module openframe_project_wrapper (por_l,
    porb_h,
    porb_l,
    resetb_h,
    resetb_l,
    vccd1,
    vdda1,
    vssa1,
    vssio,
    vccd2,
    vddio,
    vssa2,
    vdda2,
    vdda,
    vssd1,
    vssd2,
    vccd,
    vssa,
    vssd,
    analog_io,
    analog_noesd_io,
    gpio_analog_en,
    gpio_analog_pol,
    gpio_analog_sel,
    gpio_dm0,
    gpio_dm1,
    gpio_dm2,
    gpio_holdover,
    gpio_ib_mode_sel,
    gpio_in,
    gpio_in_h,
    gpio_inp_dis,
    gpio_loopback_one,
    gpio_loopback_zero,
    gpio_oeb,
    gpio_out,
    gpio_slow_sel,
    gpio_vtrip_sel,
    mask_rev);
 input por_l;
 input porb_h;
 input porb_l;
 input resetb_h;
 input resetb_l;
 input vccd1;
 input vdda1;
 input vssa1;
 input vssio;
 input vccd2;
 input vddio;
 input vssa2;
 input vdda2;
 input vdda;
 input vssd1;
 input vssd2;
 input vccd;
 input vssa;
 input vssd;
 inout [43:0] analog_io;
 inout [43:0] analog_noesd_io;
 output [43:0] gpio_analog_en;
 output [43:0] gpio_analog_pol;
 output [43:0] gpio_analog_sel;
 output [43:0] gpio_dm0;
 output [43:0] gpio_dm1;
 output [43:0] gpio_dm2;
 output [43:0] gpio_holdover;
 output [43:0] gpio_ib_mode_sel;
 input [43:0] gpio_in;
 input [43:0] gpio_in_h;
 output [43:0] gpio_inp_dis;
 input [43:0] gpio_loopback_one;
 input [43:0] gpio_loopback_zero;
 output [43:0] gpio_oeb;
 output [43:0] gpio_out;
 output [43:0] gpio_slow_sel;
 output [43:0] gpio_vtrip_sel;
 input [31:0] mask_rev;

 wire \gpio[0].gpio_I.gpio_analog_en ;
 wire \gpio[0].gpio_I.gpio_dm0 ;
 wire \top_I.branch[0].block[0].um_I.ana[0] ;
 wire \top_I.branch[0].block[0].um_I.ana[1] ;
 wire \top_I.branch[0].block[0].um_I.ana[2] ;
 wire \top_I.branch[0].block[0].um_I.ana[3] ;
 wire \top_I.branch[0].block[0].um_I.ana[4] ;
 wire \top_I.branch[0].block[0].um_I.ana[5] ;
 wire \top_I.branch[0].block[0].um_I.ana[6] ;
 wire \top_I.branch[0].block[0].um_I.ana[7] ;
 wire \top_I.branch[0].block[0].um_I.clk ;
 wire \top_I.branch[0].block[0].um_I.ena ;
 wire \top_I.branch[0].block[0].um_I.iw[10] ;
 wire \top_I.branch[0].block[0].um_I.iw[11] ;
 wire \top_I.branch[0].block[0].um_I.iw[12] ;
 wire \top_I.branch[0].block[0].um_I.iw[13] ;
 wire \top_I.branch[0].block[0].um_I.iw[14] ;
 wire \top_I.branch[0].block[0].um_I.iw[15] ;
 wire \top_I.branch[0].block[0].um_I.iw[16] ;
 wire \top_I.branch[0].block[0].um_I.iw[17] ;
 wire \top_I.branch[0].block[0].um_I.iw[1] ;
 wire \top_I.branch[0].block[0].um_I.iw[2] ;
 wire \top_I.branch[0].block[0].um_I.iw[3] ;
 wire \top_I.branch[0].block[0].um_I.iw[4] ;
 wire \top_I.branch[0].block[0].um_I.iw[5] ;
 wire \top_I.branch[0].block[0].um_I.iw[6] ;
 wire \top_I.branch[0].block[0].um_I.iw[7] ;
 wire \top_I.branch[0].block[0].um_I.iw[8] ;
 wire \top_I.branch[0].block[0].um_I.iw[9] ;
 wire \top_I.branch[0].block[0].um_I.k_zero ;
 wire \top_I.branch[0].block[0].um_I.ow[0] ;
 wire \top_I.branch[0].block[0].um_I.ow[10] ;
 wire \top_I.branch[0].block[0].um_I.ow[11] ;
 wire \top_I.branch[0].block[0].um_I.ow[12] ;
 wire \top_I.branch[0].block[0].um_I.ow[13] ;
 wire \top_I.branch[0].block[0].um_I.ow[14] ;
 wire \top_I.branch[0].block[0].um_I.ow[15] ;
 wire \top_I.branch[0].block[0].um_I.ow[16] ;
 wire \top_I.branch[0].block[0].um_I.ow[17] ;
 wire \top_I.branch[0].block[0].um_I.ow[18] ;
 wire \top_I.branch[0].block[0].um_I.ow[19] ;
 wire \top_I.branch[0].block[0].um_I.ow[1] ;
 wire \top_I.branch[0].block[0].um_I.ow[20] ;
 wire \top_I.branch[0].block[0].um_I.ow[21] ;
 wire \top_I.branch[0].block[0].um_I.ow[22] ;
 wire \top_I.branch[0].block[0].um_I.ow[23] ;
 wire \top_I.branch[0].block[0].um_I.ow[2] ;
 wire \top_I.branch[0].block[0].um_I.ow[3] ;
 wire \top_I.branch[0].block[0].um_I.ow[4] ;
 wire \top_I.branch[0].block[0].um_I.ow[5] ;
 wire \top_I.branch[0].block[0].um_I.ow[6] ;
 wire \top_I.branch[0].block[0].um_I.ow[7] ;
 wire \top_I.branch[0].block[0].um_I.ow[8] ;
 wire \top_I.branch[0].block[0].um_I.ow[9] ;
 wire \top_I.branch[0].block[0].um_I.pg_vdd ;
 wire \top_I.branch[0].block[10].um_I.ana[0] ;
 wire \top_I.branch[0].block[10].um_I.ana[1] ;
 wire \top_I.branch[0].block[10].um_I.ana[2] ;
 wire \top_I.branch[0].block[10].um_I.ana[3] ;
 wire \top_I.branch[0].block[10].um_I.ana[4] ;
 wire \top_I.branch[0].block[10].um_I.ana[5] ;
 wire \top_I.branch[0].block[10].um_I.ana[6] ;
 wire \top_I.branch[0].block[10].um_I.ana[7] ;
 wire \top_I.branch[0].block[10].um_I.clk ;
 wire \top_I.branch[0].block[10].um_I.ena ;
 wire \top_I.branch[0].block[10].um_I.iw[10] ;
 wire \top_I.branch[0].block[10].um_I.iw[11] ;
 wire \top_I.branch[0].block[10].um_I.iw[12] ;
 wire \top_I.branch[0].block[10].um_I.iw[13] ;
 wire \top_I.branch[0].block[10].um_I.iw[14] ;
 wire \top_I.branch[0].block[10].um_I.iw[15] ;
 wire \top_I.branch[0].block[10].um_I.iw[16] ;
 wire \top_I.branch[0].block[10].um_I.iw[17] ;
 wire \top_I.branch[0].block[10].um_I.iw[1] ;
 wire \top_I.branch[0].block[10].um_I.iw[2] ;
 wire \top_I.branch[0].block[10].um_I.iw[3] ;
 wire \top_I.branch[0].block[10].um_I.iw[4] ;
 wire \top_I.branch[0].block[10].um_I.iw[5] ;
 wire \top_I.branch[0].block[10].um_I.iw[6] ;
 wire \top_I.branch[0].block[10].um_I.iw[7] ;
 wire \top_I.branch[0].block[10].um_I.iw[8] ;
 wire \top_I.branch[0].block[10].um_I.iw[9] ;
 wire \top_I.branch[0].block[10].um_I.k_zero ;
 wire \top_I.branch[0].block[10].um_I.pg_vdd ;
 wire \top_I.branch[0].block[11].um_I.ana[0] ;
 wire \top_I.branch[0].block[11].um_I.ana[1] ;
 wire \top_I.branch[0].block[11].um_I.ana[2] ;
 wire \top_I.branch[0].block[11].um_I.ana[3] ;
 wire \top_I.branch[0].block[11].um_I.ana[4] ;
 wire \top_I.branch[0].block[11].um_I.ana[5] ;
 wire \top_I.branch[0].block[11].um_I.ana[6] ;
 wire \top_I.branch[0].block[11].um_I.ana[7] ;
 wire \top_I.branch[0].block[11].um_I.clk ;
 wire \top_I.branch[0].block[11].um_I.ena ;
 wire \top_I.branch[0].block[11].um_I.iw[10] ;
 wire \top_I.branch[0].block[11].um_I.iw[11] ;
 wire \top_I.branch[0].block[11].um_I.iw[12] ;
 wire \top_I.branch[0].block[11].um_I.iw[13] ;
 wire \top_I.branch[0].block[11].um_I.iw[14] ;
 wire \top_I.branch[0].block[11].um_I.iw[15] ;
 wire \top_I.branch[0].block[11].um_I.iw[16] ;
 wire \top_I.branch[0].block[11].um_I.iw[17] ;
 wire \top_I.branch[0].block[11].um_I.iw[1] ;
 wire \top_I.branch[0].block[11].um_I.iw[2] ;
 wire \top_I.branch[0].block[11].um_I.iw[3] ;
 wire \top_I.branch[0].block[11].um_I.iw[4] ;
 wire \top_I.branch[0].block[11].um_I.iw[5] ;
 wire \top_I.branch[0].block[11].um_I.iw[6] ;
 wire \top_I.branch[0].block[11].um_I.iw[7] ;
 wire \top_I.branch[0].block[11].um_I.iw[8] ;
 wire \top_I.branch[0].block[11].um_I.iw[9] ;
 wire \top_I.branch[0].block[11].um_I.k_zero ;
 wire \top_I.branch[0].block[11].um_I.pg_vdd ;
 wire \top_I.branch[0].block[12].um_I.ana[0] ;
 wire \top_I.branch[0].block[12].um_I.ana[1] ;
 wire \top_I.branch[0].block[12].um_I.ana[2] ;
 wire \top_I.branch[0].block[12].um_I.ana[3] ;
 wire \top_I.branch[0].block[12].um_I.ana[4] ;
 wire \top_I.branch[0].block[12].um_I.ana[5] ;
 wire \top_I.branch[0].block[12].um_I.ana[6] ;
 wire \top_I.branch[0].block[12].um_I.ana[7] ;
 wire \top_I.branch[0].block[12].um_I.clk ;
 wire \top_I.branch[0].block[12].um_I.ena ;
 wire \top_I.branch[0].block[12].um_I.iw[10] ;
 wire \top_I.branch[0].block[12].um_I.iw[11] ;
 wire \top_I.branch[0].block[12].um_I.iw[12] ;
 wire \top_I.branch[0].block[12].um_I.iw[13] ;
 wire \top_I.branch[0].block[12].um_I.iw[14] ;
 wire \top_I.branch[0].block[12].um_I.iw[15] ;
 wire \top_I.branch[0].block[12].um_I.iw[16] ;
 wire \top_I.branch[0].block[12].um_I.iw[17] ;
 wire \top_I.branch[0].block[12].um_I.iw[1] ;
 wire \top_I.branch[0].block[12].um_I.iw[2] ;
 wire \top_I.branch[0].block[12].um_I.iw[3] ;
 wire \top_I.branch[0].block[12].um_I.iw[4] ;
 wire \top_I.branch[0].block[12].um_I.iw[5] ;
 wire \top_I.branch[0].block[12].um_I.iw[6] ;
 wire \top_I.branch[0].block[12].um_I.iw[7] ;
 wire \top_I.branch[0].block[12].um_I.iw[8] ;
 wire \top_I.branch[0].block[12].um_I.iw[9] ;
 wire \top_I.branch[0].block[12].um_I.k_zero ;
 wire \top_I.branch[0].block[12].um_I.pg_vdd ;
 wire \top_I.branch[0].block[13].um_I.ana[0] ;
 wire \top_I.branch[0].block[13].um_I.ana[1] ;
 wire \top_I.branch[0].block[13].um_I.ana[2] ;
 wire \top_I.branch[0].block[13].um_I.ana[3] ;
 wire \top_I.branch[0].block[13].um_I.ana[4] ;
 wire \top_I.branch[0].block[13].um_I.ana[5] ;
 wire \top_I.branch[0].block[13].um_I.ana[6] ;
 wire \top_I.branch[0].block[13].um_I.ana[7] ;
 wire \top_I.branch[0].block[13].um_I.clk ;
 wire \top_I.branch[0].block[13].um_I.ena ;
 wire \top_I.branch[0].block[13].um_I.iw[10] ;
 wire \top_I.branch[0].block[13].um_I.iw[11] ;
 wire \top_I.branch[0].block[13].um_I.iw[12] ;
 wire \top_I.branch[0].block[13].um_I.iw[13] ;
 wire \top_I.branch[0].block[13].um_I.iw[14] ;
 wire \top_I.branch[0].block[13].um_I.iw[15] ;
 wire \top_I.branch[0].block[13].um_I.iw[16] ;
 wire \top_I.branch[0].block[13].um_I.iw[17] ;
 wire \top_I.branch[0].block[13].um_I.iw[1] ;
 wire \top_I.branch[0].block[13].um_I.iw[2] ;
 wire \top_I.branch[0].block[13].um_I.iw[3] ;
 wire \top_I.branch[0].block[13].um_I.iw[4] ;
 wire \top_I.branch[0].block[13].um_I.iw[5] ;
 wire \top_I.branch[0].block[13].um_I.iw[6] ;
 wire \top_I.branch[0].block[13].um_I.iw[7] ;
 wire \top_I.branch[0].block[13].um_I.iw[8] ;
 wire \top_I.branch[0].block[13].um_I.iw[9] ;
 wire \top_I.branch[0].block[13].um_I.k_zero ;
 wire \top_I.branch[0].block[13].um_I.pg_vdd ;
 wire \top_I.branch[0].block[14].um_I.ana[0] ;
 wire \top_I.branch[0].block[14].um_I.ana[1] ;
 wire \top_I.branch[0].block[14].um_I.ana[2] ;
 wire \top_I.branch[0].block[14].um_I.ana[3] ;
 wire \top_I.branch[0].block[14].um_I.ana[4] ;
 wire \top_I.branch[0].block[14].um_I.ana[5] ;
 wire \top_I.branch[0].block[14].um_I.ana[6] ;
 wire \top_I.branch[0].block[14].um_I.ana[7] ;
 wire \top_I.branch[0].block[14].um_I.clk ;
 wire \top_I.branch[0].block[14].um_I.ena ;
 wire \top_I.branch[0].block[14].um_I.iw[10] ;
 wire \top_I.branch[0].block[14].um_I.iw[11] ;
 wire \top_I.branch[0].block[14].um_I.iw[12] ;
 wire \top_I.branch[0].block[14].um_I.iw[13] ;
 wire \top_I.branch[0].block[14].um_I.iw[14] ;
 wire \top_I.branch[0].block[14].um_I.iw[15] ;
 wire \top_I.branch[0].block[14].um_I.iw[16] ;
 wire \top_I.branch[0].block[14].um_I.iw[17] ;
 wire \top_I.branch[0].block[14].um_I.iw[1] ;
 wire \top_I.branch[0].block[14].um_I.iw[2] ;
 wire \top_I.branch[0].block[14].um_I.iw[3] ;
 wire \top_I.branch[0].block[14].um_I.iw[4] ;
 wire \top_I.branch[0].block[14].um_I.iw[5] ;
 wire \top_I.branch[0].block[14].um_I.iw[6] ;
 wire \top_I.branch[0].block[14].um_I.iw[7] ;
 wire \top_I.branch[0].block[14].um_I.iw[8] ;
 wire \top_I.branch[0].block[14].um_I.iw[9] ;
 wire \top_I.branch[0].block[14].um_I.k_zero ;
 wire \top_I.branch[0].block[14].um_I.pg_vdd ;
 wire \top_I.branch[0].block[15].um_I.ana[0] ;
 wire \top_I.branch[0].block[15].um_I.ana[1] ;
 wire \top_I.branch[0].block[15].um_I.ana[2] ;
 wire \top_I.branch[0].block[15].um_I.ana[3] ;
 wire \top_I.branch[0].block[15].um_I.ana[4] ;
 wire \top_I.branch[0].block[15].um_I.ana[5] ;
 wire \top_I.branch[0].block[15].um_I.ana[6] ;
 wire \top_I.branch[0].block[15].um_I.ana[7] ;
 wire \top_I.branch[0].block[15].um_I.clk ;
 wire \top_I.branch[0].block[15].um_I.ena ;
 wire \top_I.branch[0].block[15].um_I.iw[10] ;
 wire \top_I.branch[0].block[15].um_I.iw[11] ;
 wire \top_I.branch[0].block[15].um_I.iw[12] ;
 wire \top_I.branch[0].block[15].um_I.iw[13] ;
 wire \top_I.branch[0].block[15].um_I.iw[14] ;
 wire \top_I.branch[0].block[15].um_I.iw[15] ;
 wire \top_I.branch[0].block[15].um_I.iw[16] ;
 wire \top_I.branch[0].block[15].um_I.iw[17] ;
 wire \top_I.branch[0].block[15].um_I.iw[1] ;
 wire \top_I.branch[0].block[15].um_I.iw[2] ;
 wire \top_I.branch[0].block[15].um_I.iw[3] ;
 wire \top_I.branch[0].block[15].um_I.iw[4] ;
 wire \top_I.branch[0].block[15].um_I.iw[5] ;
 wire \top_I.branch[0].block[15].um_I.iw[6] ;
 wire \top_I.branch[0].block[15].um_I.iw[7] ;
 wire \top_I.branch[0].block[15].um_I.iw[8] ;
 wire \top_I.branch[0].block[15].um_I.iw[9] ;
 wire \top_I.branch[0].block[15].um_I.k_zero ;
 wire \top_I.branch[0].block[15].um_I.pg_vdd ;
 wire \top_I.branch[0].block[1].um_I.ana[0] ;
 wire \top_I.branch[0].block[1].um_I.ana[1] ;
 wire \top_I.branch[0].block[1].um_I.ana[2] ;
 wire \top_I.branch[0].block[1].um_I.ana[3] ;
 wire \top_I.branch[0].block[1].um_I.ana[4] ;
 wire \top_I.branch[0].block[1].um_I.ana[5] ;
 wire \top_I.branch[0].block[1].um_I.ana[6] ;
 wire \top_I.branch[0].block[1].um_I.ana[7] ;
 wire \top_I.branch[0].block[1].um_I.clk ;
 wire \top_I.branch[0].block[1].um_I.ena ;
 wire \top_I.branch[0].block[1].um_I.iw[10] ;
 wire \top_I.branch[0].block[1].um_I.iw[11] ;
 wire \top_I.branch[0].block[1].um_I.iw[12] ;
 wire \top_I.branch[0].block[1].um_I.iw[13] ;
 wire \top_I.branch[0].block[1].um_I.iw[14] ;
 wire \top_I.branch[0].block[1].um_I.iw[15] ;
 wire \top_I.branch[0].block[1].um_I.iw[16] ;
 wire \top_I.branch[0].block[1].um_I.iw[17] ;
 wire \top_I.branch[0].block[1].um_I.iw[1] ;
 wire \top_I.branch[0].block[1].um_I.iw[2] ;
 wire \top_I.branch[0].block[1].um_I.iw[3] ;
 wire \top_I.branch[0].block[1].um_I.iw[4] ;
 wire \top_I.branch[0].block[1].um_I.iw[5] ;
 wire \top_I.branch[0].block[1].um_I.iw[6] ;
 wire \top_I.branch[0].block[1].um_I.iw[7] ;
 wire \top_I.branch[0].block[1].um_I.iw[8] ;
 wire \top_I.branch[0].block[1].um_I.iw[9] ;
 wire \top_I.branch[0].block[1].um_I.k_zero ;
 wire \top_I.branch[0].block[1].um_I.ow[0] ;
 wire \top_I.branch[0].block[1].um_I.ow[10] ;
 wire \top_I.branch[0].block[1].um_I.ow[11] ;
 wire \top_I.branch[0].block[1].um_I.ow[12] ;
 wire \top_I.branch[0].block[1].um_I.ow[13] ;
 wire \top_I.branch[0].block[1].um_I.ow[14] ;
 wire \top_I.branch[0].block[1].um_I.ow[15] ;
 wire \top_I.branch[0].block[1].um_I.ow[16] ;
 wire \top_I.branch[0].block[1].um_I.ow[17] ;
 wire \top_I.branch[0].block[1].um_I.ow[18] ;
 wire \top_I.branch[0].block[1].um_I.ow[19] ;
 wire \top_I.branch[0].block[1].um_I.ow[1] ;
 wire \top_I.branch[0].block[1].um_I.ow[20] ;
 wire \top_I.branch[0].block[1].um_I.ow[21] ;
 wire \top_I.branch[0].block[1].um_I.ow[22] ;
 wire \top_I.branch[0].block[1].um_I.ow[23] ;
 wire \top_I.branch[0].block[1].um_I.ow[2] ;
 wire \top_I.branch[0].block[1].um_I.ow[3] ;
 wire \top_I.branch[0].block[1].um_I.ow[4] ;
 wire \top_I.branch[0].block[1].um_I.ow[5] ;
 wire \top_I.branch[0].block[1].um_I.ow[6] ;
 wire \top_I.branch[0].block[1].um_I.ow[7] ;
 wire \top_I.branch[0].block[1].um_I.ow[8] ;
 wire \top_I.branch[0].block[1].um_I.ow[9] ;
 wire \top_I.branch[0].block[1].um_I.pg_vdd ;
 wire \top_I.branch[0].block[2].um_I.ana[0] ;
 wire \top_I.branch[0].block[2].um_I.ana[1] ;
 wire \top_I.branch[0].block[2].um_I.ana[2] ;
 wire \top_I.branch[0].block[2].um_I.ana[3] ;
 wire \top_I.branch[0].block[2].um_I.ana[4] ;
 wire \top_I.branch[0].block[2].um_I.ana[5] ;
 wire \top_I.branch[0].block[2].um_I.ana[6] ;
 wire \top_I.branch[0].block[2].um_I.ana[7] ;
 wire \top_I.branch[0].block[2].um_I.clk ;
 wire \top_I.branch[0].block[2].um_I.ena ;
 wire \top_I.branch[0].block[2].um_I.iw[10] ;
 wire \top_I.branch[0].block[2].um_I.iw[11] ;
 wire \top_I.branch[0].block[2].um_I.iw[12] ;
 wire \top_I.branch[0].block[2].um_I.iw[13] ;
 wire \top_I.branch[0].block[2].um_I.iw[14] ;
 wire \top_I.branch[0].block[2].um_I.iw[15] ;
 wire \top_I.branch[0].block[2].um_I.iw[16] ;
 wire \top_I.branch[0].block[2].um_I.iw[17] ;
 wire \top_I.branch[0].block[2].um_I.iw[1] ;
 wire \top_I.branch[0].block[2].um_I.iw[2] ;
 wire \top_I.branch[0].block[2].um_I.iw[3] ;
 wire \top_I.branch[0].block[2].um_I.iw[4] ;
 wire \top_I.branch[0].block[2].um_I.iw[5] ;
 wire \top_I.branch[0].block[2].um_I.iw[6] ;
 wire \top_I.branch[0].block[2].um_I.iw[7] ;
 wire \top_I.branch[0].block[2].um_I.iw[8] ;
 wire \top_I.branch[0].block[2].um_I.iw[9] ;
 wire \top_I.branch[0].block[2].um_I.k_zero ;
 wire \top_I.branch[0].block[2].um_I.pg_vdd ;
 wire \top_I.branch[0].block[3].um_I.ana[0] ;
 wire \top_I.branch[0].block[3].um_I.ana[1] ;
 wire \top_I.branch[0].block[3].um_I.ana[2] ;
 wire \top_I.branch[0].block[3].um_I.ana[3] ;
 wire \top_I.branch[0].block[3].um_I.ana[4] ;
 wire \top_I.branch[0].block[3].um_I.ana[5] ;
 wire \top_I.branch[0].block[3].um_I.ana[6] ;
 wire \top_I.branch[0].block[3].um_I.ana[7] ;
 wire \top_I.branch[0].block[3].um_I.clk ;
 wire \top_I.branch[0].block[3].um_I.ena ;
 wire \top_I.branch[0].block[3].um_I.iw[10] ;
 wire \top_I.branch[0].block[3].um_I.iw[11] ;
 wire \top_I.branch[0].block[3].um_I.iw[12] ;
 wire \top_I.branch[0].block[3].um_I.iw[13] ;
 wire \top_I.branch[0].block[3].um_I.iw[14] ;
 wire \top_I.branch[0].block[3].um_I.iw[15] ;
 wire \top_I.branch[0].block[3].um_I.iw[16] ;
 wire \top_I.branch[0].block[3].um_I.iw[17] ;
 wire \top_I.branch[0].block[3].um_I.iw[1] ;
 wire \top_I.branch[0].block[3].um_I.iw[2] ;
 wire \top_I.branch[0].block[3].um_I.iw[3] ;
 wire \top_I.branch[0].block[3].um_I.iw[4] ;
 wire \top_I.branch[0].block[3].um_I.iw[5] ;
 wire \top_I.branch[0].block[3].um_I.iw[6] ;
 wire \top_I.branch[0].block[3].um_I.iw[7] ;
 wire \top_I.branch[0].block[3].um_I.iw[8] ;
 wire \top_I.branch[0].block[3].um_I.iw[9] ;
 wire \top_I.branch[0].block[3].um_I.k_zero ;
 wire \top_I.branch[0].block[3].um_I.pg_vdd ;
 wire \top_I.branch[0].block[4].um_I.ana[0] ;
 wire \top_I.branch[0].block[4].um_I.ana[1] ;
 wire \top_I.branch[0].block[4].um_I.ana[2] ;
 wire \top_I.branch[0].block[4].um_I.ana[3] ;
 wire \top_I.branch[0].block[4].um_I.ana[4] ;
 wire \top_I.branch[0].block[4].um_I.ana[5] ;
 wire \top_I.branch[0].block[4].um_I.ana[6] ;
 wire \top_I.branch[0].block[4].um_I.ana[7] ;
 wire \top_I.branch[0].block[4].um_I.clk ;
 wire \top_I.branch[0].block[4].um_I.ena ;
 wire \top_I.branch[0].block[4].um_I.iw[10] ;
 wire \top_I.branch[0].block[4].um_I.iw[11] ;
 wire \top_I.branch[0].block[4].um_I.iw[12] ;
 wire \top_I.branch[0].block[4].um_I.iw[13] ;
 wire \top_I.branch[0].block[4].um_I.iw[14] ;
 wire \top_I.branch[0].block[4].um_I.iw[15] ;
 wire \top_I.branch[0].block[4].um_I.iw[16] ;
 wire \top_I.branch[0].block[4].um_I.iw[17] ;
 wire \top_I.branch[0].block[4].um_I.iw[1] ;
 wire \top_I.branch[0].block[4].um_I.iw[2] ;
 wire \top_I.branch[0].block[4].um_I.iw[3] ;
 wire \top_I.branch[0].block[4].um_I.iw[4] ;
 wire \top_I.branch[0].block[4].um_I.iw[5] ;
 wire \top_I.branch[0].block[4].um_I.iw[6] ;
 wire \top_I.branch[0].block[4].um_I.iw[7] ;
 wire \top_I.branch[0].block[4].um_I.iw[8] ;
 wire \top_I.branch[0].block[4].um_I.iw[9] ;
 wire \top_I.branch[0].block[4].um_I.k_zero ;
 wire \top_I.branch[0].block[4].um_I.pg_vdd ;
 wire \top_I.branch[0].block[5].um_I.ana[0] ;
 wire \top_I.branch[0].block[5].um_I.ana[1] ;
 wire \top_I.branch[0].block[5].um_I.ana[2] ;
 wire \top_I.branch[0].block[5].um_I.ana[3] ;
 wire \top_I.branch[0].block[5].um_I.ana[4] ;
 wire \top_I.branch[0].block[5].um_I.ana[5] ;
 wire \top_I.branch[0].block[5].um_I.ana[6] ;
 wire \top_I.branch[0].block[5].um_I.ana[7] ;
 wire \top_I.branch[0].block[5].um_I.clk ;
 wire \top_I.branch[0].block[5].um_I.ena ;
 wire \top_I.branch[0].block[5].um_I.iw[10] ;
 wire \top_I.branch[0].block[5].um_I.iw[11] ;
 wire \top_I.branch[0].block[5].um_I.iw[12] ;
 wire \top_I.branch[0].block[5].um_I.iw[13] ;
 wire \top_I.branch[0].block[5].um_I.iw[14] ;
 wire \top_I.branch[0].block[5].um_I.iw[15] ;
 wire \top_I.branch[0].block[5].um_I.iw[16] ;
 wire \top_I.branch[0].block[5].um_I.iw[17] ;
 wire \top_I.branch[0].block[5].um_I.iw[1] ;
 wire \top_I.branch[0].block[5].um_I.iw[2] ;
 wire \top_I.branch[0].block[5].um_I.iw[3] ;
 wire \top_I.branch[0].block[5].um_I.iw[4] ;
 wire \top_I.branch[0].block[5].um_I.iw[5] ;
 wire \top_I.branch[0].block[5].um_I.iw[6] ;
 wire \top_I.branch[0].block[5].um_I.iw[7] ;
 wire \top_I.branch[0].block[5].um_I.iw[8] ;
 wire \top_I.branch[0].block[5].um_I.iw[9] ;
 wire \top_I.branch[0].block[5].um_I.k_zero ;
 wire \top_I.branch[0].block[5].um_I.pg_vdd ;
 wire \top_I.branch[0].block[6].um_I.ana[0] ;
 wire \top_I.branch[0].block[6].um_I.ana[1] ;
 wire \top_I.branch[0].block[6].um_I.ana[2] ;
 wire \top_I.branch[0].block[6].um_I.ana[3] ;
 wire \top_I.branch[0].block[6].um_I.ana[4] ;
 wire \top_I.branch[0].block[6].um_I.ana[5] ;
 wire \top_I.branch[0].block[6].um_I.ana[6] ;
 wire \top_I.branch[0].block[6].um_I.ana[7] ;
 wire \top_I.branch[0].block[6].um_I.clk ;
 wire \top_I.branch[0].block[6].um_I.ena ;
 wire \top_I.branch[0].block[6].um_I.iw[10] ;
 wire \top_I.branch[0].block[6].um_I.iw[11] ;
 wire \top_I.branch[0].block[6].um_I.iw[12] ;
 wire \top_I.branch[0].block[6].um_I.iw[13] ;
 wire \top_I.branch[0].block[6].um_I.iw[14] ;
 wire \top_I.branch[0].block[6].um_I.iw[15] ;
 wire \top_I.branch[0].block[6].um_I.iw[16] ;
 wire \top_I.branch[0].block[6].um_I.iw[17] ;
 wire \top_I.branch[0].block[6].um_I.iw[1] ;
 wire \top_I.branch[0].block[6].um_I.iw[2] ;
 wire \top_I.branch[0].block[6].um_I.iw[3] ;
 wire \top_I.branch[0].block[6].um_I.iw[4] ;
 wire \top_I.branch[0].block[6].um_I.iw[5] ;
 wire \top_I.branch[0].block[6].um_I.iw[6] ;
 wire \top_I.branch[0].block[6].um_I.iw[7] ;
 wire \top_I.branch[0].block[6].um_I.iw[8] ;
 wire \top_I.branch[0].block[6].um_I.iw[9] ;
 wire \top_I.branch[0].block[6].um_I.k_zero ;
 wire \top_I.branch[0].block[6].um_I.pg_vdd ;
 wire \top_I.branch[0].block[7].um_I.ana[0] ;
 wire \top_I.branch[0].block[7].um_I.ana[1] ;
 wire \top_I.branch[0].block[7].um_I.ana[2] ;
 wire \top_I.branch[0].block[7].um_I.ana[3] ;
 wire \top_I.branch[0].block[7].um_I.ana[4] ;
 wire \top_I.branch[0].block[7].um_I.ana[5] ;
 wire \top_I.branch[0].block[7].um_I.ana[6] ;
 wire \top_I.branch[0].block[7].um_I.ana[7] ;
 wire \top_I.branch[0].block[7].um_I.clk ;
 wire \top_I.branch[0].block[7].um_I.ena ;
 wire \top_I.branch[0].block[7].um_I.iw[10] ;
 wire \top_I.branch[0].block[7].um_I.iw[11] ;
 wire \top_I.branch[0].block[7].um_I.iw[12] ;
 wire \top_I.branch[0].block[7].um_I.iw[13] ;
 wire \top_I.branch[0].block[7].um_I.iw[14] ;
 wire \top_I.branch[0].block[7].um_I.iw[15] ;
 wire \top_I.branch[0].block[7].um_I.iw[16] ;
 wire \top_I.branch[0].block[7].um_I.iw[17] ;
 wire \top_I.branch[0].block[7].um_I.iw[1] ;
 wire \top_I.branch[0].block[7].um_I.iw[2] ;
 wire \top_I.branch[0].block[7].um_I.iw[3] ;
 wire \top_I.branch[0].block[7].um_I.iw[4] ;
 wire \top_I.branch[0].block[7].um_I.iw[5] ;
 wire \top_I.branch[0].block[7].um_I.iw[6] ;
 wire \top_I.branch[0].block[7].um_I.iw[7] ;
 wire \top_I.branch[0].block[7].um_I.iw[8] ;
 wire \top_I.branch[0].block[7].um_I.iw[9] ;
 wire \top_I.branch[0].block[7].um_I.k_zero ;
 wire \top_I.branch[0].block[7].um_I.pg_vdd ;
 wire \top_I.branch[0].block[8].um_I.ana[0] ;
 wire \top_I.branch[0].block[8].um_I.ana[1] ;
 wire \top_I.branch[0].block[8].um_I.ana[2] ;
 wire \top_I.branch[0].block[8].um_I.ana[3] ;
 wire \top_I.branch[0].block[8].um_I.ana[4] ;
 wire \top_I.branch[0].block[8].um_I.ana[5] ;
 wire \top_I.branch[0].block[8].um_I.ana[6] ;
 wire \top_I.branch[0].block[8].um_I.ana[7] ;
 wire \top_I.branch[0].block[8].um_I.clk ;
 wire \top_I.branch[0].block[8].um_I.ena ;
 wire \top_I.branch[0].block[8].um_I.iw[10] ;
 wire \top_I.branch[0].block[8].um_I.iw[11] ;
 wire \top_I.branch[0].block[8].um_I.iw[12] ;
 wire \top_I.branch[0].block[8].um_I.iw[13] ;
 wire \top_I.branch[0].block[8].um_I.iw[14] ;
 wire \top_I.branch[0].block[8].um_I.iw[15] ;
 wire \top_I.branch[0].block[8].um_I.iw[16] ;
 wire \top_I.branch[0].block[8].um_I.iw[17] ;
 wire \top_I.branch[0].block[8].um_I.iw[1] ;
 wire \top_I.branch[0].block[8].um_I.iw[2] ;
 wire \top_I.branch[0].block[8].um_I.iw[3] ;
 wire \top_I.branch[0].block[8].um_I.iw[4] ;
 wire \top_I.branch[0].block[8].um_I.iw[5] ;
 wire \top_I.branch[0].block[8].um_I.iw[6] ;
 wire \top_I.branch[0].block[8].um_I.iw[7] ;
 wire \top_I.branch[0].block[8].um_I.iw[8] ;
 wire \top_I.branch[0].block[8].um_I.iw[9] ;
 wire \top_I.branch[0].block[8].um_I.k_zero ;
 wire \top_I.branch[0].block[8].um_I.pg_vdd ;
 wire \top_I.branch[0].block[9].um_I.ana[0] ;
 wire \top_I.branch[0].block[9].um_I.ana[1] ;
 wire \top_I.branch[0].block[9].um_I.ana[2] ;
 wire \top_I.branch[0].block[9].um_I.ana[3] ;
 wire \top_I.branch[0].block[9].um_I.ana[4] ;
 wire \top_I.branch[0].block[9].um_I.ana[5] ;
 wire \top_I.branch[0].block[9].um_I.ana[6] ;
 wire \top_I.branch[0].block[9].um_I.ana[7] ;
 wire \top_I.branch[0].block[9].um_I.clk ;
 wire \top_I.branch[0].block[9].um_I.ena ;
 wire \top_I.branch[0].block[9].um_I.iw[10] ;
 wire \top_I.branch[0].block[9].um_I.iw[11] ;
 wire \top_I.branch[0].block[9].um_I.iw[12] ;
 wire \top_I.branch[0].block[9].um_I.iw[13] ;
 wire \top_I.branch[0].block[9].um_I.iw[14] ;
 wire \top_I.branch[0].block[9].um_I.iw[15] ;
 wire \top_I.branch[0].block[9].um_I.iw[16] ;
 wire \top_I.branch[0].block[9].um_I.iw[17] ;
 wire \top_I.branch[0].block[9].um_I.iw[1] ;
 wire \top_I.branch[0].block[9].um_I.iw[2] ;
 wire \top_I.branch[0].block[9].um_I.iw[3] ;
 wire \top_I.branch[0].block[9].um_I.iw[4] ;
 wire \top_I.branch[0].block[9].um_I.iw[5] ;
 wire \top_I.branch[0].block[9].um_I.iw[6] ;
 wire \top_I.branch[0].block[9].um_I.iw[7] ;
 wire \top_I.branch[0].block[9].um_I.iw[8] ;
 wire \top_I.branch[0].block[9].um_I.iw[9] ;
 wire \top_I.branch[0].block[9].um_I.k_zero ;
 wire \top_I.branch[0].block[9].um_I.pg_vdd ;
 wire \top_I.branch[0].l_addr[0] ;
 wire \top_I.branch[0].l_k_one ;
 wire \top_I.branch[0].l_spine_iw[0] ;
 wire \top_I.branch[0].l_spine_iw[10] ;
 wire \top_I.branch[0].l_spine_iw[11] ;
 wire \top_I.branch[0].l_spine_iw[12] ;
 wire \top_I.branch[0].l_spine_iw[13] ;
 wire \top_I.branch[0].l_spine_iw[14] ;
 wire \top_I.branch[0].l_spine_iw[15] ;
 wire \top_I.branch[0].l_spine_iw[16] ;
 wire \top_I.branch[0].l_spine_iw[17] ;
 wire \top_I.branch[0].l_spine_iw[18] ;
 wire \top_I.branch[0].l_spine_iw[19] ;
 wire \top_I.branch[0].l_spine_iw[1] ;
 wire \top_I.branch[0].l_spine_iw[20] ;
 wire \top_I.branch[0].l_spine_iw[21] ;
 wire \top_I.branch[0].l_spine_iw[22] ;
 wire \top_I.branch[0].l_spine_iw[23] ;
 wire \top_I.branch[0].l_spine_iw[24] ;
 wire \top_I.branch[0].l_spine_iw[25] ;
 wire \top_I.branch[0].l_spine_iw[26] ;
 wire \top_I.branch[0].l_spine_iw[27] ;
 wire \top_I.branch[0].l_spine_iw[28] ;
 wire \top_I.branch[0].l_spine_iw[29] ;
 wire \top_I.branch[0].l_spine_iw[2] ;
 wire \top_I.branch[0].l_spine_iw[3] ;
 wire \top_I.branch[0].l_spine_iw[4] ;
 wire \top_I.branch[0].l_spine_iw[5] ;
 wire \top_I.branch[0].l_spine_iw[6] ;
 wire \top_I.branch[0].l_spine_iw[7] ;
 wire \top_I.branch[0].l_spine_iw[8] ;
 wire \top_I.branch[0].l_spine_iw[9] ;
 wire \top_I.branch[0].l_spine_ow[0] ;
 wire \top_I.branch[0].l_spine_ow[10] ;
 wire \top_I.branch[0].l_spine_ow[11] ;
 wire \top_I.branch[0].l_spine_ow[12] ;
 wire \top_I.branch[0].l_spine_ow[13] ;
 wire \top_I.branch[0].l_spine_ow[14] ;
 wire \top_I.branch[0].l_spine_ow[15] ;
 wire \top_I.branch[0].l_spine_ow[16] ;
 wire \top_I.branch[0].l_spine_ow[17] ;
 wire \top_I.branch[0].l_spine_ow[18] ;
 wire \top_I.branch[0].l_spine_ow[19] ;
 wire \top_I.branch[0].l_spine_ow[1] ;
 wire \top_I.branch[0].l_spine_ow[20] ;
 wire \top_I.branch[0].l_spine_ow[21] ;
 wire \top_I.branch[0].l_spine_ow[22] ;
 wire \top_I.branch[0].l_spine_ow[23] ;
 wire \top_I.branch[0].l_spine_ow[24] ;
 wire \top_I.branch[0].l_spine_ow[25] ;
 wire \top_I.branch[0].l_spine_ow[2] ;
 wire \top_I.branch[0].l_spine_ow[3] ;
 wire \top_I.branch[0].l_spine_ow[4] ;
 wire \top_I.branch[0].l_spine_ow[5] ;
 wire \top_I.branch[0].l_spine_ow[6] ;
 wire \top_I.branch[0].l_spine_ow[7] ;
 wire \top_I.branch[0].l_spine_ow[8] ;
 wire \top_I.branch[0].l_spine_ow[9] ;
 wire \top_I.branch[10].block[0].um_I.ana[0] ;
 wire \top_I.branch[10].block[0].um_I.ana[1] ;
 wire \top_I.branch[10].block[0].um_I.ana[2] ;
 wire \top_I.branch[10].block[0].um_I.ana[3] ;
 wire \top_I.branch[10].block[0].um_I.ana[4] ;
 wire \top_I.branch[10].block[0].um_I.ana[5] ;
 wire \top_I.branch[10].block[0].um_I.ana[6] ;
 wire \top_I.branch[10].block[0].um_I.ana[7] ;
 wire \top_I.branch[10].block[0].um_I.clk ;
 wire \top_I.branch[10].block[0].um_I.ena ;
 wire \top_I.branch[10].block[0].um_I.iw[10] ;
 wire \top_I.branch[10].block[0].um_I.iw[11] ;
 wire \top_I.branch[10].block[0].um_I.iw[12] ;
 wire \top_I.branch[10].block[0].um_I.iw[13] ;
 wire \top_I.branch[10].block[0].um_I.iw[14] ;
 wire \top_I.branch[10].block[0].um_I.iw[15] ;
 wire \top_I.branch[10].block[0].um_I.iw[16] ;
 wire \top_I.branch[10].block[0].um_I.iw[17] ;
 wire \top_I.branch[10].block[0].um_I.iw[1] ;
 wire \top_I.branch[10].block[0].um_I.iw[2] ;
 wire \top_I.branch[10].block[0].um_I.iw[3] ;
 wire \top_I.branch[10].block[0].um_I.iw[4] ;
 wire \top_I.branch[10].block[0].um_I.iw[5] ;
 wire \top_I.branch[10].block[0].um_I.iw[6] ;
 wire \top_I.branch[10].block[0].um_I.iw[7] ;
 wire \top_I.branch[10].block[0].um_I.iw[8] ;
 wire \top_I.branch[10].block[0].um_I.iw[9] ;
 wire \top_I.branch[10].block[0].um_I.k_zero ;
 wire \top_I.branch[10].block[0].um_I.pg_vdd ;
 wire \top_I.branch[10].block[10].um_I.ana[0] ;
 wire \top_I.branch[10].block[10].um_I.ana[1] ;
 wire \top_I.branch[10].block[10].um_I.ana[2] ;
 wire \top_I.branch[10].block[10].um_I.ana[3] ;
 wire \top_I.branch[10].block[10].um_I.ana[4] ;
 wire \top_I.branch[10].block[10].um_I.ana[5] ;
 wire \top_I.branch[10].block[10].um_I.ana[6] ;
 wire \top_I.branch[10].block[10].um_I.ana[7] ;
 wire \top_I.branch[10].block[10].um_I.clk ;
 wire \top_I.branch[10].block[10].um_I.ena ;
 wire \top_I.branch[10].block[10].um_I.iw[10] ;
 wire \top_I.branch[10].block[10].um_I.iw[11] ;
 wire \top_I.branch[10].block[10].um_I.iw[12] ;
 wire \top_I.branch[10].block[10].um_I.iw[13] ;
 wire \top_I.branch[10].block[10].um_I.iw[14] ;
 wire \top_I.branch[10].block[10].um_I.iw[15] ;
 wire \top_I.branch[10].block[10].um_I.iw[16] ;
 wire \top_I.branch[10].block[10].um_I.iw[17] ;
 wire \top_I.branch[10].block[10].um_I.iw[1] ;
 wire \top_I.branch[10].block[10].um_I.iw[2] ;
 wire \top_I.branch[10].block[10].um_I.iw[3] ;
 wire \top_I.branch[10].block[10].um_I.iw[4] ;
 wire \top_I.branch[10].block[10].um_I.iw[5] ;
 wire \top_I.branch[10].block[10].um_I.iw[6] ;
 wire \top_I.branch[10].block[10].um_I.iw[7] ;
 wire \top_I.branch[10].block[10].um_I.iw[8] ;
 wire \top_I.branch[10].block[10].um_I.iw[9] ;
 wire \top_I.branch[10].block[10].um_I.k_zero ;
 wire \top_I.branch[10].block[10].um_I.pg_vdd ;
 wire \top_I.branch[10].block[11].um_I.ana[0] ;
 wire \top_I.branch[10].block[11].um_I.ana[1] ;
 wire \top_I.branch[10].block[11].um_I.ana[2] ;
 wire \top_I.branch[10].block[11].um_I.ana[3] ;
 wire \top_I.branch[10].block[11].um_I.ana[4] ;
 wire \top_I.branch[10].block[11].um_I.ana[5] ;
 wire \top_I.branch[10].block[11].um_I.ana[6] ;
 wire \top_I.branch[10].block[11].um_I.ana[7] ;
 wire \top_I.branch[10].block[11].um_I.clk ;
 wire \top_I.branch[10].block[11].um_I.ena ;
 wire \top_I.branch[10].block[11].um_I.iw[10] ;
 wire \top_I.branch[10].block[11].um_I.iw[11] ;
 wire \top_I.branch[10].block[11].um_I.iw[12] ;
 wire \top_I.branch[10].block[11].um_I.iw[13] ;
 wire \top_I.branch[10].block[11].um_I.iw[14] ;
 wire \top_I.branch[10].block[11].um_I.iw[15] ;
 wire \top_I.branch[10].block[11].um_I.iw[16] ;
 wire \top_I.branch[10].block[11].um_I.iw[17] ;
 wire \top_I.branch[10].block[11].um_I.iw[1] ;
 wire \top_I.branch[10].block[11].um_I.iw[2] ;
 wire \top_I.branch[10].block[11].um_I.iw[3] ;
 wire \top_I.branch[10].block[11].um_I.iw[4] ;
 wire \top_I.branch[10].block[11].um_I.iw[5] ;
 wire \top_I.branch[10].block[11].um_I.iw[6] ;
 wire \top_I.branch[10].block[11].um_I.iw[7] ;
 wire \top_I.branch[10].block[11].um_I.iw[8] ;
 wire \top_I.branch[10].block[11].um_I.iw[9] ;
 wire \top_I.branch[10].block[11].um_I.k_zero ;
 wire \top_I.branch[10].block[11].um_I.pg_vdd ;
 wire \top_I.branch[10].block[12].um_I.ana[0] ;
 wire \top_I.branch[10].block[12].um_I.ana[1] ;
 wire \top_I.branch[10].block[12].um_I.ana[2] ;
 wire \top_I.branch[10].block[12].um_I.ana[3] ;
 wire \top_I.branch[10].block[12].um_I.ana[4] ;
 wire \top_I.branch[10].block[12].um_I.ana[5] ;
 wire \top_I.branch[10].block[12].um_I.ana[6] ;
 wire \top_I.branch[10].block[12].um_I.ana[7] ;
 wire \top_I.branch[10].block[12].um_I.clk ;
 wire \top_I.branch[10].block[12].um_I.ena ;
 wire \top_I.branch[10].block[12].um_I.iw[10] ;
 wire \top_I.branch[10].block[12].um_I.iw[11] ;
 wire \top_I.branch[10].block[12].um_I.iw[12] ;
 wire \top_I.branch[10].block[12].um_I.iw[13] ;
 wire \top_I.branch[10].block[12].um_I.iw[14] ;
 wire \top_I.branch[10].block[12].um_I.iw[15] ;
 wire \top_I.branch[10].block[12].um_I.iw[16] ;
 wire \top_I.branch[10].block[12].um_I.iw[17] ;
 wire \top_I.branch[10].block[12].um_I.iw[1] ;
 wire \top_I.branch[10].block[12].um_I.iw[2] ;
 wire \top_I.branch[10].block[12].um_I.iw[3] ;
 wire \top_I.branch[10].block[12].um_I.iw[4] ;
 wire \top_I.branch[10].block[12].um_I.iw[5] ;
 wire \top_I.branch[10].block[12].um_I.iw[6] ;
 wire \top_I.branch[10].block[12].um_I.iw[7] ;
 wire \top_I.branch[10].block[12].um_I.iw[8] ;
 wire \top_I.branch[10].block[12].um_I.iw[9] ;
 wire \top_I.branch[10].block[12].um_I.k_zero ;
 wire \top_I.branch[10].block[12].um_I.pg_vdd ;
 wire \top_I.branch[10].block[13].um_I.ana[0] ;
 wire \top_I.branch[10].block[13].um_I.ana[1] ;
 wire \top_I.branch[10].block[13].um_I.ana[2] ;
 wire \top_I.branch[10].block[13].um_I.ana[3] ;
 wire \top_I.branch[10].block[13].um_I.ana[4] ;
 wire \top_I.branch[10].block[13].um_I.ana[5] ;
 wire \top_I.branch[10].block[13].um_I.ana[6] ;
 wire \top_I.branch[10].block[13].um_I.ana[7] ;
 wire \top_I.branch[10].block[13].um_I.clk ;
 wire \top_I.branch[10].block[13].um_I.ena ;
 wire \top_I.branch[10].block[13].um_I.iw[10] ;
 wire \top_I.branch[10].block[13].um_I.iw[11] ;
 wire \top_I.branch[10].block[13].um_I.iw[12] ;
 wire \top_I.branch[10].block[13].um_I.iw[13] ;
 wire \top_I.branch[10].block[13].um_I.iw[14] ;
 wire \top_I.branch[10].block[13].um_I.iw[15] ;
 wire \top_I.branch[10].block[13].um_I.iw[16] ;
 wire \top_I.branch[10].block[13].um_I.iw[17] ;
 wire \top_I.branch[10].block[13].um_I.iw[1] ;
 wire \top_I.branch[10].block[13].um_I.iw[2] ;
 wire \top_I.branch[10].block[13].um_I.iw[3] ;
 wire \top_I.branch[10].block[13].um_I.iw[4] ;
 wire \top_I.branch[10].block[13].um_I.iw[5] ;
 wire \top_I.branch[10].block[13].um_I.iw[6] ;
 wire \top_I.branch[10].block[13].um_I.iw[7] ;
 wire \top_I.branch[10].block[13].um_I.iw[8] ;
 wire \top_I.branch[10].block[13].um_I.iw[9] ;
 wire \top_I.branch[10].block[13].um_I.k_zero ;
 wire \top_I.branch[10].block[13].um_I.pg_vdd ;
 wire \top_I.branch[10].block[14].um_I.ana[0] ;
 wire \top_I.branch[10].block[14].um_I.ana[1] ;
 wire \top_I.branch[10].block[14].um_I.ana[2] ;
 wire \top_I.branch[10].block[14].um_I.ana[3] ;
 wire \top_I.branch[10].block[14].um_I.ana[4] ;
 wire \top_I.branch[10].block[14].um_I.ana[5] ;
 wire \top_I.branch[10].block[14].um_I.ana[6] ;
 wire \top_I.branch[10].block[14].um_I.ana[7] ;
 wire \top_I.branch[10].block[14].um_I.clk ;
 wire \top_I.branch[10].block[14].um_I.ena ;
 wire \top_I.branch[10].block[14].um_I.iw[10] ;
 wire \top_I.branch[10].block[14].um_I.iw[11] ;
 wire \top_I.branch[10].block[14].um_I.iw[12] ;
 wire \top_I.branch[10].block[14].um_I.iw[13] ;
 wire \top_I.branch[10].block[14].um_I.iw[14] ;
 wire \top_I.branch[10].block[14].um_I.iw[15] ;
 wire \top_I.branch[10].block[14].um_I.iw[16] ;
 wire \top_I.branch[10].block[14].um_I.iw[17] ;
 wire \top_I.branch[10].block[14].um_I.iw[1] ;
 wire \top_I.branch[10].block[14].um_I.iw[2] ;
 wire \top_I.branch[10].block[14].um_I.iw[3] ;
 wire \top_I.branch[10].block[14].um_I.iw[4] ;
 wire \top_I.branch[10].block[14].um_I.iw[5] ;
 wire \top_I.branch[10].block[14].um_I.iw[6] ;
 wire \top_I.branch[10].block[14].um_I.iw[7] ;
 wire \top_I.branch[10].block[14].um_I.iw[8] ;
 wire \top_I.branch[10].block[14].um_I.iw[9] ;
 wire \top_I.branch[10].block[14].um_I.k_zero ;
 wire \top_I.branch[10].block[14].um_I.pg_vdd ;
 wire \top_I.branch[10].block[15].um_I.ana[0] ;
 wire \top_I.branch[10].block[15].um_I.ana[1] ;
 wire \top_I.branch[10].block[15].um_I.ana[2] ;
 wire \top_I.branch[10].block[15].um_I.ana[3] ;
 wire \top_I.branch[10].block[15].um_I.ana[4] ;
 wire \top_I.branch[10].block[15].um_I.ana[5] ;
 wire \top_I.branch[10].block[15].um_I.ana[6] ;
 wire \top_I.branch[10].block[15].um_I.ana[7] ;
 wire \top_I.branch[10].block[15].um_I.clk ;
 wire \top_I.branch[10].block[15].um_I.ena ;
 wire \top_I.branch[10].block[15].um_I.iw[10] ;
 wire \top_I.branch[10].block[15].um_I.iw[11] ;
 wire \top_I.branch[10].block[15].um_I.iw[12] ;
 wire \top_I.branch[10].block[15].um_I.iw[13] ;
 wire \top_I.branch[10].block[15].um_I.iw[14] ;
 wire \top_I.branch[10].block[15].um_I.iw[15] ;
 wire \top_I.branch[10].block[15].um_I.iw[16] ;
 wire \top_I.branch[10].block[15].um_I.iw[17] ;
 wire \top_I.branch[10].block[15].um_I.iw[1] ;
 wire \top_I.branch[10].block[15].um_I.iw[2] ;
 wire \top_I.branch[10].block[15].um_I.iw[3] ;
 wire \top_I.branch[10].block[15].um_I.iw[4] ;
 wire \top_I.branch[10].block[15].um_I.iw[5] ;
 wire \top_I.branch[10].block[15].um_I.iw[6] ;
 wire \top_I.branch[10].block[15].um_I.iw[7] ;
 wire \top_I.branch[10].block[15].um_I.iw[8] ;
 wire \top_I.branch[10].block[15].um_I.iw[9] ;
 wire \top_I.branch[10].block[15].um_I.k_zero ;
 wire \top_I.branch[10].block[15].um_I.pg_vdd ;
 wire \top_I.branch[10].block[1].um_I.ana[0] ;
 wire \top_I.branch[10].block[1].um_I.ana[1] ;
 wire \top_I.branch[10].block[1].um_I.ana[2] ;
 wire \top_I.branch[10].block[1].um_I.ana[3] ;
 wire \top_I.branch[10].block[1].um_I.ana[4] ;
 wire \top_I.branch[10].block[1].um_I.ana[5] ;
 wire \top_I.branch[10].block[1].um_I.ana[6] ;
 wire \top_I.branch[10].block[1].um_I.ana[7] ;
 wire \top_I.branch[10].block[1].um_I.clk ;
 wire \top_I.branch[10].block[1].um_I.ena ;
 wire \top_I.branch[10].block[1].um_I.iw[10] ;
 wire \top_I.branch[10].block[1].um_I.iw[11] ;
 wire \top_I.branch[10].block[1].um_I.iw[12] ;
 wire \top_I.branch[10].block[1].um_I.iw[13] ;
 wire \top_I.branch[10].block[1].um_I.iw[14] ;
 wire \top_I.branch[10].block[1].um_I.iw[15] ;
 wire \top_I.branch[10].block[1].um_I.iw[16] ;
 wire \top_I.branch[10].block[1].um_I.iw[17] ;
 wire \top_I.branch[10].block[1].um_I.iw[1] ;
 wire \top_I.branch[10].block[1].um_I.iw[2] ;
 wire \top_I.branch[10].block[1].um_I.iw[3] ;
 wire \top_I.branch[10].block[1].um_I.iw[4] ;
 wire \top_I.branch[10].block[1].um_I.iw[5] ;
 wire \top_I.branch[10].block[1].um_I.iw[6] ;
 wire \top_I.branch[10].block[1].um_I.iw[7] ;
 wire \top_I.branch[10].block[1].um_I.iw[8] ;
 wire \top_I.branch[10].block[1].um_I.iw[9] ;
 wire \top_I.branch[10].block[1].um_I.k_zero ;
 wire \top_I.branch[10].block[1].um_I.pg_vdd ;
 wire \top_I.branch[10].block[2].um_I.ana[0] ;
 wire \top_I.branch[10].block[2].um_I.ana[1] ;
 wire \top_I.branch[10].block[2].um_I.ana[2] ;
 wire \top_I.branch[10].block[2].um_I.ana[3] ;
 wire \top_I.branch[10].block[2].um_I.ana[4] ;
 wire \top_I.branch[10].block[2].um_I.ana[5] ;
 wire \top_I.branch[10].block[2].um_I.ana[6] ;
 wire \top_I.branch[10].block[2].um_I.ana[7] ;
 wire \top_I.branch[10].block[2].um_I.clk ;
 wire \top_I.branch[10].block[2].um_I.ena ;
 wire \top_I.branch[10].block[2].um_I.iw[10] ;
 wire \top_I.branch[10].block[2].um_I.iw[11] ;
 wire \top_I.branch[10].block[2].um_I.iw[12] ;
 wire \top_I.branch[10].block[2].um_I.iw[13] ;
 wire \top_I.branch[10].block[2].um_I.iw[14] ;
 wire \top_I.branch[10].block[2].um_I.iw[15] ;
 wire \top_I.branch[10].block[2].um_I.iw[16] ;
 wire \top_I.branch[10].block[2].um_I.iw[17] ;
 wire \top_I.branch[10].block[2].um_I.iw[1] ;
 wire \top_I.branch[10].block[2].um_I.iw[2] ;
 wire \top_I.branch[10].block[2].um_I.iw[3] ;
 wire \top_I.branch[10].block[2].um_I.iw[4] ;
 wire \top_I.branch[10].block[2].um_I.iw[5] ;
 wire \top_I.branch[10].block[2].um_I.iw[6] ;
 wire \top_I.branch[10].block[2].um_I.iw[7] ;
 wire \top_I.branch[10].block[2].um_I.iw[8] ;
 wire \top_I.branch[10].block[2].um_I.iw[9] ;
 wire \top_I.branch[10].block[2].um_I.k_zero ;
 wire \top_I.branch[10].block[2].um_I.pg_vdd ;
 wire \top_I.branch[10].block[3].um_I.ana[0] ;
 wire \top_I.branch[10].block[3].um_I.ana[1] ;
 wire \top_I.branch[10].block[3].um_I.ana[2] ;
 wire \top_I.branch[10].block[3].um_I.ana[3] ;
 wire \top_I.branch[10].block[3].um_I.ana[4] ;
 wire \top_I.branch[10].block[3].um_I.ana[5] ;
 wire \top_I.branch[10].block[3].um_I.ana[6] ;
 wire \top_I.branch[10].block[3].um_I.ana[7] ;
 wire \top_I.branch[10].block[3].um_I.clk ;
 wire \top_I.branch[10].block[3].um_I.ena ;
 wire \top_I.branch[10].block[3].um_I.iw[10] ;
 wire \top_I.branch[10].block[3].um_I.iw[11] ;
 wire \top_I.branch[10].block[3].um_I.iw[12] ;
 wire \top_I.branch[10].block[3].um_I.iw[13] ;
 wire \top_I.branch[10].block[3].um_I.iw[14] ;
 wire \top_I.branch[10].block[3].um_I.iw[15] ;
 wire \top_I.branch[10].block[3].um_I.iw[16] ;
 wire \top_I.branch[10].block[3].um_I.iw[17] ;
 wire \top_I.branch[10].block[3].um_I.iw[1] ;
 wire \top_I.branch[10].block[3].um_I.iw[2] ;
 wire \top_I.branch[10].block[3].um_I.iw[3] ;
 wire \top_I.branch[10].block[3].um_I.iw[4] ;
 wire \top_I.branch[10].block[3].um_I.iw[5] ;
 wire \top_I.branch[10].block[3].um_I.iw[6] ;
 wire \top_I.branch[10].block[3].um_I.iw[7] ;
 wire \top_I.branch[10].block[3].um_I.iw[8] ;
 wire \top_I.branch[10].block[3].um_I.iw[9] ;
 wire \top_I.branch[10].block[3].um_I.k_zero ;
 wire \top_I.branch[10].block[3].um_I.pg_vdd ;
 wire \top_I.branch[10].block[4].um_I.ana[0] ;
 wire \top_I.branch[10].block[4].um_I.ana[1] ;
 wire \top_I.branch[10].block[4].um_I.ana[2] ;
 wire \top_I.branch[10].block[4].um_I.ana[3] ;
 wire \top_I.branch[10].block[4].um_I.ana[4] ;
 wire \top_I.branch[10].block[4].um_I.ana[5] ;
 wire \top_I.branch[10].block[4].um_I.ana[6] ;
 wire \top_I.branch[10].block[4].um_I.ana[7] ;
 wire \top_I.branch[10].block[4].um_I.clk ;
 wire \top_I.branch[10].block[4].um_I.ena ;
 wire \top_I.branch[10].block[4].um_I.iw[10] ;
 wire \top_I.branch[10].block[4].um_I.iw[11] ;
 wire \top_I.branch[10].block[4].um_I.iw[12] ;
 wire \top_I.branch[10].block[4].um_I.iw[13] ;
 wire \top_I.branch[10].block[4].um_I.iw[14] ;
 wire \top_I.branch[10].block[4].um_I.iw[15] ;
 wire \top_I.branch[10].block[4].um_I.iw[16] ;
 wire \top_I.branch[10].block[4].um_I.iw[17] ;
 wire \top_I.branch[10].block[4].um_I.iw[1] ;
 wire \top_I.branch[10].block[4].um_I.iw[2] ;
 wire \top_I.branch[10].block[4].um_I.iw[3] ;
 wire \top_I.branch[10].block[4].um_I.iw[4] ;
 wire \top_I.branch[10].block[4].um_I.iw[5] ;
 wire \top_I.branch[10].block[4].um_I.iw[6] ;
 wire \top_I.branch[10].block[4].um_I.iw[7] ;
 wire \top_I.branch[10].block[4].um_I.iw[8] ;
 wire \top_I.branch[10].block[4].um_I.iw[9] ;
 wire \top_I.branch[10].block[4].um_I.k_zero ;
 wire \top_I.branch[10].block[4].um_I.pg_vdd ;
 wire \top_I.branch[10].block[5].um_I.ana[0] ;
 wire \top_I.branch[10].block[5].um_I.ana[1] ;
 wire \top_I.branch[10].block[5].um_I.ana[2] ;
 wire \top_I.branch[10].block[5].um_I.ana[3] ;
 wire \top_I.branch[10].block[5].um_I.ana[4] ;
 wire \top_I.branch[10].block[5].um_I.ana[5] ;
 wire \top_I.branch[10].block[5].um_I.ana[6] ;
 wire \top_I.branch[10].block[5].um_I.ana[7] ;
 wire \top_I.branch[10].block[5].um_I.clk ;
 wire \top_I.branch[10].block[5].um_I.ena ;
 wire \top_I.branch[10].block[5].um_I.iw[10] ;
 wire \top_I.branch[10].block[5].um_I.iw[11] ;
 wire \top_I.branch[10].block[5].um_I.iw[12] ;
 wire \top_I.branch[10].block[5].um_I.iw[13] ;
 wire \top_I.branch[10].block[5].um_I.iw[14] ;
 wire \top_I.branch[10].block[5].um_I.iw[15] ;
 wire \top_I.branch[10].block[5].um_I.iw[16] ;
 wire \top_I.branch[10].block[5].um_I.iw[17] ;
 wire \top_I.branch[10].block[5].um_I.iw[1] ;
 wire \top_I.branch[10].block[5].um_I.iw[2] ;
 wire \top_I.branch[10].block[5].um_I.iw[3] ;
 wire \top_I.branch[10].block[5].um_I.iw[4] ;
 wire \top_I.branch[10].block[5].um_I.iw[5] ;
 wire \top_I.branch[10].block[5].um_I.iw[6] ;
 wire \top_I.branch[10].block[5].um_I.iw[7] ;
 wire \top_I.branch[10].block[5].um_I.iw[8] ;
 wire \top_I.branch[10].block[5].um_I.iw[9] ;
 wire \top_I.branch[10].block[5].um_I.k_zero ;
 wire \top_I.branch[10].block[5].um_I.pg_vdd ;
 wire \top_I.branch[10].block[6].um_I.ana[0] ;
 wire \top_I.branch[10].block[6].um_I.ana[1] ;
 wire \top_I.branch[10].block[6].um_I.ana[2] ;
 wire \top_I.branch[10].block[6].um_I.ana[3] ;
 wire \top_I.branch[10].block[6].um_I.ana[4] ;
 wire \top_I.branch[10].block[6].um_I.ana[5] ;
 wire \top_I.branch[10].block[6].um_I.ana[6] ;
 wire \top_I.branch[10].block[6].um_I.ana[7] ;
 wire \top_I.branch[10].block[6].um_I.clk ;
 wire \top_I.branch[10].block[6].um_I.ena ;
 wire \top_I.branch[10].block[6].um_I.iw[10] ;
 wire \top_I.branch[10].block[6].um_I.iw[11] ;
 wire \top_I.branch[10].block[6].um_I.iw[12] ;
 wire \top_I.branch[10].block[6].um_I.iw[13] ;
 wire \top_I.branch[10].block[6].um_I.iw[14] ;
 wire \top_I.branch[10].block[6].um_I.iw[15] ;
 wire \top_I.branch[10].block[6].um_I.iw[16] ;
 wire \top_I.branch[10].block[6].um_I.iw[17] ;
 wire \top_I.branch[10].block[6].um_I.iw[1] ;
 wire \top_I.branch[10].block[6].um_I.iw[2] ;
 wire \top_I.branch[10].block[6].um_I.iw[3] ;
 wire \top_I.branch[10].block[6].um_I.iw[4] ;
 wire \top_I.branch[10].block[6].um_I.iw[5] ;
 wire \top_I.branch[10].block[6].um_I.iw[6] ;
 wire \top_I.branch[10].block[6].um_I.iw[7] ;
 wire \top_I.branch[10].block[6].um_I.iw[8] ;
 wire \top_I.branch[10].block[6].um_I.iw[9] ;
 wire \top_I.branch[10].block[6].um_I.k_zero ;
 wire \top_I.branch[10].block[6].um_I.pg_vdd ;
 wire \top_I.branch[10].block[7].um_I.ana[0] ;
 wire \top_I.branch[10].block[7].um_I.ana[1] ;
 wire \top_I.branch[10].block[7].um_I.ana[2] ;
 wire \top_I.branch[10].block[7].um_I.ana[3] ;
 wire \top_I.branch[10].block[7].um_I.ana[4] ;
 wire \top_I.branch[10].block[7].um_I.ana[5] ;
 wire \top_I.branch[10].block[7].um_I.ana[6] ;
 wire \top_I.branch[10].block[7].um_I.ana[7] ;
 wire \top_I.branch[10].block[7].um_I.clk ;
 wire \top_I.branch[10].block[7].um_I.ena ;
 wire \top_I.branch[10].block[7].um_I.iw[10] ;
 wire \top_I.branch[10].block[7].um_I.iw[11] ;
 wire \top_I.branch[10].block[7].um_I.iw[12] ;
 wire \top_I.branch[10].block[7].um_I.iw[13] ;
 wire \top_I.branch[10].block[7].um_I.iw[14] ;
 wire \top_I.branch[10].block[7].um_I.iw[15] ;
 wire \top_I.branch[10].block[7].um_I.iw[16] ;
 wire \top_I.branch[10].block[7].um_I.iw[17] ;
 wire \top_I.branch[10].block[7].um_I.iw[1] ;
 wire \top_I.branch[10].block[7].um_I.iw[2] ;
 wire \top_I.branch[10].block[7].um_I.iw[3] ;
 wire \top_I.branch[10].block[7].um_I.iw[4] ;
 wire \top_I.branch[10].block[7].um_I.iw[5] ;
 wire \top_I.branch[10].block[7].um_I.iw[6] ;
 wire \top_I.branch[10].block[7].um_I.iw[7] ;
 wire \top_I.branch[10].block[7].um_I.iw[8] ;
 wire \top_I.branch[10].block[7].um_I.iw[9] ;
 wire \top_I.branch[10].block[7].um_I.k_zero ;
 wire \top_I.branch[10].block[7].um_I.pg_vdd ;
 wire \top_I.branch[10].block[8].um_I.ana[0] ;
 wire \top_I.branch[10].block[8].um_I.ana[1] ;
 wire \top_I.branch[10].block[8].um_I.ana[2] ;
 wire \top_I.branch[10].block[8].um_I.ana[3] ;
 wire \top_I.branch[10].block[8].um_I.ana[4] ;
 wire \top_I.branch[10].block[8].um_I.ana[5] ;
 wire \top_I.branch[10].block[8].um_I.ana[6] ;
 wire \top_I.branch[10].block[8].um_I.ana[7] ;
 wire \top_I.branch[10].block[8].um_I.clk ;
 wire \top_I.branch[10].block[8].um_I.ena ;
 wire \top_I.branch[10].block[8].um_I.iw[10] ;
 wire \top_I.branch[10].block[8].um_I.iw[11] ;
 wire \top_I.branch[10].block[8].um_I.iw[12] ;
 wire \top_I.branch[10].block[8].um_I.iw[13] ;
 wire \top_I.branch[10].block[8].um_I.iw[14] ;
 wire \top_I.branch[10].block[8].um_I.iw[15] ;
 wire \top_I.branch[10].block[8].um_I.iw[16] ;
 wire \top_I.branch[10].block[8].um_I.iw[17] ;
 wire \top_I.branch[10].block[8].um_I.iw[1] ;
 wire \top_I.branch[10].block[8].um_I.iw[2] ;
 wire \top_I.branch[10].block[8].um_I.iw[3] ;
 wire \top_I.branch[10].block[8].um_I.iw[4] ;
 wire \top_I.branch[10].block[8].um_I.iw[5] ;
 wire \top_I.branch[10].block[8].um_I.iw[6] ;
 wire \top_I.branch[10].block[8].um_I.iw[7] ;
 wire \top_I.branch[10].block[8].um_I.iw[8] ;
 wire \top_I.branch[10].block[8].um_I.iw[9] ;
 wire \top_I.branch[10].block[8].um_I.k_zero ;
 wire \top_I.branch[10].block[8].um_I.pg_vdd ;
 wire \top_I.branch[10].block[9].um_I.ana[0] ;
 wire \top_I.branch[10].block[9].um_I.ana[1] ;
 wire \top_I.branch[10].block[9].um_I.ana[2] ;
 wire \top_I.branch[10].block[9].um_I.ana[3] ;
 wire \top_I.branch[10].block[9].um_I.ana[4] ;
 wire \top_I.branch[10].block[9].um_I.ana[5] ;
 wire \top_I.branch[10].block[9].um_I.ana[6] ;
 wire \top_I.branch[10].block[9].um_I.ana[7] ;
 wire \top_I.branch[10].block[9].um_I.clk ;
 wire \top_I.branch[10].block[9].um_I.ena ;
 wire \top_I.branch[10].block[9].um_I.iw[10] ;
 wire \top_I.branch[10].block[9].um_I.iw[11] ;
 wire \top_I.branch[10].block[9].um_I.iw[12] ;
 wire \top_I.branch[10].block[9].um_I.iw[13] ;
 wire \top_I.branch[10].block[9].um_I.iw[14] ;
 wire \top_I.branch[10].block[9].um_I.iw[15] ;
 wire \top_I.branch[10].block[9].um_I.iw[16] ;
 wire \top_I.branch[10].block[9].um_I.iw[17] ;
 wire \top_I.branch[10].block[9].um_I.iw[1] ;
 wire \top_I.branch[10].block[9].um_I.iw[2] ;
 wire \top_I.branch[10].block[9].um_I.iw[3] ;
 wire \top_I.branch[10].block[9].um_I.iw[4] ;
 wire \top_I.branch[10].block[9].um_I.iw[5] ;
 wire \top_I.branch[10].block[9].um_I.iw[6] ;
 wire \top_I.branch[10].block[9].um_I.iw[7] ;
 wire \top_I.branch[10].block[9].um_I.iw[8] ;
 wire \top_I.branch[10].block[9].um_I.iw[9] ;
 wire \top_I.branch[10].block[9].um_I.k_zero ;
 wire \top_I.branch[10].block[9].um_I.pg_vdd ;
 wire \top_I.branch[10].l_addr[0] ;
 wire \top_I.branch[10].l_addr[1] ;
 wire \top_I.branch[11].block[0].um_I.ana[0] ;
 wire \top_I.branch[11].block[0].um_I.ana[1] ;
 wire \top_I.branch[11].block[0].um_I.ana[2] ;
 wire \top_I.branch[11].block[0].um_I.ana[3] ;
 wire \top_I.branch[11].block[0].um_I.ana[4] ;
 wire \top_I.branch[11].block[0].um_I.ana[5] ;
 wire \top_I.branch[11].block[0].um_I.ana[6] ;
 wire \top_I.branch[11].block[0].um_I.ana[7] ;
 wire \top_I.branch[11].block[0].um_I.clk ;
 wire \top_I.branch[11].block[0].um_I.ena ;
 wire \top_I.branch[11].block[0].um_I.iw[10] ;
 wire \top_I.branch[11].block[0].um_I.iw[11] ;
 wire \top_I.branch[11].block[0].um_I.iw[12] ;
 wire \top_I.branch[11].block[0].um_I.iw[13] ;
 wire \top_I.branch[11].block[0].um_I.iw[14] ;
 wire \top_I.branch[11].block[0].um_I.iw[15] ;
 wire \top_I.branch[11].block[0].um_I.iw[16] ;
 wire \top_I.branch[11].block[0].um_I.iw[17] ;
 wire \top_I.branch[11].block[0].um_I.iw[1] ;
 wire \top_I.branch[11].block[0].um_I.iw[2] ;
 wire \top_I.branch[11].block[0].um_I.iw[3] ;
 wire \top_I.branch[11].block[0].um_I.iw[4] ;
 wire \top_I.branch[11].block[0].um_I.iw[5] ;
 wire \top_I.branch[11].block[0].um_I.iw[6] ;
 wire \top_I.branch[11].block[0].um_I.iw[7] ;
 wire \top_I.branch[11].block[0].um_I.iw[8] ;
 wire \top_I.branch[11].block[0].um_I.iw[9] ;
 wire \top_I.branch[11].block[0].um_I.k_zero ;
 wire \top_I.branch[11].block[0].um_I.pg_vdd ;
 wire \top_I.branch[11].block[10].um_I.ana[0] ;
 wire \top_I.branch[11].block[10].um_I.ana[1] ;
 wire \top_I.branch[11].block[10].um_I.ana[2] ;
 wire \top_I.branch[11].block[10].um_I.ana[3] ;
 wire \top_I.branch[11].block[10].um_I.ana[4] ;
 wire \top_I.branch[11].block[10].um_I.ana[5] ;
 wire \top_I.branch[11].block[10].um_I.ana[6] ;
 wire \top_I.branch[11].block[10].um_I.ana[7] ;
 wire \top_I.branch[11].block[10].um_I.clk ;
 wire \top_I.branch[11].block[10].um_I.ena ;
 wire \top_I.branch[11].block[10].um_I.iw[10] ;
 wire \top_I.branch[11].block[10].um_I.iw[11] ;
 wire \top_I.branch[11].block[10].um_I.iw[12] ;
 wire \top_I.branch[11].block[10].um_I.iw[13] ;
 wire \top_I.branch[11].block[10].um_I.iw[14] ;
 wire \top_I.branch[11].block[10].um_I.iw[15] ;
 wire \top_I.branch[11].block[10].um_I.iw[16] ;
 wire \top_I.branch[11].block[10].um_I.iw[17] ;
 wire \top_I.branch[11].block[10].um_I.iw[1] ;
 wire \top_I.branch[11].block[10].um_I.iw[2] ;
 wire \top_I.branch[11].block[10].um_I.iw[3] ;
 wire \top_I.branch[11].block[10].um_I.iw[4] ;
 wire \top_I.branch[11].block[10].um_I.iw[5] ;
 wire \top_I.branch[11].block[10].um_I.iw[6] ;
 wire \top_I.branch[11].block[10].um_I.iw[7] ;
 wire \top_I.branch[11].block[10].um_I.iw[8] ;
 wire \top_I.branch[11].block[10].um_I.iw[9] ;
 wire \top_I.branch[11].block[10].um_I.k_zero ;
 wire \top_I.branch[11].block[10].um_I.pg_vdd ;
 wire \top_I.branch[11].block[11].um_I.ana[0] ;
 wire \top_I.branch[11].block[11].um_I.ana[1] ;
 wire \top_I.branch[11].block[11].um_I.ana[2] ;
 wire \top_I.branch[11].block[11].um_I.ana[3] ;
 wire \top_I.branch[11].block[11].um_I.ana[4] ;
 wire \top_I.branch[11].block[11].um_I.ana[5] ;
 wire \top_I.branch[11].block[11].um_I.ana[6] ;
 wire \top_I.branch[11].block[11].um_I.ana[7] ;
 wire \top_I.branch[11].block[11].um_I.clk ;
 wire \top_I.branch[11].block[11].um_I.ena ;
 wire \top_I.branch[11].block[11].um_I.iw[10] ;
 wire \top_I.branch[11].block[11].um_I.iw[11] ;
 wire \top_I.branch[11].block[11].um_I.iw[12] ;
 wire \top_I.branch[11].block[11].um_I.iw[13] ;
 wire \top_I.branch[11].block[11].um_I.iw[14] ;
 wire \top_I.branch[11].block[11].um_I.iw[15] ;
 wire \top_I.branch[11].block[11].um_I.iw[16] ;
 wire \top_I.branch[11].block[11].um_I.iw[17] ;
 wire \top_I.branch[11].block[11].um_I.iw[1] ;
 wire \top_I.branch[11].block[11].um_I.iw[2] ;
 wire \top_I.branch[11].block[11].um_I.iw[3] ;
 wire \top_I.branch[11].block[11].um_I.iw[4] ;
 wire \top_I.branch[11].block[11].um_I.iw[5] ;
 wire \top_I.branch[11].block[11].um_I.iw[6] ;
 wire \top_I.branch[11].block[11].um_I.iw[7] ;
 wire \top_I.branch[11].block[11].um_I.iw[8] ;
 wire \top_I.branch[11].block[11].um_I.iw[9] ;
 wire \top_I.branch[11].block[11].um_I.k_zero ;
 wire \top_I.branch[11].block[11].um_I.pg_vdd ;
 wire \top_I.branch[11].block[12].um_I.ana[0] ;
 wire \top_I.branch[11].block[12].um_I.ana[1] ;
 wire \top_I.branch[11].block[12].um_I.ana[2] ;
 wire \top_I.branch[11].block[12].um_I.ana[3] ;
 wire \top_I.branch[11].block[12].um_I.ana[4] ;
 wire \top_I.branch[11].block[12].um_I.ana[5] ;
 wire \top_I.branch[11].block[12].um_I.ana[6] ;
 wire \top_I.branch[11].block[12].um_I.ana[7] ;
 wire \top_I.branch[11].block[12].um_I.clk ;
 wire \top_I.branch[11].block[12].um_I.ena ;
 wire \top_I.branch[11].block[12].um_I.iw[10] ;
 wire \top_I.branch[11].block[12].um_I.iw[11] ;
 wire \top_I.branch[11].block[12].um_I.iw[12] ;
 wire \top_I.branch[11].block[12].um_I.iw[13] ;
 wire \top_I.branch[11].block[12].um_I.iw[14] ;
 wire \top_I.branch[11].block[12].um_I.iw[15] ;
 wire \top_I.branch[11].block[12].um_I.iw[16] ;
 wire \top_I.branch[11].block[12].um_I.iw[17] ;
 wire \top_I.branch[11].block[12].um_I.iw[1] ;
 wire \top_I.branch[11].block[12].um_I.iw[2] ;
 wire \top_I.branch[11].block[12].um_I.iw[3] ;
 wire \top_I.branch[11].block[12].um_I.iw[4] ;
 wire \top_I.branch[11].block[12].um_I.iw[5] ;
 wire \top_I.branch[11].block[12].um_I.iw[6] ;
 wire \top_I.branch[11].block[12].um_I.iw[7] ;
 wire \top_I.branch[11].block[12].um_I.iw[8] ;
 wire \top_I.branch[11].block[12].um_I.iw[9] ;
 wire \top_I.branch[11].block[12].um_I.k_zero ;
 wire \top_I.branch[11].block[12].um_I.pg_vdd ;
 wire \top_I.branch[11].block[13].um_I.ana[0] ;
 wire \top_I.branch[11].block[13].um_I.ana[1] ;
 wire \top_I.branch[11].block[13].um_I.ana[2] ;
 wire \top_I.branch[11].block[13].um_I.ana[3] ;
 wire \top_I.branch[11].block[13].um_I.ana[4] ;
 wire \top_I.branch[11].block[13].um_I.ana[5] ;
 wire \top_I.branch[11].block[13].um_I.ana[6] ;
 wire \top_I.branch[11].block[13].um_I.ana[7] ;
 wire \top_I.branch[11].block[13].um_I.clk ;
 wire \top_I.branch[11].block[13].um_I.ena ;
 wire \top_I.branch[11].block[13].um_I.iw[10] ;
 wire \top_I.branch[11].block[13].um_I.iw[11] ;
 wire \top_I.branch[11].block[13].um_I.iw[12] ;
 wire \top_I.branch[11].block[13].um_I.iw[13] ;
 wire \top_I.branch[11].block[13].um_I.iw[14] ;
 wire \top_I.branch[11].block[13].um_I.iw[15] ;
 wire \top_I.branch[11].block[13].um_I.iw[16] ;
 wire \top_I.branch[11].block[13].um_I.iw[17] ;
 wire \top_I.branch[11].block[13].um_I.iw[1] ;
 wire \top_I.branch[11].block[13].um_I.iw[2] ;
 wire \top_I.branch[11].block[13].um_I.iw[3] ;
 wire \top_I.branch[11].block[13].um_I.iw[4] ;
 wire \top_I.branch[11].block[13].um_I.iw[5] ;
 wire \top_I.branch[11].block[13].um_I.iw[6] ;
 wire \top_I.branch[11].block[13].um_I.iw[7] ;
 wire \top_I.branch[11].block[13].um_I.iw[8] ;
 wire \top_I.branch[11].block[13].um_I.iw[9] ;
 wire \top_I.branch[11].block[13].um_I.k_zero ;
 wire \top_I.branch[11].block[13].um_I.pg_vdd ;
 wire \top_I.branch[11].block[14].um_I.ana[0] ;
 wire \top_I.branch[11].block[14].um_I.ana[1] ;
 wire \top_I.branch[11].block[14].um_I.ana[2] ;
 wire \top_I.branch[11].block[14].um_I.ana[3] ;
 wire \top_I.branch[11].block[14].um_I.ana[4] ;
 wire \top_I.branch[11].block[14].um_I.ana[5] ;
 wire \top_I.branch[11].block[14].um_I.ana[6] ;
 wire \top_I.branch[11].block[14].um_I.ana[7] ;
 wire \top_I.branch[11].block[14].um_I.clk ;
 wire \top_I.branch[11].block[14].um_I.ena ;
 wire \top_I.branch[11].block[14].um_I.iw[10] ;
 wire \top_I.branch[11].block[14].um_I.iw[11] ;
 wire \top_I.branch[11].block[14].um_I.iw[12] ;
 wire \top_I.branch[11].block[14].um_I.iw[13] ;
 wire \top_I.branch[11].block[14].um_I.iw[14] ;
 wire \top_I.branch[11].block[14].um_I.iw[15] ;
 wire \top_I.branch[11].block[14].um_I.iw[16] ;
 wire \top_I.branch[11].block[14].um_I.iw[17] ;
 wire \top_I.branch[11].block[14].um_I.iw[1] ;
 wire \top_I.branch[11].block[14].um_I.iw[2] ;
 wire \top_I.branch[11].block[14].um_I.iw[3] ;
 wire \top_I.branch[11].block[14].um_I.iw[4] ;
 wire \top_I.branch[11].block[14].um_I.iw[5] ;
 wire \top_I.branch[11].block[14].um_I.iw[6] ;
 wire \top_I.branch[11].block[14].um_I.iw[7] ;
 wire \top_I.branch[11].block[14].um_I.iw[8] ;
 wire \top_I.branch[11].block[14].um_I.iw[9] ;
 wire \top_I.branch[11].block[14].um_I.k_zero ;
 wire \top_I.branch[11].block[14].um_I.pg_vdd ;
 wire \top_I.branch[11].block[15].um_I.ana[0] ;
 wire \top_I.branch[11].block[15].um_I.ana[1] ;
 wire \top_I.branch[11].block[15].um_I.ana[2] ;
 wire \top_I.branch[11].block[15].um_I.ana[3] ;
 wire \top_I.branch[11].block[15].um_I.ana[4] ;
 wire \top_I.branch[11].block[15].um_I.ana[5] ;
 wire \top_I.branch[11].block[15].um_I.ana[6] ;
 wire \top_I.branch[11].block[15].um_I.ana[7] ;
 wire \top_I.branch[11].block[15].um_I.clk ;
 wire \top_I.branch[11].block[15].um_I.ena ;
 wire \top_I.branch[11].block[15].um_I.iw[10] ;
 wire \top_I.branch[11].block[15].um_I.iw[11] ;
 wire \top_I.branch[11].block[15].um_I.iw[12] ;
 wire \top_I.branch[11].block[15].um_I.iw[13] ;
 wire \top_I.branch[11].block[15].um_I.iw[14] ;
 wire \top_I.branch[11].block[15].um_I.iw[15] ;
 wire \top_I.branch[11].block[15].um_I.iw[16] ;
 wire \top_I.branch[11].block[15].um_I.iw[17] ;
 wire \top_I.branch[11].block[15].um_I.iw[1] ;
 wire \top_I.branch[11].block[15].um_I.iw[2] ;
 wire \top_I.branch[11].block[15].um_I.iw[3] ;
 wire \top_I.branch[11].block[15].um_I.iw[4] ;
 wire \top_I.branch[11].block[15].um_I.iw[5] ;
 wire \top_I.branch[11].block[15].um_I.iw[6] ;
 wire \top_I.branch[11].block[15].um_I.iw[7] ;
 wire \top_I.branch[11].block[15].um_I.iw[8] ;
 wire \top_I.branch[11].block[15].um_I.iw[9] ;
 wire \top_I.branch[11].block[15].um_I.k_zero ;
 wire \top_I.branch[11].block[15].um_I.pg_vdd ;
 wire \top_I.branch[11].block[1].um_I.ana[0] ;
 wire \top_I.branch[11].block[1].um_I.ana[1] ;
 wire \top_I.branch[11].block[1].um_I.ana[2] ;
 wire \top_I.branch[11].block[1].um_I.ana[3] ;
 wire \top_I.branch[11].block[1].um_I.ana[4] ;
 wire \top_I.branch[11].block[1].um_I.ana[5] ;
 wire \top_I.branch[11].block[1].um_I.ana[6] ;
 wire \top_I.branch[11].block[1].um_I.ana[7] ;
 wire \top_I.branch[11].block[1].um_I.clk ;
 wire \top_I.branch[11].block[1].um_I.ena ;
 wire \top_I.branch[11].block[1].um_I.iw[10] ;
 wire \top_I.branch[11].block[1].um_I.iw[11] ;
 wire \top_I.branch[11].block[1].um_I.iw[12] ;
 wire \top_I.branch[11].block[1].um_I.iw[13] ;
 wire \top_I.branch[11].block[1].um_I.iw[14] ;
 wire \top_I.branch[11].block[1].um_I.iw[15] ;
 wire \top_I.branch[11].block[1].um_I.iw[16] ;
 wire \top_I.branch[11].block[1].um_I.iw[17] ;
 wire \top_I.branch[11].block[1].um_I.iw[1] ;
 wire \top_I.branch[11].block[1].um_I.iw[2] ;
 wire \top_I.branch[11].block[1].um_I.iw[3] ;
 wire \top_I.branch[11].block[1].um_I.iw[4] ;
 wire \top_I.branch[11].block[1].um_I.iw[5] ;
 wire \top_I.branch[11].block[1].um_I.iw[6] ;
 wire \top_I.branch[11].block[1].um_I.iw[7] ;
 wire \top_I.branch[11].block[1].um_I.iw[8] ;
 wire \top_I.branch[11].block[1].um_I.iw[9] ;
 wire \top_I.branch[11].block[1].um_I.k_zero ;
 wire \top_I.branch[11].block[1].um_I.pg_vdd ;
 wire \top_I.branch[11].block[2].um_I.ana[0] ;
 wire \top_I.branch[11].block[2].um_I.ana[1] ;
 wire \top_I.branch[11].block[2].um_I.ana[2] ;
 wire \top_I.branch[11].block[2].um_I.ana[3] ;
 wire \top_I.branch[11].block[2].um_I.ana[4] ;
 wire \top_I.branch[11].block[2].um_I.ana[5] ;
 wire \top_I.branch[11].block[2].um_I.ana[6] ;
 wire \top_I.branch[11].block[2].um_I.ana[7] ;
 wire \top_I.branch[11].block[2].um_I.clk ;
 wire \top_I.branch[11].block[2].um_I.ena ;
 wire \top_I.branch[11].block[2].um_I.iw[10] ;
 wire \top_I.branch[11].block[2].um_I.iw[11] ;
 wire \top_I.branch[11].block[2].um_I.iw[12] ;
 wire \top_I.branch[11].block[2].um_I.iw[13] ;
 wire \top_I.branch[11].block[2].um_I.iw[14] ;
 wire \top_I.branch[11].block[2].um_I.iw[15] ;
 wire \top_I.branch[11].block[2].um_I.iw[16] ;
 wire \top_I.branch[11].block[2].um_I.iw[17] ;
 wire \top_I.branch[11].block[2].um_I.iw[1] ;
 wire \top_I.branch[11].block[2].um_I.iw[2] ;
 wire \top_I.branch[11].block[2].um_I.iw[3] ;
 wire \top_I.branch[11].block[2].um_I.iw[4] ;
 wire \top_I.branch[11].block[2].um_I.iw[5] ;
 wire \top_I.branch[11].block[2].um_I.iw[6] ;
 wire \top_I.branch[11].block[2].um_I.iw[7] ;
 wire \top_I.branch[11].block[2].um_I.iw[8] ;
 wire \top_I.branch[11].block[2].um_I.iw[9] ;
 wire \top_I.branch[11].block[2].um_I.k_zero ;
 wire \top_I.branch[11].block[2].um_I.pg_vdd ;
 wire \top_I.branch[11].block[3].um_I.ana[0] ;
 wire \top_I.branch[11].block[3].um_I.ana[1] ;
 wire \top_I.branch[11].block[3].um_I.ana[2] ;
 wire \top_I.branch[11].block[3].um_I.ana[3] ;
 wire \top_I.branch[11].block[3].um_I.ana[4] ;
 wire \top_I.branch[11].block[3].um_I.ana[5] ;
 wire \top_I.branch[11].block[3].um_I.ana[6] ;
 wire \top_I.branch[11].block[3].um_I.ana[7] ;
 wire \top_I.branch[11].block[3].um_I.clk ;
 wire \top_I.branch[11].block[3].um_I.ena ;
 wire \top_I.branch[11].block[3].um_I.iw[10] ;
 wire \top_I.branch[11].block[3].um_I.iw[11] ;
 wire \top_I.branch[11].block[3].um_I.iw[12] ;
 wire \top_I.branch[11].block[3].um_I.iw[13] ;
 wire \top_I.branch[11].block[3].um_I.iw[14] ;
 wire \top_I.branch[11].block[3].um_I.iw[15] ;
 wire \top_I.branch[11].block[3].um_I.iw[16] ;
 wire \top_I.branch[11].block[3].um_I.iw[17] ;
 wire \top_I.branch[11].block[3].um_I.iw[1] ;
 wire \top_I.branch[11].block[3].um_I.iw[2] ;
 wire \top_I.branch[11].block[3].um_I.iw[3] ;
 wire \top_I.branch[11].block[3].um_I.iw[4] ;
 wire \top_I.branch[11].block[3].um_I.iw[5] ;
 wire \top_I.branch[11].block[3].um_I.iw[6] ;
 wire \top_I.branch[11].block[3].um_I.iw[7] ;
 wire \top_I.branch[11].block[3].um_I.iw[8] ;
 wire \top_I.branch[11].block[3].um_I.iw[9] ;
 wire \top_I.branch[11].block[3].um_I.k_zero ;
 wire \top_I.branch[11].block[3].um_I.pg_vdd ;
 wire \top_I.branch[11].block[4].um_I.ana[0] ;
 wire \top_I.branch[11].block[4].um_I.ana[1] ;
 wire \top_I.branch[11].block[4].um_I.ana[2] ;
 wire \top_I.branch[11].block[4].um_I.ana[3] ;
 wire \top_I.branch[11].block[4].um_I.ana[4] ;
 wire \top_I.branch[11].block[4].um_I.ana[5] ;
 wire \top_I.branch[11].block[4].um_I.ana[6] ;
 wire \top_I.branch[11].block[4].um_I.ana[7] ;
 wire \top_I.branch[11].block[4].um_I.clk ;
 wire \top_I.branch[11].block[4].um_I.ena ;
 wire \top_I.branch[11].block[4].um_I.iw[10] ;
 wire \top_I.branch[11].block[4].um_I.iw[11] ;
 wire \top_I.branch[11].block[4].um_I.iw[12] ;
 wire \top_I.branch[11].block[4].um_I.iw[13] ;
 wire \top_I.branch[11].block[4].um_I.iw[14] ;
 wire \top_I.branch[11].block[4].um_I.iw[15] ;
 wire \top_I.branch[11].block[4].um_I.iw[16] ;
 wire \top_I.branch[11].block[4].um_I.iw[17] ;
 wire \top_I.branch[11].block[4].um_I.iw[1] ;
 wire \top_I.branch[11].block[4].um_I.iw[2] ;
 wire \top_I.branch[11].block[4].um_I.iw[3] ;
 wire \top_I.branch[11].block[4].um_I.iw[4] ;
 wire \top_I.branch[11].block[4].um_I.iw[5] ;
 wire \top_I.branch[11].block[4].um_I.iw[6] ;
 wire \top_I.branch[11].block[4].um_I.iw[7] ;
 wire \top_I.branch[11].block[4].um_I.iw[8] ;
 wire \top_I.branch[11].block[4].um_I.iw[9] ;
 wire \top_I.branch[11].block[4].um_I.k_zero ;
 wire \top_I.branch[11].block[4].um_I.pg_vdd ;
 wire \top_I.branch[11].block[5].um_I.ana[0] ;
 wire \top_I.branch[11].block[5].um_I.ana[1] ;
 wire \top_I.branch[11].block[5].um_I.ana[2] ;
 wire \top_I.branch[11].block[5].um_I.ana[3] ;
 wire \top_I.branch[11].block[5].um_I.ana[4] ;
 wire \top_I.branch[11].block[5].um_I.ana[5] ;
 wire \top_I.branch[11].block[5].um_I.ana[6] ;
 wire \top_I.branch[11].block[5].um_I.ana[7] ;
 wire \top_I.branch[11].block[5].um_I.clk ;
 wire \top_I.branch[11].block[5].um_I.ena ;
 wire \top_I.branch[11].block[5].um_I.iw[10] ;
 wire \top_I.branch[11].block[5].um_I.iw[11] ;
 wire \top_I.branch[11].block[5].um_I.iw[12] ;
 wire \top_I.branch[11].block[5].um_I.iw[13] ;
 wire \top_I.branch[11].block[5].um_I.iw[14] ;
 wire \top_I.branch[11].block[5].um_I.iw[15] ;
 wire \top_I.branch[11].block[5].um_I.iw[16] ;
 wire \top_I.branch[11].block[5].um_I.iw[17] ;
 wire \top_I.branch[11].block[5].um_I.iw[1] ;
 wire \top_I.branch[11].block[5].um_I.iw[2] ;
 wire \top_I.branch[11].block[5].um_I.iw[3] ;
 wire \top_I.branch[11].block[5].um_I.iw[4] ;
 wire \top_I.branch[11].block[5].um_I.iw[5] ;
 wire \top_I.branch[11].block[5].um_I.iw[6] ;
 wire \top_I.branch[11].block[5].um_I.iw[7] ;
 wire \top_I.branch[11].block[5].um_I.iw[8] ;
 wire \top_I.branch[11].block[5].um_I.iw[9] ;
 wire \top_I.branch[11].block[5].um_I.k_zero ;
 wire \top_I.branch[11].block[5].um_I.pg_vdd ;
 wire \top_I.branch[11].block[6].um_I.ana[0] ;
 wire \top_I.branch[11].block[6].um_I.ana[1] ;
 wire \top_I.branch[11].block[6].um_I.ana[2] ;
 wire \top_I.branch[11].block[6].um_I.ana[3] ;
 wire \top_I.branch[11].block[6].um_I.ana[4] ;
 wire \top_I.branch[11].block[6].um_I.ana[5] ;
 wire \top_I.branch[11].block[6].um_I.ana[6] ;
 wire \top_I.branch[11].block[6].um_I.ana[7] ;
 wire \top_I.branch[11].block[6].um_I.clk ;
 wire \top_I.branch[11].block[6].um_I.ena ;
 wire \top_I.branch[11].block[6].um_I.iw[10] ;
 wire \top_I.branch[11].block[6].um_I.iw[11] ;
 wire \top_I.branch[11].block[6].um_I.iw[12] ;
 wire \top_I.branch[11].block[6].um_I.iw[13] ;
 wire \top_I.branch[11].block[6].um_I.iw[14] ;
 wire \top_I.branch[11].block[6].um_I.iw[15] ;
 wire \top_I.branch[11].block[6].um_I.iw[16] ;
 wire \top_I.branch[11].block[6].um_I.iw[17] ;
 wire \top_I.branch[11].block[6].um_I.iw[1] ;
 wire \top_I.branch[11].block[6].um_I.iw[2] ;
 wire \top_I.branch[11].block[6].um_I.iw[3] ;
 wire \top_I.branch[11].block[6].um_I.iw[4] ;
 wire \top_I.branch[11].block[6].um_I.iw[5] ;
 wire \top_I.branch[11].block[6].um_I.iw[6] ;
 wire \top_I.branch[11].block[6].um_I.iw[7] ;
 wire \top_I.branch[11].block[6].um_I.iw[8] ;
 wire \top_I.branch[11].block[6].um_I.iw[9] ;
 wire \top_I.branch[11].block[6].um_I.k_zero ;
 wire \top_I.branch[11].block[6].um_I.pg_vdd ;
 wire \top_I.branch[11].block[7].um_I.ana[0] ;
 wire \top_I.branch[11].block[7].um_I.ana[1] ;
 wire \top_I.branch[11].block[7].um_I.ana[2] ;
 wire \top_I.branch[11].block[7].um_I.ana[3] ;
 wire \top_I.branch[11].block[7].um_I.ana[4] ;
 wire \top_I.branch[11].block[7].um_I.ana[5] ;
 wire \top_I.branch[11].block[7].um_I.ana[6] ;
 wire \top_I.branch[11].block[7].um_I.ana[7] ;
 wire \top_I.branch[11].block[7].um_I.clk ;
 wire \top_I.branch[11].block[7].um_I.ena ;
 wire \top_I.branch[11].block[7].um_I.iw[10] ;
 wire \top_I.branch[11].block[7].um_I.iw[11] ;
 wire \top_I.branch[11].block[7].um_I.iw[12] ;
 wire \top_I.branch[11].block[7].um_I.iw[13] ;
 wire \top_I.branch[11].block[7].um_I.iw[14] ;
 wire \top_I.branch[11].block[7].um_I.iw[15] ;
 wire \top_I.branch[11].block[7].um_I.iw[16] ;
 wire \top_I.branch[11].block[7].um_I.iw[17] ;
 wire \top_I.branch[11].block[7].um_I.iw[1] ;
 wire \top_I.branch[11].block[7].um_I.iw[2] ;
 wire \top_I.branch[11].block[7].um_I.iw[3] ;
 wire \top_I.branch[11].block[7].um_I.iw[4] ;
 wire \top_I.branch[11].block[7].um_I.iw[5] ;
 wire \top_I.branch[11].block[7].um_I.iw[6] ;
 wire \top_I.branch[11].block[7].um_I.iw[7] ;
 wire \top_I.branch[11].block[7].um_I.iw[8] ;
 wire \top_I.branch[11].block[7].um_I.iw[9] ;
 wire \top_I.branch[11].block[7].um_I.k_zero ;
 wire \top_I.branch[11].block[7].um_I.pg_vdd ;
 wire \top_I.branch[11].block[8].um_I.ana[0] ;
 wire \top_I.branch[11].block[8].um_I.ana[1] ;
 wire \top_I.branch[11].block[8].um_I.ana[2] ;
 wire \top_I.branch[11].block[8].um_I.ana[3] ;
 wire \top_I.branch[11].block[8].um_I.ana[4] ;
 wire \top_I.branch[11].block[8].um_I.ana[5] ;
 wire \top_I.branch[11].block[8].um_I.ana[6] ;
 wire \top_I.branch[11].block[8].um_I.ana[7] ;
 wire \top_I.branch[11].block[8].um_I.clk ;
 wire \top_I.branch[11].block[8].um_I.ena ;
 wire \top_I.branch[11].block[8].um_I.iw[10] ;
 wire \top_I.branch[11].block[8].um_I.iw[11] ;
 wire \top_I.branch[11].block[8].um_I.iw[12] ;
 wire \top_I.branch[11].block[8].um_I.iw[13] ;
 wire \top_I.branch[11].block[8].um_I.iw[14] ;
 wire \top_I.branch[11].block[8].um_I.iw[15] ;
 wire \top_I.branch[11].block[8].um_I.iw[16] ;
 wire \top_I.branch[11].block[8].um_I.iw[17] ;
 wire \top_I.branch[11].block[8].um_I.iw[1] ;
 wire \top_I.branch[11].block[8].um_I.iw[2] ;
 wire \top_I.branch[11].block[8].um_I.iw[3] ;
 wire \top_I.branch[11].block[8].um_I.iw[4] ;
 wire \top_I.branch[11].block[8].um_I.iw[5] ;
 wire \top_I.branch[11].block[8].um_I.iw[6] ;
 wire \top_I.branch[11].block[8].um_I.iw[7] ;
 wire \top_I.branch[11].block[8].um_I.iw[8] ;
 wire \top_I.branch[11].block[8].um_I.iw[9] ;
 wire \top_I.branch[11].block[8].um_I.k_zero ;
 wire \top_I.branch[11].block[8].um_I.pg_vdd ;
 wire \top_I.branch[11].block[9].um_I.ana[0] ;
 wire \top_I.branch[11].block[9].um_I.ana[1] ;
 wire \top_I.branch[11].block[9].um_I.ana[2] ;
 wire \top_I.branch[11].block[9].um_I.ana[3] ;
 wire \top_I.branch[11].block[9].um_I.ana[4] ;
 wire \top_I.branch[11].block[9].um_I.ana[5] ;
 wire \top_I.branch[11].block[9].um_I.ana[6] ;
 wire \top_I.branch[11].block[9].um_I.ana[7] ;
 wire \top_I.branch[11].block[9].um_I.clk ;
 wire \top_I.branch[11].block[9].um_I.ena ;
 wire \top_I.branch[11].block[9].um_I.iw[10] ;
 wire \top_I.branch[11].block[9].um_I.iw[11] ;
 wire \top_I.branch[11].block[9].um_I.iw[12] ;
 wire \top_I.branch[11].block[9].um_I.iw[13] ;
 wire \top_I.branch[11].block[9].um_I.iw[14] ;
 wire \top_I.branch[11].block[9].um_I.iw[15] ;
 wire \top_I.branch[11].block[9].um_I.iw[16] ;
 wire \top_I.branch[11].block[9].um_I.iw[17] ;
 wire \top_I.branch[11].block[9].um_I.iw[1] ;
 wire \top_I.branch[11].block[9].um_I.iw[2] ;
 wire \top_I.branch[11].block[9].um_I.iw[3] ;
 wire \top_I.branch[11].block[9].um_I.iw[4] ;
 wire \top_I.branch[11].block[9].um_I.iw[5] ;
 wire \top_I.branch[11].block[9].um_I.iw[6] ;
 wire \top_I.branch[11].block[9].um_I.iw[7] ;
 wire \top_I.branch[11].block[9].um_I.iw[8] ;
 wire \top_I.branch[11].block[9].um_I.iw[9] ;
 wire \top_I.branch[11].block[9].um_I.k_zero ;
 wire \top_I.branch[11].block[9].um_I.pg_vdd ;
 wire \top_I.branch[11].l_addr[0] ;
 wire \top_I.branch[11].l_addr[1] ;
 wire \top_I.branch[11].l_spine_iw[0] ;
 wire \top_I.branch[11].l_spine_iw[10] ;
 wire \top_I.branch[11].l_spine_iw[11] ;
 wire \top_I.branch[11].l_spine_iw[12] ;
 wire \top_I.branch[11].l_spine_iw[13] ;
 wire \top_I.branch[11].l_spine_iw[14] ;
 wire \top_I.branch[11].l_spine_iw[15] ;
 wire \top_I.branch[11].l_spine_iw[16] ;
 wire \top_I.branch[11].l_spine_iw[17] ;
 wire \top_I.branch[11].l_spine_iw[18] ;
 wire \top_I.branch[11].l_spine_iw[19] ;
 wire \top_I.branch[11].l_spine_iw[1] ;
 wire \top_I.branch[11].l_spine_iw[20] ;
 wire \top_I.branch[11].l_spine_iw[21] ;
 wire \top_I.branch[11].l_spine_iw[22] ;
 wire \top_I.branch[11].l_spine_iw[23] ;
 wire \top_I.branch[11].l_spine_iw[24] ;
 wire \top_I.branch[11].l_spine_iw[25] ;
 wire \top_I.branch[11].l_spine_iw[26] ;
 wire \top_I.branch[11].l_spine_iw[27] ;
 wire \top_I.branch[11].l_spine_iw[28] ;
 wire \top_I.branch[11].l_spine_iw[29] ;
 wire \top_I.branch[11].l_spine_iw[2] ;
 wire \top_I.branch[11].l_spine_iw[3] ;
 wire \top_I.branch[11].l_spine_iw[4] ;
 wire \top_I.branch[11].l_spine_iw[5] ;
 wire \top_I.branch[11].l_spine_iw[6] ;
 wire \top_I.branch[11].l_spine_iw[7] ;
 wire \top_I.branch[11].l_spine_iw[8] ;
 wire \top_I.branch[11].l_spine_iw[9] ;
 wire \top_I.branch[11].l_spine_ow[0] ;
 wire \top_I.branch[11].l_spine_ow[10] ;
 wire \top_I.branch[11].l_spine_ow[11] ;
 wire \top_I.branch[11].l_spine_ow[12] ;
 wire \top_I.branch[11].l_spine_ow[13] ;
 wire \top_I.branch[11].l_spine_ow[14] ;
 wire \top_I.branch[11].l_spine_ow[15] ;
 wire \top_I.branch[11].l_spine_ow[16] ;
 wire \top_I.branch[11].l_spine_ow[17] ;
 wire \top_I.branch[11].l_spine_ow[18] ;
 wire \top_I.branch[11].l_spine_ow[19] ;
 wire \top_I.branch[11].l_spine_ow[1] ;
 wire \top_I.branch[11].l_spine_ow[20] ;
 wire \top_I.branch[11].l_spine_ow[21] ;
 wire \top_I.branch[11].l_spine_ow[22] ;
 wire \top_I.branch[11].l_spine_ow[23] ;
 wire \top_I.branch[11].l_spine_ow[24] ;
 wire \top_I.branch[11].l_spine_ow[25] ;
 wire \top_I.branch[11].l_spine_ow[2] ;
 wire \top_I.branch[11].l_spine_ow[3] ;
 wire \top_I.branch[11].l_spine_ow[4] ;
 wire \top_I.branch[11].l_spine_ow[5] ;
 wire \top_I.branch[11].l_spine_ow[6] ;
 wire \top_I.branch[11].l_spine_ow[7] ;
 wire \top_I.branch[11].l_spine_ow[8] ;
 wire \top_I.branch[11].l_spine_ow[9] ;
 wire \top_I.branch[12].block[0].um_I.ana[0] ;
 wire \top_I.branch[12].block[0].um_I.ana[1] ;
 wire \top_I.branch[12].block[0].um_I.ana[2] ;
 wire \top_I.branch[12].block[0].um_I.ana[3] ;
 wire \top_I.branch[12].block[0].um_I.ana[4] ;
 wire \top_I.branch[12].block[0].um_I.ana[5] ;
 wire \top_I.branch[12].block[0].um_I.ana[6] ;
 wire \top_I.branch[12].block[0].um_I.ana[7] ;
 wire \top_I.branch[12].block[0].um_I.clk ;
 wire \top_I.branch[12].block[0].um_I.ena ;
 wire \top_I.branch[12].block[0].um_I.iw[10] ;
 wire \top_I.branch[12].block[0].um_I.iw[11] ;
 wire \top_I.branch[12].block[0].um_I.iw[12] ;
 wire \top_I.branch[12].block[0].um_I.iw[13] ;
 wire \top_I.branch[12].block[0].um_I.iw[14] ;
 wire \top_I.branch[12].block[0].um_I.iw[15] ;
 wire \top_I.branch[12].block[0].um_I.iw[16] ;
 wire \top_I.branch[12].block[0].um_I.iw[17] ;
 wire \top_I.branch[12].block[0].um_I.iw[1] ;
 wire \top_I.branch[12].block[0].um_I.iw[2] ;
 wire \top_I.branch[12].block[0].um_I.iw[3] ;
 wire \top_I.branch[12].block[0].um_I.iw[4] ;
 wire \top_I.branch[12].block[0].um_I.iw[5] ;
 wire \top_I.branch[12].block[0].um_I.iw[6] ;
 wire \top_I.branch[12].block[0].um_I.iw[7] ;
 wire \top_I.branch[12].block[0].um_I.iw[8] ;
 wire \top_I.branch[12].block[0].um_I.iw[9] ;
 wire \top_I.branch[12].block[0].um_I.k_zero ;
 wire \top_I.branch[12].block[0].um_I.pg_vdd ;
 wire \top_I.branch[12].block[10].um_I.ana[0] ;
 wire \top_I.branch[12].block[10].um_I.ana[1] ;
 wire \top_I.branch[12].block[10].um_I.ana[2] ;
 wire \top_I.branch[12].block[10].um_I.ana[3] ;
 wire \top_I.branch[12].block[10].um_I.ana[4] ;
 wire \top_I.branch[12].block[10].um_I.ana[5] ;
 wire \top_I.branch[12].block[10].um_I.ana[6] ;
 wire \top_I.branch[12].block[10].um_I.ana[7] ;
 wire \top_I.branch[12].block[10].um_I.clk ;
 wire \top_I.branch[12].block[10].um_I.ena ;
 wire \top_I.branch[12].block[10].um_I.iw[10] ;
 wire \top_I.branch[12].block[10].um_I.iw[11] ;
 wire \top_I.branch[12].block[10].um_I.iw[12] ;
 wire \top_I.branch[12].block[10].um_I.iw[13] ;
 wire \top_I.branch[12].block[10].um_I.iw[14] ;
 wire \top_I.branch[12].block[10].um_I.iw[15] ;
 wire \top_I.branch[12].block[10].um_I.iw[16] ;
 wire \top_I.branch[12].block[10].um_I.iw[17] ;
 wire \top_I.branch[12].block[10].um_I.iw[1] ;
 wire \top_I.branch[12].block[10].um_I.iw[2] ;
 wire \top_I.branch[12].block[10].um_I.iw[3] ;
 wire \top_I.branch[12].block[10].um_I.iw[4] ;
 wire \top_I.branch[12].block[10].um_I.iw[5] ;
 wire \top_I.branch[12].block[10].um_I.iw[6] ;
 wire \top_I.branch[12].block[10].um_I.iw[7] ;
 wire \top_I.branch[12].block[10].um_I.iw[8] ;
 wire \top_I.branch[12].block[10].um_I.iw[9] ;
 wire \top_I.branch[12].block[10].um_I.k_zero ;
 wire \top_I.branch[12].block[10].um_I.pg_vdd ;
 wire \top_I.branch[12].block[11].um_I.ana[0] ;
 wire \top_I.branch[12].block[11].um_I.ana[1] ;
 wire \top_I.branch[12].block[11].um_I.ana[2] ;
 wire \top_I.branch[12].block[11].um_I.ana[3] ;
 wire \top_I.branch[12].block[11].um_I.ana[4] ;
 wire \top_I.branch[12].block[11].um_I.ana[5] ;
 wire \top_I.branch[12].block[11].um_I.ana[6] ;
 wire \top_I.branch[12].block[11].um_I.ana[7] ;
 wire \top_I.branch[12].block[11].um_I.clk ;
 wire \top_I.branch[12].block[11].um_I.ena ;
 wire \top_I.branch[12].block[11].um_I.iw[10] ;
 wire \top_I.branch[12].block[11].um_I.iw[11] ;
 wire \top_I.branch[12].block[11].um_I.iw[12] ;
 wire \top_I.branch[12].block[11].um_I.iw[13] ;
 wire \top_I.branch[12].block[11].um_I.iw[14] ;
 wire \top_I.branch[12].block[11].um_I.iw[15] ;
 wire \top_I.branch[12].block[11].um_I.iw[16] ;
 wire \top_I.branch[12].block[11].um_I.iw[17] ;
 wire \top_I.branch[12].block[11].um_I.iw[1] ;
 wire \top_I.branch[12].block[11].um_I.iw[2] ;
 wire \top_I.branch[12].block[11].um_I.iw[3] ;
 wire \top_I.branch[12].block[11].um_I.iw[4] ;
 wire \top_I.branch[12].block[11].um_I.iw[5] ;
 wire \top_I.branch[12].block[11].um_I.iw[6] ;
 wire \top_I.branch[12].block[11].um_I.iw[7] ;
 wire \top_I.branch[12].block[11].um_I.iw[8] ;
 wire \top_I.branch[12].block[11].um_I.iw[9] ;
 wire \top_I.branch[12].block[11].um_I.k_zero ;
 wire \top_I.branch[12].block[11].um_I.pg_vdd ;
 wire \top_I.branch[12].block[12].um_I.ana[0] ;
 wire \top_I.branch[12].block[12].um_I.ana[1] ;
 wire \top_I.branch[12].block[12].um_I.ana[2] ;
 wire \top_I.branch[12].block[12].um_I.ana[3] ;
 wire \top_I.branch[12].block[12].um_I.ana[4] ;
 wire \top_I.branch[12].block[12].um_I.ana[5] ;
 wire \top_I.branch[12].block[12].um_I.ana[6] ;
 wire \top_I.branch[12].block[12].um_I.ana[7] ;
 wire \top_I.branch[12].block[12].um_I.clk ;
 wire \top_I.branch[12].block[12].um_I.ena ;
 wire \top_I.branch[12].block[12].um_I.iw[10] ;
 wire \top_I.branch[12].block[12].um_I.iw[11] ;
 wire \top_I.branch[12].block[12].um_I.iw[12] ;
 wire \top_I.branch[12].block[12].um_I.iw[13] ;
 wire \top_I.branch[12].block[12].um_I.iw[14] ;
 wire \top_I.branch[12].block[12].um_I.iw[15] ;
 wire \top_I.branch[12].block[12].um_I.iw[16] ;
 wire \top_I.branch[12].block[12].um_I.iw[17] ;
 wire \top_I.branch[12].block[12].um_I.iw[1] ;
 wire \top_I.branch[12].block[12].um_I.iw[2] ;
 wire \top_I.branch[12].block[12].um_I.iw[3] ;
 wire \top_I.branch[12].block[12].um_I.iw[4] ;
 wire \top_I.branch[12].block[12].um_I.iw[5] ;
 wire \top_I.branch[12].block[12].um_I.iw[6] ;
 wire \top_I.branch[12].block[12].um_I.iw[7] ;
 wire \top_I.branch[12].block[12].um_I.iw[8] ;
 wire \top_I.branch[12].block[12].um_I.iw[9] ;
 wire \top_I.branch[12].block[12].um_I.k_zero ;
 wire \top_I.branch[12].block[12].um_I.pg_vdd ;
 wire \top_I.branch[12].block[13].um_I.ana[0] ;
 wire \top_I.branch[12].block[13].um_I.ana[1] ;
 wire \top_I.branch[12].block[13].um_I.ana[2] ;
 wire \top_I.branch[12].block[13].um_I.ana[3] ;
 wire \top_I.branch[12].block[13].um_I.ana[4] ;
 wire \top_I.branch[12].block[13].um_I.ana[5] ;
 wire \top_I.branch[12].block[13].um_I.ana[6] ;
 wire \top_I.branch[12].block[13].um_I.ana[7] ;
 wire \top_I.branch[12].block[13].um_I.clk ;
 wire \top_I.branch[12].block[13].um_I.ena ;
 wire \top_I.branch[12].block[13].um_I.iw[10] ;
 wire \top_I.branch[12].block[13].um_I.iw[11] ;
 wire \top_I.branch[12].block[13].um_I.iw[12] ;
 wire \top_I.branch[12].block[13].um_I.iw[13] ;
 wire \top_I.branch[12].block[13].um_I.iw[14] ;
 wire \top_I.branch[12].block[13].um_I.iw[15] ;
 wire \top_I.branch[12].block[13].um_I.iw[16] ;
 wire \top_I.branch[12].block[13].um_I.iw[17] ;
 wire \top_I.branch[12].block[13].um_I.iw[1] ;
 wire \top_I.branch[12].block[13].um_I.iw[2] ;
 wire \top_I.branch[12].block[13].um_I.iw[3] ;
 wire \top_I.branch[12].block[13].um_I.iw[4] ;
 wire \top_I.branch[12].block[13].um_I.iw[5] ;
 wire \top_I.branch[12].block[13].um_I.iw[6] ;
 wire \top_I.branch[12].block[13].um_I.iw[7] ;
 wire \top_I.branch[12].block[13].um_I.iw[8] ;
 wire \top_I.branch[12].block[13].um_I.iw[9] ;
 wire \top_I.branch[12].block[13].um_I.k_zero ;
 wire \top_I.branch[12].block[13].um_I.pg_vdd ;
 wire \top_I.branch[12].block[14].um_I.ana[0] ;
 wire \top_I.branch[12].block[14].um_I.ana[1] ;
 wire \top_I.branch[12].block[14].um_I.ana[2] ;
 wire \top_I.branch[12].block[14].um_I.ana[3] ;
 wire \top_I.branch[12].block[14].um_I.ana[4] ;
 wire \top_I.branch[12].block[14].um_I.ana[5] ;
 wire \top_I.branch[12].block[14].um_I.ana[6] ;
 wire \top_I.branch[12].block[14].um_I.ana[7] ;
 wire \top_I.branch[12].block[14].um_I.clk ;
 wire \top_I.branch[12].block[14].um_I.ena ;
 wire \top_I.branch[12].block[14].um_I.iw[10] ;
 wire \top_I.branch[12].block[14].um_I.iw[11] ;
 wire \top_I.branch[12].block[14].um_I.iw[12] ;
 wire \top_I.branch[12].block[14].um_I.iw[13] ;
 wire \top_I.branch[12].block[14].um_I.iw[14] ;
 wire \top_I.branch[12].block[14].um_I.iw[15] ;
 wire \top_I.branch[12].block[14].um_I.iw[16] ;
 wire \top_I.branch[12].block[14].um_I.iw[17] ;
 wire \top_I.branch[12].block[14].um_I.iw[1] ;
 wire \top_I.branch[12].block[14].um_I.iw[2] ;
 wire \top_I.branch[12].block[14].um_I.iw[3] ;
 wire \top_I.branch[12].block[14].um_I.iw[4] ;
 wire \top_I.branch[12].block[14].um_I.iw[5] ;
 wire \top_I.branch[12].block[14].um_I.iw[6] ;
 wire \top_I.branch[12].block[14].um_I.iw[7] ;
 wire \top_I.branch[12].block[14].um_I.iw[8] ;
 wire \top_I.branch[12].block[14].um_I.iw[9] ;
 wire \top_I.branch[12].block[14].um_I.k_zero ;
 wire \top_I.branch[12].block[14].um_I.pg_vdd ;
 wire \top_I.branch[12].block[15].um_I.ana[0] ;
 wire \top_I.branch[12].block[15].um_I.ana[1] ;
 wire \top_I.branch[12].block[15].um_I.ana[2] ;
 wire \top_I.branch[12].block[15].um_I.ana[3] ;
 wire \top_I.branch[12].block[15].um_I.ana[4] ;
 wire \top_I.branch[12].block[15].um_I.ana[5] ;
 wire \top_I.branch[12].block[15].um_I.ana[6] ;
 wire \top_I.branch[12].block[15].um_I.ana[7] ;
 wire \top_I.branch[12].block[15].um_I.clk ;
 wire \top_I.branch[12].block[15].um_I.ena ;
 wire \top_I.branch[12].block[15].um_I.iw[10] ;
 wire \top_I.branch[12].block[15].um_I.iw[11] ;
 wire \top_I.branch[12].block[15].um_I.iw[12] ;
 wire \top_I.branch[12].block[15].um_I.iw[13] ;
 wire \top_I.branch[12].block[15].um_I.iw[14] ;
 wire \top_I.branch[12].block[15].um_I.iw[15] ;
 wire \top_I.branch[12].block[15].um_I.iw[16] ;
 wire \top_I.branch[12].block[15].um_I.iw[17] ;
 wire \top_I.branch[12].block[15].um_I.iw[1] ;
 wire \top_I.branch[12].block[15].um_I.iw[2] ;
 wire \top_I.branch[12].block[15].um_I.iw[3] ;
 wire \top_I.branch[12].block[15].um_I.iw[4] ;
 wire \top_I.branch[12].block[15].um_I.iw[5] ;
 wire \top_I.branch[12].block[15].um_I.iw[6] ;
 wire \top_I.branch[12].block[15].um_I.iw[7] ;
 wire \top_I.branch[12].block[15].um_I.iw[8] ;
 wire \top_I.branch[12].block[15].um_I.iw[9] ;
 wire \top_I.branch[12].block[15].um_I.k_zero ;
 wire \top_I.branch[12].block[15].um_I.pg_vdd ;
 wire \top_I.branch[12].block[1].um_I.ana[0] ;
 wire \top_I.branch[12].block[1].um_I.ana[1] ;
 wire \top_I.branch[12].block[1].um_I.ana[2] ;
 wire \top_I.branch[12].block[1].um_I.ana[3] ;
 wire \top_I.branch[12].block[1].um_I.ana[4] ;
 wire \top_I.branch[12].block[1].um_I.ana[5] ;
 wire \top_I.branch[12].block[1].um_I.ana[6] ;
 wire \top_I.branch[12].block[1].um_I.ana[7] ;
 wire \top_I.branch[12].block[1].um_I.clk ;
 wire \top_I.branch[12].block[1].um_I.ena ;
 wire \top_I.branch[12].block[1].um_I.iw[10] ;
 wire \top_I.branch[12].block[1].um_I.iw[11] ;
 wire \top_I.branch[12].block[1].um_I.iw[12] ;
 wire \top_I.branch[12].block[1].um_I.iw[13] ;
 wire \top_I.branch[12].block[1].um_I.iw[14] ;
 wire \top_I.branch[12].block[1].um_I.iw[15] ;
 wire \top_I.branch[12].block[1].um_I.iw[16] ;
 wire \top_I.branch[12].block[1].um_I.iw[17] ;
 wire \top_I.branch[12].block[1].um_I.iw[1] ;
 wire \top_I.branch[12].block[1].um_I.iw[2] ;
 wire \top_I.branch[12].block[1].um_I.iw[3] ;
 wire \top_I.branch[12].block[1].um_I.iw[4] ;
 wire \top_I.branch[12].block[1].um_I.iw[5] ;
 wire \top_I.branch[12].block[1].um_I.iw[6] ;
 wire \top_I.branch[12].block[1].um_I.iw[7] ;
 wire \top_I.branch[12].block[1].um_I.iw[8] ;
 wire \top_I.branch[12].block[1].um_I.iw[9] ;
 wire \top_I.branch[12].block[1].um_I.k_zero ;
 wire \top_I.branch[12].block[1].um_I.pg_vdd ;
 wire \top_I.branch[12].block[2].um_I.ana[0] ;
 wire \top_I.branch[12].block[2].um_I.ana[1] ;
 wire \top_I.branch[12].block[2].um_I.ana[2] ;
 wire \top_I.branch[12].block[2].um_I.ana[3] ;
 wire \top_I.branch[12].block[2].um_I.ana[4] ;
 wire \top_I.branch[12].block[2].um_I.ana[5] ;
 wire \top_I.branch[12].block[2].um_I.ana[6] ;
 wire \top_I.branch[12].block[2].um_I.ana[7] ;
 wire \top_I.branch[12].block[2].um_I.clk ;
 wire \top_I.branch[12].block[2].um_I.ena ;
 wire \top_I.branch[12].block[2].um_I.iw[10] ;
 wire \top_I.branch[12].block[2].um_I.iw[11] ;
 wire \top_I.branch[12].block[2].um_I.iw[12] ;
 wire \top_I.branch[12].block[2].um_I.iw[13] ;
 wire \top_I.branch[12].block[2].um_I.iw[14] ;
 wire \top_I.branch[12].block[2].um_I.iw[15] ;
 wire \top_I.branch[12].block[2].um_I.iw[16] ;
 wire \top_I.branch[12].block[2].um_I.iw[17] ;
 wire \top_I.branch[12].block[2].um_I.iw[1] ;
 wire \top_I.branch[12].block[2].um_I.iw[2] ;
 wire \top_I.branch[12].block[2].um_I.iw[3] ;
 wire \top_I.branch[12].block[2].um_I.iw[4] ;
 wire \top_I.branch[12].block[2].um_I.iw[5] ;
 wire \top_I.branch[12].block[2].um_I.iw[6] ;
 wire \top_I.branch[12].block[2].um_I.iw[7] ;
 wire \top_I.branch[12].block[2].um_I.iw[8] ;
 wire \top_I.branch[12].block[2].um_I.iw[9] ;
 wire \top_I.branch[12].block[2].um_I.k_zero ;
 wire \top_I.branch[12].block[2].um_I.pg_vdd ;
 wire \top_I.branch[12].block[3].um_I.ana[0] ;
 wire \top_I.branch[12].block[3].um_I.ana[1] ;
 wire \top_I.branch[12].block[3].um_I.ana[2] ;
 wire \top_I.branch[12].block[3].um_I.ana[3] ;
 wire \top_I.branch[12].block[3].um_I.ana[4] ;
 wire \top_I.branch[12].block[3].um_I.ana[5] ;
 wire \top_I.branch[12].block[3].um_I.ana[6] ;
 wire \top_I.branch[12].block[3].um_I.ana[7] ;
 wire \top_I.branch[12].block[3].um_I.clk ;
 wire \top_I.branch[12].block[3].um_I.ena ;
 wire \top_I.branch[12].block[3].um_I.iw[10] ;
 wire \top_I.branch[12].block[3].um_I.iw[11] ;
 wire \top_I.branch[12].block[3].um_I.iw[12] ;
 wire \top_I.branch[12].block[3].um_I.iw[13] ;
 wire \top_I.branch[12].block[3].um_I.iw[14] ;
 wire \top_I.branch[12].block[3].um_I.iw[15] ;
 wire \top_I.branch[12].block[3].um_I.iw[16] ;
 wire \top_I.branch[12].block[3].um_I.iw[17] ;
 wire \top_I.branch[12].block[3].um_I.iw[1] ;
 wire \top_I.branch[12].block[3].um_I.iw[2] ;
 wire \top_I.branch[12].block[3].um_I.iw[3] ;
 wire \top_I.branch[12].block[3].um_I.iw[4] ;
 wire \top_I.branch[12].block[3].um_I.iw[5] ;
 wire \top_I.branch[12].block[3].um_I.iw[6] ;
 wire \top_I.branch[12].block[3].um_I.iw[7] ;
 wire \top_I.branch[12].block[3].um_I.iw[8] ;
 wire \top_I.branch[12].block[3].um_I.iw[9] ;
 wire \top_I.branch[12].block[3].um_I.k_zero ;
 wire \top_I.branch[12].block[3].um_I.pg_vdd ;
 wire \top_I.branch[12].block[4].um_I.ana[0] ;
 wire \top_I.branch[12].block[4].um_I.ana[1] ;
 wire \top_I.branch[12].block[4].um_I.ana[2] ;
 wire \top_I.branch[12].block[4].um_I.ana[3] ;
 wire \top_I.branch[12].block[4].um_I.ana[4] ;
 wire \top_I.branch[12].block[4].um_I.ana[5] ;
 wire \top_I.branch[12].block[4].um_I.ana[6] ;
 wire \top_I.branch[12].block[4].um_I.ana[7] ;
 wire \top_I.branch[12].block[4].um_I.clk ;
 wire \top_I.branch[12].block[4].um_I.ena ;
 wire \top_I.branch[12].block[4].um_I.iw[10] ;
 wire \top_I.branch[12].block[4].um_I.iw[11] ;
 wire \top_I.branch[12].block[4].um_I.iw[12] ;
 wire \top_I.branch[12].block[4].um_I.iw[13] ;
 wire \top_I.branch[12].block[4].um_I.iw[14] ;
 wire \top_I.branch[12].block[4].um_I.iw[15] ;
 wire \top_I.branch[12].block[4].um_I.iw[16] ;
 wire \top_I.branch[12].block[4].um_I.iw[17] ;
 wire \top_I.branch[12].block[4].um_I.iw[1] ;
 wire \top_I.branch[12].block[4].um_I.iw[2] ;
 wire \top_I.branch[12].block[4].um_I.iw[3] ;
 wire \top_I.branch[12].block[4].um_I.iw[4] ;
 wire \top_I.branch[12].block[4].um_I.iw[5] ;
 wire \top_I.branch[12].block[4].um_I.iw[6] ;
 wire \top_I.branch[12].block[4].um_I.iw[7] ;
 wire \top_I.branch[12].block[4].um_I.iw[8] ;
 wire \top_I.branch[12].block[4].um_I.iw[9] ;
 wire \top_I.branch[12].block[4].um_I.k_zero ;
 wire \top_I.branch[12].block[4].um_I.pg_vdd ;
 wire \top_I.branch[12].block[5].um_I.ana[0] ;
 wire \top_I.branch[12].block[5].um_I.ana[1] ;
 wire \top_I.branch[12].block[5].um_I.ana[2] ;
 wire \top_I.branch[12].block[5].um_I.ana[3] ;
 wire \top_I.branch[12].block[5].um_I.ana[4] ;
 wire \top_I.branch[12].block[5].um_I.ana[5] ;
 wire \top_I.branch[12].block[5].um_I.ana[6] ;
 wire \top_I.branch[12].block[5].um_I.ana[7] ;
 wire \top_I.branch[12].block[5].um_I.clk ;
 wire \top_I.branch[12].block[5].um_I.ena ;
 wire \top_I.branch[12].block[5].um_I.iw[10] ;
 wire \top_I.branch[12].block[5].um_I.iw[11] ;
 wire \top_I.branch[12].block[5].um_I.iw[12] ;
 wire \top_I.branch[12].block[5].um_I.iw[13] ;
 wire \top_I.branch[12].block[5].um_I.iw[14] ;
 wire \top_I.branch[12].block[5].um_I.iw[15] ;
 wire \top_I.branch[12].block[5].um_I.iw[16] ;
 wire \top_I.branch[12].block[5].um_I.iw[17] ;
 wire \top_I.branch[12].block[5].um_I.iw[1] ;
 wire \top_I.branch[12].block[5].um_I.iw[2] ;
 wire \top_I.branch[12].block[5].um_I.iw[3] ;
 wire \top_I.branch[12].block[5].um_I.iw[4] ;
 wire \top_I.branch[12].block[5].um_I.iw[5] ;
 wire \top_I.branch[12].block[5].um_I.iw[6] ;
 wire \top_I.branch[12].block[5].um_I.iw[7] ;
 wire \top_I.branch[12].block[5].um_I.iw[8] ;
 wire \top_I.branch[12].block[5].um_I.iw[9] ;
 wire \top_I.branch[12].block[5].um_I.k_zero ;
 wire \top_I.branch[12].block[5].um_I.pg_vdd ;
 wire \top_I.branch[12].block[6].um_I.ana[0] ;
 wire \top_I.branch[12].block[6].um_I.ana[1] ;
 wire \top_I.branch[12].block[6].um_I.ana[2] ;
 wire \top_I.branch[12].block[6].um_I.ana[3] ;
 wire \top_I.branch[12].block[6].um_I.ana[4] ;
 wire \top_I.branch[12].block[6].um_I.ana[5] ;
 wire \top_I.branch[12].block[6].um_I.ana[6] ;
 wire \top_I.branch[12].block[6].um_I.ana[7] ;
 wire \top_I.branch[12].block[6].um_I.clk ;
 wire \top_I.branch[12].block[6].um_I.ena ;
 wire \top_I.branch[12].block[6].um_I.iw[10] ;
 wire \top_I.branch[12].block[6].um_I.iw[11] ;
 wire \top_I.branch[12].block[6].um_I.iw[12] ;
 wire \top_I.branch[12].block[6].um_I.iw[13] ;
 wire \top_I.branch[12].block[6].um_I.iw[14] ;
 wire \top_I.branch[12].block[6].um_I.iw[15] ;
 wire \top_I.branch[12].block[6].um_I.iw[16] ;
 wire \top_I.branch[12].block[6].um_I.iw[17] ;
 wire \top_I.branch[12].block[6].um_I.iw[1] ;
 wire \top_I.branch[12].block[6].um_I.iw[2] ;
 wire \top_I.branch[12].block[6].um_I.iw[3] ;
 wire \top_I.branch[12].block[6].um_I.iw[4] ;
 wire \top_I.branch[12].block[6].um_I.iw[5] ;
 wire \top_I.branch[12].block[6].um_I.iw[6] ;
 wire \top_I.branch[12].block[6].um_I.iw[7] ;
 wire \top_I.branch[12].block[6].um_I.iw[8] ;
 wire \top_I.branch[12].block[6].um_I.iw[9] ;
 wire \top_I.branch[12].block[6].um_I.k_zero ;
 wire \top_I.branch[12].block[6].um_I.pg_vdd ;
 wire \top_I.branch[12].block[7].um_I.ana[0] ;
 wire \top_I.branch[12].block[7].um_I.ana[1] ;
 wire \top_I.branch[12].block[7].um_I.ana[2] ;
 wire \top_I.branch[12].block[7].um_I.ana[3] ;
 wire \top_I.branch[12].block[7].um_I.ana[4] ;
 wire \top_I.branch[12].block[7].um_I.ana[5] ;
 wire \top_I.branch[12].block[7].um_I.ana[6] ;
 wire \top_I.branch[12].block[7].um_I.ana[7] ;
 wire \top_I.branch[12].block[7].um_I.clk ;
 wire \top_I.branch[12].block[7].um_I.ena ;
 wire \top_I.branch[12].block[7].um_I.iw[10] ;
 wire \top_I.branch[12].block[7].um_I.iw[11] ;
 wire \top_I.branch[12].block[7].um_I.iw[12] ;
 wire \top_I.branch[12].block[7].um_I.iw[13] ;
 wire \top_I.branch[12].block[7].um_I.iw[14] ;
 wire \top_I.branch[12].block[7].um_I.iw[15] ;
 wire \top_I.branch[12].block[7].um_I.iw[16] ;
 wire \top_I.branch[12].block[7].um_I.iw[17] ;
 wire \top_I.branch[12].block[7].um_I.iw[1] ;
 wire \top_I.branch[12].block[7].um_I.iw[2] ;
 wire \top_I.branch[12].block[7].um_I.iw[3] ;
 wire \top_I.branch[12].block[7].um_I.iw[4] ;
 wire \top_I.branch[12].block[7].um_I.iw[5] ;
 wire \top_I.branch[12].block[7].um_I.iw[6] ;
 wire \top_I.branch[12].block[7].um_I.iw[7] ;
 wire \top_I.branch[12].block[7].um_I.iw[8] ;
 wire \top_I.branch[12].block[7].um_I.iw[9] ;
 wire \top_I.branch[12].block[7].um_I.k_zero ;
 wire \top_I.branch[12].block[7].um_I.pg_vdd ;
 wire \top_I.branch[12].block[8].um_I.ana[0] ;
 wire \top_I.branch[12].block[8].um_I.ana[1] ;
 wire \top_I.branch[12].block[8].um_I.ana[2] ;
 wire \top_I.branch[12].block[8].um_I.ana[3] ;
 wire \top_I.branch[12].block[8].um_I.ana[4] ;
 wire \top_I.branch[12].block[8].um_I.ana[5] ;
 wire \top_I.branch[12].block[8].um_I.ana[6] ;
 wire \top_I.branch[12].block[8].um_I.ana[7] ;
 wire \top_I.branch[12].block[8].um_I.clk ;
 wire \top_I.branch[12].block[8].um_I.ena ;
 wire \top_I.branch[12].block[8].um_I.iw[10] ;
 wire \top_I.branch[12].block[8].um_I.iw[11] ;
 wire \top_I.branch[12].block[8].um_I.iw[12] ;
 wire \top_I.branch[12].block[8].um_I.iw[13] ;
 wire \top_I.branch[12].block[8].um_I.iw[14] ;
 wire \top_I.branch[12].block[8].um_I.iw[15] ;
 wire \top_I.branch[12].block[8].um_I.iw[16] ;
 wire \top_I.branch[12].block[8].um_I.iw[17] ;
 wire \top_I.branch[12].block[8].um_I.iw[1] ;
 wire \top_I.branch[12].block[8].um_I.iw[2] ;
 wire \top_I.branch[12].block[8].um_I.iw[3] ;
 wire \top_I.branch[12].block[8].um_I.iw[4] ;
 wire \top_I.branch[12].block[8].um_I.iw[5] ;
 wire \top_I.branch[12].block[8].um_I.iw[6] ;
 wire \top_I.branch[12].block[8].um_I.iw[7] ;
 wire \top_I.branch[12].block[8].um_I.iw[8] ;
 wire \top_I.branch[12].block[8].um_I.iw[9] ;
 wire \top_I.branch[12].block[8].um_I.k_zero ;
 wire \top_I.branch[12].block[8].um_I.pg_vdd ;
 wire \top_I.branch[12].block[9].um_I.ana[0] ;
 wire \top_I.branch[12].block[9].um_I.ana[1] ;
 wire \top_I.branch[12].block[9].um_I.ana[2] ;
 wire \top_I.branch[12].block[9].um_I.ana[3] ;
 wire \top_I.branch[12].block[9].um_I.ana[4] ;
 wire \top_I.branch[12].block[9].um_I.ana[5] ;
 wire \top_I.branch[12].block[9].um_I.ana[6] ;
 wire \top_I.branch[12].block[9].um_I.ana[7] ;
 wire \top_I.branch[12].block[9].um_I.clk ;
 wire \top_I.branch[12].block[9].um_I.ena ;
 wire \top_I.branch[12].block[9].um_I.iw[10] ;
 wire \top_I.branch[12].block[9].um_I.iw[11] ;
 wire \top_I.branch[12].block[9].um_I.iw[12] ;
 wire \top_I.branch[12].block[9].um_I.iw[13] ;
 wire \top_I.branch[12].block[9].um_I.iw[14] ;
 wire \top_I.branch[12].block[9].um_I.iw[15] ;
 wire \top_I.branch[12].block[9].um_I.iw[16] ;
 wire \top_I.branch[12].block[9].um_I.iw[17] ;
 wire \top_I.branch[12].block[9].um_I.iw[1] ;
 wire \top_I.branch[12].block[9].um_I.iw[2] ;
 wire \top_I.branch[12].block[9].um_I.iw[3] ;
 wire \top_I.branch[12].block[9].um_I.iw[4] ;
 wire \top_I.branch[12].block[9].um_I.iw[5] ;
 wire \top_I.branch[12].block[9].um_I.iw[6] ;
 wire \top_I.branch[12].block[9].um_I.iw[7] ;
 wire \top_I.branch[12].block[9].um_I.iw[8] ;
 wire \top_I.branch[12].block[9].um_I.iw[9] ;
 wire \top_I.branch[12].block[9].um_I.k_zero ;
 wire \top_I.branch[12].block[9].um_I.pg_vdd ;
 wire \top_I.branch[12].l_addr[0] ;
 wire \top_I.branch[12].l_addr[1] ;
 wire \top_I.branch[13].block[0].um_I.ana[0] ;
 wire \top_I.branch[13].block[0].um_I.ana[1] ;
 wire \top_I.branch[13].block[0].um_I.ana[2] ;
 wire \top_I.branch[13].block[0].um_I.ana[3] ;
 wire \top_I.branch[13].block[0].um_I.ana[4] ;
 wire \top_I.branch[13].block[0].um_I.ana[5] ;
 wire \top_I.branch[13].block[0].um_I.ana[6] ;
 wire \top_I.branch[13].block[0].um_I.ana[7] ;
 wire \top_I.branch[13].block[0].um_I.clk ;
 wire \top_I.branch[13].block[0].um_I.ena ;
 wire \top_I.branch[13].block[0].um_I.iw[10] ;
 wire \top_I.branch[13].block[0].um_I.iw[11] ;
 wire \top_I.branch[13].block[0].um_I.iw[12] ;
 wire \top_I.branch[13].block[0].um_I.iw[13] ;
 wire \top_I.branch[13].block[0].um_I.iw[14] ;
 wire \top_I.branch[13].block[0].um_I.iw[15] ;
 wire \top_I.branch[13].block[0].um_I.iw[16] ;
 wire \top_I.branch[13].block[0].um_I.iw[17] ;
 wire \top_I.branch[13].block[0].um_I.iw[1] ;
 wire \top_I.branch[13].block[0].um_I.iw[2] ;
 wire \top_I.branch[13].block[0].um_I.iw[3] ;
 wire \top_I.branch[13].block[0].um_I.iw[4] ;
 wire \top_I.branch[13].block[0].um_I.iw[5] ;
 wire \top_I.branch[13].block[0].um_I.iw[6] ;
 wire \top_I.branch[13].block[0].um_I.iw[7] ;
 wire \top_I.branch[13].block[0].um_I.iw[8] ;
 wire \top_I.branch[13].block[0].um_I.iw[9] ;
 wire \top_I.branch[13].block[0].um_I.k_zero ;
 wire \top_I.branch[13].block[0].um_I.pg_vdd ;
 wire \top_I.branch[13].block[10].um_I.ana[0] ;
 wire \top_I.branch[13].block[10].um_I.ana[1] ;
 wire \top_I.branch[13].block[10].um_I.ana[2] ;
 wire \top_I.branch[13].block[10].um_I.ana[3] ;
 wire \top_I.branch[13].block[10].um_I.ana[4] ;
 wire \top_I.branch[13].block[10].um_I.ana[5] ;
 wire \top_I.branch[13].block[10].um_I.ana[6] ;
 wire \top_I.branch[13].block[10].um_I.ana[7] ;
 wire \top_I.branch[13].block[10].um_I.clk ;
 wire \top_I.branch[13].block[10].um_I.ena ;
 wire \top_I.branch[13].block[10].um_I.iw[10] ;
 wire \top_I.branch[13].block[10].um_I.iw[11] ;
 wire \top_I.branch[13].block[10].um_I.iw[12] ;
 wire \top_I.branch[13].block[10].um_I.iw[13] ;
 wire \top_I.branch[13].block[10].um_I.iw[14] ;
 wire \top_I.branch[13].block[10].um_I.iw[15] ;
 wire \top_I.branch[13].block[10].um_I.iw[16] ;
 wire \top_I.branch[13].block[10].um_I.iw[17] ;
 wire \top_I.branch[13].block[10].um_I.iw[1] ;
 wire \top_I.branch[13].block[10].um_I.iw[2] ;
 wire \top_I.branch[13].block[10].um_I.iw[3] ;
 wire \top_I.branch[13].block[10].um_I.iw[4] ;
 wire \top_I.branch[13].block[10].um_I.iw[5] ;
 wire \top_I.branch[13].block[10].um_I.iw[6] ;
 wire \top_I.branch[13].block[10].um_I.iw[7] ;
 wire \top_I.branch[13].block[10].um_I.iw[8] ;
 wire \top_I.branch[13].block[10].um_I.iw[9] ;
 wire \top_I.branch[13].block[10].um_I.k_zero ;
 wire \top_I.branch[13].block[10].um_I.pg_vdd ;
 wire \top_I.branch[13].block[11].um_I.ana[0] ;
 wire \top_I.branch[13].block[11].um_I.ana[1] ;
 wire \top_I.branch[13].block[11].um_I.ana[2] ;
 wire \top_I.branch[13].block[11].um_I.ana[3] ;
 wire \top_I.branch[13].block[11].um_I.ana[4] ;
 wire \top_I.branch[13].block[11].um_I.ana[5] ;
 wire \top_I.branch[13].block[11].um_I.ana[6] ;
 wire \top_I.branch[13].block[11].um_I.ana[7] ;
 wire \top_I.branch[13].block[11].um_I.clk ;
 wire \top_I.branch[13].block[11].um_I.ena ;
 wire \top_I.branch[13].block[11].um_I.iw[10] ;
 wire \top_I.branch[13].block[11].um_I.iw[11] ;
 wire \top_I.branch[13].block[11].um_I.iw[12] ;
 wire \top_I.branch[13].block[11].um_I.iw[13] ;
 wire \top_I.branch[13].block[11].um_I.iw[14] ;
 wire \top_I.branch[13].block[11].um_I.iw[15] ;
 wire \top_I.branch[13].block[11].um_I.iw[16] ;
 wire \top_I.branch[13].block[11].um_I.iw[17] ;
 wire \top_I.branch[13].block[11].um_I.iw[1] ;
 wire \top_I.branch[13].block[11].um_I.iw[2] ;
 wire \top_I.branch[13].block[11].um_I.iw[3] ;
 wire \top_I.branch[13].block[11].um_I.iw[4] ;
 wire \top_I.branch[13].block[11].um_I.iw[5] ;
 wire \top_I.branch[13].block[11].um_I.iw[6] ;
 wire \top_I.branch[13].block[11].um_I.iw[7] ;
 wire \top_I.branch[13].block[11].um_I.iw[8] ;
 wire \top_I.branch[13].block[11].um_I.iw[9] ;
 wire \top_I.branch[13].block[11].um_I.k_zero ;
 wire \top_I.branch[13].block[11].um_I.pg_vdd ;
 wire \top_I.branch[13].block[12].um_I.ana[0] ;
 wire \top_I.branch[13].block[12].um_I.ana[1] ;
 wire \top_I.branch[13].block[12].um_I.ana[2] ;
 wire \top_I.branch[13].block[12].um_I.ana[3] ;
 wire \top_I.branch[13].block[12].um_I.ana[4] ;
 wire \top_I.branch[13].block[12].um_I.ana[5] ;
 wire \top_I.branch[13].block[12].um_I.ana[6] ;
 wire \top_I.branch[13].block[12].um_I.ana[7] ;
 wire \top_I.branch[13].block[12].um_I.clk ;
 wire \top_I.branch[13].block[12].um_I.ena ;
 wire \top_I.branch[13].block[12].um_I.iw[10] ;
 wire \top_I.branch[13].block[12].um_I.iw[11] ;
 wire \top_I.branch[13].block[12].um_I.iw[12] ;
 wire \top_I.branch[13].block[12].um_I.iw[13] ;
 wire \top_I.branch[13].block[12].um_I.iw[14] ;
 wire \top_I.branch[13].block[12].um_I.iw[15] ;
 wire \top_I.branch[13].block[12].um_I.iw[16] ;
 wire \top_I.branch[13].block[12].um_I.iw[17] ;
 wire \top_I.branch[13].block[12].um_I.iw[1] ;
 wire \top_I.branch[13].block[12].um_I.iw[2] ;
 wire \top_I.branch[13].block[12].um_I.iw[3] ;
 wire \top_I.branch[13].block[12].um_I.iw[4] ;
 wire \top_I.branch[13].block[12].um_I.iw[5] ;
 wire \top_I.branch[13].block[12].um_I.iw[6] ;
 wire \top_I.branch[13].block[12].um_I.iw[7] ;
 wire \top_I.branch[13].block[12].um_I.iw[8] ;
 wire \top_I.branch[13].block[12].um_I.iw[9] ;
 wire \top_I.branch[13].block[12].um_I.k_zero ;
 wire \top_I.branch[13].block[12].um_I.pg_vdd ;
 wire \top_I.branch[13].block[13].um_I.ana[0] ;
 wire \top_I.branch[13].block[13].um_I.ana[1] ;
 wire \top_I.branch[13].block[13].um_I.ana[2] ;
 wire \top_I.branch[13].block[13].um_I.ana[3] ;
 wire \top_I.branch[13].block[13].um_I.ana[4] ;
 wire \top_I.branch[13].block[13].um_I.ana[5] ;
 wire \top_I.branch[13].block[13].um_I.ana[6] ;
 wire \top_I.branch[13].block[13].um_I.ana[7] ;
 wire \top_I.branch[13].block[13].um_I.clk ;
 wire \top_I.branch[13].block[13].um_I.ena ;
 wire \top_I.branch[13].block[13].um_I.iw[10] ;
 wire \top_I.branch[13].block[13].um_I.iw[11] ;
 wire \top_I.branch[13].block[13].um_I.iw[12] ;
 wire \top_I.branch[13].block[13].um_I.iw[13] ;
 wire \top_I.branch[13].block[13].um_I.iw[14] ;
 wire \top_I.branch[13].block[13].um_I.iw[15] ;
 wire \top_I.branch[13].block[13].um_I.iw[16] ;
 wire \top_I.branch[13].block[13].um_I.iw[17] ;
 wire \top_I.branch[13].block[13].um_I.iw[1] ;
 wire \top_I.branch[13].block[13].um_I.iw[2] ;
 wire \top_I.branch[13].block[13].um_I.iw[3] ;
 wire \top_I.branch[13].block[13].um_I.iw[4] ;
 wire \top_I.branch[13].block[13].um_I.iw[5] ;
 wire \top_I.branch[13].block[13].um_I.iw[6] ;
 wire \top_I.branch[13].block[13].um_I.iw[7] ;
 wire \top_I.branch[13].block[13].um_I.iw[8] ;
 wire \top_I.branch[13].block[13].um_I.iw[9] ;
 wire \top_I.branch[13].block[13].um_I.k_zero ;
 wire \top_I.branch[13].block[13].um_I.pg_vdd ;
 wire \top_I.branch[13].block[14].um_I.ana[0] ;
 wire \top_I.branch[13].block[14].um_I.ana[1] ;
 wire \top_I.branch[13].block[14].um_I.ana[2] ;
 wire \top_I.branch[13].block[14].um_I.ana[3] ;
 wire \top_I.branch[13].block[14].um_I.ana[4] ;
 wire \top_I.branch[13].block[14].um_I.ana[5] ;
 wire \top_I.branch[13].block[14].um_I.ana[6] ;
 wire \top_I.branch[13].block[14].um_I.ana[7] ;
 wire \top_I.branch[13].block[14].um_I.clk ;
 wire \top_I.branch[13].block[14].um_I.ena ;
 wire \top_I.branch[13].block[14].um_I.iw[10] ;
 wire \top_I.branch[13].block[14].um_I.iw[11] ;
 wire \top_I.branch[13].block[14].um_I.iw[12] ;
 wire \top_I.branch[13].block[14].um_I.iw[13] ;
 wire \top_I.branch[13].block[14].um_I.iw[14] ;
 wire \top_I.branch[13].block[14].um_I.iw[15] ;
 wire \top_I.branch[13].block[14].um_I.iw[16] ;
 wire \top_I.branch[13].block[14].um_I.iw[17] ;
 wire \top_I.branch[13].block[14].um_I.iw[1] ;
 wire \top_I.branch[13].block[14].um_I.iw[2] ;
 wire \top_I.branch[13].block[14].um_I.iw[3] ;
 wire \top_I.branch[13].block[14].um_I.iw[4] ;
 wire \top_I.branch[13].block[14].um_I.iw[5] ;
 wire \top_I.branch[13].block[14].um_I.iw[6] ;
 wire \top_I.branch[13].block[14].um_I.iw[7] ;
 wire \top_I.branch[13].block[14].um_I.iw[8] ;
 wire \top_I.branch[13].block[14].um_I.iw[9] ;
 wire \top_I.branch[13].block[14].um_I.k_zero ;
 wire \top_I.branch[13].block[14].um_I.pg_vdd ;
 wire \top_I.branch[13].block[15].um_I.ana[0] ;
 wire \top_I.branch[13].block[15].um_I.ana[1] ;
 wire \top_I.branch[13].block[15].um_I.ana[2] ;
 wire \top_I.branch[13].block[15].um_I.ana[3] ;
 wire \top_I.branch[13].block[15].um_I.ana[4] ;
 wire \top_I.branch[13].block[15].um_I.ana[5] ;
 wire \top_I.branch[13].block[15].um_I.ana[6] ;
 wire \top_I.branch[13].block[15].um_I.ana[7] ;
 wire \top_I.branch[13].block[15].um_I.clk ;
 wire \top_I.branch[13].block[15].um_I.ena ;
 wire \top_I.branch[13].block[15].um_I.iw[10] ;
 wire \top_I.branch[13].block[15].um_I.iw[11] ;
 wire \top_I.branch[13].block[15].um_I.iw[12] ;
 wire \top_I.branch[13].block[15].um_I.iw[13] ;
 wire \top_I.branch[13].block[15].um_I.iw[14] ;
 wire \top_I.branch[13].block[15].um_I.iw[15] ;
 wire \top_I.branch[13].block[15].um_I.iw[16] ;
 wire \top_I.branch[13].block[15].um_I.iw[17] ;
 wire \top_I.branch[13].block[15].um_I.iw[1] ;
 wire \top_I.branch[13].block[15].um_I.iw[2] ;
 wire \top_I.branch[13].block[15].um_I.iw[3] ;
 wire \top_I.branch[13].block[15].um_I.iw[4] ;
 wire \top_I.branch[13].block[15].um_I.iw[5] ;
 wire \top_I.branch[13].block[15].um_I.iw[6] ;
 wire \top_I.branch[13].block[15].um_I.iw[7] ;
 wire \top_I.branch[13].block[15].um_I.iw[8] ;
 wire \top_I.branch[13].block[15].um_I.iw[9] ;
 wire \top_I.branch[13].block[15].um_I.k_zero ;
 wire \top_I.branch[13].block[15].um_I.pg_vdd ;
 wire \top_I.branch[13].block[1].um_I.ana[0] ;
 wire \top_I.branch[13].block[1].um_I.ana[1] ;
 wire \top_I.branch[13].block[1].um_I.ana[2] ;
 wire \top_I.branch[13].block[1].um_I.ana[3] ;
 wire \top_I.branch[13].block[1].um_I.ana[4] ;
 wire \top_I.branch[13].block[1].um_I.ana[5] ;
 wire \top_I.branch[13].block[1].um_I.ana[6] ;
 wire \top_I.branch[13].block[1].um_I.ana[7] ;
 wire \top_I.branch[13].block[1].um_I.clk ;
 wire \top_I.branch[13].block[1].um_I.ena ;
 wire \top_I.branch[13].block[1].um_I.iw[10] ;
 wire \top_I.branch[13].block[1].um_I.iw[11] ;
 wire \top_I.branch[13].block[1].um_I.iw[12] ;
 wire \top_I.branch[13].block[1].um_I.iw[13] ;
 wire \top_I.branch[13].block[1].um_I.iw[14] ;
 wire \top_I.branch[13].block[1].um_I.iw[15] ;
 wire \top_I.branch[13].block[1].um_I.iw[16] ;
 wire \top_I.branch[13].block[1].um_I.iw[17] ;
 wire \top_I.branch[13].block[1].um_I.iw[1] ;
 wire \top_I.branch[13].block[1].um_I.iw[2] ;
 wire \top_I.branch[13].block[1].um_I.iw[3] ;
 wire \top_I.branch[13].block[1].um_I.iw[4] ;
 wire \top_I.branch[13].block[1].um_I.iw[5] ;
 wire \top_I.branch[13].block[1].um_I.iw[6] ;
 wire \top_I.branch[13].block[1].um_I.iw[7] ;
 wire \top_I.branch[13].block[1].um_I.iw[8] ;
 wire \top_I.branch[13].block[1].um_I.iw[9] ;
 wire \top_I.branch[13].block[1].um_I.k_zero ;
 wire \top_I.branch[13].block[1].um_I.pg_vdd ;
 wire \top_I.branch[13].block[2].um_I.ana[0] ;
 wire \top_I.branch[13].block[2].um_I.ana[1] ;
 wire \top_I.branch[13].block[2].um_I.ana[2] ;
 wire \top_I.branch[13].block[2].um_I.ana[3] ;
 wire \top_I.branch[13].block[2].um_I.ana[4] ;
 wire \top_I.branch[13].block[2].um_I.ana[5] ;
 wire \top_I.branch[13].block[2].um_I.ana[6] ;
 wire \top_I.branch[13].block[2].um_I.ana[7] ;
 wire \top_I.branch[13].block[2].um_I.clk ;
 wire \top_I.branch[13].block[2].um_I.ena ;
 wire \top_I.branch[13].block[2].um_I.iw[10] ;
 wire \top_I.branch[13].block[2].um_I.iw[11] ;
 wire \top_I.branch[13].block[2].um_I.iw[12] ;
 wire \top_I.branch[13].block[2].um_I.iw[13] ;
 wire \top_I.branch[13].block[2].um_I.iw[14] ;
 wire \top_I.branch[13].block[2].um_I.iw[15] ;
 wire \top_I.branch[13].block[2].um_I.iw[16] ;
 wire \top_I.branch[13].block[2].um_I.iw[17] ;
 wire \top_I.branch[13].block[2].um_I.iw[1] ;
 wire \top_I.branch[13].block[2].um_I.iw[2] ;
 wire \top_I.branch[13].block[2].um_I.iw[3] ;
 wire \top_I.branch[13].block[2].um_I.iw[4] ;
 wire \top_I.branch[13].block[2].um_I.iw[5] ;
 wire \top_I.branch[13].block[2].um_I.iw[6] ;
 wire \top_I.branch[13].block[2].um_I.iw[7] ;
 wire \top_I.branch[13].block[2].um_I.iw[8] ;
 wire \top_I.branch[13].block[2].um_I.iw[9] ;
 wire \top_I.branch[13].block[2].um_I.k_zero ;
 wire \top_I.branch[13].block[2].um_I.pg_vdd ;
 wire \top_I.branch[13].block[3].um_I.ana[0] ;
 wire \top_I.branch[13].block[3].um_I.ana[1] ;
 wire \top_I.branch[13].block[3].um_I.ana[2] ;
 wire \top_I.branch[13].block[3].um_I.ana[3] ;
 wire \top_I.branch[13].block[3].um_I.ana[4] ;
 wire \top_I.branch[13].block[3].um_I.ana[5] ;
 wire \top_I.branch[13].block[3].um_I.ana[6] ;
 wire \top_I.branch[13].block[3].um_I.ana[7] ;
 wire \top_I.branch[13].block[3].um_I.clk ;
 wire \top_I.branch[13].block[3].um_I.ena ;
 wire \top_I.branch[13].block[3].um_I.iw[10] ;
 wire \top_I.branch[13].block[3].um_I.iw[11] ;
 wire \top_I.branch[13].block[3].um_I.iw[12] ;
 wire \top_I.branch[13].block[3].um_I.iw[13] ;
 wire \top_I.branch[13].block[3].um_I.iw[14] ;
 wire \top_I.branch[13].block[3].um_I.iw[15] ;
 wire \top_I.branch[13].block[3].um_I.iw[16] ;
 wire \top_I.branch[13].block[3].um_I.iw[17] ;
 wire \top_I.branch[13].block[3].um_I.iw[1] ;
 wire \top_I.branch[13].block[3].um_I.iw[2] ;
 wire \top_I.branch[13].block[3].um_I.iw[3] ;
 wire \top_I.branch[13].block[3].um_I.iw[4] ;
 wire \top_I.branch[13].block[3].um_I.iw[5] ;
 wire \top_I.branch[13].block[3].um_I.iw[6] ;
 wire \top_I.branch[13].block[3].um_I.iw[7] ;
 wire \top_I.branch[13].block[3].um_I.iw[8] ;
 wire \top_I.branch[13].block[3].um_I.iw[9] ;
 wire \top_I.branch[13].block[3].um_I.k_zero ;
 wire \top_I.branch[13].block[3].um_I.pg_vdd ;
 wire \top_I.branch[13].block[4].um_I.ana[0] ;
 wire \top_I.branch[13].block[4].um_I.ana[1] ;
 wire \top_I.branch[13].block[4].um_I.ana[2] ;
 wire \top_I.branch[13].block[4].um_I.ana[3] ;
 wire \top_I.branch[13].block[4].um_I.ana[4] ;
 wire \top_I.branch[13].block[4].um_I.ana[5] ;
 wire \top_I.branch[13].block[4].um_I.ana[6] ;
 wire \top_I.branch[13].block[4].um_I.ana[7] ;
 wire \top_I.branch[13].block[4].um_I.clk ;
 wire \top_I.branch[13].block[4].um_I.ena ;
 wire \top_I.branch[13].block[4].um_I.iw[10] ;
 wire \top_I.branch[13].block[4].um_I.iw[11] ;
 wire \top_I.branch[13].block[4].um_I.iw[12] ;
 wire \top_I.branch[13].block[4].um_I.iw[13] ;
 wire \top_I.branch[13].block[4].um_I.iw[14] ;
 wire \top_I.branch[13].block[4].um_I.iw[15] ;
 wire \top_I.branch[13].block[4].um_I.iw[16] ;
 wire \top_I.branch[13].block[4].um_I.iw[17] ;
 wire \top_I.branch[13].block[4].um_I.iw[1] ;
 wire \top_I.branch[13].block[4].um_I.iw[2] ;
 wire \top_I.branch[13].block[4].um_I.iw[3] ;
 wire \top_I.branch[13].block[4].um_I.iw[4] ;
 wire \top_I.branch[13].block[4].um_I.iw[5] ;
 wire \top_I.branch[13].block[4].um_I.iw[6] ;
 wire \top_I.branch[13].block[4].um_I.iw[7] ;
 wire \top_I.branch[13].block[4].um_I.iw[8] ;
 wire \top_I.branch[13].block[4].um_I.iw[9] ;
 wire \top_I.branch[13].block[4].um_I.k_zero ;
 wire \top_I.branch[13].block[4].um_I.pg_vdd ;
 wire \top_I.branch[13].block[5].um_I.ana[0] ;
 wire \top_I.branch[13].block[5].um_I.ana[1] ;
 wire \top_I.branch[13].block[5].um_I.ana[2] ;
 wire \top_I.branch[13].block[5].um_I.ana[3] ;
 wire \top_I.branch[13].block[5].um_I.ana[4] ;
 wire \top_I.branch[13].block[5].um_I.ana[5] ;
 wire \top_I.branch[13].block[5].um_I.ana[6] ;
 wire \top_I.branch[13].block[5].um_I.ana[7] ;
 wire \top_I.branch[13].block[5].um_I.clk ;
 wire \top_I.branch[13].block[5].um_I.ena ;
 wire \top_I.branch[13].block[5].um_I.iw[10] ;
 wire \top_I.branch[13].block[5].um_I.iw[11] ;
 wire \top_I.branch[13].block[5].um_I.iw[12] ;
 wire \top_I.branch[13].block[5].um_I.iw[13] ;
 wire \top_I.branch[13].block[5].um_I.iw[14] ;
 wire \top_I.branch[13].block[5].um_I.iw[15] ;
 wire \top_I.branch[13].block[5].um_I.iw[16] ;
 wire \top_I.branch[13].block[5].um_I.iw[17] ;
 wire \top_I.branch[13].block[5].um_I.iw[1] ;
 wire \top_I.branch[13].block[5].um_I.iw[2] ;
 wire \top_I.branch[13].block[5].um_I.iw[3] ;
 wire \top_I.branch[13].block[5].um_I.iw[4] ;
 wire \top_I.branch[13].block[5].um_I.iw[5] ;
 wire \top_I.branch[13].block[5].um_I.iw[6] ;
 wire \top_I.branch[13].block[5].um_I.iw[7] ;
 wire \top_I.branch[13].block[5].um_I.iw[8] ;
 wire \top_I.branch[13].block[5].um_I.iw[9] ;
 wire \top_I.branch[13].block[5].um_I.k_zero ;
 wire \top_I.branch[13].block[5].um_I.pg_vdd ;
 wire \top_I.branch[13].block[6].um_I.ana[0] ;
 wire \top_I.branch[13].block[6].um_I.ana[1] ;
 wire \top_I.branch[13].block[6].um_I.ana[2] ;
 wire \top_I.branch[13].block[6].um_I.ana[3] ;
 wire \top_I.branch[13].block[6].um_I.ana[4] ;
 wire \top_I.branch[13].block[6].um_I.ana[5] ;
 wire \top_I.branch[13].block[6].um_I.ana[6] ;
 wire \top_I.branch[13].block[6].um_I.ana[7] ;
 wire \top_I.branch[13].block[6].um_I.clk ;
 wire \top_I.branch[13].block[6].um_I.ena ;
 wire \top_I.branch[13].block[6].um_I.iw[10] ;
 wire \top_I.branch[13].block[6].um_I.iw[11] ;
 wire \top_I.branch[13].block[6].um_I.iw[12] ;
 wire \top_I.branch[13].block[6].um_I.iw[13] ;
 wire \top_I.branch[13].block[6].um_I.iw[14] ;
 wire \top_I.branch[13].block[6].um_I.iw[15] ;
 wire \top_I.branch[13].block[6].um_I.iw[16] ;
 wire \top_I.branch[13].block[6].um_I.iw[17] ;
 wire \top_I.branch[13].block[6].um_I.iw[1] ;
 wire \top_I.branch[13].block[6].um_I.iw[2] ;
 wire \top_I.branch[13].block[6].um_I.iw[3] ;
 wire \top_I.branch[13].block[6].um_I.iw[4] ;
 wire \top_I.branch[13].block[6].um_I.iw[5] ;
 wire \top_I.branch[13].block[6].um_I.iw[6] ;
 wire \top_I.branch[13].block[6].um_I.iw[7] ;
 wire \top_I.branch[13].block[6].um_I.iw[8] ;
 wire \top_I.branch[13].block[6].um_I.iw[9] ;
 wire \top_I.branch[13].block[6].um_I.k_zero ;
 wire \top_I.branch[13].block[6].um_I.pg_vdd ;
 wire \top_I.branch[13].block[7].um_I.ana[0] ;
 wire \top_I.branch[13].block[7].um_I.ana[1] ;
 wire \top_I.branch[13].block[7].um_I.ana[2] ;
 wire \top_I.branch[13].block[7].um_I.ana[3] ;
 wire \top_I.branch[13].block[7].um_I.ana[4] ;
 wire \top_I.branch[13].block[7].um_I.ana[5] ;
 wire \top_I.branch[13].block[7].um_I.ana[6] ;
 wire \top_I.branch[13].block[7].um_I.ana[7] ;
 wire \top_I.branch[13].block[7].um_I.clk ;
 wire \top_I.branch[13].block[7].um_I.ena ;
 wire \top_I.branch[13].block[7].um_I.iw[10] ;
 wire \top_I.branch[13].block[7].um_I.iw[11] ;
 wire \top_I.branch[13].block[7].um_I.iw[12] ;
 wire \top_I.branch[13].block[7].um_I.iw[13] ;
 wire \top_I.branch[13].block[7].um_I.iw[14] ;
 wire \top_I.branch[13].block[7].um_I.iw[15] ;
 wire \top_I.branch[13].block[7].um_I.iw[16] ;
 wire \top_I.branch[13].block[7].um_I.iw[17] ;
 wire \top_I.branch[13].block[7].um_I.iw[1] ;
 wire \top_I.branch[13].block[7].um_I.iw[2] ;
 wire \top_I.branch[13].block[7].um_I.iw[3] ;
 wire \top_I.branch[13].block[7].um_I.iw[4] ;
 wire \top_I.branch[13].block[7].um_I.iw[5] ;
 wire \top_I.branch[13].block[7].um_I.iw[6] ;
 wire \top_I.branch[13].block[7].um_I.iw[7] ;
 wire \top_I.branch[13].block[7].um_I.iw[8] ;
 wire \top_I.branch[13].block[7].um_I.iw[9] ;
 wire \top_I.branch[13].block[7].um_I.k_zero ;
 wire \top_I.branch[13].block[7].um_I.pg_vdd ;
 wire \top_I.branch[13].block[8].um_I.ana[0] ;
 wire \top_I.branch[13].block[8].um_I.ana[1] ;
 wire \top_I.branch[13].block[8].um_I.ana[2] ;
 wire \top_I.branch[13].block[8].um_I.ana[3] ;
 wire \top_I.branch[13].block[8].um_I.ana[4] ;
 wire \top_I.branch[13].block[8].um_I.ana[5] ;
 wire \top_I.branch[13].block[8].um_I.ana[6] ;
 wire \top_I.branch[13].block[8].um_I.ana[7] ;
 wire \top_I.branch[13].block[8].um_I.clk ;
 wire \top_I.branch[13].block[8].um_I.ena ;
 wire \top_I.branch[13].block[8].um_I.iw[10] ;
 wire \top_I.branch[13].block[8].um_I.iw[11] ;
 wire \top_I.branch[13].block[8].um_I.iw[12] ;
 wire \top_I.branch[13].block[8].um_I.iw[13] ;
 wire \top_I.branch[13].block[8].um_I.iw[14] ;
 wire \top_I.branch[13].block[8].um_I.iw[15] ;
 wire \top_I.branch[13].block[8].um_I.iw[16] ;
 wire \top_I.branch[13].block[8].um_I.iw[17] ;
 wire \top_I.branch[13].block[8].um_I.iw[1] ;
 wire \top_I.branch[13].block[8].um_I.iw[2] ;
 wire \top_I.branch[13].block[8].um_I.iw[3] ;
 wire \top_I.branch[13].block[8].um_I.iw[4] ;
 wire \top_I.branch[13].block[8].um_I.iw[5] ;
 wire \top_I.branch[13].block[8].um_I.iw[6] ;
 wire \top_I.branch[13].block[8].um_I.iw[7] ;
 wire \top_I.branch[13].block[8].um_I.iw[8] ;
 wire \top_I.branch[13].block[8].um_I.iw[9] ;
 wire \top_I.branch[13].block[8].um_I.k_zero ;
 wire \top_I.branch[13].block[8].um_I.pg_vdd ;
 wire \top_I.branch[13].block[9].um_I.ana[0] ;
 wire \top_I.branch[13].block[9].um_I.ana[1] ;
 wire \top_I.branch[13].block[9].um_I.ana[2] ;
 wire \top_I.branch[13].block[9].um_I.ana[3] ;
 wire \top_I.branch[13].block[9].um_I.ana[4] ;
 wire \top_I.branch[13].block[9].um_I.ana[5] ;
 wire \top_I.branch[13].block[9].um_I.ana[6] ;
 wire \top_I.branch[13].block[9].um_I.ana[7] ;
 wire \top_I.branch[13].block[9].um_I.clk ;
 wire \top_I.branch[13].block[9].um_I.ena ;
 wire \top_I.branch[13].block[9].um_I.iw[10] ;
 wire \top_I.branch[13].block[9].um_I.iw[11] ;
 wire \top_I.branch[13].block[9].um_I.iw[12] ;
 wire \top_I.branch[13].block[9].um_I.iw[13] ;
 wire \top_I.branch[13].block[9].um_I.iw[14] ;
 wire \top_I.branch[13].block[9].um_I.iw[15] ;
 wire \top_I.branch[13].block[9].um_I.iw[16] ;
 wire \top_I.branch[13].block[9].um_I.iw[17] ;
 wire \top_I.branch[13].block[9].um_I.iw[1] ;
 wire \top_I.branch[13].block[9].um_I.iw[2] ;
 wire \top_I.branch[13].block[9].um_I.iw[3] ;
 wire \top_I.branch[13].block[9].um_I.iw[4] ;
 wire \top_I.branch[13].block[9].um_I.iw[5] ;
 wire \top_I.branch[13].block[9].um_I.iw[6] ;
 wire \top_I.branch[13].block[9].um_I.iw[7] ;
 wire \top_I.branch[13].block[9].um_I.iw[8] ;
 wire \top_I.branch[13].block[9].um_I.iw[9] ;
 wire \top_I.branch[13].block[9].um_I.k_zero ;
 wire \top_I.branch[13].block[9].um_I.pg_vdd ;
 wire \top_I.branch[13].l_addr[0] ;
 wire \top_I.branch[13].l_addr[1] ;
 wire \top_I.branch[14].block[0].um_I.ana[0] ;
 wire \top_I.branch[14].block[0].um_I.ana[1] ;
 wire \top_I.branch[14].block[0].um_I.ana[2] ;
 wire \top_I.branch[14].block[0].um_I.ana[3] ;
 wire \top_I.branch[14].block[0].um_I.ana[4] ;
 wire \top_I.branch[14].block[0].um_I.ana[5] ;
 wire \top_I.branch[14].block[0].um_I.ana[6] ;
 wire \top_I.branch[14].block[0].um_I.ana[7] ;
 wire \top_I.branch[14].block[0].um_I.clk ;
 wire \top_I.branch[14].block[0].um_I.ena ;
 wire \top_I.branch[14].block[0].um_I.iw[10] ;
 wire \top_I.branch[14].block[0].um_I.iw[11] ;
 wire \top_I.branch[14].block[0].um_I.iw[12] ;
 wire \top_I.branch[14].block[0].um_I.iw[13] ;
 wire \top_I.branch[14].block[0].um_I.iw[14] ;
 wire \top_I.branch[14].block[0].um_I.iw[15] ;
 wire \top_I.branch[14].block[0].um_I.iw[16] ;
 wire \top_I.branch[14].block[0].um_I.iw[17] ;
 wire \top_I.branch[14].block[0].um_I.iw[1] ;
 wire \top_I.branch[14].block[0].um_I.iw[2] ;
 wire \top_I.branch[14].block[0].um_I.iw[3] ;
 wire \top_I.branch[14].block[0].um_I.iw[4] ;
 wire \top_I.branch[14].block[0].um_I.iw[5] ;
 wire \top_I.branch[14].block[0].um_I.iw[6] ;
 wire \top_I.branch[14].block[0].um_I.iw[7] ;
 wire \top_I.branch[14].block[0].um_I.iw[8] ;
 wire \top_I.branch[14].block[0].um_I.iw[9] ;
 wire \top_I.branch[14].block[0].um_I.k_zero ;
 wire \top_I.branch[14].block[0].um_I.pg_vdd ;
 wire \top_I.branch[14].block[10].um_I.ana[0] ;
 wire \top_I.branch[14].block[10].um_I.ana[1] ;
 wire \top_I.branch[14].block[10].um_I.ana[2] ;
 wire \top_I.branch[14].block[10].um_I.ana[3] ;
 wire \top_I.branch[14].block[10].um_I.ana[4] ;
 wire \top_I.branch[14].block[10].um_I.ana[5] ;
 wire \top_I.branch[14].block[10].um_I.ana[6] ;
 wire \top_I.branch[14].block[10].um_I.ana[7] ;
 wire \top_I.branch[14].block[10].um_I.clk ;
 wire \top_I.branch[14].block[10].um_I.ena ;
 wire \top_I.branch[14].block[10].um_I.iw[10] ;
 wire \top_I.branch[14].block[10].um_I.iw[11] ;
 wire \top_I.branch[14].block[10].um_I.iw[12] ;
 wire \top_I.branch[14].block[10].um_I.iw[13] ;
 wire \top_I.branch[14].block[10].um_I.iw[14] ;
 wire \top_I.branch[14].block[10].um_I.iw[15] ;
 wire \top_I.branch[14].block[10].um_I.iw[16] ;
 wire \top_I.branch[14].block[10].um_I.iw[17] ;
 wire \top_I.branch[14].block[10].um_I.iw[1] ;
 wire \top_I.branch[14].block[10].um_I.iw[2] ;
 wire \top_I.branch[14].block[10].um_I.iw[3] ;
 wire \top_I.branch[14].block[10].um_I.iw[4] ;
 wire \top_I.branch[14].block[10].um_I.iw[5] ;
 wire \top_I.branch[14].block[10].um_I.iw[6] ;
 wire \top_I.branch[14].block[10].um_I.iw[7] ;
 wire \top_I.branch[14].block[10].um_I.iw[8] ;
 wire \top_I.branch[14].block[10].um_I.iw[9] ;
 wire \top_I.branch[14].block[10].um_I.k_zero ;
 wire \top_I.branch[14].block[10].um_I.pg_vdd ;
 wire \top_I.branch[14].block[11].um_I.ana[0] ;
 wire \top_I.branch[14].block[11].um_I.ana[1] ;
 wire \top_I.branch[14].block[11].um_I.ana[2] ;
 wire \top_I.branch[14].block[11].um_I.ana[3] ;
 wire \top_I.branch[14].block[11].um_I.ana[4] ;
 wire \top_I.branch[14].block[11].um_I.ana[5] ;
 wire \top_I.branch[14].block[11].um_I.ana[6] ;
 wire \top_I.branch[14].block[11].um_I.ana[7] ;
 wire \top_I.branch[14].block[11].um_I.clk ;
 wire \top_I.branch[14].block[11].um_I.ena ;
 wire \top_I.branch[14].block[11].um_I.iw[10] ;
 wire \top_I.branch[14].block[11].um_I.iw[11] ;
 wire \top_I.branch[14].block[11].um_I.iw[12] ;
 wire \top_I.branch[14].block[11].um_I.iw[13] ;
 wire \top_I.branch[14].block[11].um_I.iw[14] ;
 wire \top_I.branch[14].block[11].um_I.iw[15] ;
 wire \top_I.branch[14].block[11].um_I.iw[16] ;
 wire \top_I.branch[14].block[11].um_I.iw[17] ;
 wire \top_I.branch[14].block[11].um_I.iw[1] ;
 wire \top_I.branch[14].block[11].um_I.iw[2] ;
 wire \top_I.branch[14].block[11].um_I.iw[3] ;
 wire \top_I.branch[14].block[11].um_I.iw[4] ;
 wire \top_I.branch[14].block[11].um_I.iw[5] ;
 wire \top_I.branch[14].block[11].um_I.iw[6] ;
 wire \top_I.branch[14].block[11].um_I.iw[7] ;
 wire \top_I.branch[14].block[11].um_I.iw[8] ;
 wire \top_I.branch[14].block[11].um_I.iw[9] ;
 wire \top_I.branch[14].block[11].um_I.k_zero ;
 wire \top_I.branch[14].block[11].um_I.pg_vdd ;
 wire \top_I.branch[14].block[12].um_I.ana[0] ;
 wire \top_I.branch[14].block[12].um_I.ana[1] ;
 wire \top_I.branch[14].block[12].um_I.ana[2] ;
 wire \top_I.branch[14].block[12].um_I.ana[3] ;
 wire \top_I.branch[14].block[12].um_I.ana[4] ;
 wire \top_I.branch[14].block[12].um_I.ana[5] ;
 wire \top_I.branch[14].block[12].um_I.ana[6] ;
 wire \top_I.branch[14].block[12].um_I.ana[7] ;
 wire \top_I.branch[14].block[12].um_I.clk ;
 wire \top_I.branch[14].block[12].um_I.ena ;
 wire \top_I.branch[14].block[12].um_I.iw[10] ;
 wire \top_I.branch[14].block[12].um_I.iw[11] ;
 wire \top_I.branch[14].block[12].um_I.iw[12] ;
 wire \top_I.branch[14].block[12].um_I.iw[13] ;
 wire \top_I.branch[14].block[12].um_I.iw[14] ;
 wire \top_I.branch[14].block[12].um_I.iw[15] ;
 wire \top_I.branch[14].block[12].um_I.iw[16] ;
 wire \top_I.branch[14].block[12].um_I.iw[17] ;
 wire \top_I.branch[14].block[12].um_I.iw[1] ;
 wire \top_I.branch[14].block[12].um_I.iw[2] ;
 wire \top_I.branch[14].block[12].um_I.iw[3] ;
 wire \top_I.branch[14].block[12].um_I.iw[4] ;
 wire \top_I.branch[14].block[12].um_I.iw[5] ;
 wire \top_I.branch[14].block[12].um_I.iw[6] ;
 wire \top_I.branch[14].block[12].um_I.iw[7] ;
 wire \top_I.branch[14].block[12].um_I.iw[8] ;
 wire \top_I.branch[14].block[12].um_I.iw[9] ;
 wire \top_I.branch[14].block[12].um_I.k_zero ;
 wire \top_I.branch[14].block[12].um_I.pg_vdd ;
 wire \top_I.branch[14].block[13].um_I.ana[0] ;
 wire \top_I.branch[14].block[13].um_I.ana[1] ;
 wire \top_I.branch[14].block[13].um_I.ana[2] ;
 wire \top_I.branch[14].block[13].um_I.ana[3] ;
 wire \top_I.branch[14].block[13].um_I.ana[4] ;
 wire \top_I.branch[14].block[13].um_I.ana[5] ;
 wire \top_I.branch[14].block[13].um_I.ana[6] ;
 wire \top_I.branch[14].block[13].um_I.ana[7] ;
 wire \top_I.branch[14].block[13].um_I.clk ;
 wire \top_I.branch[14].block[13].um_I.ena ;
 wire \top_I.branch[14].block[13].um_I.iw[10] ;
 wire \top_I.branch[14].block[13].um_I.iw[11] ;
 wire \top_I.branch[14].block[13].um_I.iw[12] ;
 wire \top_I.branch[14].block[13].um_I.iw[13] ;
 wire \top_I.branch[14].block[13].um_I.iw[14] ;
 wire \top_I.branch[14].block[13].um_I.iw[15] ;
 wire \top_I.branch[14].block[13].um_I.iw[16] ;
 wire \top_I.branch[14].block[13].um_I.iw[17] ;
 wire \top_I.branch[14].block[13].um_I.iw[1] ;
 wire \top_I.branch[14].block[13].um_I.iw[2] ;
 wire \top_I.branch[14].block[13].um_I.iw[3] ;
 wire \top_I.branch[14].block[13].um_I.iw[4] ;
 wire \top_I.branch[14].block[13].um_I.iw[5] ;
 wire \top_I.branch[14].block[13].um_I.iw[6] ;
 wire \top_I.branch[14].block[13].um_I.iw[7] ;
 wire \top_I.branch[14].block[13].um_I.iw[8] ;
 wire \top_I.branch[14].block[13].um_I.iw[9] ;
 wire \top_I.branch[14].block[13].um_I.k_zero ;
 wire \top_I.branch[14].block[13].um_I.pg_vdd ;
 wire \top_I.branch[14].block[14].um_I.ana[0] ;
 wire \top_I.branch[14].block[14].um_I.ana[1] ;
 wire \top_I.branch[14].block[14].um_I.ana[2] ;
 wire \top_I.branch[14].block[14].um_I.ana[3] ;
 wire \top_I.branch[14].block[14].um_I.ana[4] ;
 wire \top_I.branch[14].block[14].um_I.ana[5] ;
 wire \top_I.branch[14].block[14].um_I.ana[6] ;
 wire \top_I.branch[14].block[14].um_I.ana[7] ;
 wire \top_I.branch[14].block[14].um_I.clk ;
 wire \top_I.branch[14].block[14].um_I.ena ;
 wire \top_I.branch[14].block[14].um_I.iw[10] ;
 wire \top_I.branch[14].block[14].um_I.iw[11] ;
 wire \top_I.branch[14].block[14].um_I.iw[12] ;
 wire \top_I.branch[14].block[14].um_I.iw[13] ;
 wire \top_I.branch[14].block[14].um_I.iw[14] ;
 wire \top_I.branch[14].block[14].um_I.iw[15] ;
 wire \top_I.branch[14].block[14].um_I.iw[16] ;
 wire \top_I.branch[14].block[14].um_I.iw[17] ;
 wire \top_I.branch[14].block[14].um_I.iw[1] ;
 wire \top_I.branch[14].block[14].um_I.iw[2] ;
 wire \top_I.branch[14].block[14].um_I.iw[3] ;
 wire \top_I.branch[14].block[14].um_I.iw[4] ;
 wire \top_I.branch[14].block[14].um_I.iw[5] ;
 wire \top_I.branch[14].block[14].um_I.iw[6] ;
 wire \top_I.branch[14].block[14].um_I.iw[7] ;
 wire \top_I.branch[14].block[14].um_I.iw[8] ;
 wire \top_I.branch[14].block[14].um_I.iw[9] ;
 wire \top_I.branch[14].block[14].um_I.k_zero ;
 wire \top_I.branch[14].block[14].um_I.pg_vdd ;
 wire \top_I.branch[14].block[15].um_I.ana[0] ;
 wire \top_I.branch[14].block[15].um_I.ana[1] ;
 wire \top_I.branch[14].block[15].um_I.ana[2] ;
 wire \top_I.branch[14].block[15].um_I.ana[3] ;
 wire \top_I.branch[14].block[15].um_I.ana[4] ;
 wire \top_I.branch[14].block[15].um_I.ana[5] ;
 wire \top_I.branch[14].block[15].um_I.ana[6] ;
 wire \top_I.branch[14].block[15].um_I.ana[7] ;
 wire \top_I.branch[14].block[15].um_I.clk ;
 wire \top_I.branch[14].block[15].um_I.ena ;
 wire \top_I.branch[14].block[15].um_I.iw[10] ;
 wire \top_I.branch[14].block[15].um_I.iw[11] ;
 wire \top_I.branch[14].block[15].um_I.iw[12] ;
 wire \top_I.branch[14].block[15].um_I.iw[13] ;
 wire \top_I.branch[14].block[15].um_I.iw[14] ;
 wire \top_I.branch[14].block[15].um_I.iw[15] ;
 wire \top_I.branch[14].block[15].um_I.iw[16] ;
 wire \top_I.branch[14].block[15].um_I.iw[17] ;
 wire \top_I.branch[14].block[15].um_I.iw[1] ;
 wire \top_I.branch[14].block[15].um_I.iw[2] ;
 wire \top_I.branch[14].block[15].um_I.iw[3] ;
 wire \top_I.branch[14].block[15].um_I.iw[4] ;
 wire \top_I.branch[14].block[15].um_I.iw[5] ;
 wire \top_I.branch[14].block[15].um_I.iw[6] ;
 wire \top_I.branch[14].block[15].um_I.iw[7] ;
 wire \top_I.branch[14].block[15].um_I.iw[8] ;
 wire \top_I.branch[14].block[15].um_I.iw[9] ;
 wire \top_I.branch[14].block[15].um_I.k_zero ;
 wire \top_I.branch[14].block[15].um_I.pg_vdd ;
 wire \top_I.branch[14].block[1].um_I.ana[0] ;
 wire \top_I.branch[14].block[1].um_I.ana[1] ;
 wire \top_I.branch[14].block[1].um_I.ana[2] ;
 wire \top_I.branch[14].block[1].um_I.ana[3] ;
 wire \top_I.branch[14].block[1].um_I.ana[4] ;
 wire \top_I.branch[14].block[1].um_I.ana[5] ;
 wire \top_I.branch[14].block[1].um_I.ana[6] ;
 wire \top_I.branch[14].block[1].um_I.ana[7] ;
 wire \top_I.branch[14].block[1].um_I.clk ;
 wire \top_I.branch[14].block[1].um_I.ena ;
 wire \top_I.branch[14].block[1].um_I.iw[10] ;
 wire \top_I.branch[14].block[1].um_I.iw[11] ;
 wire \top_I.branch[14].block[1].um_I.iw[12] ;
 wire \top_I.branch[14].block[1].um_I.iw[13] ;
 wire \top_I.branch[14].block[1].um_I.iw[14] ;
 wire \top_I.branch[14].block[1].um_I.iw[15] ;
 wire \top_I.branch[14].block[1].um_I.iw[16] ;
 wire \top_I.branch[14].block[1].um_I.iw[17] ;
 wire \top_I.branch[14].block[1].um_I.iw[1] ;
 wire \top_I.branch[14].block[1].um_I.iw[2] ;
 wire \top_I.branch[14].block[1].um_I.iw[3] ;
 wire \top_I.branch[14].block[1].um_I.iw[4] ;
 wire \top_I.branch[14].block[1].um_I.iw[5] ;
 wire \top_I.branch[14].block[1].um_I.iw[6] ;
 wire \top_I.branch[14].block[1].um_I.iw[7] ;
 wire \top_I.branch[14].block[1].um_I.iw[8] ;
 wire \top_I.branch[14].block[1].um_I.iw[9] ;
 wire \top_I.branch[14].block[1].um_I.k_zero ;
 wire \top_I.branch[14].block[1].um_I.pg_vdd ;
 wire \top_I.branch[14].block[2].um_I.ana[0] ;
 wire \top_I.branch[14].block[2].um_I.ana[1] ;
 wire \top_I.branch[14].block[2].um_I.ana[2] ;
 wire \top_I.branch[14].block[2].um_I.ana[3] ;
 wire \top_I.branch[14].block[2].um_I.ana[4] ;
 wire \top_I.branch[14].block[2].um_I.ana[5] ;
 wire \top_I.branch[14].block[2].um_I.ana[6] ;
 wire \top_I.branch[14].block[2].um_I.ana[7] ;
 wire \top_I.branch[14].block[2].um_I.clk ;
 wire \top_I.branch[14].block[2].um_I.ena ;
 wire \top_I.branch[14].block[2].um_I.iw[10] ;
 wire \top_I.branch[14].block[2].um_I.iw[11] ;
 wire \top_I.branch[14].block[2].um_I.iw[12] ;
 wire \top_I.branch[14].block[2].um_I.iw[13] ;
 wire \top_I.branch[14].block[2].um_I.iw[14] ;
 wire \top_I.branch[14].block[2].um_I.iw[15] ;
 wire \top_I.branch[14].block[2].um_I.iw[16] ;
 wire \top_I.branch[14].block[2].um_I.iw[17] ;
 wire \top_I.branch[14].block[2].um_I.iw[1] ;
 wire \top_I.branch[14].block[2].um_I.iw[2] ;
 wire \top_I.branch[14].block[2].um_I.iw[3] ;
 wire \top_I.branch[14].block[2].um_I.iw[4] ;
 wire \top_I.branch[14].block[2].um_I.iw[5] ;
 wire \top_I.branch[14].block[2].um_I.iw[6] ;
 wire \top_I.branch[14].block[2].um_I.iw[7] ;
 wire \top_I.branch[14].block[2].um_I.iw[8] ;
 wire \top_I.branch[14].block[2].um_I.iw[9] ;
 wire \top_I.branch[14].block[2].um_I.k_zero ;
 wire \top_I.branch[14].block[2].um_I.pg_vdd ;
 wire \top_I.branch[14].block[3].um_I.ana[0] ;
 wire \top_I.branch[14].block[3].um_I.ana[1] ;
 wire \top_I.branch[14].block[3].um_I.ana[2] ;
 wire \top_I.branch[14].block[3].um_I.ana[3] ;
 wire \top_I.branch[14].block[3].um_I.ana[4] ;
 wire \top_I.branch[14].block[3].um_I.ana[5] ;
 wire \top_I.branch[14].block[3].um_I.ana[6] ;
 wire \top_I.branch[14].block[3].um_I.ana[7] ;
 wire \top_I.branch[14].block[3].um_I.clk ;
 wire \top_I.branch[14].block[3].um_I.ena ;
 wire \top_I.branch[14].block[3].um_I.iw[10] ;
 wire \top_I.branch[14].block[3].um_I.iw[11] ;
 wire \top_I.branch[14].block[3].um_I.iw[12] ;
 wire \top_I.branch[14].block[3].um_I.iw[13] ;
 wire \top_I.branch[14].block[3].um_I.iw[14] ;
 wire \top_I.branch[14].block[3].um_I.iw[15] ;
 wire \top_I.branch[14].block[3].um_I.iw[16] ;
 wire \top_I.branch[14].block[3].um_I.iw[17] ;
 wire \top_I.branch[14].block[3].um_I.iw[1] ;
 wire \top_I.branch[14].block[3].um_I.iw[2] ;
 wire \top_I.branch[14].block[3].um_I.iw[3] ;
 wire \top_I.branch[14].block[3].um_I.iw[4] ;
 wire \top_I.branch[14].block[3].um_I.iw[5] ;
 wire \top_I.branch[14].block[3].um_I.iw[6] ;
 wire \top_I.branch[14].block[3].um_I.iw[7] ;
 wire \top_I.branch[14].block[3].um_I.iw[8] ;
 wire \top_I.branch[14].block[3].um_I.iw[9] ;
 wire \top_I.branch[14].block[3].um_I.k_zero ;
 wire \top_I.branch[14].block[3].um_I.pg_vdd ;
 wire \top_I.branch[14].block[4].um_I.ana[0] ;
 wire \top_I.branch[14].block[4].um_I.ana[1] ;
 wire \top_I.branch[14].block[4].um_I.ana[2] ;
 wire \top_I.branch[14].block[4].um_I.ana[3] ;
 wire \top_I.branch[14].block[4].um_I.ana[4] ;
 wire \top_I.branch[14].block[4].um_I.ana[5] ;
 wire \top_I.branch[14].block[4].um_I.ana[6] ;
 wire \top_I.branch[14].block[4].um_I.ana[7] ;
 wire \top_I.branch[14].block[4].um_I.clk ;
 wire \top_I.branch[14].block[4].um_I.ena ;
 wire \top_I.branch[14].block[4].um_I.iw[10] ;
 wire \top_I.branch[14].block[4].um_I.iw[11] ;
 wire \top_I.branch[14].block[4].um_I.iw[12] ;
 wire \top_I.branch[14].block[4].um_I.iw[13] ;
 wire \top_I.branch[14].block[4].um_I.iw[14] ;
 wire \top_I.branch[14].block[4].um_I.iw[15] ;
 wire \top_I.branch[14].block[4].um_I.iw[16] ;
 wire \top_I.branch[14].block[4].um_I.iw[17] ;
 wire \top_I.branch[14].block[4].um_I.iw[1] ;
 wire \top_I.branch[14].block[4].um_I.iw[2] ;
 wire \top_I.branch[14].block[4].um_I.iw[3] ;
 wire \top_I.branch[14].block[4].um_I.iw[4] ;
 wire \top_I.branch[14].block[4].um_I.iw[5] ;
 wire \top_I.branch[14].block[4].um_I.iw[6] ;
 wire \top_I.branch[14].block[4].um_I.iw[7] ;
 wire \top_I.branch[14].block[4].um_I.iw[8] ;
 wire \top_I.branch[14].block[4].um_I.iw[9] ;
 wire \top_I.branch[14].block[4].um_I.k_zero ;
 wire \top_I.branch[14].block[4].um_I.pg_vdd ;
 wire \top_I.branch[14].block[5].um_I.ana[0] ;
 wire \top_I.branch[14].block[5].um_I.ana[1] ;
 wire \top_I.branch[14].block[5].um_I.ana[2] ;
 wire \top_I.branch[14].block[5].um_I.ana[3] ;
 wire \top_I.branch[14].block[5].um_I.ana[4] ;
 wire \top_I.branch[14].block[5].um_I.ana[5] ;
 wire \top_I.branch[14].block[5].um_I.ana[6] ;
 wire \top_I.branch[14].block[5].um_I.ana[7] ;
 wire \top_I.branch[14].block[5].um_I.clk ;
 wire \top_I.branch[14].block[5].um_I.ena ;
 wire \top_I.branch[14].block[5].um_I.iw[10] ;
 wire \top_I.branch[14].block[5].um_I.iw[11] ;
 wire \top_I.branch[14].block[5].um_I.iw[12] ;
 wire \top_I.branch[14].block[5].um_I.iw[13] ;
 wire \top_I.branch[14].block[5].um_I.iw[14] ;
 wire \top_I.branch[14].block[5].um_I.iw[15] ;
 wire \top_I.branch[14].block[5].um_I.iw[16] ;
 wire \top_I.branch[14].block[5].um_I.iw[17] ;
 wire \top_I.branch[14].block[5].um_I.iw[1] ;
 wire \top_I.branch[14].block[5].um_I.iw[2] ;
 wire \top_I.branch[14].block[5].um_I.iw[3] ;
 wire \top_I.branch[14].block[5].um_I.iw[4] ;
 wire \top_I.branch[14].block[5].um_I.iw[5] ;
 wire \top_I.branch[14].block[5].um_I.iw[6] ;
 wire \top_I.branch[14].block[5].um_I.iw[7] ;
 wire \top_I.branch[14].block[5].um_I.iw[8] ;
 wire \top_I.branch[14].block[5].um_I.iw[9] ;
 wire \top_I.branch[14].block[5].um_I.k_zero ;
 wire \top_I.branch[14].block[5].um_I.pg_vdd ;
 wire \top_I.branch[14].block[6].um_I.ana[0] ;
 wire \top_I.branch[14].block[6].um_I.ana[1] ;
 wire \top_I.branch[14].block[6].um_I.ana[2] ;
 wire \top_I.branch[14].block[6].um_I.ana[3] ;
 wire \top_I.branch[14].block[6].um_I.ana[4] ;
 wire \top_I.branch[14].block[6].um_I.ana[5] ;
 wire \top_I.branch[14].block[6].um_I.ana[6] ;
 wire \top_I.branch[14].block[6].um_I.ana[7] ;
 wire \top_I.branch[14].block[6].um_I.clk ;
 wire \top_I.branch[14].block[6].um_I.ena ;
 wire \top_I.branch[14].block[6].um_I.iw[10] ;
 wire \top_I.branch[14].block[6].um_I.iw[11] ;
 wire \top_I.branch[14].block[6].um_I.iw[12] ;
 wire \top_I.branch[14].block[6].um_I.iw[13] ;
 wire \top_I.branch[14].block[6].um_I.iw[14] ;
 wire \top_I.branch[14].block[6].um_I.iw[15] ;
 wire \top_I.branch[14].block[6].um_I.iw[16] ;
 wire \top_I.branch[14].block[6].um_I.iw[17] ;
 wire \top_I.branch[14].block[6].um_I.iw[1] ;
 wire \top_I.branch[14].block[6].um_I.iw[2] ;
 wire \top_I.branch[14].block[6].um_I.iw[3] ;
 wire \top_I.branch[14].block[6].um_I.iw[4] ;
 wire \top_I.branch[14].block[6].um_I.iw[5] ;
 wire \top_I.branch[14].block[6].um_I.iw[6] ;
 wire \top_I.branch[14].block[6].um_I.iw[7] ;
 wire \top_I.branch[14].block[6].um_I.iw[8] ;
 wire \top_I.branch[14].block[6].um_I.iw[9] ;
 wire \top_I.branch[14].block[6].um_I.k_zero ;
 wire \top_I.branch[14].block[6].um_I.pg_vdd ;
 wire \top_I.branch[14].block[7].um_I.ana[0] ;
 wire \top_I.branch[14].block[7].um_I.ana[1] ;
 wire \top_I.branch[14].block[7].um_I.ana[2] ;
 wire \top_I.branch[14].block[7].um_I.ana[3] ;
 wire \top_I.branch[14].block[7].um_I.ana[4] ;
 wire \top_I.branch[14].block[7].um_I.ana[5] ;
 wire \top_I.branch[14].block[7].um_I.ana[6] ;
 wire \top_I.branch[14].block[7].um_I.ana[7] ;
 wire \top_I.branch[14].block[7].um_I.clk ;
 wire \top_I.branch[14].block[7].um_I.ena ;
 wire \top_I.branch[14].block[7].um_I.iw[10] ;
 wire \top_I.branch[14].block[7].um_I.iw[11] ;
 wire \top_I.branch[14].block[7].um_I.iw[12] ;
 wire \top_I.branch[14].block[7].um_I.iw[13] ;
 wire \top_I.branch[14].block[7].um_I.iw[14] ;
 wire \top_I.branch[14].block[7].um_I.iw[15] ;
 wire \top_I.branch[14].block[7].um_I.iw[16] ;
 wire \top_I.branch[14].block[7].um_I.iw[17] ;
 wire \top_I.branch[14].block[7].um_I.iw[1] ;
 wire \top_I.branch[14].block[7].um_I.iw[2] ;
 wire \top_I.branch[14].block[7].um_I.iw[3] ;
 wire \top_I.branch[14].block[7].um_I.iw[4] ;
 wire \top_I.branch[14].block[7].um_I.iw[5] ;
 wire \top_I.branch[14].block[7].um_I.iw[6] ;
 wire \top_I.branch[14].block[7].um_I.iw[7] ;
 wire \top_I.branch[14].block[7].um_I.iw[8] ;
 wire \top_I.branch[14].block[7].um_I.iw[9] ;
 wire \top_I.branch[14].block[7].um_I.k_zero ;
 wire \top_I.branch[14].block[7].um_I.pg_vdd ;
 wire \top_I.branch[14].block[8].um_I.ana[0] ;
 wire \top_I.branch[14].block[8].um_I.ana[1] ;
 wire \top_I.branch[14].block[8].um_I.ana[2] ;
 wire \top_I.branch[14].block[8].um_I.ana[3] ;
 wire \top_I.branch[14].block[8].um_I.ana[4] ;
 wire \top_I.branch[14].block[8].um_I.ana[5] ;
 wire \top_I.branch[14].block[8].um_I.ana[6] ;
 wire \top_I.branch[14].block[8].um_I.ana[7] ;
 wire \top_I.branch[14].block[8].um_I.clk ;
 wire \top_I.branch[14].block[8].um_I.ena ;
 wire \top_I.branch[14].block[8].um_I.iw[10] ;
 wire \top_I.branch[14].block[8].um_I.iw[11] ;
 wire \top_I.branch[14].block[8].um_I.iw[12] ;
 wire \top_I.branch[14].block[8].um_I.iw[13] ;
 wire \top_I.branch[14].block[8].um_I.iw[14] ;
 wire \top_I.branch[14].block[8].um_I.iw[15] ;
 wire \top_I.branch[14].block[8].um_I.iw[16] ;
 wire \top_I.branch[14].block[8].um_I.iw[17] ;
 wire \top_I.branch[14].block[8].um_I.iw[1] ;
 wire \top_I.branch[14].block[8].um_I.iw[2] ;
 wire \top_I.branch[14].block[8].um_I.iw[3] ;
 wire \top_I.branch[14].block[8].um_I.iw[4] ;
 wire \top_I.branch[14].block[8].um_I.iw[5] ;
 wire \top_I.branch[14].block[8].um_I.iw[6] ;
 wire \top_I.branch[14].block[8].um_I.iw[7] ;
 wire \top_I.branch[14].block[8].um_I.iw[8] ;
 wire \top_I.branch[14].block[8].um_I.iw[9] ;
 wire \top_I.branch[14].block[8].um_I.k_zero ;
 wire \top_I.branch[14].block[8].um_I.pg_vdd ;
 wire \top_I.branch[14].block[9].um_I.ana[0] ;
 wire \top_I.branch[14].block[9].um_I.ana[1] ;
 wire \top_I.branch[14].block[9].um_I.ana[2] ;
 wire \top_I.branch[14].block[9].um_I.ana[3] ;
 wire \top_I.branch[14].block[9].um_I.ana[4] ;
 wire \top_I.branch[14].block[9].um_I.ana[5] ;
 wire \top_I.branch[14].block[9].um_I.ana[6] ;
 wire \top_I.branch[14].block[9].um_I.ana[7] ;
 wire \top_I.branch[14].block[9].um_I.clk ;
 wire \top_I.branch[14].block[9].um_I.ena ;
 wire \top_I.branch[14].block[9].um_I.iw[10] ;
 wire \top_I.branch[14].block[9].um_I.iw[11] ;
 wire \top_I.branch[14].block[9].um_I.iw[12] ;
 wire \top_I.branch[14].block[9].um_I.iw[13] ;
 wire \top_I.branch[14].block[9].um_I.iw[14] ;
 wire \top_I.branch[14].block[9].um_I.iw[15] ;
 wire \top_I.branch[14].block[9].um_I.iw[16] ;
 wire \top_I.branch[14].block[9].um_I.iw[17] ;
 wire \top_I.branch[14].block[9].um_I.iw[1] ;
 wire \top_I.branch[14].block[9].um_I.iw[2] ;
 wire \top_I.branch[14].block[9].um_I.iw[3] ;
 wire \top_I.branch[14].block[9].um_I.iw[4] ;
 wire \top_I.branch[14].block[9].um_I.iw[5] ;
 wire \top_I.branch[14].block[9].um_I.iw[6] ;
 wire \top_I.branch[14].block[9].um_I.iw[7] ;
 wire \top_I.branch[14].block[9].um_I.iw[8] ;
 wire \top_I.branch[14].block[9].um_I.iw[9] ;
 wire \top_I.branch[14].block[9].um_I.k_zero ;
 wire \top_I.branch[14].block[9].um_I.pg_vdd ;
 wire \top_I.branch[14].l_addr[0] ;
 wire \top_I.branch[14].l_addr[3] ;
 wire \top_I.branch[15].block[0].um_I.ana[0] ;
 wire \top_I.branch[15].block[0].um_I.ana[1] ;
 wire \top_I.branch[15].block[0].um_I.ana[2] ;
 wire \top_I.branch[15].block[0].um_I.ana[3] ;
 wire \top_I.branch[15].block[0].um_I.ana[4] ;
 wire \top_I.branch[15].block[0].um_I.ana[5] ;
 wire \top_I.branch[15].block[0].um_I.ana[6] ;
 wire \top_I.branch[15].block[0].um_I.ana[7] ;
 wire \top_I.branch[15].block[0].um_I.clk ;
 wire \top_I.branch[15].block[0].um_I.ena ;
 wire \top_I.branch[15].block[0].um_I.iw[10] ;
 wire \top_I.branch[15].block[0].um_I.iw[11] ;
 wire \top_I.branch[15].block[0].um_I.iw[12] ;
 wire \top_I.branch[15].block[0].um_I.iw[13] ;
 wire \top_I.branch[15].block[0].um_I.iw[14] ;
 wire \top_I.branch[15].block[0].um_I.iw[15] ;
 wire \top_I.branch[15].block[0].um_I.iw[16] ;
 wire \top_I.branch[15].block[0].um_I.iw[17] ;
 wire \top_I.branch[15].block[0].um_I.iw[1] ;
 wire \top_I.branch[15].block[0].um_I.iw[2] ;
 wire \top_I.branch[15].block[0].um_I.iw[3] ;
 wire \top_I.branch[15].block[0].um_I.iw[4] ;
 wire \top_I.branch[15].block[0].um_I.iw[5] ;
 wire \top_I.branch[15].block[0].um_I.iw[6] ;
 wire \top_I.branch[15].block[0].um_I.iw[7] ;
 wire \top_I.branch[15].block[0].um_I.iw[8] ;
 wire \top_I.branch[15].block[0].um_I.iw[9] ;
 wire \top_I.branch[15].block[0].um_I.k_zero ;
 wire \top_I.branch[15].block[0].um_I.pg_vdd ;
 wire \top_I.branch[15].block[10].um_I.ana[0] ;
 wire \top_I.branch[15].block[10].um_I.ana[1] ;
 wire \top_I.branch[15].block[10].um_I.ana[2] ;
 wire \top_I.branch[15].block[10].um_I.ana[3] ;
 wire \top_I.branch[15].block[10].um_I.ana[4] ;
 wire \top_I.branch[15].block[10].um_I.ana[5] ;
 wire \top_I.branch[15].block[10].um_I.ana[6] ;
 wire \top_I.branch[15].block[10].um_I.ana[7] ;
 wire \top_I.branch[15].block[10].um_I.clk ;
 wire \top_I.branch[15].block[10].um_I.ena ;
 wire \top_I.branch[15].block[10].um_I.iw[10] ;
 wire \top_I.branch[15].block[10].um_I.iw[11] ;
 wire \top_I.branch[15].block[10].um_I.iw[12] ;
 wire \top_I.branch[15].block[10].um_I.iw[13] ;
 wire \top_I.branch[15].block[10].um_I.iw[14] ;
 wire \top_I.branch[15].block[10].um_I.iw[15] ;
 wire \top_I.branch[15].block[10].um_I.iw[16] ;
 wire \top_I.branch[15].block[10].um_I.iw[17] ;
 wire \top_I.branch[15].block[10].um_I.iw[1] ;
 wire \top_I.branch[15].block[10].um_I.iw[2] ;
 wire \top_I.branch[15].block[10].um_I.iw[3] ;
 wire \top_I.branch[15].block[10].um_I.iw[4] ;
 wire \top_I.branch[15].block[10].um_I.iw[5] ;
 wire \top_I.branch[15].block[10].um_I.iw[6] ;
 wire \top_I.branch[15].block[10].um_I.iw[7] ;
 wire \top_I.branch[15].block[10].um_I.iw[8] ;
 wire \top_I.branch[15].block[10].um_I.iw[9] ;
 wire \top_I.branch[15].block[10].um_I.k_zero ;
 wire \top_I.branch[15].block[10].um_I.pg_vdd ;
 wire \top_I.branch[15].block[11].um_I.ana[0] ;
 wire \top_I.branch[15].block[11].um_I.ana[1] ;
 wire \top_I.branch[15].block[11].um_I.ana[2] ;
 wire \top_I.branch[15].block[11].um_I.ana[3] ;
 wire \top_I.branch[15].block[11].um_I.ana[4] ;
 wire \top_I.branch[15].block[11].um_I.ana[5] ;
 wire \top_I.branch[15].block[11].um_I.ana[6] ;
 wire \top_I.branch[15].block[11].um_I.ana[7] ;
 wire \top_I.branch[15].block[11].um_I.clk ;
 wire \top_I.branch[15].block[11].um_I.ena ;
 wire \top_I.branch[15].block[11].um_I.iw[10] ;
 wire \top_I.branch[15].block[11].um_I.iw[11] ;
 wire \top_I.branch[15].block[11].um_I.iw[12] ;
 wire \top_I.branch[15].block[11].um_I.iw[13] ;
 wire \top_I.branch[15].block[11].um_I.iw[14] ;
 wire \top_I.branch[15].block[11].um_I.iw[15] ;
 wire \top_I.branch[15].block[11].um_I.iw[16] ;
 wire \top_I.branch[15].block[11].um_I.iw[17] ;
 wire \top_I.branch[15].block[11].um_I.iw[1] ;
 wire \top_I.branch[15].block[11].um_I.iw[2] ;
 wire \top_I.branch[15].block[11].um_I.iw[3] ;
 wire \top_I.branch[15].block[11].um_I.iw[4] ;
 wire \top_I.branch[15].block[11].um_I.iw[5] ;
 wire \top_I.branch[15].block[11].um_I.iw[6] ;
 wire \top_I.branch[15].block[11].um_I.iw[7] ;
 wire \top_I.branch[15].block[11].um_I.iw[8] ;
 wire \top_I.branch[15].block[11].um_I.iw[9] ;
 wire \top_I.branch[15].block[11].um_I.k_zero ;
 wire \top_I.branch[15].block[11].um_I.pg_vdd ;
 wire \top_I.branch[15].block[12].um_I.ana[0] ;
 wire \top_I.branch[15].block[12].um_I.ana[1] ;
 wire \top_I.branch[15].block[12].um_I.ana[2] ;
 wire \top_I.branch[15].block[12].um_I.ana[3] ;
 wire \top_I.branch[15].block[12].um_I.ana[4] ;
 wire \top_I.branch[15].block[12].um_I.ana[5] ;
 wire \top_I.branch[15].block[12].um_I.ana[6] ;
 wire \top_I.branch[15].block[12].um_I.ana[7] ;
 wire \top_I.branch[15].block[12].um_I.clk ;
 wire \top_I.branch[15].block[12].um_I.ena ;
 wire \top_I.branch[15].block[12].um_I.iw[10] ;
 wire \top_I.branch[15].block[12].um_I.iw[11] ;
 wire \top_I.branch[15].block[12].um_I.iw[12] ;
 wire \top_I.branch[15].block[12].um_I.iw[13] ;
 wire \top_I.branch[15].block[12].um_I.iw[14] ;
 wire \top_I.branch[15].block[12].um_I.iw[15] ;
 wire \top_I.branch[15].block[12].um_I.iw[16] ;
 wire \top_I.branch[15].block[12].um_I.iw[17] ;
 wire \top_I.branch[15].block[12].um_I.iw[1] ;
 wire \top_I.branch[15].block[12].um_I.iw[2] ;
 wire \top_I.branch[15].block[12].um_I.iw[3] ;
 wire \top_I.branch[15].block[12].um_I.iw[4] ;
 wire \top_I.branch[15].block[12].um_I.iw[5] ;
 wire \top_I.branch[15].block[12].um_I.iw[6] ;
 wire \top_I.branch[15].block[12].um_I.iw[7] ;
 wire \top_I.branch[15].block[12].um_I.iw[8] ;
 wire \top_I.branch[15].block[12].um_I.iw[9] ;
 wire \top_I.branch[15].block[12].um_I.k_zero ;
 wire \top_I.branch[15].block[12].um_I.pg_vdd ;
 wire \top_I.branch[15].block[13].um_I.ana[0] ;
 wire \top_I.branch[15].block[13].um_I.ana[1] ;
 wire \top_I.branch[15].block[13].um_I.ana[2] ;
 wire \top_I.branch[15].block[13].um_I.ana[3] ;
 wire \top_I.branch[15].block[13].um_I.ana[4] ;
 wire \top_I.branch[15].block[13].um_I.ana[5] ;
 wire \top_I.branch[15].block[13].um_I.ana[6] ;
 wire \top_I.branch[15].block[13].um_I.ana[7] ;
 wire \top_I.branch[15].block[13].um_I.clk ;
 wire \top_I.branch[15].block[13].um_I.ena ;
 wire \top_I.branch[15].block[13].um_I.iw[10] ;
 wire \top_I.branch[15].block[13].um_I.iw[11] ;
 wire \top_I.branch[15].block[13].um_I.iw[12] ;
 wire \top_I.branch[15].block[13].um_I.iw[13] ;
 wire \top_I.branch[15].block[13].um_I.iw[14] ;
 wire \top_I.branch[15].block[13].um_I.iw[15] ;
 wire \top_I.branch[15].block[13].um_I.iw[16] ;
 wire \top_I.branch[15].block[13].um_I.iw[17] ;
 wire \top_I.branch[15].block[13].um_I.iw[1] ;
 wire \top_I.branch[15].block[13].um_I.iw[2] ;
 wire \top_I.branch[15].block[13].um_I.iw[3] ;
 wire \top_I.branch[15].block[13].um_I.iw[4] ;
 wire \top_I.branch[15].block[13].um_I.iw[5] ;
 wire \top_I.branch[15].block[13].um_I.iw[6] ;
 wire \top_I.branch[15].block[13].um_I.iw[7] ;
 wire \top_I.branch[15].block[13].um_I.iw[8] ;
 wire \top_I.branch[15].block[13].um_I.iw[9] ;
 wire \top_I.branch[15].block[13].um_I.k_zero ;
 wire \top_I.branch[15].block[13].um_I.pg_vdd ;
 wire \top_I.branch[15].block[14].um_I.ana[0] ;
 wire \top_I.branch[15].block[14].um_I.ana[1] ;
 wire \top_I.branch[15].block[14].um_I.ana[2] ;
 wire \top_I.branch[15].block[14].um_I.ana[3] ;
 wire \top_I.branch[15].block[14].um_I.ana[4] ;
 wire \top_I.branch[15].block[14].um_I.ana[5] ;
 wire \top_I.branch[15].block[14].um_I.ana[6] ;
 wire \top_I.branch[15].block[14].um_I.ana[7] ;
 wire \top_I.branch[15].block[14].um_I.clk ;
 wire \top_I.branch[15].block[14].um_I.ena ;
 wire \top_I.branch[15].block[14].um_I.iw[10] ;
 wire \top_I.branch[15].block[14].um_I.iw[11] ;
 wire \top_I.branch[15].block[14].um_I.iw[12] ;
 wire \top_I.branch[15].block[14].um_I.iw[13] ;
 wire \top_I.branch[15].block[14].um_I.iw[14] ;
 wire \top_I.branch[15].block[14].um_I.iw[15] ;
 wire \top_I.branch[15].block[14].um_I.iw[16] ;
 wire \top_I.branch[15].block[14].um_I.iw[17] ;
 wire \top_I.branch[15].block[14].um_I.iw[1] ;
 wire \top_I.branch[15].block[14].um_I.iw[2] ;
 wire \top_I.branch[15].block[14].um_I.iw[3] ;
 wire \top_I.branch[15].block[14].um_I.iw[4] ;
 wire \top_I.branch[15].block[14].um_I.iw[5] ;
 wire \top_I.branch[15].block[14].um_I.iw[6] ;
 wire \top_I.branch[15].block[14].um_I.iw[7] ;
 wire \top_I.branch[15].block[14].um_I.iw[8] ;
 wire \top_I.branch[15].block[14].um_I.iw[9] ;
 wire \top_I.branch[15].block[14].um_I.k_zero ;
 wire \top_I.branch[15].block[14].um_I.pg_vdd ;
 wire \top_I.branch[15].block[15].um_I.ana[0] ;
 wire \top_I.branch[15].block[15].um_I.ana[1] ;
 wire \top_I.branch[15].block[15].um_I.ana[2] ;
 wire \top_I.branch[15].block[15].um_I.ana[3] ;
 wire \top_I.branch[15].block[15].um_I.ana[4] ;
 wire \top_I.branch[15].block[15].um_I.ana[5] ;
 wire \top_I.branch[15].block[15].um_I.ana[6] ;
 wire \top_I.branch[15].block[15].um_I.ana[7] ;
 wire \top_I.branch[15].block[15].um_I.clk ;
 wire \top_I.branch[15].block[15].um_I.ena ;
 wire \top_I.branch[15].block[15].um_I.iw[10] ;
 wire \top_I.branch[15].block[15].um_I.iw[11] ;
 wire \top_I.branch[15].block[15].um_I.iw[12] ;
 wire \top_I.branch[15].block[15].um_I.iw[13] ;
 wire \top_I.branch[15].block[15].um_I.iw[14] ;
 wire \top_I.branch[15].block[15].um_I.iw[15] ;
 wire \top_I.branch[15].block[15].um_I.iw[16] ;
 wire \top_I.branch[15].block[15].um_I.iw[17] ;
 wire \top_I.branch[15].block[15].um_I.iw[1] ;
 wire \top_I.branch[15].block[15].um_I.iw[2] ;
 wire \top_I.branch[15].block[15].um_I.iw[3] ;
 wire \top_I.branch[15].block[15].um_I.iw[4] ;
 wire \top_I.branch[15].block[15].um_I.iw[5] ;
 wire \top_I.branch[15].block[15].um_I.iw[6] ;
 wire \top_I.branch[15].block[15].um_I.iw[7] ;
 wire \top_I.branch[15].block[15].um_I.iw[8] ;
 wire \top_I.branch[15].block[15].um_I.iw[9] ;
 wire \top_I.branch[15].block[15].um_I.k_zero ;
 wire \top_I.branch[15].block[15].um_I.pg_vdd ;
 wire \top_I.branch[15].block[1].um_I.ana[0] ;
 wire \top_I.branch[15].block[1].um_I.ana[1] ;
 wire \top_I.branch[15].block[1].um_I.ana[2] ;
 wire \top_I.branch[15].block[1].um_I.ana[3] ;
 wire \top_I.branch[15].block[1].um_I.ana[4] ;
 wire \top_I.branch[15].block[1].um_I.ana[5] ;
 wire \top_I.branch[15].block[1].um_I.ana[6] ;
 wire \top_I.branch[15].block[1].um_I.ana[7] ;
 wire \top_I.branch[15].block[1].um_I.clk ;
 wire \top_I.branch[15].block[1].um_I.ena ;
 wire \top_I.branch[15].block[1].um_I.iw[10] ;
 wire \top_I.branch[15].block[1].um_I.iw[11] ;
 wire \top_I.branch[15].block[1].um_I.iw[12] ;
 wire \top_I.branch[15].block[1].um_I.iw[13] ;
 wire \top_I.branch[15].block[1].um_I.iw[14] ;
 wire \top_I.branch[15].block[1].um_I.iw[15] ;
 wire \top_I.branch[15].block[1].um_I.iw[16] ;
 wire \top_I.branch[15].block[1].um_I.iw[17] ;
 wire \top_I.branch[15].block[1].um_I.iw[1] ;
 wire \top_I.branch[15].block[1].um_I.iw[2] ;
 wire \top_I.branch[15].block[1].um_I.iw[3] ;
 wire \top_I.branch[15].block[1].um_I.iw[4] ;
 wire \top_I.branch[15].block[1].um_I.iw[5] ;
 wire \top_I.branch[15].block[1].um_I.iw[6] ;
 wire \top_I.branch[15].block[1].um_I.iw[7] ;
 wire \top_I.branch[15].block[1].um_I.iw[8] ;
 wire \top_I.branch[15].block[1].um_I.iw[9] ;
 wire \top_I.branch[15].block[1].um_I.k_zero ;
 wire \top_I.branch[15].block[1].um_I.pg_vdd ;
 wire \top_I.branch[15].block[2].um_I.ana[0] ;
 wire \top_I.branch[15].block[2].um_I.ana[1] ;
 wire \top_I.branch[15].block[2].um_I.ana[2] ;
 wire \top_I.branch[15].block[2].um_I.ana[3] ;
 wire \top_I.branch[15].block[2].um_I.ana[4] ;
 wire \top_I.branch[15].block[2].um_I.ana[5] ;
 wire \top_I.branch[15].block[2].um_I.ana[6] ;
 wire \top_I.branch[15].block[2].um_I.ana[7] ;
 wire \top_I.branch[15].block[2].um_I.clk ;
 wire \top_I.branch[15].block[2].um_I.ena ;
 wire \top_I.branch[15].block[2].um_I.iw[10] ;
 wire \top_I.branch[15].block[2].um_I.iw[11] ;
 wire \top_I.branch[15].block[2].um_I.iw[12] ;
 wire \top_I.branch[15].block[2].um_I.iw[13] ;
 wire \top_I.branch[15].block[2].um_I.iw[14] ;
 wire \top_I.branch[15].block[2].um_I.iw[15] ;
 wire \top_I.branch[15].block[2].um_I.iw[16] ;
 wire \top_I.branch[15].block[2].um_I.iw[17] ;
 wire \top_I.branch[15].block[2].um_I.iw[1] ;
 wire \top_I.branch[15].block[2].um_I.iw[2] ;
 wire \top_I.branch[15].block[2].um_I.iw[3] ;
 wire \top_I.branch[15].block[2].um_I.iw[4] ;
 wire \top_I.branch[15].block[2].um_I.iw[5] ;
 wire \top_I.branch[15].block[2].um_I.iw[6] ;
 wire \top_I.branch[15].block[2].um_I.iw[7] ;
 wire \top_I.branch[15].block[2].um_I.iw[8] ;
 wire \top_I.branch[15].block[2].um_I.iw[9] ;
 wire \top_I.branch[15].block[2].um_I.k_zero ;
 wire \top_I.branch[15].block[2].um_I.pg_vdd ;
 wire \top_I.branch[15].block[3].um_I.ana[0] ;
 wire \top_I.branch[15].block[3].um_I.ana[1] ;
 wire \top_I.branch[15].block[3].um_I.ana[2] ;
 wire \top_I.branch[15].block[3].um_I.ana[3] ;
 wire \top_I.branch[15].block[3].um_I.ana[4] ;
 wire \top_I.branch[15].block[3].um_I.ana[5] ;
 wire \top_I.branch[15].block[3].um_I.ana[6] ;
 wire \top_I.branch[15].block[3].um_I.ana[7] ;
 wire \top_I.branch[15].block[3].um_I.clk ;
 wire \top_I.branch[15].block[3].um_I.ena ;
 wire \top_I.branch[15].block[3].um_I.iw[10] ;
 wire \top_I.branch[15].block[3].um_I.iw[11] ;
 wire \top_I.branch[15].block[3].um_I.iw[12] ;
 wire \top_I.branch[15].block[3].um_I.iw[13] ;
 wire \top_I.branch[15].block[3].um_I.iw[14] ;
 wire \top_I.branch[15].block[3].um_I.iw[15] ;
 wire \top_I.branch[15].block[3].um_I.iw[16] ;
 wire \top_I.branch[15].block[3].um_I.iw[17] ;
 wire \top_I.branch[15].block[3].um_I.iw[1] ;
 wire \top_I.branch[15].block[3].um_I.iw[2] ;
 wire \top_I.branch[15].block[3].um_I.iw[3] ;
 wire \top_I.branch[15].block[3].um_I.iw[4] ;
 wire \top_I.branch[15].block[3].um_I.iw[5] ;
 wire \top_I.branch[15].block[3].um_I.iw[6] ;
 wire \top_I.branch[15].block[3].um_I.iw[7] ;
 wire \top_I.branch[15].block[3].um_I.iw[8] ;
 wire \top_I.branch[15].block[3].um_I.iw[9] ;
 wire \top_I.branch[15].block[3].um_I.k_zero ;
 wire \top_I.branch[15].block[3].um_I.pg_vdd ;
 wire \top_I.branch[15].block[4].um_I.ana[0] ;
 wire \top_I.branch[15].block[4].um_I.ana[1] ;
 wire \top_I.branch[15].block[4].um_I.ana[2] ;
 wire \top_I.branch[15].block[4].um_I.ana[3] ;
 wire \top_I.branch[15].block[4].um_I.ana[4] ;
 wire \top_I.branch[15].block[4].um_I.ana[5] ;
 wire \top_I.branch[15].block[4].um_I.ana[6] ;
 wire \top_I.branch[15].block[4].um_I.ana[7] ;
 wire \top_I.branch[15].block[4].um_I.clk ;
 wire \top_I.branch[15].block[4].um_I.ena ;
 wire \top_I.branch[15].block[4].um_I.iw[10] ;
 wire \top_I.branch[15].block[4].um_I.iw[11] ;
 wire \top_I.branch[15].block[4].um_I.iw[12] ;
 wire \top_I.branch[15].block[4].um_I.iw[13] ;
 wire \top_I.branch[15].block[4].um_I.iw[14] ;
 wire \top_I.branch[15].block[4].um_I.iw[15] ;
 wire \top_I.branch[15].block[4].um_I.iw[16] ;
 wire \top_I.branch[15].block[4].um_I.iw[17] ;
 wire \top_I.branch[15].block[4].um_I.iw[1] ;
 wire \top_I.branch[15].block[4].um_I.iw[2] ;
 wire \top_I.branch[15].block[4].um_I.iw[3] ;
 wire \top_I.branch[15].block[4].um_I.iw[4] ;
 wire \top_I.branch[15].block[4].um_I.iw[5] ;
 wire \top_I.branch[15].block[4].um_I.iw[6] ;
 wire \top_I.branch[15].block[4].um_I.iw[7] ;
 wire \top_I.branch[15].block[4].um_I.iw[8] ;
 wire \top_I.branch[15].block[4].um_I.iw[9] ;
 wire \top_I.branch[15].block[4].um_I.k_zero ;
 wire \top_I.branch[15].block[4].um_I.pg_vdd ;
 wire \top_I.branch[15].block[5].um_I.ana[0] ;
 wire \top_I.branch[15].block[5].um_I.ana[1] ;
 wire \top_I.branch[15].block[5].um_I.ana[2] ;
 wire \top_I.branch[15].block[5].um_I.ana[3] ;
 wire \top_I.branch[15].block[5].um_I.ana[4] ;
 wire \top_I.branch[15].block[5].um_I.ana[5] ;
 wire \top_I.branch[15].block[5].um_I.ana[6] ;
 wire \top_I.branch[15].block[5].um_I.ana[7] ;
 wire \top_I.branch[15].block[5].um_I.clk ;
 wire \top_I.branch[15].block[5].um_I.ena ;
 wire \top_I.branch[15].block[5].um_I.iw[10] ;
 wire \top_I.branch[15].block[5].um_I.iw[11] ;
 wire \top_I.branch[15].block[5].um_I.iw[12] ;
 wire \top_I.branch[15].block[5].um_I.iw[13] ;
 wire \top_I.branch[15].block[5].um_I.iw[14] ;
 wire \top_I.branch[15].block[5].um_I.iw[15] ;
 wire \top_I.branch[15].block[5].um_I.iw[16] ;
 wire \top_I.branch[15].block[5].um_I.iw[17] ;
 wire \top_I.branch[15].block[5].um_I.iw[1] ;
 wire \top_I.branch[15].block[5].um_I.iw[2] ;
 wire \top_I.branch[15].block[5].um_I.iw[3] ;
 wire \top_I.branch[15].block[5].um_I.iw[4] ;
 wire \top_I.branch[15].block[5].um_I.iw[5] ;
 wire \top_I.branch[15].block[5].um_I.iw[6] ;
 wire \top_I.branch[15].block[5].um_I.iw[7] ;
 wire \top_I.branch[15].block[5].um_I.iw[8] ;
 wire \top_I.branch[15].block[5].um_I.iw[9] ;
 wire \top_I.branch[15].block[5].um_I.k_zero ;
 wire \top_I.branch[15].block[5].um_I.pg_vdd ;
 wire \top_I.branch[15].block[6].um_I.ana[0] ;
 wire \top_I.branch[15].block[6].um_I.ana[1] ;
 wire \top_I.branch[15].block[6].um_I.ana[2] ;
 wire \top_I.branch[15].block[6].um_I.ana[3] ;
 wire \top_I.branch[15].block[6].um_I.ana[4] ;
 wire \top_I.branch[15].block[6].um_I.ana[5] ;
 wire \top_I.branch[15].block[6].um_I.ana[6] ;
 wire \top_I.branch[15].block[6].um_I.ana[7] ;
 wire \top_I.branch[15].block[6].um_I.clk ;
 wire \top_I.branch[15].block[6].um_I.ena ;
 wire \top_I.branch[15].block[6].um_I.iw[10] ;
 wire \top_I.branch[15].block[6].um_I.iw[11] ;
 wire \top_I.branch[15].block[6].um_I.iw[12] ;
 wire \top_I.branch[15].block[6].um_I.iw[13] ;
 wire \top_I.branch[15].block[6].um_I.iw[14] ;
 wire \top_I.branch[15].block[6].um_I.iw[15] ;
 wire \top_I.branch[15].block[6].um_I.iw[16] ;
 wire \top_I.branch[15].block[6].um_I.iw[17] ;
 wire \top_I.branch[15].block[6].um_I.iw[1] ;
 wire \top_I.branch[15].block[6].um_I.iw[2] ;
 wire \top_I.branch[15].block[6].um_I.iw[3] ;
 wire \top_I.branch[15].block[6].um_I.iw[4] ;
 wire \top_I.branch[15].block[6].um_I.iw[5] ;
 wire \top_I.branch[15].block[6].um_I.iw[6] ;
 wire \top_I.branch[15].block[6].um_I.iw[7] ;
 wire \top_I.branch[15].block[6].um_I.iw[8] ;
 wire \top_I.branch[15].block[6].um_I.iw[9] ;
 wire \top_I.branch[15].block[6].um_I.k_zero ;
 wire \top_I.branch[15].block[6].um_I.pg_vdd ;
 wire \top_I.branch[15].block[7].um_I.ana[0] ;
 wire \top_I.branch[15].block[7].um_I.ana[1] ;
 wire \top_I.branch[15].block[7].um_I.ana[2] ;
 wire \top_I.branch[15].block[7].um_I.ana[3] ;
 wire \top_I.branch[15].block[7].um_I.ana[4] ;
 wire \top_I.branch[15].block[7].um_I.ana[5] ;
 wire \top_I.branch[15].block[7].um_I.ana[6] ;
 wire \top_I.branch[15].block[7].um_I.ana[7] ;
 wire \top_I.branch[15].block[7].um_I.clk ;
 wire \top_I.branch[15].block[7].um_I.ena ;
 wire \top_I.branch[15].block[7].um_I.iw[10] ;
 wire \top_I.branch[15].block[7].um_I.iw[11] ;
 wire \top_I.branch[15].block[7].um_I.iw[12] ;
 wire \top_I.branch[15].block[7].um_I.iw[13] ;
 wire \top_I.branch[15].block[7].um_I.iw[14] ;
 wire \top_I.branch[15].block[7].um_I.iw[15] ;
 wire \top_I.branch[15].block[7].um_I.iw[16] ;
 wire \top_I.branch[15].block[7].um_I.iw[17] ;
 wire \top_I.branch[15].block[7].um_I.iw[1] ;
 wire \top_I.branch[15].block[7].um_I.iw[2] ;
 wire \top_I.branch[15].block[7].um_I.iw[3] ;
 wire \top_I.branch[15].block[7].um_I.iw[4] ;
 wire \top_I.branch[15].block[7].um_I.iw[5] ;
 wire \top_I.branch[15].block[7].um_I.iw[6] ;
 wire \top_I.branch[15].block[7].um_I.iw[7] ;
 wire \top_I.branch[15].block[7].um_I.iw[8] ;
 wire \top_I.branch[15].block[7].um_I.iw[9] ;
 wire \top_I.branch[15].block[7].um_I.k_zero ;
 wire \top_I.branch[15].block[7].um_I.pg_vdd ;
 wire \top_I.branch[15].block[8].um_I.ana[0] ;
 wire \top_I.branch[15].block[8].um_I.ana[1] ;
 wire \top_I.branch[15].block[8].um_I.ana[2] ;
 wire \top_I.branch[15].block[8].um_I.ana[3] ;
 wire \top_I.branch[15].block[8].um_I.ana[4] ;
 wire \top_I.branch[15].block[8].um_I.ana[5] ;
 wire \top_I.branch[15].block[8].um_I.ana[6] ;
 wire \top_I.branch[15].block[8].um_I.ana[7] ;
 wire \top_I.branch[15].block[8].um_I.clk ;
 wire \top_I.branch[15].block[8].um_I.ena ;
 wire \top_I.branch[15].block[8].um_I.iw[10] ;
 wire \top_I.branch[15].block[8].um_I.iw[11] ;
 wire \top_I.branch[15].block[8].um_I.iw[12] ;
 wire \top_I.branch[15].block[8].um_I.iw[13] ;
 wire \top_I.branch[15].block[8].um_I.iw[14] ;
 wire \top_I.branch[15].block[8].um_I.iw[15] ;
 wire \top_I.branch[15].block[8].um_I.iw[16] ;
 wire \top_I.branch[15].block[8].um_I.iw[17] ;
 wire \top_I.branch[15].block[8].um_I.iw[1] ;
 wire \top_I.branch[15].block[8].um_I.iw[2] ;
 wire \top_I.branch[15].block[8].um_I.iw[3] ;
 wire \top_I.branch[15].block[8].um_I.iw[4] ;
 wire \top_I.branch[15].block[8].um_I.iw[5] ;
 wire \top_I.branch[15].block[8].um_I.iw[6] ;
 wire \top_I.branch[15].block[8].um_I.iw[7] ;
 wire \top_I.branch[15].block[8].um_I.iw[8] ;
 wire \top_I.branch[15].block[8].um_I.iw[9] ;
 wire \top_I.branch[15].block[8].um_I.k_zero ;
 wire \top_I.branch[15].block[8].um_I.pg_vdd ;
 wire \top_I.branch[15].block[9].um_I.ana[0] ;
 wire \top_I.branch[15].block[9].um_I.ana[1] ;
 wire \top_I.branch[15].block[9].um_I.ana[2] ;
 wire \top_I.branch[15].block[9].um_I.ana[3] ;
 wire \top_I.branch[15].block[9].um_I.ana[4] ;
 wire \top_I.branch[15].block[9].um_I.ana[5] ;
 wire \top_I.branch[15].block[9].um_I.ana[6] ;
 wire \top_I.branch[15].block[9].um_I.ana[7] ;
 wire \top_I.branch[15].block[9].um_I.clk ;
 wire \top_I.branch[15].block[9].um_I.ena ;
 wire \top_I.branch[15].block[9].um_I.iw[10] ;
 wire \top_I.branch[15].block[9].um_I.iw[11] ;
 wire \top_I.branch[15].block[9].um_I.iw[12] ;
 wire \top_I.branch[15].block[9].um_I.iw[13] ;
 wire \top_I.branch[15].block[9].um_I.iw[14] ;
 wire \top_I.branch[15].block[9].um_I.iw[15] ;
 wire \top_I.branch[15].block[9].um_I.iw[16] ;
 wire \top_I.branch[15].block[9].um_I.iw[17] ;
 wire \top_I.branch[15].block[9].um_I.iw[1] ;
 wire \top_I.branch[15].block[9].um_I.iw[2] ;
 wire \top_I.branch[15].block[9].um_I.iw[3] ;
 wire \top_I.branch[15].block[9].um_I.iw[4] ;
 wire \top_I.branch[15].block[9].um_I.iw[5] ;
 wire \top_I.branch[15].block[9].um_I.iw[6] ;
 wire \top_I.branch[15].block[9].um_I.iw[7] ;
 wire \top_I.branch[15].block[9].um_I.iw[8] ;
 wire \top_I.branch[15].block[9].um_I.iw[9] ;
 wire \top_I.branch[15].block[9].um_I.k_zero ;
 wire \top_I.branch[15].block[9].um_I.pg_vdd ;
 wire \top_I.branch[15].l_addr[0] ;
 wire \top_I.branch[15].l_addr[3] ;
 wire \top_I.branch[16].block[0].um_I.ana[0] ;
 wire \top_I.branch[16].block[0].um_I.ana[1] ;
 wire \top_I.branch[16].block[0].um_I.ana[2] ;
 wire \top_I.branch[16].block[0].um_I.ana[3] ;
 wire \top_I.branch[16].block[0].um_I.ana[4] ;
 wire \top_I.branch[16].block[0].um_I.ana[5] ;
 wire \top_I.branch[16].block[0].um_I.ana[6] ;
 wire \top_I.branch[16].block[0].um_I.ana[7] ;
 wire \top_I.branch[16].block[0].um_I.clk ;
 wire \top_I.branch[16].block[0].um_I.ena ;
 wire \top_I.branch[16].block[0].um_I.iw[10] ;
 wire \top_I.branch[16].block[0].um_I.iw[11] ;
 wire \top_I.branch[16].block[0].um_I.iw[12] ;
 wire \top_I.branch[16].block[0].um_I.iw[13] ;
 wire \top_I.branch[16].block[0].um_I.iw[14] ;
 wire \top_I.branch[16].block[0].um_I.iw[15] ;
 wire \top_I.branch[16].block[0].um_I.iw[16] ;
 wire \top_I.branch[16].block[0].um_I.iw[17] ;
 wire \top_I.branch[16].block[0].um_I.iw[1] ;
 wire \top_I.branch[16].block[0].um_I.iw[2] ;
 wire \top_I.branch[16].block[0].um_I.iw[3] ;
 wire \top_I.branch[16].block[0].um_I.iw[4] ;
 wire \top_I.branch[16].block[0].um_I.iw[5] ;
 wire \top_I.branch[16].block[0].um_I.iw[6] ;
 wire \top_I.branch[16].block[0].um_I.iw[7] ;
 wire \top_I.branch[16].block[0].um_I.iw[8] ;
 wire \top_I.branch[16].block[0].um_I.iw[9] ;
 wire \top_I.branch[16].block[0].um_I.k_zero ;
 wire \top_I.branch[16].block[0].um_I.pg_vdd ;
 wire \top_I.branch[16].block[10].um_I.ana[0] ;
 wire \top_I.branch[16].block[10].um_I.ana[1] ;
 wire \top_I.branch[16].block[10].um_I.ana[2] ;
 wire \top_I.branch[16].block[10].um_I.ana[3] ;
 wire \top_I.branch[16].block[10].um_I.ana[4] ;
 wire \top_I.branch[16].block[10].um_I.ana[5] ;
 wire \top_I.branch[16].block[10].um_I.ana[6] ;
 wire \top_I.branch[16].block[10].um_I.ana[7] ;
 wire \top_I.branch[16].block[10].um_I.clk ;
 wire \top_I.branch[16].block[10].um_I.ena ;
 wire \top_I.branch[16].block[10].um_I.iw[10] ;
 wire \top_I.branch[16].block[10].um_I.iw[11] ;
 wire \top_I.branch[16].block[10].um_I.iw[12] ;
 wire \top_I.branch[16].block[10].um_I.iw[13] ;
 wire \top_I.branch[16].block[10].um_I.iw[14] ;
 wire \top_I.branch[16].block[10].um_I.iw[15] ;
 wire \top_I.branch[16].block[10].um_I.iw[16] ;
 wire \top_I.branch[16].block[10].um_I.iw[17] ;
 wire \top_I.branch[16].block[10].um_I.iw[1] ;
 wire \top_I.branch[16].block[10].um_I.iw[2] ;
 wire \top_I.branch[16].block[10].um_I.iw[3] ;
 wire \top_I.branch[16].block[10].um_I.iw[4] ;
 wire \top_I.branch[16].block[10].um_I.iw[5] ;
 wire \top_I.branch[16].block[10].um_I.iw[6] ;
 wire \top_I.branch[16].block[10].um_I.iw[7] ;
 wire \top_I.branch[16].block[10].um_I.iw[8] ;
 wire \top_I.branch[16].block[10].um_I.iw[9] ;
 wire \top_I.branch[16].block[10].um_I.k_zero ;
 wire \top_I.branch[16].block[10].um_I.pg_vdd ;
 wire \top_I.branch[16].block[11].um_I.ana[0] ;
 wire \top_I.branch[16].block[11].um_I.ana[1] ;
 wire \top_I.branch[16].block[11].um_I.ana[2] ;
 wire \top_I.branch[16].block[11].um_I.ana[3] ;
 wire \top_I.branch[16].block[11].um_I.ana[4] ;
 wire \top_I.branch[16].block[11].um_I.ana[5] ;
 wire \top_I.branch[16].block[11].um_I.ana[6] ;
 wire \top_I.branch[16].block[11].um_I.ana[7] ;
 wire \top_I.branch[16].block[11].um_I.clk ;
 wire \top_I.branch[16].block[11].um_I.ena ;
 wire \top_I.branch[16].block[11].um_I.iw[10] ;
 wire \top_I.branch[16].block[11].um_I.iw[11] ;
 wire \top_I.branch[16].block[11].um_I.iw[12] ;
 wire \top_I.branch[16].block[11].um_I.iw[13] ;
 wire \top_I.branch[16].block[11].um_I.iw[14] ;
 wire \top_I.branch[16].block[11].um_I.iw[15] ;
 wire \top_I.branch[16].block[11].um_I.iw[16] ;
 wire \top_I.branch[16].block[11].um_I.iw[17] ;
 wire \top_I.branch[16].block[11].um_I.iw[1] ;
 wire \top_I.branch[16].block[11].um_I.iw[2] ;
 wire \top_I.branch[16].block[11].um_I.iw[3] ;
 wire \top_I.branch[16].block[11].um_I.iw[4] ;
 wire \top_I.branch[16].block[11].um_I.iw[5] ;
 wire \top_I.branch[16].block[11].um_I.iw[6] ;
 wire \top_I.branch[16].block[11].um_I.iw[7] ;
 wire \top_I.branch[16].block[11].um_I.iw[8] ;
 wire \top_I.branch[16].block[11].um_I.iw[9] ;
 wire \top_I.branch[16].block[11].um_I.k_zero ;
 wire \top_I.branch[16].block[11].um_I.pg_vdd ;
 wire \top_I.branch[16].block[12].um_I.ana[0] ;
 wire \top_I.branch[16].block[12].um_I.ana[1] ;
 wire \top_I.branch[16].block[12].um_I.ana[2] ;
 wire \top_I.branch[16].block[12].um_I.ana[3] ;
 wire \top_I.branch[16].block[12].um_I.ana[4] ;
 wire \top_I.branch[16].block[12].um_I.ana[5] ;
 wire \top_I.branch[16].block[12].um_I.ana[6] ;
 wire \top_I.branch[16].block[12].um_I.ana[7] ;
 wire \top_I.branch[16].block[12].um_I.clk ;
 wire \top_I.branch[16].block[12].um_I.ena ;
 wire \top_I.branch[16].block[12].um_I.iw[10] ;
 wire \top_I.branch[16].block[12].um_I.iw[11] ;
 wire \top_I.branch[16].block[12].um_I.iw[12] ;
 wire \top_I.branch[16].block[12].um_I.iw[13] ;
 wire \top_I.branch[16].block[12].um_I.iw[14] ;
 wire \top_I.branch[16].block[12].um_I.iw[15] ;
 wire \top_I.branch[16].block[12].um_I.iw[16] ;
 wire \top_I.branch[16].block[12].um_I.iw[17] ;
 wire \top_I.branch[16].block[12].um_I.iw[1] ;
 wire \top_I.branch[16].block[12].um_I.iw[2] ;
 wire \top_I.branch[16].block[12].um_I.iw[3] ;
 wire \top_I.branch[16].block[12].um_I.iw[4] ;
 wire \top_I.branch[16].block[12].um_I.iw[5] ;
 wire \top_I.branch[16].block[12].um_I.iw[6] ;
 wire \top_I.branch[16].block[12].um_I.iw[7] ;
 wire \top_I.branch[16].block[12].um_I.iw[8] ;
 wire \top_I.branch[16].block[12].um_I.iw[9] ;
 wire \top_I.branch[16].block[12].um_I.k_zero ;
 wire \top_I.branch[16].block[12].um_I.pg_vdd ;
 wire \top_I.branch[16].block[13].um_I.ana[0] ;
 wire \top_I.branch[16].block[13].um_I.ana[1] ;
 wire \top_I.branch[16].block[13].um_I.ana[2] ;
 wire \top_I.branch[16].block[13].um_I.ana[3] ;
 wire \top_I.branch[16].block[13].um_I.ana[4] ;
 wire \top_I.branch[16].block[13].um_I.ana[5] ;
 wire \top_I.branch[16].block[13].um_I.ana[6] ;
 wire \top_I.branch[16].block[13].um_I.ana[7] ;
 wire \top_I.branch[16].block[13].um_I.clk ;
 wire \top_I.branch[16].block[13].um_I.ena ;
 wire \top_I.branch[16].block[13].um_I.iw[10] ;
 wire \top_I.branch[16].block[13].um_I.iw[11] ;
 wire \top_I.branch[16].block[13].um_I.iw[12] ;
 wire \top_I.branch[16].block[13].um_I.iw[13] ;
 wire \top_I.branch[16].block[13].um_I.iw[14] ;
 wire \top_I.branch[16].block[13].um_I.iw[15] ;
 wire \top_I.branch[16].block[13].um_I.iw[16] ;
 wire \top_I.branch[16].block[13].um_I.iw[17] ;
 wire \top_I.branch[16].block[13].um_I.iw[1] ;
 wire \top_I.branch[16].block[13].um_I.iw[2] ;
 wire \top_I.branch[16].block[13].um_I.iw[3] ;
 wire \top_I.branch[16].block[13].um_I.iw[4] ;
 wire \top_I.branch[16].block[13].um_I.iw[5] ;
 wire \top_I.branch[16].block[13].um_I.iw[6] ;
 wire \top_I.branch[16].block[13].um_I.iw[7] ;
 wire \top_I.branch[16].block[13].um_I.iw[8] ;
 wire \top_I.branch[16].block[13].um_I.iw[9] ;
 wire \top_I.branch[16].block[13].um_I.k_zero ;
 wire \top_I.branch[16].block[13].um_I.pg_vdd ;
 wire \top_I.branch[16].block[14].um_I.ana[0] ;
 wire \top_I.branch[16].block[14].um_I.ana[1] ;
 wire \top_I.branch[16].block[14].um_I.ana[2] ;
 wire \top_I.branch[16].block[14].um_I.ana[3] ;
 wire \top_I.branch[16].block[14].um_I.ana[4] ;
 wire \top_I.branch[16].block[14].um_I.ana[5] ;
 wire \top_I.branch[16].block[14].um_I.ana[6] ;
 wire \top_I.branch[16].block[14].um_I.ana[7] ;
 wire \top_I.branch[16].block[14].um_I.clk ;
 wire \top_I.branch[16].block[14].um_I.ena ;
 wire \top_I.branch[16].block[14].um_I.iw[10] ;
 wire \top_I.branch[16].block[14].um_I.iw[11] ;
 wire \top_I.branch[16].block[14].um_I.iw[12] ;
 wire \top_I.branch[16].block[14].um_I.iw[13] ;
 wire \top_I.branch[16].block[14].um_I.iw[14] ;
 wire \top_I.branch[16].block[14].um_I.iw[15] ;
 wire \top_I.branch[16].block[14].um_I.iw[16] ;
 wire \top_I.branch[16].block[14].um_I.iw[17] ;
 wire \top_I.branch[16].block[14].um_I.iw[1] ;
 wire \top_I.branch[16].block[14].um_I.iw[2] ;
 wire \top_I.branch[16].block[14].um_I.iw[3] ;
 wire \top_I.branch[16].block[14].um_I.iw[4] ;
 wire \top_I.branch[16].block[14].um_I.iw[5] ;
 wire \top_I.branch[16].block[14].um_I.iw[6] ;
 wire \top_I.branch[16].block[14].um_I.iw[7] ;
 wire \top_I.branch[16].block[14].um_I.iw[8] ;
 wire \top_I.branch[16].block[14].um_I.iw[9] ;
 wire \top_I.branch[16].block[14].um_I.k_zero ;
 wire \top_I.branch[16].block[14].um_I.pg_vdd ;
 wire \top_I.branch[16].block[15].um_I.ana[0] ;
 wire \top_I.branch[16].block[15].um_I.ana[1] ;
 wire \top_I.branch[16].block[15].um_I.ana[2] ;
 wire \top_I.branch[16].block[15].um_I.ana[3] ;
 wire \top_I.branch[16].block[15].um_I.ana[4] ;
 wire \top_I.branch[16].block[15].um_I.ana[5] ;
 wire \top_I.branch[16].block[15].um_I.ana[6] ;
 wire \top_I.branch[16].block[15].um_I.ana[7] ;
 wire \top_I.branch[16].block[15].um_I.clk ;
 wire \top_I.branch[16].block[15].um_I.ena ;
 wire \top_I.branch[16].block[15].um_I.iw[10] ;
 wire \top_I.branch[16].block[15].um_I.iw[11] ;
 wire \top_I.branch[16].block[15].um_I.iw[12] ;
 wire \top_I.branch[16].block[15].um_I.iw[13] ;
 wire \top_I.branch[16].block[15].um_I.iw[14] ;
 wire \top_I.branch[16].block[15].um_I.iw[15] ;
 wire \top_I.branch[16].block[15].um_I.iw[16] ;
 wire \top_I.branch[16].block[15].um_I.iw[17] ;
 wire \top_I.branch[16].block[15].um_I.iw[1] ;
 wire \top_I.branch[16].block[15].um_I.iw[2] ;
 wire \top_I.branch[16].block[15].um_I.iw[3] ;
 wire \top_I.branch[16].block[15].um_I.iw[4] ;
 wire \top_I.branch[16].block[15].um_I.iw[5] ;
 wire \top_I.branch[16].block[15].um_I.iw[6] ;
 wire \top_I.branch[16].block[15].um_I.iw[7] ;
 wire \top_I.branch[16].block[15].um_I.iw[8] ;
 wire \top_I.branch[16].block[15].um_I.iw[9] ;
 wire \top_I.branch[16].block[15].um_I.k_zero ;
 wire \top_I.branch[16].block[15].um_I.pg_vdd ;
 wire \top_I.branch[16].block[1].um_I.ana[0] ;
 wire \top_I.branch[16].block[1].um_I.ana[1] ;
 wire \top_I.branch[16].block[1].um_I.ana[2] ;
 wire \top_I.branch[16].block[1].um_I.ana[3] ;
 wire \top_I.branch[16].block[1].um_I.ana[4] ;
 wire \top_I.branch[16].block[1].um_I.ana[5] ;
 wire \top_I.branch[16].block[1].um_I.ana[6] ;
 wire \top_I.branch[16].block[1].um_I.ana[7] ;
 wire \top_I.branch[16].block[1].um_I.clk ;
 wire \top_I.branch[16].block[1].um_I.ena ;
 wire \top_I.branch[16].block[1].um_I.iw[10] ;
 wire \top_I.branch[16].block[1].um_I.iw[11] ;
 wire \top_I.branch[16].block[1].um_I.iw[12] ;
 wire \top_I.branch[16].block[1].um_I.iw[13] ;
 wire \top_I.branch[16].block[1].um_I.iw[14] ;
 wire \top_I.branch[16].block[1].um_I.iw[15] ;
 wire \top_I.branch[16].block[1].um_I.iw[16] ;
 wire \top_I.branch[16].block[1].um_I.iw[17] ;
 wire \top_I.branch[16].block[1].um_I.iw[1] ;
 wire \top_I.branch[16].block[1].um_I.iw[2] ;
 wire \top_I.branch[16].block[1].um_I.iw[3] ;
 wire \top_I.branch[16].block[1].um_I.iw[4] ;
 wire \top_I.branch[16].block[1].um_I.iw[5] ;
 wire \top_I.branch[16].block[1].um_I.iw[6] ;
 wire \top_I.branch[16].block[1].um_I.iw[7] ;
 wire \top_I.branch[16].block[1].um_I.iw[8] ;
 wire \top_I.branch[16].block[1].um_I.iw[9] ;
 wire \top_I.branch[16].block[1].um_I.k_zero ;
 wire \top_I.branch[16].block[1].um_I.pg_vdd ;
 wire \top_I.branch[16].block[2].um_I.ana[0] ;
 wire \top_I.branch[16].block[2].um_I.ana[1] ;
 wire \top_I.branch[16].block[2].um_I.ana[2] ;
 wire \top_I.branch[16].block[2].um_I.ana[3] ;
 wire \top_I.branch[16].block[2].um_I.ana[4] ;
 wire \top_I.branch[16].block[2].um_I.ana[5] ;
 wire \top_I.branch[16].block[2].um_I.ana[6] ;
 wire \top_I.branch[16].block[2].um_I.ana[7] ;
 wire \top_I.branch[16].block[2].um_I.clk ;
 wire \top_I.branch[16].block[2].um_I.ena ;
 wire \top_I.branch[16].block[2].um_I.iw[10] ;
 wire \top_I.branch[16].block[2].um_I.iw[11] ;
 wire \top_I.branch[16].block[2].um_I.iw[12] ;
 wire \top_I.branch[16].block[2].um_I.iw[13] ;
 wire \top_I.branch[16].block[2].um_I.iw[14] ;
 wire \top_I.branch[16].block[2].um_I.iw[15] ;
 wire \top_I.branch[16].block[2].um_I.iw[16] ;
 wire \top_I.branch[16].block[2].um_I.iw[17] ;
 wire \top_I.branch[16].block[2].um_I.iw[1] ;
 wire \top_I.branch[16].block[2].um_I.iw[2] ;
 wire \top_I.branch[16].block[2].um_I.iw[3] ;
 wire \top_I.branch[16].block[2].um_I.iw[4] ;
 wire \top_I.branch[16].block[2].um_I.iw[5] ;
 wire \top_I.branch[16].block[2].um_I.iw[6] ;
 wire \top_I.branch[16].block[2].um_I.iw[7] ;
 wire \top_I.branch[16].block[2].um_I.iw[8] ;
 wire \top_I.branch[16].block[2].um_I.iw[9] ;
 wire \top_I.branch[16].block[2].um_I.k_zero ;
 wire \top_I.branch[16].block[2].um_I.pg_vdd ;
 wire \top_I.branch[16].block[3].um_I.ana[0] ;
 wire \top_I.branch[16].block[3].um_I.ana[1] ;
 wire \top_I.branch[16].block[3].um_I.ana[2] ;
 wire \top_I.branch[16].block[3].um_I.ana[3] ;
 wire \top_I.branch[16].block[3].um_I.ana[4] ;
 wire \top_I.branch[16].block[3].um_I.ana[5] ;
 wire \top_I.branch[16].block[3].um_I.ana[6] ;
 wire \top_I.branch[16].block[3].um_I.ana[7] ;
 wire \top_I.branch[16].block[3].um_I.clk ;
 wire \top_I.branch[16].block[3].um_I.ena ;
 wire \top_I.branch[16].block[3].um_I.iw[10] ;
 wire \top_I.branch[16].block[3].um_I.iw[11] ;
 wire \top_I.branch[16].block[3].um_I.iw[12] ;
 wire \top_I.branch[16].block[3].um_I.iw[13] ;
 wire \top_I.branch[16].block[3].um_I.iw[14] ;
 wire \top_I.branch[16].block[3].um_I.iw[15] ;
 wire \top_I.branch[16].block[3].um_I.iw[16] ;
 wire \top_I.branch[16].block[3].um_I.iw[17] ;
 wire \top_I.branch[16].block[3].um_I.iw[1] ;
 wire \top_I.branch[16].block[3].um_I.iw[2] ;
 wire \top_I.branch[16].block[3].um_I.iw[3] ;
 wire \top_I.branch[16].block[3].um_I.iw[4] ;
 wire \top_I.branch[16].block[3].um_I.iw[5] ;
 wire \top_I.branch[16].block[3].um_I.iw[6] ;
 wire \top_I.branch[16].block[3].um_I.iw[7] ;
 wire \top_I.branch[16].block[3].um_I.iw[8] ;
 wire \top_I.branch[16].block[3].um_I.iw[9] ;
 wire \top_I.branch[16].block[3].um_I.k_zero ;
 wire \top_I.branch[16].block[3].um_I.pg_vdd ;
 wire \top_I.branch[16].block[4].um_I.ana[0] ;
 wire \top_I.branch[16].block[4].um_I.ana[1] ;
 wire \top_I.branch[16].block[4].um_I.ana[2] ;
 wire \top_I.branch[16].block[4].um_I.ana[3] ;
 wire \top_I.branch[16].block[4].um_I.ana[4] ;
 wire \top_I.branch[16].block[4].um_I.ana[5] ;
 wire \top_I.branch[16].block[4].um_I.ana[6] ;
 wire \top_I.branch[16].block[4].um_I.ana[7] ;
 wire \top_I.branch[16].block[4].um_I.clk ;
 wire \top_I.branch[16].block[4].um_I.ena ;
 wire \top_I.branch[16].block[4].um_I.iw[10] ;
 wire \top_I.branch[16].block[4].um_I.iw[11] ;
 wire \top_I.branch[16].block[4].um_I.iw[12] ;
 wire \top_I.branch[16].block[4].um_I.iw[13] ;
 wire \top_I.branch[16].block[4].um_I.iw[14] ;
 wire \top_I.branch[16].block[4].um_I.iw[15] ;
 wire \top_I.branch[16].block[4].um_I.iw[16] ;
 wire \top_I.branch[16].block[4].um_I.iw[17] ;
 wire \top_I.branch[16].block[4].um_I.iw[1] ;
 wire \top_I.branch[16].block[4].um_I.iw[2] ;
 wire \top_I.branch[16].block[4].um_I.iw[3] ;
 wire \top_I.branch[16].block[4].um_I.iw[4] ;
 wire \top_I.branch[16].block[4].um_I.iw[5] ;
 wire \top_I.branch[16].block[4].um_I.iw[6] ;
 wire \top_I.branch[16].block[4].um_I.iw[7] ;
 wire \top_I.branch[16].block[4].um_I.iw[8] ;
 wire \top_I.branch[16].block[4].um_I.iw[9] ;
 wire \top_I.branch[16].block[4].um_I.k_zero ;
 wire \top_I.branch[16].block[4].um_I.pg_vdd ;
 wire \top_I.branch[16].block[5].um_I.ana[0] ;
 wire \top_I.branch[16].block[5].um_I.ana[1] ;
 wire \top_I.branch[16].block[5].um_I.ana[2] ;
 wire \top_I.branch[16].block[5].um_I.ana[3] ;
 wire \top_I.branch[16].block[5].um_I.ana[4] ;
 wire \top_I.branch[16].block[5].um_I.ana[5] ;
 wire \top_I.branch[16].block[5].um_I.ana[6] ;
 wire \top_I.branch[16].block[5].um_I.ana[7] ;
 wire \top_I.branch[16].block[5].um_I.clk ;
 wire \top_I.branch[16].block[5].um_I.ena ;
 wire \top_I.branch[16].block[5].um_I.iw[10] ;
 wire \top_I.branch[16].block[5].um_I.iw[11] ;
 wire \top_I.branch[16].block[5].um_I.iw[12] ;
 wire \top_I.branch[16].block[5].um_I.iw[13] ;
 wire \top_I.branch[16].block[5].um_I.iw[14] ;
 wire \top_I.branch[16].block[5].um_I.iw[15] ;
 wire \top_I.branch[16].block[5].um_I.iw[16] ;
 wire \top_I.branch[16].block[5].um_I.iw[17] ;
 wire \top_I.branch[16].block[5].um_I.iw[1] ;
 wire \top_I.branch[16].block[5].um_I.iw[2] ;
 wire \top_I.branch[16].block[5].um_I.iw[3] ;
 wire \top_I.branch[16].block[5].um_I.iw[4] ;
 wire \top_I.branch[16].block[5].um_I.iw[5] ;
 wire \top_I.branch[16].block[5].um_I.iw[6] ;
 wire \top_I.branch[16].block[5].um_I.iw[7] ;
 wire \top_I.branch[16].block[5].um_I.iw[8] ;
 wire \top_I.branch[16].block[5].um_I.iw[9] ;
 wire \top_I.branch[16].block[5].um_I.k_zero ;
 wire \top_I.branch[16].block[5].um_I.pg_vdd ;
 wire \top_I.branch[16].block[6].um_I.ana[0] ;
 wire \top_I.branch[16].block[6].um_I.ana[1] ;
 wire \top_I.branch[16].block[6].um_I.ana[2] ;
 wire \top_I.branch[16].block[6].um_I.ana[3] ;
 wire \top_I.branch[16].block[6].um_I.ana[4] ;
 wire \top_I.branch[16].block[6].um_I.ana[5] ;
 wire \top_I.branch[16].block[6].um_I.ana[6] ;
 wire \top_I.branch[16].block[6].um_I.ana[7] ;
 wire \top_I.branch[16].block[6].um_I.clk ;
 wire \top_I.branch[16].block[6].um_I.ena ;
 wire \top_I.branch[16].block[6].um_I.iw[10] ;
 wire \top_I.branch[16].block[6].um_I.iw[11] ;
 wire \top_I.branch[16].block[6].um_I.iw[12] ;
 wire \top_I.branch[16].block[6].um_I.iw[13] ;
 wire \top_I.branch[16].block[6].um_I.iw[14] ;
 wire \top_I.branch[16].block[6].um_I.iw[15] ;
 wire \top_I.branch[16].block[6].um_I.iw[16] ;
 wire \top_I.branch[16].block[6].um_I.iw[17] ;
 wire \top_I.branch[16].block[6].um_I.iw[1] ;
 wire \top_I.branch[16].block[6].um_I.iw[2] ;
 wire \top_I.branch[16].block[6].um_I.iw[3] ;
 wire \top_I.branch[16].block[6].um_I.iw[4] ;
 wire \top_I.branch[16].block[6].um_I.iw[5] ;
 wire \top_I.branch[16].block[6].um_I.iw[6] ;
 wire \top_I.branch[16].block[6].um_I.iw[7] ;
 wire \top_I.branch[16].block[6].um_I.iw[8] ;
 wire \top_I.branch[16].block[6].um_I.iw[9] ;
 wire \top_I.branch[16].block[6].um_I.k_zero ;
 wire \top_I.branch[16].block[6].um_I.pg_vdd ;
 wire \top_I.branch[16].block[7].um_I.ana[0] ;
 wire \top_I.branch[16].block[7].um_I.ana[1] ;
 wire \top_I.branch[16].block[7].um_I.ana[2] ;
 wire \top_I.branch[16].block[7].um_I.ana[3] ;
 wire \top_I.branch[16].block[7].um_I.ana[4] ;
 wire \top_I.branch[16].block[7].um_I.ana[5] ;
 wire \top_I.branch[16].block[7].um_I.ana[6] ;
 wire \top_I.branch[16].block[7].um_I.ana[7] ;
 wire \top_I.branch[16].block[7].um_I.clk ;
 wire \top_I.branch[16].block[7].um_I.ena ;
 wire \top_I.branch[16].block[7].um_I.iw[10] ;
 wire \top_I.branch[16].block[7].um_I.iw[11] ;
 wire \top_I.branch[16].block[7].um_I.iw[12] ;
 wire \top_I.branch[16].block[7].um_I.iw[13] ;
 wire \top_I.branch[16].block[7].um_I.iw[14] ;
 wire \top_I.branch[16].block[7].um_I.iw[15] ;
 wire \top_I.branch[16].block[7].um_I.iw[16] ;
 wire \top_I.branch[16].block[7].um_I.iw[17] ;
 wire \top_I.branch[16].block[7].um_I.iw[1] ;
 wire \top_I.branch[16].block[7].um_I.iw[2] ;
 wire \top_I.branch[16].block[7].um_I.iw[3] ;
 wire \top_I.branch[16].block[7].um_I.iw[4] ;
 wire \top_I.branch[16].block[7].um_I.iw[5] ;
 wire \top_I.branch[16].block[7].um_I.iw[6] ;
 wire \top_I.branch[16].block[7].um_I.iw[7] ;
 wire \top_I.branch[16].block[7].um_I.iw[8] ;
 wire \top_I.branch[16].block[7].um_I.iw[9] ;
 wire \top_I.branch[16].block[7].um_I.k_zero ;
 wire \top_I.branch[16].block[7].um_I.pg_vdd ;
 wire \top_I.branch[16].block[8].um_I.ana[0] ;
 wire \top_I.branch[16].block[8].um_I.ana[1] ;
 wire \top_I.branch[16].block[8].um_I.ana[2] ;
 wire \top_I.branch[16].block[8].um_I.ana[3] ;
 wire \top_I.branch[16].block[8].um_I.ana[4] ;
 wire \top_I.branch[16].block[8].um_I.ana[5] ;
 wire \top_I.branch[16].block[8].um_I.ana[6] ;
 wire \top_I.branch[16].block[8].um_I.ana[7] ;
 wire \top_I.branch[16].block[8].um_I.clk ;
 wire \top_I.branch[16].block[8].um_I.ena ;
 wire \top_I.branch[16].block[8].um_I.iw[10] ;
 wire \top_I.branch[16].block[8].um_I.iw[11] ;
 wire \top_I.branch[16].block[8].um_I.iw[12] ;
 wire \top_I.branch[16].block[8].um_I.iw[13] ;
 wire \top_I.branch[16].block[8].um_I.iw[14] ;
 wire \top_I.branch[16].block[8].um_I.iw[15] ;
 wire \top_I.branch[16].block[8].um_I.iw[16] ;
 wire \top_I.branch[16].block[8].um_I.iw[17] ;
 wire \top_I.branch[16].block[8].um_I.iw[1] ;
 wire \top_I.branch[16].block[8].um_I.iw[2] ;
 wire \top_I.branch[16].block[8].um_I.iw[3] ;
 wire \top_I.branch[16].block[8].um_I.iw[4] ;
 wire \top_I.branch[16].block[8].um_I.iw[5] ;
 wire \top_I.branch[16].block[8].um_I.iw[6] ;
 wire \top_I.branch[16].block[8].um_I.iw[7] ;
 wire \top_I.branch[16].block[8].um_I.iw[8] ;
 wire \top_I.branch[16].block[8].um_I.iw[9] ;
 wire \top_I.branch[16].block[8].um_I.k_zero ;
 wire \top_I.branch[16].block[8].um_I.pg_vdd ;
 wire \top_I.branch[16].block[9].um_I.ana[0] ;
 wire \top_I.branch[16].block[9].um_I.ana[1] ;
 wire \top_I.branch[16].block[9].um_I.ana[2] ;
 wire \top_I.branch[16].block[9].um_I.ana[3] ;
 wire \top_I.branch[16].block[9].um_I.ana[4] ;
 wire \top_I.branch[16].block[9].um_I.ana[5] ;
 wire \top_I.branch[16].block[9].um_I.ana[6] ;
 wire \top_I.branch[16].block[9].um_I.ana[7] ;
 wire \top_I.branch[16].block[9].um_I.clk ;
 wire \top_I.branch[16].block[9].um_I.ena ;
 wire \top_I.branch[16].block[9].um_I.iw[10] ;
 wire \top_I.branch[16].block[9].um_I.iw[11] ;
 wire \top_I.branch[16].block[9].um_I.iw[12] ;
 wire \top_I.branch[16].block[9].um_I.iw[13] ;
 wire \top_I.branch[16].block[9].um_I.iw[14] ;
 wire \top_I.branch[16].block[9].um_I.iw[15] ;
 wire \top_I.branch[16].block[9].um_I.iw[16] ;
 wire \top_I.branch[16].block[9].um_I.iw[17] ;
 wire \top_I.branch[16].block[9].um_I.iw[1] ;
 wire \top_I.branch[16].block[9].um_I.iw[2] ;
 wire \top_I.branch[16].block[9].um_I.iw[3] ;
 wire \top_I.branch[16].block[9].um_I.iw[4] ;
 wire \top_I.branch[16].block[9].um_I.iw[5] ;
 wire \top_I.branch[16].block[9].um_I.iw[6] ;
 wire \top_I.branch[16].block[9].um_I.iw[7] ;
 wire \top_I.branch[16].block[9].um_I.iw[8] ;
 wire \top_I.branch[16].block[9].um_I.iw[9] ;
 wire \top_I.branch[16].block[9].um_I.k_zero ;
 wire \top_I.branch[16].block[9].um_I.pg_vdd ;
 wire \top_I.branch[16].l_addr[0] ;
 wire \top_I.branch[16].l_addr[3] ;
 wire \top_I.branch[17].block[0].um_I.ana[0] ;
 wire \top_I.branch[17].block[0].um_I.ana[1] ;
 wire \top_I.branch[17].block[0].um_I.ana[2] ;
 wire \top_I.branch[17].block[0].um_I.ana[3] ;
 wire \top_I.branch[17].block[0].um_I.ana[4] ;
 wire \top_I.branch[17].block[0].um_I.ana[5] ;
 wire \top_I.branch[17].block[0].um_I.ana[6] ;
 wire \top_I.branch[17].block[0].um_I.ana[7] ;
 wire \top_I.branch[17].block[0].um_I.clk ;
 wire \top_I.branch[17].block[0].um_I.ena ;
 wire \top_I.branch[17].block[0].um_I.iw[10] ;
 wire \top_I.branch[17].block[0].um_I.iw[11] ;
 wire \top_I.branch[17].block[0].um_I.iw[12] ;
 wire \top_I.branch[17].block[0].um_I.iw[13] ;
 wire \top_I.branch[17].block[0].um_I.iw[14] ;
 wire \top_I.branch[17].block[0].um_I.iw[15] ;
 wire \top_I.branch[17].block[0].um_I.iw[16] ;
 wire \top_I.branch[17].block[0].um_I.iw[17] ;
 wire \top_I.branch[17].block[0].um_I.iw[1] ;
 wire \top_I.branch[17].block[0].um_I.iw[2] ;
 wire \top_I.branch[17].block[0].um_I.iw[3] ;
 wire \top_I.branch[17].block[0].um_I.iw[4] ;
 wire \top_I.branch[17].block[0].um_I.iw[5] ;
 wire \top_I.branch[17].block[0].um_I.iw[6] ;
 wire \top_I.branch[17].block[0].um_I.iw[7] ;
 wire \top_I.branch[17].block[0].um_I.iw[8] ;
 wire \top_I.branch[17].block[0].um_I.iw[9] ;
 wire \top_I.branch[17].block[0].um_I.k_zero ;
 wire \top_I.branch[17].block[0].um_I.pg_vdd ;
 wire \top_I.branch[17].block[10].um_I.ana[0] ;
 wire \top_I.branch[17].block[10].um_I.ana[1] ;
 wire \top_I.branch[17].block[10].um_I.ana[2] ;
 wire \top_I.branch[17].block[10].um_I.ana[3] ;
 wire \top_I.branch[17].block[10].um_I.ana[4] ;
 wire \top_I.branch[17].block[10].um_I.ana[5] ;
 wire \top_I.branch[17].block[10].um_I.ana[6] ;
 wire \top_I.branch[17].block[10].um_I.ana[7] ;
 wire \top_I.branch[17].block[10].um_I.clk ;
 wire \top_I.branch[17].block[10].um_I.ena ;
 wire \top_I.branch[17].block[10].um_I.iw[10] ;
 wire \top_I.branch[17].block[10].um_I.iw[11] ;
 wire \top_I.branch[17].block[10].um_I.iw[12] ;
 wire \top_I.branch[17].block[10].um_I.iw[13] ;
 wire \top_I.branch[17].block[10].um_I.iw[14] ;
 wire \top_I.branch[17].block[10].um_I.iw[15] ;
 wire \top_I.branch[17].block[10].um_I.iw[16] ;
 wire \top_I.branch[17].block[10].um_I.iw[17] ;
 wire \top_I.branch[17].block[10].um_I.iw[1] ;
 wire \top_I.branch[17].block[10].um_I.iw[2] ;
 wire \top_I.branch[17].block[10].um_I.iw[3] ;
 wire \top_I.branch[17].block[10].um_I.iw[4] ;
 wire \top_I.branch[17].block[10].um_I.iw[5] ;
 wire \top_I.branch[17].block[10].um_I.iw[6] ;
 wire \top_I.branch[17].block[10].um_I.iw[7] ;
 wire \top_I.branch[17].block[10].um_I.iw[8] ;
 wire \top_I.branch[17].block[10].um_I.iw[9] ;
 wire \top_I.branch[17].block[10].um_I.k_zero ;
 wire \top_I.branch[17].block[10].um_I.pg_vdd ;
 wire \top_I.branch[17].block[11].um_I.ana[0] ;
 wire \top_I.branch[17].block[11].um_I.ana[1] ;
 wire \top_I.branch[17].block[11].um_I.ana[2] ;
 wire \top_I.branch[17].block[11].um_I.ana[3] ;
 wire \top_I.branch[17].block[11].um_I.ana[4] ;
 wire \top_I.branch[17].block[11].um_I.ana[5] ;
 wire \top_I.branch[17].block[11].um_I.ana[6] ;
 wire \top_I.branch[17].block[11].um_I.ana[7] ;
 wire \top_I.branch[17].block[11].um_I.clk ;
 wire \top_I.branch[17].block[11].um_I.ena ;
 wire \top_I.branch[17].block[11].um_I.iw[10] ;
 wire \top_I.branch[17].block[11].um_I.iw[11] ;
 wire \top_I.branch[17].block[11].um_I.iw[12] ;
 wire \top_I.branch[17].block[11].um_I.iw[13] ;
 wire \top_I.branch[17].block[11].um_I.iw[14] ;
 wire \top_I.branch[17].block[11].um_I.iw[15] ;
 wire \top_I.branch[17].block[11].um_I.iw[16] ;
 wire \top_I.branch[17].block[11].um_I.iw[17] ;
 wire \top_I.branch[17].block[11].um_I.iw[1] ;
 wire \top_I.branch[17].block[11].um_I.iw[2] ;
 wire \top_I.branch[17].block[11].um_I.iw[3] ;
 wire \top_I.branch[17].block[11].um_I.iw[4] ;
 wire \top_I.branch[17].block[11].um_I.iw[5] ;
 wire \top_I.branch[17].block[11].um_I.iw[6] ;
 wire \top_I.branch[17].block[11].um_I.iw[7] ;
 wire \top_I.branch[17].block[11].um_I.iw[8] ;
 wire \top_I.branch[17].block[11].um_I.iw[9] ;
 wire \top_I.branch[17].block[11].um_I.k_zero ;
 wire \top_I.branch[17].block[11].um_I.pg_vdd ;
 wire \top_I.branch[17].block[12].um_I.ana[0] ;
 wire \top_I.branch[17].block[12].um_I.ana[1] ;
 wire \top_I.branch[17].block[12].um_I.ana[2] ;
 wire \top_I.branch[17].block[12].um_I.ana[3] ;
 wire \top_I.branch[17].block[12].um_I.ana[4] ;
 wire \top_I.branch[17].block[12].um_I.ana[5] ;
 wire \top_I.branch[17].block[12].um_I.ana[6] ;
 wire \top_I.branch[17].block[12].um_I.ana[7] ;
 wire \top_I.branch[17].block[12].um_I.clk ;
 wire \top_I.branch[17].block[12].um_I.ena ;
 wire \top_I.branch[17].block[12].um_I.iw[10] ;
 wire \top_I.branch[17].block[12].um_I.iw[11] ;
 wire \top_I.branch[17].block[12].um_I.iw[12] ;
 wire \top_I.branch[17].block[12].um_I.iw[13] ;
 wire \top_I.branch[17].block[12].um_I.iw[14] ;
 wire \top_I.branch[17].block[12].um_I.iw[15] ;
 wire \top_I.branch[17].block[12].um_I.iw[16] ;
 wire \top_I.branch[17].block[12].um_I.iw[17] ;
 wire \top_I.branch[17].block[12].um_I.iw[1] ;
 wire \top_I.branch[17].block[12].um_I.iw[2] ;
 wire \top_I.branch[17].block[12].um_I.iw[3] ;
 wire \top_I.branch[17].block[12].um_I.iw[4] ;
 wire \top_I.branch[17].block[12].um_I.iw[5] ;
 wire \top_I.branch[17].block[12].um_I.iw[6] ;
 wire \top_I.branch[17].block[12].um_I.iw[7] ;
 wire \top_I.branch[17].block[12].um_I.iw[8] ;
 wire \top_I.branch[17].block[12].um_I.iw[9] ;
 wire \top_I.branch[17].block[12].um_I.k_zero ;
 wire \top_I.branch[17].block[12].um_I.pg_vdd ;
 wire \top_I.branch[17].block[13].um_I.ana[0] ;
 wire \top_I.branch[17].block[13].um_I.ana[1] ;
 wire \top_I.branch[17].block[13].um_I.ana[2] ;
 wire \top_I.branch[17].block[13].um_I.ana[3] ;
 wire \top_I.branch[17].block[13].um_I.ana[4] ;
 wire \top_I.branch[17].block[13].um_I.ana[5] ;
 wire \top_I.branch[17].block[13].um_I.ana[6] ;
 wire \top_I.branch[17].block[13].um_I.ana[7] ;
 wire \top_I.branch[17].block[13].um_I.clk ;
 wire \top_I.branch[17].block[13].um_I.ena ;
 wire \top_I.branch[17].block[13].um_I.iw[10] ;
 wire \top_I.branch[17].block[13].um_I.iw[11] ;
 wire \top_I.branch[17].block[13].um_I.iw[12] ;
 wire \top_I.branch[17].block[13].um_I.iw[13] ;
 wire \top_I.branch[17].block[13].um_I.iw[14] ;
 wire \top_I.branch[17].block[13].um_I.iw[15] ;
 wire \top_I.branch[17].block[13].um_I.iw[16] ;
 wire \top_I.branch[17].block[13].um_I.iw[17] ;
 wire \top_I.branch[17].block[13].um_I.iw[1] ;
 wire \top_I.branch[17].block[13].um_I.iw[2] ;
 wire \top_I.branch[17].block[13].um_I.iw[3] ;
 wire \top_I.branch[17].block[13].um_I.iw[4] ;
 wire \top_I.branch[17].block[13].um_I.iw[5] ;
 wire \top_I.branch[17].block[13].um_I.iw[6] ;
 wire \top_I.branch[17].block[13].um_I.iw[7] ;
 wire \top_I.branch[17].block[13].um_I.iw[8] ;
 wire \top_I.branch[17].block[13].um_I.iw[9] ;
 wire \top_I.branch[17].block[13].um_I.k_zero ;
 wire \top_I.branch[17].block[13].um_I.pg_vdd ;
 wire \top_I.branch[17].block[14].um_I.ana[0] ;
 wire \top_I.branch[17].block[14].um_I.ana[1] ;
 wire \top_I.branch[17].block[14].um_I.ana[2] ;
 wire \top_I.branch[17].block[14].um_I.ana[3] ;
 wire \top_I.branch[17].block[14].um_I.ana[4] ;
 wire \top_I.branch[17].block[14].um_I.ana[5] ;
 wire \top_I.branch[17].block[14].um_I.ana[6] ;
 wire \top_I.branch[17].block[14].um_I.ana[7] ;
 wire \top_I.branch[17].block[14].um_I.clk ;
 wire \top_I.branch[17].block[14].um_I.ena ;
 wire \top_I.branch[17].block[14].um_I.iw[10] ;
 wire \top_I.branch[17].block[14].um_I.iw[11] ;
 wire \top_I.branch[17].block[14].um_I.iw[12] ;
 wire \top_I.branch[17].block[14].um_I.iw[13] ;
 wire \top_I.branch[17].block[14].um_I.iw[14] ;
 wire \top_I.branch[17].block[14].um_I.iw[15] ;
 wire \top_I.branch[17].block[14].um_I.iw[16] ;
 wire \top_I.branch[17].block[14].um_I.iw[17] ;
 wire \top_I.branch[17].block[14].um_I.iw[1] ;
 wire \top_I.branch[17].block[14].um_I.iw[2] ;
 wire \top_I.branch[17].block[14].um_I.iw[3] ;
 wire \top_I.branch[17].block[14].um_I.iw[4] ;
 wire \top_I.branch[17].block[14].um_I.iw[5] ;
 wire \top_I.branch[17].block[14].um_I.iw[6] ;
 wire \top_I.branch[17].block[14].um_I.iw[7] ;
 wire \top_I.branch[17].block[14].um_I.iw[8] ;
 wire \top_I.branch[17].block[14].um_I.iw[9] ;
 wire \top_I.branch[17].block[14].um_I.k_zero ;
 wire \top_I.branch[17].block[14].um_I.pg_vdd ;
 wire \top_I.branch[17].block[15].um_I.ana[0] ;
 wire \top_I.branch[17].block[15].um_I.ana[1] ;
 wire \top_I.branch[17].block[15].um_I.ana[2] ;
 wire \top_I.branch[17].block[15].um_I.ana[3] ;
 wire \top_I.branch[17].block[15].um_I.ana[4] ;
 wire \top_I.branch[17].block[15].um_I.ana[5] ;
 wire \top_I.branch[17].block[15].um_I.ana[6] ;
 wire \top_I.branch[17].block[15].um_I.ana[7] ;
 wire \top_I.branch[17].block[15].um_I.clk ;
 wire \top_I.branch[17].block[15].um_I.ena ;
 wire \top_I.branch[17].block[15].um_I.iw[10] ;
 wire \top_I.branch[17].block[15].um_I.iw[11] ;
 wire \top_I.branch[17].block[15].um_I.iw[12] ;
 wire \top_I.branch[17].block[15].um_I.iw[13] ;
 wire \top_I.branch[17].block[15].um_I.iw[14] ;
 wire \top_I.branch[17].block[15].um_I.iw[15] ;
 wire \top_I.branch[17].block[15].um_I.iw[16] ;
 wire \top_I.branch[17].block[15].um_I.iw[17] ;
 wire \top_I.branch[17].block[15].um_I.iw[1] ;
 wire \top_I.branch[17].block[15].um_I.iw[2] ;
 wire \top_I.branch[17].block[15].um_I.iw[3] ;
 wire \top_I.branch[17].block[15].um_I.iw[4] ;
 wire \top_I.branch[17].block[15].um_I.iw[5] ;
 wire \top_I.branch[17].block[15].um_I.iw[6] ;
 wire \top_I.branch[17].block[15].um_I.iw[7] ;
 wire \top_I.branch[17].block[15].um_I.iw[8] ;
 wire \top_I.branch[17].block[15].um_I.iw[9] ;
 wire \top_I.branch[17].block[15].um_I.k_zero ;
 wire \top_I.branch[17].block[15].um_I.pg_vdd ;
 wire \top_I.branch[17].block[1].um_I.ana[0] ;
 wire \top_I.branch[17].block[1].um_I.ana[1] ;
 wire \top_I.branch[17].block[1].um_I.ana[2] ;
 wire \top_I.branch[17].block[1].um_I.ana[3] ;
 wire \top_I.branch[17].block[1].um_I.ana[4] ;
 wire \top_I.branch[17].block[1].um_I.ana[5] ;
 wire \top_I.branch[17].block[1].um_I.ana[6] ;
 wire \top_I.branch[17].block[1].um_I.ana[7] ;
 wire \top_I.branch[17].block[1].um_I.clk ;
 wire \top_I.branch[17].block[1].um_I.ena ;
 wire \top_I.branch[17].block[1].um_I.iw[10] ;
 wire \top_I.branch[17].block[1].um_I.iw[11] ;
 wire \top_I.branch[17].block[1].um_I.iw[12] ;
 wire \top_I.branch[17].block[1].um_I.iw[13] ;
 wire \top_I.branch[17].block[1].um_I.iw[14] ;
 wire \top_I.branch[17].block[1].um_I.iw[15] ;
 wire \top_I.branch[17].block[1].um_I.iw[16] ;
 wire \top_I.branch[17].block[1].um_I.iw[17] ;
 wire \top_I.branch[17].block[1].um_I.iw[1] ;
 wire \top_I.branch[17].block[1].um_I.iw[2] ;
 wire \top_I.branch[17].block[1].um_I.iw[3] ;
 wire \top_I.branch[17].block[1].um_I.iw[4] ;
 wire \top_I.branch[17].block[1].um_I.iw[5] ;
 wire \top_I.branch[17].block[1].um_I.iw[6] ;
 wire \top_I.branch[17].block[1].um_I.iw[7] ;
 wire \top_I.branch[17].block[1].um_I.iw[8] ;
 wire \top_I.branch[17].block[1].um_I.iw[9] ;
 wire \top_I.branch[17].block[1].um_I.k_zero ;
 wire \top_I.branch[17].block[1].um_I.pg_vdd ;
 wire \top_I.branch[17].block[2].um_I.ana[0] ;
 wire \top_I.branch[17].block[2].um_I.ana[1] ;
 wire \top_I.branch[17].block[2].um_I.ana[2] ;
 wire \top_I.branch[17].block[2].um_I.ana[3] ;
 wire \top_I.branch[17].block[2].um_I.ana[4] ;
 wire \top_I.branch[17].block[2].um_I.ana[5] ;
 wire \top_I.branch[17].block[2].um_I.ana[6] ;
 wire \top_I.branch[17].block[2].um_I.ana[7] ;
 wire \top_I.branch[17].block[2].um_I.clk ;
 wire \top_I.branch[17].block[2].um_I.ena ;
 wire \top_I.branch[17].block[2].um_I.iw[10] ;
 wire \top_I.branch[17].block[2].um_I.iw[11] ;
 wire \top_I.branch[17].block[2].um_I.iw[12] ;
 wire \top_I.branch[17].block[2].um_I.iw[13] ;
 wire \top_I.branch[17].block[2].um_I.iw[14] ;
 wire \top_I.branch[17].block[2].um_I.iw[15] ;
 wire \top_I.branch[17].block[2].um_I.iw[16] ;
 wire \top_I.branch[17].block[2].um_I.iw[17] ;
 wire \top_I.branch[17].block[2].um_I.iw[1] ;
 wire \top_I.branch[17].block[2].um_I.iw[2] ;
 wire \top_I.branch[17].block[2].um_I.iw[3] ;
 wire \top_I.branch[17].block[2].um_I.iw[4] ;
 wire \top_I.branch[17].block[2].um_I.iw[5] ;
 wire \top_I.branch[17].block[2].um_I.iw[6] ;
 wire \top_I.branch[17].block[2].um_I.iw[7] ;
 wire \top_I.branch[17].block[2].um_I.iw[8] ;
 wire \top_I.branch[17].block[2].um_I.iw[9] ;
 wire \top_I.branch[17].block[2].um_I.k_zero ;
 wire \top_I.branch[17].block[2].um_I.pg_vdd ;
 wire \top_I.branch[17].block[3].um_I.ana[0] ;
 wire \top_I.branch[17].block[3].um_I.ana[1] ;
 wire \top_I.branch[17].block[3].um_I.ana[2] ;
 wire \top_I.branch[17].block[3].um_I.ana[3] ;
 wire \top_I.branch[17].block[3].um_I.ana[4] ;
 wire \top_I.branch[17].block[3].um_I.ana[5] ;
 wire \top_I.branch[17].block[3].um_I.ana[6] ;
 wire \top_I.branch[17].block[3].um_I.ana[7] ;
 wire \top_I.branch[17].block[3].um_I.clk ;
 wire \top_I.branch[17].block[3].um_I.ena ;
 wire \top_I.branch[17].block[3].um_I.iw[10] ;
 wire \top_I.branch[17].block[3].um_I.iw[11] ;
 wire \top_I.branch[17].block[3].um_I.iw[12] ;
 wire \top_I.branch[17].block[3].um_I.iw[13] ;
 wire \top_I.branch[17].block[3].um_I.iw[14] ;
 wire \top_I.branch[17].block[3].um_I.iw[15] ;
 wire \top_I.branch[17].block[3].um_I.iw[16] ;
 wire \top_I.branch[17].block[3].um_I.iw[17] ;
 wire \top_I.branch[17].block[3].um_I.iw[1] ;
 wire \top_I.branch[17].block[3].um_I.iw[2] ;
 wire \top_I.branch[17].block[3].um_I.iw[3] ;
 wire \top_I.branch[17].block[3].um_I.iw[4] ;
 wire \top_I.branch[17].block[3].um_I.iw[5] ;
 wire \top_I.branch[17].block[3].um_I.iw[6] ;
 wire \top_I.branch[17].block[3].um_I.iw[7] ;
 wire \top_I.branch[17].block[3].um_I.iw[8] ;
 wire \top_I.branch[17].block[3].um_I.iw[9] ;
 wire \top_I.branch[17].block[3].um_I.k_zero ;
 wire \top_I.branch[17].block[3].um_I.pg_vdd ;
 wire \top_I.branch[17].block[4].um_I.ana[0] ;
 wire \top_I.branch[17].block[4].um_I.ana[1] ;
 wire \top_I.branch[17].block[4].um_I.ana[2] ;
 wire \top_I.branch[17].block[4].um_I.ana[3] ;
 wire \top_I.branch[17].block[4].um_I.ana[4] ;
 wire \top_I.branch[17].block[4].um_I.ana[5] ;
 wire \top_I.branch[17].block[4].um_I.ana[6] ;
 wire \top_I.branch[17].block[4].um_I.ana[7] ;
 wire \top_I.branch[17].block[4].um_I.clk ;
 wire \top_I.branch[17].block[4].um_I.ena ;
 wire \top_I.branch[17].block[4].um_I.iw[10] ;
 wire \top_I.branch[17].block[4].um_I.iw[11] ;
 wire \top_I.branch[17].block[4].um_I.iw[12] ;
 wire \top_I.branch[17].block[4].um_I.iw[13] ;
 wire \top_I.branch[17].block[4].um_I.iw[14] ;
 wire \top_I.branch[17].block[4].um_I.iw[15] ;
 wire \top_I.branch[17].block[4].um_I.iw[16] ;
 wire \top_I.branch[17].block[4].um_I.iw[17] ;
 wire \top_I.branch[17].block[4].um_I.iw[1] ;
 wire \top_I.branch[17].block[4].um_I.iw[2] ;
 wire \top_I.branch[17].block[4].um_I.iw[3] ;
 wire \top_I.branch[17].block[4].um_I.iw[4] ;
 wire \top_I.branch[17].block[4].um_I.iw[5] ;
 wire \top_I.branch[17].block[4].um_I.iw[6] ;
 wire \top_I.branch[17].block[4].um_I.iw[7] ;
 wire \top_I.branch[17].block[4].um_I.iw[8] ;
 wire \top_I.branch[17].block[4].um_I.iw[9] ;
 wire \top_I.branch[17].block[4].um_I.k_zero ;
 wire \top_I.branch[17].block[4].um_I.pg_vdd ;
 wire \top_I.branch[17].block[5].um_I.ana[0] ;
 wire \top_I.branch[17].block[5].um_I.ana[1] ;
 wire \top_I.branch[17].block[5].um_I.ana[2] ;
 wire \top_I.branch[17].block[5].um_I.ana[3] ;
 wire \top_I.branch[17].block[5].um_I.ana[4] ;
 wire \top_I.branch[17].block[5].um_I.ana[5] ;
 wire \top_I.branch[17].block[5].um_I.ana[6] ;
 wire \top_I.branch[17].block[5].um_I.ana[7] ;
 wire \top_I.branch[17].block[5].um_I.clk ;
 wire \top_I.branch[17].block[5].um_I.ena ;
 wire \top_I.branch[17].block[5].um_I.iw[10] ;
 wire \top_I.branch[17].block[5].um_I.iw[11] ;
 wire \top_I.branch[17].block[5].um_I.iw[12] ;
 wire \top_I.branch[17].block[5].um_I.iw[13] ;
 wire \top_I.branch[17].block[5].um_I.iw[14] ;
 wire \top_I.branch[17].block[5].um_I.iw[15] ;
 wire \top_I.branch[17].block[5].um_I.iw[16] ;
 wire \top_I.branch[17].block[5].um_I.iw[17] ;
 wire \top_I.branch[17].block[5].um_I.iw[1] ;
 wire \top_I.branch[17].block[5].um_I.iw[2] ;
 wire \top_I.branch[17].block[5].um_I.iw[3] ;
 wire \top_I.branch[17].block[5].um_I.iw[4] ;
 wire \top_I.branch[17].block[5].um_I.iw[5] ;
 wire \top_I.branch[17].block[5].um_I.iw[6] ;
 wire \top_I.branch[17].block[5].um_I.iw[7] ;
 wire \top_I.branch[17].block[5].um_I.iw[8] ;
 wire \top_I.branch[17].block[5].um_I.iw[9] ;
 wire \top_I.branch[17].block[5].um_I.k_zero ;
 wire \top_I.branch[17].block[5].um_I.pg_vdd ;
 wire \top_I.branch[17].block[6].um_I.ana[0] ;
 wire \top_I.branch[17].block[6].um_I.ana[1] ;
 wire \top_I.branch[17].block[6].um_I.ana[2] ;
 wire \top_I.branch[17].block[6].um_I.ana[3] ;
 wire \top_I.branch[17].block[6].um_I.ana[4] ;
 wire \top_I.branch[17].block[6].um_I.ana[5] ;
 wire \top_I.branch[17].block[6].um_I.ana[6] ;
 wire \top_I.branch[17].block[6].um_I.ana[7] ;
 wire \top_I.branch[17].block[6].um_I.clk ;
 wire \top_I.branch[17].block[6].um_I.ena ;
 wire \top_I.branch[17].block[6].um_I.iw[10] ;
 wire \top_I.branch[17].block[6].um_I.iw[11] ;
 wire \top_I.branch[17].block[6].um_I.iw[12] ;
 wire \top_I.branch[17].block[6].um_I.iw[13] ;
 wire \top_I.branch[17].block[6].um_I.iw[14] ;
 wire \top_I.branch[17].block[6].um_I.iw[15] ;
 wire \top_I.branch[17].block[6].um_I.iw[16] ;
 wire \top_I.branch[17].block[6].um_I.iw[17] ;
 wire \top_I.branch[17].block[6].um_I.iw[1] ;
 wire \top_I.branch[17].block[6].um_I.iw[2] ;
 wire \top_I.branch[17].block[6].um_I.iw[3] ;
 wire \top_I.branch[17].block[6].um_I.iw[4] ;
 wire \top_I.branch[17].block[6].um_I.iw[5] ;
 wire \top_I.branch[17].block[6].um_I.iw[6] ;
 wire \top_I.branch[17].block[6].um_I.iw[7] ;
 wire \top_I.branch[17].block[6].um_I.iw[8] ;
 wire \top_I.branch[17].block[6].um_I.iw[9] ;
 wire \top_I.branch[17].block[6].um_I.k_zero ;
 wire \top_I.branch[17].block[6].um_I.pg_vdd ;
 wire \top_I.branch[17].block[7].um_I.ana[0] ;
 wire \top_I.branch[17].block[7].um_I.ana[1] ;
 wire \top_I.branch[17].block[7].um_I.ana[2] ;
 wire \top_I.branch[17].block[7].um_I.ana[3] ;
 wire \top_I.branch[17].block[7].um_I.ana[4] ;
 wire \top_I.branch[17].block[7].um_I.ana[5] ;
 wire \top_I.branch[17].block[7].um_I.ana[6] ;
 wire \top_I.branch[17].block[7].um_I.ana[7] ;
 wire \top_I.branch[17].block[7].um_I.clk ;
 wire \top_I.branch[17].block[7].um_I.ena ;
 wire \top_I.branch[17].block[7].um_I.iw[10] ;
 wire \top_I.branch[17].block[7].um_I.iw[11] ;
 wire \top_I.branch[17].block[7].um_I.iw[12] ;
 wire \top_I.branch[17].block[7].um_I.iw[13] ;
 wire \top_I.branch[17].block[7].um_I.iw[14] ;
 wire \top_I.branch[17].block[7].um_I.iw[15] ;
 wire \top_I.branch[17].block[7].um_I.iw[16] ;
 wire \top_I.branch[17].block[7].um_I.iw[17] ;
 wire \top_I.branch[17].block[7].um_I.iw[1] ;
 wire \top_I.branch[17].block[7].um_I.iw[2] ;
 wire \top_I.branch[17].block[7].um_I.iw[3] ;
 wire \top_I.branch[17].block[7].um_I.iw[4] ;
 wire \top_I.branch[17].block[7].um_I.iw[5] ;
 wire \top_I.branch[17].block[7].um_I.iw[6] ;
 wire \top_I.branch[17].block[7].um_I.iw[7] ;
 wire \top_I.branch[17].block[7].um_I.iw[8] ;
 wire \top_I.branch[17].block[7].um_I.iw[9] ;
 wire \top_I.branch[17].block[7].um_I.k_zero ;
 wire \top_I.branch[17].block[7].um_I.pg_vdd ;
 wire \top_I.branch[17].block[8].um_I.ana[0] ;
 wire \top_I.branch[17].block[8].um_I.ana[1] ;
 wire \top_I.branch[17].block[8].um_I.ana[2] ;
 wire \top_I.branch[17].block[8].um_I.ana[3] ;
 wire \top_I.branch[17].block[8].um_I.ana[4] ;
 wire \top_I.branch[17].block[8].um_I.ana[5] ;
 wire \top_I.branch[17].block[8].um_I.ana[6] ;
 wire \top_I.branch[17].block[8].um_I.ana[7] ;
 wire \top_I.branch[17].block[8].um_I.clk ;
 wire \top_I.branch[17].block[8].um_I.ena ;
 wire \top_I.branch[17].block[8].um_I.iw[10] ;
 wire \top_I.branch[17].block[8].um_I.iw[11] ;
 wire \top_I.branch[17].block[8].um_I.iw[12] ;
 wire \top_I.branch[17].block[8].um_I.iw[13] ;
 wire \top_I.branch[17].block[8].um_I.iw[14] ;
 wire \top_I.branch[17].block[8].um_I.iw[15] ;
 wire \top_I.branch[17].block[8].um_I.iw[16] ;
 wire \top_I.branch[17].block[8].um_I.iw[17] ;
 wire \top_I.branch[17].block[8].um_I.iw[1] ;
 wire \top_I.branch[17].block[8].um_I.iw[2] ;
 wire \top_I.branch[17].block[8].um_I.iw[3] ;
 wire \top_I.branch[17].block[8].um_I.iw[4] ;
 wire \top_I.branch[17].block[8].um_I.iw[5] ;
 wire \top_I.branch[17].block[8].um_I.iw[6] ;
 wire \top_I.branch[17].block[8].um_I.iw[7] ;
 wire \top_I.branch[17].block[8].um_I.iw[8] ;
 wire \top_I.branch[17].block[8].um_I.iw[9] ;
 wire \top_I.branch[17].block[8].um_I.k_zero ;
 wire \top_I.branch[17].block[8].um_I.pg_vdd ;
 wire \top_I.branch[17].block[9].um_I.ana[0] ;
 wire \top_I.branch[17].block[9].um_I.ana[1] ;
 wire \top_I.branch[17].block[9].um_I.ana[2] ;
 wire \top_I.branch[17].block[9].um_I.ana[3] ;
 wire \top_I.branch[17].block[9].um_I.ana[4] ;
 wire \top_I.branch[17].block[9].um_I.ana[5] ;
 wire \top_I.branch[17].block[9].um_I.ana[6] ;
 wire \top_I.branch[17].block[9].um_I.ana[7] ;
 wire \top_I.branch[17].block[9].um_I.clk ;
 wire \top_I.branch[17].block[9].um_I.ena ;
 wire \top_I.branch[17].block[9].um_I.iw[10] ;
 wire \top_I.branch[17].block[9].um_I.iw[11] ;
 wire \top_I.branch[17].block[9].um_I.iw[12] ;
 wire \top_I.branch[17].block[9].um_I.iw[13] ;
 wire \top_I.branch[17].block[9].um_I.iw[14] ;
 wire \top_I.branch[17].block[9].um_I.iw[15] ;
 wire \top_I.branch[17].block[9].um_I.iw[16] ;
 wire \top_I.branch[17].block[9].um_I.iw[17] ;
 wire \top_I.branch[17].block[9].um_I.iw[1] ;
 wire \top_I.branch[17].block[9].um_I.iw[2] ;
 wire \top_I.branch[17].block[9].um_I.iw[3] ;
 wire \top_I.branch[17].block[9].um_I.iw[4] ;
 wire \top_I.branch[17].block[9].um_I.iw[5] ;
 wire \top_I.branch[17].block[9].um_I.iw[6] ;
 wire \top_I.branch[17].block[9].um_I.iw[7] ;
 wire \top_I.branch[17].block[9].um_I.iw[8] ;
 wire \top_I.branch[17].block[9].um_I.iw[9] ;
 wire \top_I.branch[17].block[9].um_I.k_zero ;
 wire \top_I.branch[17].block[9].um_I.pg_vdd ;
 wire \top_I.branch[17].l_addr[0] ;
 wire \top_I.branch[17].l_addr[3] ;
 wire \top_I.branch[18].block[0].um_I.ana[0] ;
 wire \top_I.branch[18].block[0].um_I.ana[1] ;
 wire \top_I.branch[18].block[0].um_I.ana[2] ;
 wire \top_I.branch[18].block[0].um_I.ana[3] ;
 wire \top_I.branch[18].block[0].um_I.ana[4] ;
 wire \top_I.branch[18].block[0].um_I.ana[5] ;
 wire \top_I.branch[18].block[0].um_I.ana[6] ;
 wire \top_I.branch[18].block[0].um_I.ana[7] ;
 wire \top_I.branch[18].block[0].um_I.clk ;
 wire \top_I.branch[18].block[0].um_I.ena ;
 wire \top_I.branch[18].block[0].um_I.iw[10] ;
 wire \top_I.branch[18].block[0].um_I.iw[11] ;
 wire \top_I.branch[18].block[0].um_I.iw[12] ;
 wire \top_I.branch[18].block[0].um_I.iw[13] ;
 wire \top_I.branch[18].block[0].um_I.iw[14] ;
 wire \top_I.branch[18].block[0].um_I.iw[15] ;
 wire \top_I.branch[18].block[0].um_I.iw[16] ;
 wire \top_I.branch[18].block[0].um_I.iw[17] ;
 wire \top_I.branch[18].block[0].um_I.iw[1] ;
 wire \top_I.branch[18].block[0].um_I.iw[2] ;
 wire \top_I.branch[18].block[0].um_I.iw[3] ;
 wire \top_I.branch[18].block[0].um_I.iw[4] ;
 wire \top_I.branch[18].block[0].um_I.iw[5] ;
 wire \top_I.branch[18].block[0].um_I.iw[6] ;
 wire \top_I.branch[18].block[0].um_I.iw[7] ;
 wire \top_I.branch[18].block[0].um_I.iw[8] ;
 wire \top_I.branch[18].block[0].um_I.iw[9] ;
 wire \top_I.branch[18].block[0].um_I.k_zero ;
 wire \top_I.branch[18].block[0].um_I.pg_vdd ;
 wire \top_I.branch[18].block[10].um_I.ana[0] ;
 wire \top_I.branch[18].block[10].um_I.ana[1] ;
 wire \top_I.branch[18].block[10].um_I.ana[2] ;
 wire \top_I.branch[18].block[10].um_I.ana[3] ;
 wire \top_I.branch[18].block[10].um_I.ana[4] ;
 wire \top_I.branch[18].block[10].um_I.ana[5] ;
 wire \top_I.branch[18].block[10].um_I.ana[6] ;
 wire \top_I.branch[18].block[10].um_I.ana[7] ;
 wire \top_I.branch[18].block[10].um_I.clk ;
 wire \top_I.branch[18].block[10].um_I.ena ;
 wire \top_I.branch[18].block[10].um_I.iw[10] ;
 wire \top_I.branch[18].block[10].um_I.iw[11] ;
 wire \top_I.branch[18].block[10].um_I.iw[12] ;
 wire \top_I.branch[18].block[10].um_I.iw[13] ;
 wire \top_I.branch[18].block[10].um_I.iw[14] ;
 wire \top_I.branch[18].block[10].um_I.iw[15] ;
 wire \top_I.branch[18].block[10].um_I.iw[16] ;
 wire \top_I.branch[18].block[10].um_I.iw[17] ;
 wire \top_I.branch[18].block[10].um_I.iw[1] ;
 wire \top_I.branch[18].block[10].um_I.iw[2] ;
 wire \top_I.branch[18].block[10].um_I.iw[3] ;
 wire \top_I.branch[18].block[10].um_I.iw[4] ;
 wire \top_I.branch[18].block[10].um_I.iw[5] ;
 wire \top_I.branch[18].block[10].um_I.iw[6] ;
 wire \top_I.branch[18].block[10].um_I.iw[7] ;
 wire \top_I.branch[18].block[10].um_I.iw[8] ;
 wire \top_I.branch[18].block[10].um_I.iw[9] ;
 wire \top_I.branch[18].block[10].um_I.k_zero ;
 wire \top_I.branch[18].block[10].um_I.pg_vdd ;
 wire \top_I.branch[18].block[11].um_I.ana[0] ;
 wire \top_I.branch[18].block[11].um_I.ana[1] ;
 wire \top_I.branch[18].block[11].um_I.ana[2] ;
 wire \top_I.branch[18].block[11].um_I.ana[3] ;
 wire \top_I.branch[18].block[11].um_I.ana[4] ;
 wire \top_I.branch[18].block[11].um_I.ana[5] ;
 wire \top_I.branch[18].block[11].um_I.ana[6] ;
 wire \top_I.branch[18].block[11].um_I.ana[7] ;
 wire \top_I.branch[18].block[11].um_I.clk ;
 wire \top_I.branch[18].block[11].um_I.ena ;
 wire \top_I.branch[18].block[11].um_I.iw[10] ;
 wire \top_I.branch[18].block[11].um_I.iw[11] ;
 wire \top_I.branch[18].block[11].um_I.iw[12] ;
 wire \top_I.branch[18].block[11].um_I.iw[13] ;
 wire \top_I.branch[18].block[11].um_I.iw[14] ;
 wire \top_I.branch[18].block[11].um_I.iw[15] ;
 wire \top_I.branch[18].block[11].um_I.iw[16] ;
 wire \top_I.branch[18].block[11].um_I.iw[17] ;
 wire \top_I.branch[18].block[11].um_I.iw[1] ;
 wire \top_I.branch[18].block[11].um_I.iw[2] ;
 wire \top_I.branch[18].block[11].um_I.iw[3] ;
 wire \top_I.branch[18].block[11].um_I.iw[4] ;
 wire \top_I.branch[18].block[11].um_I.iw[5] ;
 wire \top_I.branch[18].block[11].um_I.iw[6] ;
 wire \top_I.branch[18].block[11].um_I.iw[7] ;
 wire \top_I.branch[18].block[11].um_I.iw[8] ;
 wire \top_I.branch[18].block[11].um_I.iw[9] ;
 wire \top_I.branch[18].block[11].um_I.k_zero ;
 wire \top_I.branch[18].block[11].um_I.pg_vdd ;
 wire \top_I.branch[18].block[12].um_I.ana[0] ;
 wire \top_I.branch[18].block[12].um_I.ana[1] ;
 wire \top_I.branch[18].block[12].um_I.ana[2] ;
 wire \top_I.branch[18].block[12].um_I.ana[3] ;
 wire \top_I.branch[18].block[12].um_I.ana[4] ;
 wire \top_I.branch[18].block[12].um_I.ana[5] ;
 wire \top_I.branch[18].block[12].um_I.ana[6] ;
 wire \top_I.branch[18].block[12].um_I.ana[7] ;
 wire \top_I.branch[18].block[12].um_I.clk ;
 wire \top_I.branch[18].block[12].um_I.ena ;
 wire \top_I.branch[18].block[12].um_I.iw[10] ;
 wire \top_I.branch[18].block[12].um_I.iw[11] ;
 wire \top_I.branch[18].block[12].um_I.iw[12] ;
 wire \top_I.branch[18].block[12].um_I.iw[13] ;
 wire \top_I.branch[18].block[12].um_I.iw[14] ;
 wire \top_I.branch[18].block[12].um_I.iw[15] ;
 wire \top_I.branch[18].block[12].um_I.iw[16] ;
 wire \top_I.branch[18].block[12].um_I.iw[17] ;
 wire \top_I.branch[18].block[12].um_I.iw[1] ;
 wire \top_I.branch[18].block[12].um_I.iw[2] ;
 wire \top_I.branch[18].block[12].um_I.iw[3] ;
 wire \top_I.branch[18].block[12].um_I.iw[4] ;
 wire \top_I.branch[18].block[12].um_I.iw[5] ;
 wire \top_I.branch[18].block[12].um_I.iw[6] ;
 wire \top_I.branch[18].block[12].um_I.iw[7] ;
 wire \top_I.branch[18].block[12].um_I.iw[8] ;
 wire \top_I.branch[18].block[12].um_I.iw[9] ;
 wire \top_I.branch[18].block[12].um_I.k_zero ;
 wire \top_I.branch[18].block[12].um_I.pg_vdd ;
 wire \top_I.branch[18].block[13].um_I.ana[0] ;
 wire \top_I.branch[18].block[13].um_I.ana[1] ;
 wire \top_I.branch[18].block[13].um_I.ana[2] ;
 wire \top_I.branch[18].block[13].um_I.ana[3] ;
 wire \top_I.branch[18].block[13].um_I.ana[4] ;
 wire \top_I.branch[18].block[13].um_I.ana[5] ;
 wire \top_I.branch[18].block[13].um_I.ana[6] ;
 wire \top_I.branch[18].block[13].um_I.ana[7] ;
 wire \top_I.branch[18].block[13].um_I.clk ;
 wire \top_I.branch[18].block[13].um_I.ena ;
 wire \top_I.branch[18].block[13].um_I.iw[10] ;
 wire \top_I.branch[18].block[13].um_I.iw[11] ;
 wire \top_I.branch[18].block[13].um_I.iw[12] ;
 wire \top_I.branch[18].block[13].um_I.iw[13] ;
 wire \top_I.branch[18].block[13].um_I.iw[14] ;
 wire \top_I.branch[18].block[13].um_I.iw[15] ;
 wire \top_I.branch[18].block[13].um_I.iw[16] ;
 wire \top_I.branch[18].block[13].um_I.iw[17] ;
 wire \top_I.branch[18].block[13].um_I.iw[1] ;
 wire \top_I.branch[18].block[13].um_I.iw[2] ;
 wire \top_I.branch[18].block[13].um_I.iw[3] ;
 wire \top_I.branch[18].block[13].um_I.iw[4] ;
 wire \top_I.branch[18].block[13].um_I.iw[5] ;
 wire \top_I.branch[18].block[13].um_I.iw[6] ;
 wire \top_I.branch[18].block[13].um_I.iw[7] ;
 wire \top_I.branch[18].block[13].um_I.iw[8] ;
 wire \top_I.branch[18].block[13].um_I.iw[9] ;
 wire \top_I.branch[18].block[13].um_I.k_zero ;
 wire \top_I.branch[18].block[13].um_I.pg_vdd ;
 wire \top_I.branch[18].block[14].um_I.ana[0] ;
 wire \top_I.branch[18].block[14].um_I.ana[1] ;
 wire \top_I.branch[18].block[14].um_I.ana[2] ;
 wire \top_I.branch[18].block[14].um_I.ana[3] ;
 wire \top_I.branch[18].block[14].um_I.ana[4] ;
 wire \top_I.branch[18].block[14].um_I.ana[5] ;
 wire \top_I.branch[18].block[14].um_I.ana[6] ;
 wire \top_I.branch[18].block[14].um_I.ana[7] ;
 wire \top_I.branch[18].block[14].um_I.clk ;
 wire \top_I.branch[18].block[14].um_I.ena ;
 wire \top_I.branch[18].block[14].um_I.iw[10] ;
 wire \top_I.branch[18].block[14].um_I.iw[11] ;
 wire \top_I.branch[18].block[14].um_I.iw[12] ;
 wire \top_I.branch[18].block[14].um_I.iw[13] ;
 wire \top_I.branch[18].block[14].um_I.iw[14] ;
 wire \top_I.branch[18].block[14].um_I.iw[15] ;
 wire \top_I.branch[18].block[14].um_I.iw[16] ;
 wire \top_I.branch[18].block[14].um_I.iw[17] ;
 wire \top_I.branch[18].block[14].um_I.iw[1] ;
 wire \top_I.branch[18].block[14].um_I.iw[2] ;
 wire \top_I.branch[18].block[14].um_I.iw[3] ;
 wire \top_I.branch[18].block[14].um_I.iw[4] ;
 wire \top_I.branch[18].block[14].um_I.iw[5] ;
 wire \top_I.branch[18].block[14].um_I.iw[6] ;
 wire \top_I.branch[18].block[14].um_I.iw[7] ;
 wire \top_I.branch[18].block[14].um_I.iw[8] ;
 wire \top_I.branch[18].block[14].um_I.iw[9] ;
 wire \top_I.branch[18].block[14].um_I.k_zero ;
 wire \top_I.branch[18].block[14].um_I.pg_vdd ;
 wire \top_I.branch[18].block[15].um_I.ana[0] ;
 wire \top_I.branch[18].block[15].um_I.ana[1] ;
 wire \top_I.branch[18].block[15].um_I.ana[2] ;
 wire \top_I.branch[18].block[15].um_I.ana[3] ;
 wire \top_I.branch[18].block[15].um_I.ana[4] ;
 wire \top_I.branch[18].block[15].um_I.ana[5] ;
 wire \top_I.branch[18].block[15].um_I.ana[6] ;
 wire \top_I.branch[18].block[15].um_I.ana[7] ;
 wire \top_I.branch[18].block[15].um_I.clk ;
 wire \top_I.branch[18].block[15].um_I.ena ;
 wire \top_I.branch[18].block[15].um_I.iw[10] ;
 wire \top_I.branch[18].block[15].um_I.iw[11] ;
 wire \top_I.branch[18].block[15].um_I.iw[12] ;
 wire \top_I.branch[18].block[15].um_I.iw[13] ;
 wire \top_I.branch[18].block[15].um_I.iw[14] ;
 wire \top_I.branch[18].block[15].um_I.iw[15] ;
 wire \top_I.branch[18].block[15].um_I.iw[16] ;
 wire \top_I.branch[18].block[15].um_I.iw[17] ;
 wire \top_I.branch[18].block[15].um_I.iw[1] ;
 wire \top_I.branch[18].block[15].um_I.iw[2] ;
 wire \top_I.branch[18].block[15].um_I.iw[3] ;
 wire \top_I.branch[18].block[15].um_I.iw[4] ;
 wire \top_I.branch[18].block[15].um_I.iw[5] ;
 wire \top_I.branch[18].block[15].um_I.iw[6] ;
 wire \top_I.branch[18].block[15].um_I.iw[7] ;
 wire \top_I.branch[18].block[15].um_I.iw[8] ;
 wire \top_I.branch[18].block[15].um_I.iw[9] ;
 wire \top_I.branch[18].block[15].um_I.k_zero ;
 wire \top_I.branch[18].block[15].um_I.pg_vdd ;
 wire \top_I.branch[18].block[1].um_I.ana[0] ;
 wire \top_I.branch[18].block[1].um_I.ana[1] ;
 wire \top_I.branch[18].block[1].um_I.ana[2] ;
 wire \top_I.branch[18].block[1].um_I.ana[3] ;
 wire \top_I.branch[18].block[1].um_I.ana[4] ;
 wire \top_I.branch[18].block[1].um_I.ana[5] ;
 wire \top_I.branch[18].block[1].um_I.ana[6] ;
 wire \top_I.branch[18].block[1].um_I.ana[7] ;
 wire \top_I.branch[18].block[1].um_I.clk ;
 wire \top_I.branch[18].block[1].um_I.ena ;
 wire \top_I.branch[18].block[1].um_I.iw[10] ;
 wire \top_I.branch[18].block[1].um_I.iw[11] ;
 wire \top_I.branch[18].block[1].um_I.iw[12] ;
 wire \top_I.branch[18].block[1].um_I.iw[13] ;
 wire \top_I.branch[18].block[1].um_I.iw[14] ;
 wire \top_I.branch[18].block[1].um_I.iw[15] ;
 wire \top_I.branch[18].block[1].um_I.iw[16] ;
 wire \top_I.branch[18].block[1].um_I.iw[17] ;
 wire \top_I.branch[18].block[1].um_I.iw[1] ;
 wire \top_I.branch[18].block[1].um_I.iw[2] ;
 wire \top_I.branch[18].block[1].um_I.iw[3] ;
 wire \top_I.branch[18].block[1].um_I.iw[4] ;
 wire \top_I.branch[18].block[1].um_I.iw[5] ;
 wire \top_I.branch[18].block[1].um_I.iw[6] ;
 wire \top_I.branch[18].block[1].um_I.iw[7] ;
 wire \top_I.branch[18].block[1].um_I.iw[8] ;
 wire \top_I.branch[18].block[1].um_I.iw[9] ;
 wire \top_I.branch[18].block[1].um_I.k_zero ;
 wire \top_I.branch[18].block[1].um_I.pg_vdd ;
 wire \top_I.branch[18].block[2].um_I.ana[0] ;
 wire \top_I.branch[18].block[2].um_I.ana[1] ;
 wire \top_I.branch[18].block[2].um_I.ana[2] ;
 wire \top_I.branch[18].block[2].um_I.ana[3] ;
 wire \top_I.branch[18].block[2].um_I.ana[4] ;
 wire \top_I.branch[18].block[2].um_I.ana[5] ;
 wire \top_I.branch[18].block[2].um_I.ana[6] ;
 wire \top_I.branch[18].block[2].um_I.ana[7] ;
 wire \top_I.branch[18].block[2].um_I.clk ;
 wire \top_I.branch[18].block[2].um_I.ena ;
 wire \top_I.branch[18].block[2].um_I.iw[10] ;
 wire \top_I.branch[18].block[2].um_I.iw[11] ;
 wire \top_I.branch[18].block[2].um_I.iw[12] ;
 wire \top_I.branch[18].block[2].um_I.iw[13] ;
 wire \top_I.branch[18].block[2].um_I.iw[14] ;
 wire \top_I.branch[18].block[2].um_I.iw[15] ;
 wire \top_I.branch[18].block[2].um_I.iw[16] ;
 wire \top_I.branch[18].block[2].um_I.iw[17] ;
 wire \top_I.branch[18].block[2].um_I.iw[1] ;
 wire \top_I.branch[18].block[2].um_I.iw[2] ;
 wire \top_I.branch[18].block[2].um_I.iw[3] ;
 wire \top_I.branch[18].block[2].um_I.iw[4] ;
 wire \top_I.branch[18].block[2].um_I.iw[5] ;
 wire \top_I.branch[18].block[2].um_I.iw[6] ;
 wire \top_I.branch[18].block[2].um_I.iw[7] ;
 wire \top_I.branch[18].block[2].um_I.iw[8] ;
 wire \top_I.branch[18].block[2].um_I.iw[9] ;
 wire \top_I.branch[18].block[2].um_I.k_zero ;
 wire \top_I.branch[18].block[2].um_I.pg_vdd ;
 wire \top_I.branch[18].block[3].um_I.ana[0] ;
 wire \top_I.branch[18].block[3].um_I.ana[1] ;
 wire \top_I.branch[18].block[3].um_I.ana[2] ;
 wire \top_I.branch[18].block[3].um_I.ana[3] ;
 wire \top_I.branch[18].block[3].um_I.ana[4] ;
 wire \top_I.branch[18].block[3].um_I.ana[5] ;
 wire \top_I.branch[18].block[3].um_I.ana[6] ;
 wire \top_I.branch[18].block[3].um_I.ana[7] ;
 wire \top_I.branch[18].block[3].um_I.clk ;
 wire \top_I.branch[18].block[3].um_I.ena ;
 wire \top_I.branch[18].block[3].um_I.iw[10] ;
 wire \top_I.branch[18].block[3].um_I.iw[11] ;
 wire \top_I.branch[18].block[3].um_I.iw[12] ;
 wire \top_I.branch[18].block[3].um_I.iw[13] ;
 wire \top_I.branch[18].block[3].um_I.iw[14] ;
 wire \top_I.branch[18].block[3].um_I.iw[15] ;
 wire \top_I.branch[18].block[3].um_I.iw[16] ;
 wire \top_I.branch[18].block[3].um_I.iw[17] ;
 wire \top_I.branch[18].block[3].um_I.iw[1] ;
 wire \top_I.branch[18].block[3].um_I.iw[2] ;
 wire \top_I.branch[18].block[3].um_I.iw[3] ;
 wire \top_I.branch[18].block[3].um_I.iw[4] ;
 wire \top_I.branch[18].block[3].um_I.iw[5] ;
 wire \top_I.branch[18].block[3].um_I.iw[6] ;
 wire \top_I.branch[18].block[3].um_I.iw[7] ;
 wire \top_I.branch[18].block[3].um_I.iw[8] ;
 wire \top_I.branch[18].block[3].um_I.iw[9] ;
 wire \top_I.branch[18].block[3].um_I.k_zero ;
 wire \top_I.branch[18].block[3].um_I.pg_vdd ;
 wire \top_I.branch[18].block[4].um_I.ana[0] ;
 wire \top_I.branch[18].block[4].um_I.ana[1] ;
 wire \top_I.branch[18].block[4].um_I.ana[2] ;
 wire \top_I.branch[18].block[4].um_I.ana[3] ;
 wire \top_I.branch[18].block[4].um_I.ana[4] ;
 wire \top_I.branch[18].block[4].um_I.ana[5] ;
 wire \top_I.branch[18].block[4].um_I.ana[6] ;
 wire \top_I.branch[18].block[4].um_I.ana[7] ;
 wire \top_I.branch[18].block[4].um_I.clk ;
 wire \top_I.branch[18].block[4].um_I.ena ;
 wire \top_I.branch[18].block[4].um_I.iw[10] ;
 wire \top_I.branch[18].block[4].um_I.iw[11] ;
 wire \top_I.branch[18].block[4].um_I.iw[12] ;
 wire \top_I.branch[18].block[4].um_I.iw[13] ;
 wire \top_I.branch[18].block[4].um_I.iw[14] ;
 wire \top_I.branch[18].block[4].um_I.iw[15] ;
 wire \top_I.branch[18].block[4].um_I.iw[16] ;
 wire \top_I.branch[18].block[4].um_I.iw[17] ;
 wire \top_I.branch[18].block[4].um_I.iw[1] ;
 wire \top_I.branch[18].block[4].um_I.iw[2] ;
 wire \top_I.branch[18].block[4].um_I.iw[3] ;
 wire \top_I.branch[18].block[4].um_I.iw[4] ;
 wire \top_I.branch[18].block[4].um_I.iw[5] ;
 wire \top_I.branch[18].block[4].um_I.iw[6] ;
 wire \top_I.branch[18].block[4].um_I.iw[7] ;
 wire \top_I.branch[18].block[4].um_I.iw[8] ;
 wire \top_I.branch[18].block[4].um_I.iw[9] ;
 wire \top_I.branch[18].block[4].um_I.k_zero ;
 wire \top_I.branch[18].block[4].um_I.pg_vdd ;
 wire \top_I.branch[18].block[5].um_I.ana[0] ;
 wire \top_I.branch[18].block[5].um_I.ana[1] ;
 wire \top_I.branch[18].block[5].um_I.ana[2] ;
 wire \top_I.branch[18].block[5].um_I.ana[3] ;
 wire \top_I.branch[18].block[5].um_I.ana[4] ;
 wire \top_I.branch[18].block[5].um_I.ana[5] ;
 wire \top_I.branch[18].block[5].um_I.ana[6] ;
 wire \top_I.branch[18].block[5].um_I.ana[7] ;
 wire \top_I.branch[18].block[5].um_I.clk ;
 wire \top_I.branch[18].block[5].um_I.ena ;
 wire \top_I.branch[18].block[5].um_I.iw[10] ;
 wire \top_I.branch[18].block[5].um_I.iw[11] ;
 wire \top_I.branch[18].block[5].um_I.iw[12] ;
 wire \top_I.branch[18].block[5].um_I.iw[13] ;
 wire \top_I.branch[18].block[5].um_I.iw[14] ;
 wire \top_I.branch[18].block[5].um_I.iw[15] ;
 wire \top_I.branch[18].block[5].um_I.iw[16] ;
 wire \top_I.branch[18].block[5].um_I.iw[17] ;
 wire \top_I.branch[18].block[5].um_I.iw[1] ;
 wire \top_I.branch[18].block[5].um_I.iw[2] ;
 wire \top_I.branch[18].block[5].um_I.iw[3] ;
 wire \top_I.branch[18].block[5].um_I.iw[4] ;
 wire \top_I.branch[18].block[5].um_I.iw[5] ;
 wire \top_I.branch[18].block[5].um_I.iw[6] ;
 wire \top_I.branch[18].block[5].um_I.iw[7] ;
 wire \top_I.branch[18].block[5].um_I.iw[8] ;
 wire \top_I.branch[18].block[5].um_I.iw[9] ;
 wire \top_I.branch[18].block[5].um_I.k_zero ;
 wire \top_I.branch[18].block[5].um_I.pg_vdd ;
 wire \top_I.branch[18].block[6].um_I.ana[0] ;
 wire \top_I.branch[18].block[6].um_I.ana[1] ;
 wire \top_I.branch[18].block[6].um_I.ana[2] ;
 wire \top_I.branch[18].block[6].um_I.ana[3] ;
 wire \top_I.branch[18].block[6].um_I.ana[4] ;
 wire \top_I.branch[18].block[6].um_I.ana[5] ;
 wire \top_I.branch[18].block[6].um_I.ana[6] ;
 wire \top_I.branch[18].block[6].um_I.ana[7] ;
 wire \top_I.branch[18].block[6].um_I.clk ;
 wire \top_I.branch[18].block[6].um_I.ena ;
 wire \top_I.branch[18].block[6].um_I.iw[10] ;
 wire \top_I.branch[18].block[6].um_I.iw[11] ;
 wire \top_I.branch[18].block[6].um_I.iw[12] ;
 wire \top_I.branch[18].block[6].um_I.iw[13] ;
 wire \top_I.branch[18].block[6].um_I.iw[14] ;
 wire \top_I.branch[18].block[6].um_I.iw[15] ;
 wire \top_I.branch[18].block[6].um_I.iw[16] ;
 wire \top_I.branch[18].block[6].um_I.iw[17] ;
 wire \top_I.branch[18].block[6].um_I.iw[1] ;
 wire \top_I.branch[18].block[6].um_I.iw[2] ;
 wire \top_I.branch[18].block[6].um_I.iw[3] ;
 wire \top_I.branch[18].block[6].um_I.iw[4] ;
 wire \top_I.branch[18].block[6].um_I.iw[5] ;
 wire \top_I.branch[18].block[6].um_I.iw[6] ;
 wire \top_I.branch[18].block[6].um_I.iw[7] ;
 wire \top_I.branch[18].block[6].um_I.iw[8] ;
 wire \top_I.branch[18].block[6].um_I.iw[9] ;
 wire \top_I.branch[18].block[6].um_I.k_zero ;
 wire \top_I.branch[18].block[6].um_I.pg_vdd ;
 wire \top_I.branch[18].block[7].um_I.ana[0] ;
 wire \top_I.branch[18].block[7].um_I.ana[1] ;
 wire \top_I.branch[18].block[7].um_I.ana[2] ;
 wire \top_I.branch[18].block[7].um_I.ana[3] ;
 wire \top_I.branch[18].block[7].um_I.ana[4] ;
 wire \top_I.branch[18].block[7].um_I.ana[5] ;
 wire \top_I.branch[18].block[7].um_I.ana[6] ;
 wire \top_I.branch[18].block[7].um_I.ana[7] ;
 wire \top_I.branch[18].block[7].um_I.clk ;
 wire \top_I.branch[18].block[7].um_I.ena ;
 wire \top_I.branch[18].block[7].um_I.iw[10] ;
 wire \top_I.branch[18].block[7].um_I.iw[11] ;
 wire \top_I.branch[18].block[7].um_I.iw[12] ;
 wire \top_I.branch[18].block[7].um_I.iw[13] ;
 wire \top_I.branch[18].block[7].um_I.iw[14] ;
 wire \top_I.branch[18].block[7].um_I.iw[15] ;
 wire \top_I.branch[18].block[7].um_I.iw[16] ;
 wire \top_I.branch[18].block[7].um_I.iw[17] ;
 wire \top_I.branch[18].block[7].um_I.iw[1] ;
 wire \top_I.branch[18].block[7].um_I.iw[2] ;
 wire \top_I.branch[18].block[7].um_I.iw[3] ;
 wire \top_I.branch[18].block[7].um_I.iw[4] ;
 wire \top_I.branch[18].block[7].um_I.iw[5] ;
 wire \top_I.branch[18].block[7].um_I.iw[6] ;
 wire \top_I.branch[18].block[7].um_I.iw[7] ;
 wire \top_I.branch[18].block[7].um_I.iw[8] ;
 wire \top_I.branch[18].block[7].um_I.iw[9] ;
 wire \top_I.branch[18].block[7].um_I.k_zero ;
 wire \top_I.branch[18].block[7].um_I.pg_vdd ;
 wire \top_I.branch[18].block[8].um_I.ana[0] ;
 wire \top_I.branch[18].block[8].um_I.ana[1] ;
 wire \top_I.branch[18].block[8].um_I.ana[2] ;
 wire \top_I.branch[18].block[8].um_I.ana[3] ;
 wire \top_I.branch[18].block[8].um_I.ana[4] ;
 wire \top_I.branch[18].block[8].um_I.ana[5] ;
 wire \top_I.branch[18].block[8].um_I.ana[6] ;
 wire \top_I.branch[18].block[8].um_I.ana[7] ;
 wire \top_I.branch[18].block[8].um_I.clk ;
 wire \top_I.branch[18].block[8].um_I.ena ;
 wire \top_I.branch[18].block[8].um_I.iw[10] ;
 wire \top_I.branch[18].block[8].um_I.iw[11] ;
 wire \top_I.branch[18].block[8].um_I.iw[12] ;
 wire \top_I.branch[18].block[8].um_I.iw[13] ;
 wire \top_I.branch[18].block[8].um_I.iw[14] ;
 wire \top_I.branch[18].block[8].um_I.iw[15] ;
 wire \top_I.branch[18].block[8].um_I.iw[16] ;
 wire \top_I.branch[18].block[8].um_I.iw[17] ;
 wire \top_I.branch[18].block[8].um_I.iw[1] ;
 wire \top_I.branch[18].block[8].um_I.iw[2] ;
 wire \top_I.branch[18].block[8].um_I.iw[3] ;
 wire \top_I.branch[18].block[8].um_I.iw[4] ;
 wire \top_I.branch[18].block[8].um_I.iw[5] ;
 wire \top_I.branch[18].block[8].um_I.iw[6] ;
 wire \top_I.branch[18].block[8].um_I.iw[7] ;
 wire \top_I.branch[18].block[8].um_I.iw[8] ;
 wire \top_I.branch[18].block[8].um_I.iw[9] ;
 wire \top_I.branch[18].block[8].um_I.k_zero ;
 wire \top_I.branch[18].block[8].um_I.pg_vdd ;
 wire \top_I.branch[18].block[9].um_I.ana[0] ;
 wire \top_I.branch[18].block[9].um_I.ana[1] ;
 wire \top_I.branch[18].block[9].um_I.ana[2] ;
 wire \top_I.branch[18].block[9].um_I.ana[3] ;
 wire \top_I.branch[18].block[9].um_I.ana[4] ;
 wire \top_I.branch[18].block[9].um_I.ana[5] ;
 wire \top_I.branch[18].block[9].um_I.ana[6] ;
 wire \top_I.branch[18].block[9].um_I.ana[7] ;
 wire \top_I.branch[18].block[9].um_I.clk ;
 wire \top_I.branch[18].block[9].um_I.ena ;
 wire \top_I.branch[18].block[9].um_I.iw[10] ;
 wire \top_I.branch[18].block[9].um_I.iw[11] ;
 wire \top_I.branch[18].block[9].um_I.iw[12] ;
 wire \top_I.branch[18].block[9].um_I.iw[13] ;
 wire \top_I.branch[18].block[9].um_I.iw[14] ;
 wire \top_I.branch[18].block[9].um_I.iw[15] ;
 wire \top_I.branch[18].block[9].um_I.iw[16] ;
 wire \top_I.branch[18].block[9].um_I.iw[17] ;
 wire \top_I.branch[18].block[9].um_I.iw[1] ;
 wire \top_I.branch[18].block[9].um_I.iw[2] ;
 wire \top_I.branch[18].block[9].um_I.iw[3] ;
 wire \top_I.branch[18].block[9].um_I.iw[4] ;
 wire \top_I.branch[18].block[9].um_I.iw[5] ;
 wire \top_I.branch[18].block[9].um_I.iw[6] ;
 wire \top_I.branch[18].block[9].um_I.iw[7] ;
 wire \top_I.branch[18].block[9].um_I.iw[8] ;
 wire \top_I.branch[18].block[9].um_I.iw[9] ;
 wire \top_I.branch[18].block[9].um_I.k_zero ;
 wire \top_I.branch[18].block[9].um_I.pg_vdd ;
 wire \top_I.branch[18].l_addr[0] ;
 wire \top_I.branch[18].l_addr[1] ;
 wire \top_I.branch[19].block[0].um_I.ana[0] ;
 wire \top_I.branch[19].block[0].um_I.ana[1] ;
 wire \top_I.branch[19].block[0].um_I.ana[2] ;
 wire \top_I.branch[19].block[0].um_I.ana[3] ;
 wire \top_I.branch[19].block[0].um_I.ana[4] ;
 wire \top_I.branch[19].block[0].um_I.ana[5] ;
 wire \top_I.branch[19].block[0].um_I.ana[6] ;
 wire \top_I.branch[19].block[0].um_I.ana[7] ;
 wire \top_I.branch[19].block[0].um_I.clk ;
 wire \top_I.branch[19].block[0].um_I.ena ;
 wire \top_I.branch[19].block[0].um_I.iw[10] ;
 wire \top_I.branch[19].block[0].um_I.iw[11] ;
 wire \top_I.branch[19].block[0].um_I.iw[12] ;
 wire \top_I.branch[19].block[0].um_I.iw[13] ;
 wire \top_I.branch[19].block[0].um_I.iw[14] ;
 wire \top_I.branch[19].block[0].um_I.iw[15] ;
 wire \top_I.branch[19].block[0].um_I.iw[16] ;
 wire \top_I.branch[19].block[0].um_I.iw[17] ;
 wire \top_I.branch[19].block[0].um_I.iw[1] ;
 wire \top_I.branch[19].block[0].um_I.iw[2] ;
 wire \top_I.branch[19].block[0].um_I.iw[3] ;
 wire \top_I.branch[19].block[0].um_I.iw[4] ;
 wire \top_I.branch[19].block[0].um_I.iw[5] ;
 wire \top_I.branch[19].block[0].um_I.iw[6] ;
 wire \top_I.branch[19].block[0].um_I.iw[7] ;
 wire \top_I.branch[19].block[0].um_I.iw[8] ;
 wire \top_I.branch[19].block[0].um_I.iw[9] ;
 wire \top_I.branch[19].block[0].um_I.k_zero ;
 wire \top_I.branch[19].block[0].um_I.pg_vdd ;
 wire \top_I.branch[19].block[10].um_I.ana[0] ;
 wire \top_I.branch[19].block[10].um_I.ana[1] ;
 wire \top_I.branch[19].block[10].um_I.ana[2] ;
 wire \top_I.branch[19].block[10].um_I.ana[3] ;
 wire \top_I.branch[19].block[10].um_I.ana[4] ;
 wire \top_I.branch[19].block[10].um_I.ana[5] ;
 wire \top_I.branch[19].block[10].um_I.ana[6] ;
 wire \top_I.branch[19].block[10].um_I.ana[7] ;
 wire \top_I.branch[19].block[10].um_I.clk ;
 wire \top_I.branch[19].block[10].um_I.ena ;
 wire \top_I.branch[19].block[10].um_I.iw[10] ;
 wire \top_I.branch[19].block[10].um_I.iw[11] ;
 wire \top_I.branch[19].block[10].um_I.iw[12] ;
 wire \top_I.branch[19].block[10].um_I.iw[13] ;
 wire \top_I.branch[19].block[10].um_I.iw[14] ;
 wire \top_I.branch[19].block[10].um_I.iw[15] ;
 wire \top_I.branch[19].block[10].um_I.iw[16] ;
 wire \top_I.branch[19].block[10].um_I.iw[17] ;
 wire \top_I.branch[19].block[10].um_I.iw[1] ;
 wire \top_I.branch[19].block[10].um_I.iw[2] ;
 wire \top_I.branch[19].block[10].um_I.iw[3] ;
 wire \top_I.branch[19].block[10].um_I.iw[4] ;
 wire \top_I.branch[19].block[10].um_I.iw[5] ;
 wire \top_I.branch[19].block[10].um_I.iw[6] ;
 wire \top_I.branch[19].block[10].um_I.iw[7] ;
 wire \top_I.branch[19].block[10].um_I.iw[8] ;
 wire \top_I.branch[19].block[10].um_I.iw[9] ;
 wire \top_I.branch[19].block[10].um_I.k_zero ;
 wire \top_I.branch[19].block[10].um_I.pg_vdd ;
 wire \top_I.branch[19].block[11].um_I.ana[0] ;
 wire \top_I.branch[19].block[11].um_I.ana[1] ;
 wire \top_I.branch[19].block[11].um_I.ana[2] ;
 wire \top_I.branch[19].block[11].um_I.ana[3] ;
 wire \top_I.branch[19].block[11].um_I.ana[4] ;
 wire \top_I.branch[19].block[11].um_I.ana[5] ;
 wire \top_I.branch[19].block[11].um_I.ana[6] ;
 wire \top_I.branch[19].block[11].um_I.ana[7] ;
 wire \top_I.branch[19].block[11].um_I.clk ;
 wire \top_I.branch[19].block[11].um_I.ena ;
 wire \top_I.branch[19].block[11].um_I.iw[10] ;
 wire \top_I.branch[19].block[11].um_I.iw[11] ;
 wire \top_I.branch[19].block[11].um_I.iw[12] ;
 wire \top_I.branch[19].block[11].um_I.iw[13] ;
 wire \top_I.branch[19].block[11].um_I.iw[14] ;
 wire \top_I.branch[19].block[11].um_I.iw[15] ;
 wire \top_I.branch[19].block[11].um_I.iw[16] ;
 wire \top_I.branch[19].block[11].um_I.iw[17] ;
 wire \top_I.branch[19].block[11].um_I.iw[1] ;
 wire \top_I.branch[19].block[11].um_I.iw[2] ;
 wire \top_I.branch[19].block[11].um_I.iw[3] ;
 wire \top_I.branch[19].block[11].um_I.iw[4] ;
 wire \top_I.branch[19].block[11].um_I.iw[5] ;
 wire \top_I.branch[19].block[11].um_I.iw[6] ;
 wire \top_I.branch[19].block[11].um_I.iw[7] ;
 wire \top_I.branch[19].block[11].um_I.iw[8] ;
 wire \top_I.branch[19].block[11].um_I.iw[9] ;
 wire \top_I.branch[19].block[11].um_I.k_zero ;
 wire \top_I.branch[19].block[11].um_I.pg_vdd ;
 wire \top_I.branch[19].block[12].um_I.ana[0] ;
 wire \top_I.branch[19].block[12].um_I.ana[1] ;
 wire \top_I.branch[19].block[12].um_I.ana[2] ;
 wire \top_I.branch[19].block[12].um_I.ana[3] ;
 wire \top_I.branch[19].block[12].um_I.ana[4] ;
 wire \top_I.branch[19].block[12].um_I.ana[5] ;
 wire \top_I.branch[19].block[12].um_I.ana[6] ;
 wire \top_I.branch[19].block[12].um_I.ana[7] ;
 wire \top_I.branch[19].block[12].um_I.clk ;
 wire \top_I.branch[19].block[12].um_I.ena ;
 wire \top_I.branch[19].block[12].um_I.iw[10] ;
 wire \top_I.branch[19].block[12].um_I.iw[11] ;
 wire \top_I.branch[19].block[12].um_I.iw[12] ;
 wire \top_I.branch[19].block[12].um_I.iw[13] ;
 wire \top_I.branch[19].block[12].um_I.iw[14] ;
 wire \top_I.branch[19].block[12].um_I.iw[15] ;
 wire \top_I.branch[19].block[12].um_I.iw[16] ;
 wire \top_I.branch[19].block[12].um_I.iw[17] ;
 wire \top_I.branch[19].block[12].um_I.iw[1] ;
 wire \top_I.branch[19].block[12].um_I.iw[2] ;
 wire \top_I.branch[19].block[12].um_I.iw[3] ;
 wire \top_I.branch[19].block[12].um_I.iw[4] ;
 wire \top_I.branch[19].block[12].um_I.iw[5] ;
 wire \top_I.branch[19].block[12].um_I.iw[6] ;
 wire \top_I.branch[19].block[12].um_I.iw[7] ;
 wire \top_I.branch[19].block[12].um_I.iw[8] ;
 wire \top_I.branch[19].block[12].um_I.iw[9] ;
 wire \top_I.branch[19].block[12].um_I.k_zero ;
 wire \top_I.branch[19].block[12].um_I.pg_vdd ;
 wire \top_I.branch[19].block[13].um_I.ana[0] ;
 wire \top_I.branch[19].block[13].um_I.ana[1] ;
 wire \top_I.branch[19].block[13].um_I.ana[2] ;
 wire \top_I.branch[19].block[13].um_I.ana[3] ;
 wire \top_I.branch[19].block[13].um_I.ana[4] ;
 wire \top_I.branch[19].block[13].um_I.ana[5] ;
 wire \top_I.branch[19].block[13].um_I.ana[6] ;
 wire \top_I.branch[19].block[13].um_I.ana[7] ;
 wire \top_I.branch[19].block[13].um_I.clk ;
 wire \top_I.branch[19].block[13].um_I.ena ;
 wire \top_I.branch[19].block[13].um_I.iw[10] ;
 wire \top_I.branch[19].block[13].um_I.iw[11] ;
 wire \top_I.branch[19].block[13].um_I.iw[12] ;
 wire \top_I.branch[19].block[13].um_I.iw[13] ;
 wire \top_I.branch[19].block[13].um_I.iw[14] ;
 wire \top_I.branch[19].block[13].um_I.iw[15] ;
 wire \top_I.branch[19].block[13].um_I.iw[16] ;
 wire \top_I.branch[19].block[13].um_I.iw[17] ;
 wire \top_I.branch[19].block[13].um_I.iw[1] ;
 wire \top_I.branch[19].block[13].um_I.iw[2] ;
 wire \top_I.branch[19].block[13].um_I.iw[3] ;
 wire \top_I.branch[19].block[13].um_I.iw[4] ;
 wire \top_I.branch[19].block[13].um_I.iw[5] ;
 wire \top_I.branch[19].block[13].um_I.iw[6] ;
 wire \top_I.branch[19].block[13].um_I.iw[7] ;
 wire \top_I.branch[19].block[13].um_I.iw[8] ;
 wire \top_I.branch[19].block[13].um_I.iw[9] ;
 wire \top_I.branch[19].block[13].um_I.k_zero ;
 wire \top_I.branch[19].block[13].um_I.pg_vdd ;
 wire \top_I.branch[19].block[14].um_I.ana[0] ;
 wire \top_I.branch[19].block[14].um_I.ana[1] ;
 wire \top_I.branch[19].block[14].um_I.ana[2] ;
 wire \top_I.branch[19].block[14].um_I.ana[3] ;
 wire \top_I.branch[19].block[14].um_I.ana[4] ;
 wire \top_I.branch[19].block[14].um_I.ana[5] ;
 wire \top_I.branch[19].block[14].um_I.ana[6] ;
 wire \top_I.branch[19].block[14].um_I.ana[7] ;
 wire \top_I.branch[19].block[14].um_I.clk ;
 wire \top_I.branch[19].block[14].um_I.ena ;
 wire \top_I.branch[19].block[14].um_I.iw[10] ;
 wire \top_I.branch[19].block[14].um_I.iw[11] ;
 wire \top_I.branch[19].block[14].um_I.iw[12] ;
 wire \top_I.branch[19].block[14].um_I.iw[13] ;
 wire \top_I.branch[19].block[14].um_I.iw[14] ;
 wire \top_I.branch[19].block[14].um_I.iw[15] ;
 wire \top_I.branch[19].block[14].um_I.iw[16] ;
 wire \top_I.branch[19].block[14].um_I.iw[17] ;
 wire \top_I.branch[19].block[14].um_I.iw[1] ;
 wire \top_I.branch[19].block[14].um_I.iw[2] ;
 wire \top_I.branch[19].block[14].um_I.iw[3] ;
 wire \top_I.branch[19].block[14].um_I.iw[4] ;
 wire \top_I.branch[19].block[14].um_I.iw[5] ;
 wire \top_I.branch[19].block[14].um_I.iw[6] ;
 wire \top_I.branch[19].block[14].um_I.iw[7] ;
 wire \top_I.branch[19].block[14].um_I.iw[8] ;
 wire \top_I.branch[19].block[14].um_I.iw[9] ;
 wire \top_I.branch[19].block[14].um_I.k_zero ;
 wire \top_I.branch[19].block[14].um_I.pg_vdd ;
 wire \top_I.branch[19].block[15].um_I.ana[0] ;
 wire \top_I.branch[19].block[15].um_I.ana[1] ;
 wire \top_I.branch[19].block[15].um_I.ana[2] ;
 wire \top_I.branch[19].block[15].um_I.ana[3] ;
 wire \top_I.branch[19].block[15].um_I.ana[4] ;
 wire \top_I.branch[19].block[15].um_I.ana[5] ;
 wire \top_I.branch[19].block[15].um_I.ana[6] ;
 wire \top_I.branch[19].block[15].um_I.ana[7] ;
 wire \top_I.branch[19].block[15].um_I.clk ;
 wire \top_I.branch[19].block[15].um_I.ena ;
 wire \top_I.branch[19].block[15].um_I.iw[10] ;
 wire \top_I.branch[19].block[15].um_I.iw[11] ;
 wire \top_I.branch[19].block[15].um_I.iw[12] ;
 wire \top_I.branch[19].block[15].um_I.iw[13] ;
 wire \top_I.branch[19].block[15].um_I.iw[14] ;
 wire \top_I.branch[19].block[15].um_I.iw[15] ;
 wire \top_I.branch[19].block[15].um_I.iw[16] ;
 wire \top_I.branch[19].block[15].um_I.iw[17] ;
 wire \top_I.branch[19].block[15].um_I.iw[1] ;
 wire \top_I.branch[19].block[15].um_I.iw[2] ;
 wire \top_I.branch[19].block[15].um_I.iw[3] ;
 wire \top_I.branch[19].block[15].um_I.iw[4] ;
 wire \top_I.branch[19].block[15].um_I.iw[5] ;
 wire \top_I.branch[19].block[15].um_I.iw[6] ;
 wire \top_I.branch[19].block[15].um_I.iw[7] ;
 wire \top_I.branch[19].block[15].um_I.iw[8] ;
 wire \top_I.branch[19].block[15].um_I.iw[9] ;
 wire \top_I.branch[19].block[15].um_I.k_zero ;
 wire \top_I.branch[19].block[15].um_I.pg_vdd ;
 wire \top_I.branch[19].block[1].um_I.ana[0] ;
 wire \top_I.branch[19].block[1].um_I.ana[1] ;
 wire \top_I.branch[19].block[1].um_I.ana[2] ;
 wire \top_I.branch[19].block[1].um_I.ana[3] ;
 wire \top_I.branch[19].block[1].um_I.ana[4] ;
 wire \top_I.branch[19].block[1].um_I.ana[5] ;
 wire \top_I.branch[19].block[1].um_I.ana[6] ;
 wire \top_I.branch[19].block[1].um_I.ana[7] ;
 wire \top_I.branch[19].block[1].um_I.clk ;
 wire \top_I.branch[19].block[1].um_I.ena ;
 wire \top_I.branch[19].block[1].um_I.iw[10] ;
 wire \top_I.branch[19].block[1].um_I.iw[11] ;
 wire \top_I.branch[19].block[1].um_I.iw[12] ;
 wire \top_I.branch[19].block[1].um_I.iw[13] ;
 wire \top_I.branch[19].block[1].um_I.iw[14] ;
 wire \top_I.branch[19].block[1].um_I.iw[15] ;
 wire \top_I.branch[19].block[1].um_I.iw[16] ;
 wire \top_I.branch[19].block[1].um_I.iw[17] ;
 wire \top_I.branch[19].block[1].um_I.iw[1] ;
 wire \top_I.branch[19].block[1].um_I.iw[2] ;
 wire \top_I.branch[19].block[1].um_I.iw[3] ;
 wire \top_I.branch[19].block[1].um_I.iw[4] ;
 wire \top_I.branch[19].block[1].um_I.iw[5] ;
 wire \top_I.branch[19].block[1].um_I.iw[6] ;
 wire \top_I.branch[19].block[1].um_I.iw[7] ;
 wire \top_I.branch[19].block[1].um_I.iw[8] ;
 wire \top_I.branch[19].block[1].um_I.iw[9] ;
 wire \top_I.branch[19].block[1].um_I.k_zero ;
 wire \top_I.branch[19].block[1].um_I.pg_vdd ;
 wire \top_I.branch[19].block[2].um_I.ana[0] ;
 wire \top_I.branch[19].block[2].um_I.ana[1] ;
 wire \top_I.branch[19].block[2].um_I.ana[2] ;
 wire \top_I.branch[19].block[2].um_I.ana[3] ;
 wire \top_I.branch[19].block[2].um_I.ana[4] ;
 wire \top_I.branch[19].block[2].um_I.ana[5] ;
 wire \top_I.branch[19].block[2].um_I.ana[6] ;
 wire \top_I.branch[19].block[2].um_I.ana[7] ;
 wire \top_I.branch[19].block[2].um_I.clk ;
 wire \top_I.branch[19].block[2].um_I.ena ;
 wire \top_I.branch[19].block[2].um_I.iw[10] ;
 wire \top_I.branch[19].block[2].um_I.iw[11] ;
 wire \top_I.branch[19].block[2].um_I.iw[12] ;
 wire \top_I.branch[19].block[2].um_I.iw[13] ;
 wire \top_I.branch[19].block[2].um_I.iw[14] ;
 wire \top_I.branch[19].block[2].um_I.iw[15] ;
 wire \top_I.branch[19].block[2].um_I.iw[16] ;
 wire \top_I.branch[19].block[2].um_I.iw[17] ;
 wire \top_I.branch[19].block[2].um_I.iw[1] ;
 wire \top_I.branch[19].block[2].um_I.iw[2] ;
 wire \top_I.branch[19].block[2].um_I.iw[3] ;
 wire \top_I.branch[19].block[2].um_I.iw[4] ;
 wire \top_I.branch[19].block[2].um_I.iw[5] ;
 wire \top_I.branch[19].block[2].um_I.iw[6] ;
 wire \top_I.branch[19].block[2].um_I.iw[7] ;
 wire \top_I.branch[19].block[2].um_I.iw[8] ;
 wire \top_I.branch[19].block[2].um_I.iw[9] ;
 wire \top_I.branch[19].block[2].um_I.k_zero ;
 wire \top_I.branch[19].block[2].um_I.pg_vdd ;
 wire \top_I.branch[19].block[3].um_I.ana[0] ;
 wire \top_I.branch[19].block[3].um_I.ana[1] ;
 wire \top_I.branch[19].block[3].um_I.ana[2] ;
 wire \top_I.branch[19].block[3].um_I.ana[3] ;
 wire \top_I.branch[19].block[3].um_I.ana[4] ;
 wire \top_I.branch[19].block[3].um_I.ana[5] ;
 wire \top_I.branch[19].block[3].um_I.ana[6] ;
 wire \top_I.branch[19].block[3].um_I.ana[7] ;
 wire \top_I.branch[19].block[3].um_I.clk ;
 wire \top_I.branch[19].block[3].um_I.ena ;
 wire \top_I.branch[19].block[3].um_I.iw[10] ;
 wire \top_I.branch[19].block[3].um_I.iw[11] ;
 wire \top_I.branch[19].block[3].um_I.iw[12] ;
 wire \top_I.branch[19].block[3].um_I.iw[13] ;
 wire \top_I.branch[19].block[3].um_I.iw[14] ;
 wire \top_I.branch[19].block[3].um_I.iw[15] ;
 wire \top_I.branch[19].block[3].um_I.iw[16] ;
 wire \top_I.branch[19].block[3].um_I.iw[17] ;
 wire \top_I.branch[19].block[3].um_I.iw[1] ;
 wire \top_I.branch[19].block[3].um_I.iw[2] ;
 wire \top_I.branch[19].block[3].um_I.iw[3] ;
 wire \top_I.branch[19].block[3].um_I.iw[4] ;
 wire \top_I.branch[19].block[3].um_I.iw[5] ;
 wire \top_I.branch[19].block[3].um_I.iw[6] ;
 wire \top_I.branch[19].block[3].um_I.iw[7] ;
 wire \top_I.branch[19].block[3].um_I.iw[8] ;
 wire \top_I.branch[19].block[3].um_I.iw[9] ;
 wire \top_I.branch[19].block[3].um_I.k_zero ;
 wire \top_I.branch[19].block[3].um_I.pg_vdd ;
 wire \top_I.branch[19].block[4].um_I.ana[0] ;
 wire \top_I.branch[19].block[4].um_I.ana[1] ;
 wire \top_I.branch[19].block[4].um_I.ana[2] ;
 wire \top_I.branch[19].block[4].um_I.ana[3] ;
 wire \top_I.branch[19].block[4].um_I.ana[4] ;
 wire \top_I.branch[19].block[4].um_I.ana[5] ;
 wire \top_I.branch[19].block[4].um_I.ana[6] ;
 wire \top_I.branch[19].block[4].um_I.ana[7] ;
 wire \top_I.branch[19].block[4].um_I.clk ;
 wire \top_I.branch[19].block[4].um_I.ena ;
 wire \top_I.branch[19].block[4].um_I.iw[10] ;
 wire \top_I.branch[19].block[4].um_I.iw[11] ;
 wire \top_I.branch[19].block[4].um_I.iw[12] ;
 wire \top_I.branch[19].block[4].um_I.iw[13] ;
 wire \top_I.branch[19].block[4].um_I.iw[14] ;
 wire \top_I.branch[19].block[4].um_I.iw[15] ;
 wire \top_I.branch[19].block[4].um_I.iw[16] ;
 wire \top_I.branch[19].block[4].um_I.iw[17] ;
 wire \top_I.branch[19].block[4].um_I.iw[1] ;
 wire \top_I.branch[19].block[4].um_I.iw[2] ;
 wire \top_I.branch[19].block[4].um_I.iw[3] ;
 wire \top_I.branch[19].block[4].um_I.iw[4] ;
 wire \top_I.branch[19].block[4].um_I.iw[5] ;
 wire \top_I.branch[19].block[4].um_I.iw[6] ;
 wire \top_I.branch[19].block[4].um_I.iw[7] ;
 wire \top_I.branch[19].block[4].um_I.iw[8] ;
 wire \top_I.branch[19].block[4].um_I.iw[9] ;
 wire \top_I.branch[19].block[4].um_I.k_zero ;
 wire \top_I.branch[19].block[4].um_I.pg_vdd ;
 wire \top_I.branch[19].block[5].um_I.ana[0] ;
 wire \top_I.branch[19].block[5].um_I.ana[1] ;
 wire \top_I.branch[19].block[5].um_I.ana[2] ;
 wire \top_I.branch[19].block[5].um_I.ana[3] ;
 wire \top_I.branch[19].block[5].um_I.ana[4] ;
 wire \top_I.branch[19].block[5].um_I.ana[5] ;
 wire \top_I.branch[19].block[5].um_I.ana[6] ;
 wire \top_I.branch[19].block[5].um_I.ana[7] ;
 wire \top_I.branch[19].block[5].um_I.clk ;
 wire \top_I.branch[19].block[5].um_I.ena ;
 wire \top_I.branch[19].block[5].um_I.iw[10] ;
 wire \top_I.branch[19].block[5].um_I.iw[11] ;
 wire \top_I.branch[19].block[5].um_I.iw[12] ;
 wire \top_I.branch[19].block[5].um_I.iw[13] ;
 wire \top_I.branch[19].block[5].um_I.iw[14] ;
 wire \top_I.branch[19].block[5].um_I.iw[15] ;
 wire \top_I.branch[19].block[5].um_I.iw[16] ;
 wire \top_I.branch[19].block[5].um_I.iw[17] ;
 wire \top_I.branch[19].block[5].um_I.iw[1] ;
 wire \top_I.branch[19].block[5].um_I.iw[2] ;
 wire \top_I.branch[19].block[5].um_I.iw[3] ;
 wire \top_I.branch[19].block[5].um_I.iw[4] ;
 wire \top_I.branch[19].block[5].um_I.iw[5] ;
 wire \top_I.branch[19].block[5].um_I.iw[6] ;
 wire \top_I.branch[19].block[5].um_I.iw[7] ;
 wire \top_I.branch[19].block[5].um_I.iw[8] ;
 wire \top_I.branch[19].block[5].um_I.iw[9] ;
 wire \top_I.branch[19].block[5].um_I.k_zero ;
 wire \top_I.branch[19].block[5].um_I.pg_vdd ;
 wire \top_I.branch[19].block[6].um_I.ana[0] ;
 wire \top_I.branch[19].block[6].um_I.ana[1] ;
 wire \top_I.branch[19].block[6].um_I.ana[2] ;
 wire \top_I.branch[19].block[6].um_I.ana[3] ;
 wire \top_I.branch[19].block[6].um_I.ana[4] ;
 wire \top_I.branch[19].block[6].um_I.ana[5] ;
 wire \top_I.branch[19].block[6].um_I.ana[6] ;
 wire \top_I.branch[19].block[6].um_I.ana[7] ;
 wire \top_I.branch[19].block[6].um_I.clk ;
 wire \top_I.branch[19].block[6].um_I.ena ;
 wire \top_I.branch[19].block[6].um_I.iw[10] ;
 wire \top_I.branch[19].block[6].um_I.iw[11] ;
 wire \top_I.branch[19].block[6].um_I.iw[12] ;
 wire \top_I.branch[19].block[6].um_I.iw[13] ;
 wire \top_I.branch[19].block[6].um_I.iw[14] ;
 wire \top_I.branch[19].block[6].um_I.iw[15] ;
 wire \top_I.branch[19].block[6].um_I.iw[16] ;
 wire \top_I.branch[19].block[6].um_I.iw[17] ;
 wire \top_I.branch[19].block[6].um_I.iw[1] ;
 wire \top_I.branch[19].block[6].um_I.iw[2] ;
 wire \top_I.branch[19].block[6].um_I.iw[3] ;
 wire \top_I.branch[19].block[6].um_I.iw[4] ;
 wire \top_I.branch[19].block[6].um_I.iw[5] ;
 wire \top_I.branch[19].block[6].um_I.iw[6] ;
 wire \top_I.branch[19].block[6].um_I.iw[7] ;
 wire \top_I.branch[19].block[6].um_I.iw[8] ;
 wire \top_I.branch[19].block[6].um_I.iw[9] ;
 wire \top_I.branch[19].block[6].um_I.k_zero ;
 wire \top_I.branch[19].block[6].um_I.pg_vdd ;
 wire \top_I.branch[19].block[7].um_I.ana[0] ;
 wire \top_I.branch[19].block[7].um_I.ana[1] ;
 wire \top_I.branch[19].block[7].um_I.ana[2] ;
 wire \top_I.branch[19].block[7].um_I.ana[3] ;
 wire \top_I.branch[19].block[7].um_I.ana[4] ;
 wire \top_I.branch[19].block[7].um_I.ana[5] ;
 wire \top_I.branch[19].block[7].um_I.ana[6] ;
 wire \top_I.branch[19].block[7].um_I.ana[7] ;
 wire \top_I.branch[19].block[7].um_I.clk ;
 wire \top_I.branch[19].block[7].um_I.ena ;
 wire \top_I.branch[19].block[7].um_I.iw[10] ;
 wire \top_I.branch[19].block[7].um_I.iw[11] ;
 wire \top_I.branch[19].block[7].um_I.iw[12] ;
 wire \top_I.branch[19].block[7].um_I.iw[13] ;
 wire \top_I.branch[19].block[7].um_I.iw[14] ;
 wire \top_I.branch[19].block[7].um_I.iw[15] ;
 wire \top_I.branch[19].block[7].um_I.iw[16] ;
 wire \top_I.branch[19].block[7].um_I.iw[17] ;
 wire \top_I.branch[19].block[7].um_I.iw[1] ;
 wire \top_I.branch[19].block[7].um_I.iw[2] ;
 wire \top_I.branch[19].block[7].um_I.iw[3] ;
 wire \top_I.branch[19].block[7].um_I.iw[4] ;
 wire \top_I.branch[19].block[7].um_I.iw[5] ;
 wire \top_I.branch[19].block[7].um_I.iw[6] ;
 wire \top_I.branch[19].block[7].um_I.iw[7] ;
 wire \top_I.branch[19].block[7].um_I.iw[8] ;
 wire \top_I.branch[19].block[7].um_I.iw[9] ;
 wire \top_I.branch[19].block[7].um_I.k_zero ;
 wire \top_I.branch[19].block[7].um_I.pg_vdd ;
 wire \top_I.branch[19].block[8].um_I.ana[0] ;
 wire \top_I.branch[19].block[8].um_I.ana[1] ;
 wire \top_I.branch[19].block[8].um_I.ana[2] ;
 wire \top_I.branch[19].block[8].um_I.ana[3] ;
 wire \top_I.branch[19].block[8].um_I.ana[4] ;
 wire \top_I.branch[19].block[8].um_I.ana[5] ;
 wire \top_I.branch[19].block[8].um_I.ana[6] ;
 wire \top_I.branch[19].block[8].um_I.ana[7] ;
 wire \top_I.branch[19].block[8].um_I.clk ;
 wire \top_I.branch[19].block[8].um_I.ena ;
 wire \top_I.branch[19].block[8].um_I.iw[10] ;
 wire \top_I.branch[19].block[8].um_I.iw[11] ;
 wire \top_I.branch[19].block[8].um_I.iw[12] ;
 wire \top_I.branch[19].block[8].um_I.iw[13] ;
 wire \top_I.branch[19].block[8].um_I.iw[14] ;
 wire \top_I.branch[19].block[8].um_I.iw[15] ;
 wire \top_I.branch[19].block[8].um_I.iw[16] ;
 wire \top_I.branch[19].block[8].um_I.iw[17] ;
 wire \top_I.branch[19].block[8].um_I.iw[1] ;
 wire \top_I.branch[19].block[8].um_I.iw[2] ;
 wire \top_I.branch[19].block[8].um_I.iw[3] ;
 wire \top_I.branch[19].block[8].um_I.iw[4] ;
 wire \top_I.branch[19].block[8].um_I.iw[5] ;
 wire \top_I.branch[19].block[8].um_I.iw[6] ;
 wire \top_I.branch[19].block[8].um_I.iw[7] ;
 wire \top_I.branch[19].block[8].um_I.iw[8] ;
 wire \top_I.branch[19].block[8].um_I.iw[9] ;
 wire \top_I.branch[19].block[8].um_I.k_zero ;
 wire \top_I.branch[19].block[8].um_I.pg_vdd ;
 wire \top_I.branch[19].block[9].um_I.ana[0] ;
 wire \top_I.branch[19].block[9].um_I.ana[1] ;
 wire \top_I.branch[19].block[9].um_I.ana[2] ;
 wire \top_I.branch[19].block[9].um_I.ana[3] ;
 wire \top_I.branch[19].block[9].um_I.ana[4] ;
 wire \top_I.branch[19].block[9].um_I.ana[5] ;
 wire \top_I.branch[19].block[9].um_I.ana[6] ;
 wire \top_I.branch[19].block[9].um_I.ana[7] ;
 wire \top_I.branch[19].block[9].um_I.clk ;
 wire \top_I.branch[19].block[9].um_I.ena ;
 wire \top_I.branch[19].block[9].um_I.iw[10] ;
 wire \top_I.branch[19].block[9].um_I.iw[11] ;
 wire \top_I.branch[19].block[9].um_I.iw[12] ;
 wire \top_I.branch[19].block[9].um_I.iw[13] ;
 wire \top_I.branch[19].block[9].um_I.iw[14] ;
 wire \top_I.branch[19].block[9].um_I.iw[15] ;
 wire \top_I.branch[19].block[9].um_I.iw[16] ;
 wire \top_I.branch[19].block[9].um_I.iw[17] ;
 wire \top_I.branch[19].block[9].um_I.iw[1] ;
 wire \top_I.branch[19].block[9].um_I.iw[2] ;
 wire \top_I.branch[19].block[9].um_I.iw[3] ;
 wire \top_I.branch[19].block[9].um_I.iw[4] ;
 wire \top_I.branch[19].block[9].um_I.iw[5] ;
 wire \top_I.branch[19].block[9].um_I.iw[6] ;
 wire \top_I.branch[19].block[9].um_I.iw[7] ;
 wire \top_I.branch[19].block[9].um_I.iw[8] ;
 wire \top_I.branch[19].block[9].um_I.iw[9] ;
 wire \top_I.branch[19].block[9].um_I.k_zero ;
 wire \top_I.branch[19].block[9].um_I.pg_vdd ;
 wire \top_I.branch[19].l_addr[0] ;
 wire \top_I.branch[19].l_addr[1] ;
 wire \top_I.branch[1].block[0].um_I.ana[0] ;
 wire \top_I.branch[1].block[0].um_I.ana[1] ;
 wire \top_I.branch[1].block[0].um_I.ana[2] ;
 wire \top_I.branch[1].block[0].um_I.ana[3] ;
 wire \top_I.branch[1].block[0].um_I.ana[4] ;
 wire \top_I.branch[1].block[0].um_I.ana[5] ;
 wire \top_I.branch[1].block[0].um_I.ana[6] ;
 wire \top_I.branch[1].block[0].um_I.ana[7] ;
 wire \top_I.branch[1].block[0].um_I.clk ;
 wire \top_I.branch[1].block[0].um_I.ena ;
 wire \top_I.branch[1].block[0].um_I.iw[10] ;
 wire \top_I.branch[1].block[0].um_I.iw[11] ;
 wire \top_I.branch[1].block[0].um_I.iw[12] ;
 wire \top_I.branch[1].block[0].um_I.iw[13] ;
 wire \top_I.branch[1].block[0].um_I.iw[14] ;
 wire \top_I.branch[1].block[0].um_I.iw[15] ;
 wire \top_I.branch[1].block[0].um_I.iw[16] ;
 wire \top_I.branch[1].block[0].um_I.iw[17] ;
 wire \top_I.branch[1].block[0].um_I.iw[1] ;
 wire \top_I.branch[1].block[0].um_I.iw[2] ;
 wire \top_I.branch[1].block[0].um_I.iw[3] ;
 wire \top_I.branch[1].block[0].um_I.iw[4] ;
 wire \top_I.branch[1].block[0].um_I.iw[5] ;
 wire \top_I.branch[1].block[0].um_I.iw[6] ;
 wire \top_I.branch[1].block[0].um_I.iw[7] ;
 wire \top_I.branch[1].block[0].um_I.iw[8] ;
 wire \top_I.branch[1].block[0].um_I.iw[9] ;
 wire \top_I.branch[1].block[0].um_I.k_zero ;
 wire \top_I.branch[1].block[0].um_I.pg_vdd ;
 wire \top_I.branch[1].block[10].um_I.ana[0] ;
 wire \top_I.branch[1].block[10].um_I.ana[1] ;
 wire \top_I.branch[1].block[10].um_I.ana[2] ;
 wire \top_I.branch[1].block[10].um_I.ana[3] ;
 wire \top_I.branch[1].block[10].um_I.ana[4] ;
 wire \top_I.branch[1].block[10].um_I.ana[5] ;
 wire \top_I.branch[1].block[10].um_I.ana[6] ;
 wire \top_I.branch[1].block[10].um_I.ana[7] ;
 wire \top_I.branch[1].block[10].um_I.clk ;
 wire \top_I.branch[1].block[10].um_I.ena ;
 wire \top_I.branch[1].block[10].um_I.iw[10] ;
 wire \top_I.branch[1].block[10].um_I.iw[11] ;
 wire \top_I.branch[1].block[10].um_I.iw[12] ;
 wire \top_I.branch[1].block[10].um_I.iw[13] ;
 wire \top_I.branch[1].block[10].um_I.iw[14] ;
 wire \top_I.branch[1].block[10].um_I.iw[15] ;
 wire \top_I.branch[1].block[10].um_I.iw[16] ;
 wire \top_I.branch[1].block[10].um_I.iw[17] ;
 wire \top_I.branch[1].block[10].um_I.iw[1] ;
 wire \top_I.branch[1].block[10].um_I.iw[2] ;
 wire \top_I.branch[1].block[10].um_I.iw[3] ;
 wire \top_I.branch[1].block[10].um_I.iw[4] ;
 wire \top_I.branch[1].block[10].um_I.iw[5] ;
 wire \top_I.branch[1].block[10].um_I.iw[6] ;
 wire \top_I.branch[1].block[10].um_I.iw[7] ;
 wire \top_I.branch[1].block[10].um_I.iw[8] ;
 wire \top_I.branch[1].block[10].um_I.iw[9] ;
 wire \top_I.branch[1].block[10].um_I.k_zero ;
 wire \top_I.branch[1].block[10].um_I.pg_vdd ;
 wire \top_I.branch[1].block[11].um_I.ana[0] ;
 wire \top_I.branch[1].block[11].um_I.ana[1] ;
 wire \top_I.branch[1].block[11].um_I.ana[2] ;
 wire \top_I.branch[1].block[11].um_I.ana[3] ;
 wire \top_I.branch[1].block[11].um_I.ana[4] ;
 wire \top_I.branch[1].block[11].um_I.ana[5] ;
 wire \top_I.branch[1].block[11].um_I.ana[6] ;
 wire \top_I.branch[1].block[11].um_I.ana[7] ;
 wire \top_I.branch[1].block[11].um_I.clk ;
 wire \top_I.branch[1].block[11].um_I.ena ;
 wire \top_I.branch[1].block[11].um_I.iw[10] ;
 wire \top_I.branch[1].block[11].um_I.iw[11] ;
 wire \top_I.branch[1].block[11].um_I.iw[12] ;
 wire \top_I.branch[1].block[11].um_I.iw[13] ;
 wire \top_I.branch[1].block[11].um_I.iw[14] ;
 wire \top_I.branch[1].block[11].um_I.iw[15] ;
 wire \top_I.branch[1].block[11].um_I.iw[16] ;
 wire \top_I.branch[1].block[11].um_I.iw[17] ;
 wire \top_I.branch[1].block[11].um_I.iw[1] ;
 wire \top_I.branch[1].block[11].um_I.iw[2] ;
 wire \top_I.branch[1].block[11].um_I.iw[3] ;
 wire \top_I.branch[1].block[11].um_I.iw[4] ;
 wire \top_I.branch[1].block[11].um_I.iw[5] ;
 wire \top_I.branch[1].block[11].um_I.iw[6] ;
 wire \top_I.branch[1].block[11].um_I.iw[7] ;
 wire \top_I.branch[1].block[11].um_I.iw[8] ;
 wire \top_I.branch[1].block[11].um_I.iw[9] ;
 wire \top_I.branch[1].block[11].um_I.k_zero ;
 wire \top_I.branch[1].block[11].um_I.pg_vdd ;
 wire \top_I.branch[1].block[12].um_I.ana[0] ;
 wire \top_I.branch[1].block[12].um_I.ana[1] ;
 wire \top_I.branch[1].block[12].um_I.ana[2] ;
 wire \top_I.branch[1].block[12].um_I.ana[3] ;
 wire \top_I.branch[1].block[12].um_I.ana[4] ;
 wire \top_I.branch[1].block[12].um_I.ana[5] ;
 wire \top_I.branch[1].block[12].um_I.ana[6] ;
 wire \top_I.branch[1].block[12].um_I.ana[7] ;
 wire \top_I.branch[1].block[12].um_I.clk ;
 wire \top_I.branch[1].block[12].um_I.ena ;
 wire \top_I.branch[1].block[12].um_I.iw[10] ;
 wire \top_I.branch[1].block[12].um_I.iw[11] ;
 wire \top_I.branch[1].block[12].um_I.iw[12] ;
 wire \top_I.branch[1].block[12].um_I.iw[13] ;
 wire \top_I.branch[1].block[12].um_I.iw[14] ;
 wire \top_I.branch[1].block[12].um_I.iw[15] ;
 wire \top_I.branch[1].block[12].um_I.iw[16] ;
 wire \top_I.branch[1].block[12].um_I.iw[17] ;
 wire \top_I.branch[1].block[12].um_I.iw[1] ;
 wire \top_I.branch[1].block[12].um_I.iw[2] ;
 wire \top_I.branch[1].block[12].um_I.iw[3] ;
 wire \top_I.branch[1].block[12].um_I.iw[4] ;
 wire \top_I.branch[1].block[12].um_I.iw[5] ;
 wire \top_I.branch[1].block[12].um_I.iw[6] ;
 wire \top_I.branch[1].block[12].um_I.iw[7] ;
 wire \top_I.branch[1].block[12].um_I.iw[8] ;
 wire \top_I.branch[1].block[12].um_I.iw[9] ;
 wire \top_I.branch[1].block[12].um_I.k_zero ;
 wire \top_I.branch[1].block[12].um_I.pg_vdd ;
 wire \top_I.branch[1].block[13].um_I.ana[0] ;
 wire \top_I.branch[1].block[13].um_I.ana[1] ;
 wire \top_I.branch[1].block[13].um_I.ana[2] ;
 wire \top_I.branch[1].block[13].um_I.ana[3] ;
 wire \top_I.branch[1].block[13].um_I.ana[4] ;
 wire \top_I.branch[1].block[13].um_I.ana[5] ;
 wire \top_I.branch[1].block[13].um_I.ana[6] ;
 wire \top_I.branch[1].block[13].um_I.ana[7] ;
 wire \top_I.branch[1].block[13].um_I.clk ;
 wire \top_I.branch[1].block[13].um_I.ena ;
 wire \top_I.branch[1].block[13].um_I.iw[10] ;
 wire \top_I.branch[1].block[13].um_I.iw[11] ;
 wire \top_I.branch[1].block[13].um_I.iw[12] ;
 wire \top_I.branch[1].block[13].um_I.iw[13] ;
 wire \top_I.branch[1].block[13].um_I.iw[14] ;
 wire \top_I.branch[1].block[13].um_I.iw[15] ;
 wire \top_I.branch[1].block[13].um_I.iw[16] ;
 wire \top_I.branch[1].block[13].um_I.iw[17] ;
 wire \top_I.branch[1].block[13].um_I.iw[1] ;
 wire \top_I.branch[1].block[13].um_I.iw[2] ;
 wire \top_I.branch[1].block[13].um_I.iw[3] ;
 wire \top_I.branch[1].block[13].um_I.iw[4] ;
 wire \top_I.branch[1].block[13].um_I.iw[5] ;
 wire \top_I.branch[1].block[13].um_I.iw[6] ;
 wire \top_I.branch[1].block[13].um_I.iw[7] ;
 wire \top_I.branch[1].block[13].um_I.iw[8] ;
 wire \top_I.branch[1].block[13].um_I.iw[9] ;
 wire \top_I.branch[1].block[13].um_I.k_zero ;
 wire \top_I.branch[1].block[13].um_I.pg_vdd ;
 wire \top_I.branch[1].block[14].um_I.ana[0] ;
 wire \top_I.branch[1].block[14].um_I.ana[1] ;
 wire \top_I.branch[1].block[14].um_I.ana[2] ;
 wire \top_I.branch[1].block[14].um_I.ana[3] ;
 wire \top_I.branch[1].block[14].um_I.ana[4] ;
 wire \top_I.branch[1].block[14].um_I.ana[5] ;
 wire \top_I.branch[1].block[14].um_I.ana[6] ;
 wire \top_I.branch[1].block[14].um_I.ana[7] ;
 wire \top_I.branch[1].block[14].um_I.clk ;
 wire \top_I.branch[1].block[14].um_I.ena ;
 wire \top_I.branch[1].block[14].um_I.iw[10] ;
 wire \top_I.branch[1].block[14].um_I.iw[11] ;
 wire \top_I.branch[1].block[14].um_I.iw[12] ;
 wire \top_I.branch[1].block[14].um_I.iw[13] ;
 wire \top_I.branch[1].block[14].um_I.iw[14] ;
 wire \top_I.branch[1].block[14].um_I.iw[15] ;
 wire \top_I.branch[1].block[14].um_I.iw[16] ;
 wire \top_I.branch[1].block[14].um_I.iw[17] ;
 wire \top_I.branch[1].block[14].um_I.iw[1] ;
 wire \top_I.branch[1].block[14].um_I.iw[2] ;
 wire \top_I.branch[1].block[14].um_I.iw[3] ;
 wire \top_I.branch[1].block[14].um_I.iw[4] ;
 wire \top_I.branch[1].block[14].um_I.iw[5] ;
 wire \top_I.branch[1].block[14].um_I.iw[6] ;
 wire \top_I.branch[1].block[14].um_I.iw[7] ;
 wire \top_I.branch[1].block[14].um_I.iw[8] ;
 wire \top_I.branch[1].block[14].um_I.iw[9] ;
 wire \top_I.branch[1].block[14].um_I.k_zero ;
 wire \top_I.branch[1].block[14].um_I.pg_vdd ;
 wire \top_I.branch[1].block[15].um_I.ana[0] ;
 wire \top_I.branch[1].block[15].um_I.ana[1] ;
 wire \top_I.branch[1].block[15].um_I.ana[2] ;
 wire \top_I.branch[1].block[15].um_I.ana[3] ;
 wire \top_I.branch[1].block[15].um_I.ana[4] ;
 wire \top_I.branch[1].block[15].um_I.ana[5] ;
 wire \top_I.branch[1].block[15].um_I.ana[6] ;
 wire \top_I.branch[1].block[15].um_I.ana[7] ;
 wire \top_I.branch[1].block[15].um_I.clk ;
 wire \top_I.branch[1].block[15].um_I.ena ;
 wire \top_I.branch[1].block[15].um_I.iw[10] ;
 wire \top_I.branch[1].block[15].um_I.iw[11] ;
 wire \top_I.branch[1].block[15].um_I.iw[12] ;
 wire \top_I.branch[1].block[15].um_I.iw[13] ;
 wire \top_I.branch[1].block[15].um_I.iw[14] ;
 wire \top_I.branch[1].block[15].um_I.iw[15] ;
 wire \top_I.branch[1].block[15].um_I.iw[16] ;
 wire \top_I.branch[1].block[15].um_I.iw[17] ;
 wire \top_I.branch[1].block[15].um_I.iw[1] ;
 wire \top_I.branch[1].block[15].um_I.iw[2] ;
 wire \top_I.branch[1].block[15].um_I.iw[3] ;
 wire \top_I.branch[1].block[15].um_I.iw[4] ;
 wire \top_I.branch[1].block[15].um_I.iw[5] ;
 wire \top_I.branch[1].block[15].um_I.iw[6] ;
 wire \top_I.branch[1].block[15].um_I.iw[7] ;
 wire \top_I.branch[1].block[15].um_I.iw[8] ;
 wire \top_I.branch[1].block[15].um_I.iw[9] ;
 wire \top_I.branch[1].block[15].um_I.k_zero ;
 wire \top_I.branch[1].block[15].um_I.pg_vdd ;
 wire \top_I.branch[1].block[1].um_I.ana[0] ;
 wire \top_I.branch[1].block[1].um_I.ana[1] ;
 wire \top_I.branch[1].block[1].um_I.ana[2] ;
 wire \top_I.branch[1].block[1].um_I.ana[3] ;
 wire \top_I.branch[1].block[1].um_I.ana[4] ;
 wire \top_I.branch[1].block[1].um_I.ana[5] ;
 wire \top_I.branch[1].block[1].um_I.ana[6] ;
 wire \top_I.branch[1].block[1].um_I.ana[7] ;
 wire \top_I.branch[1].block[1].um_I.clk ;
 wire \top_I.branch[1].block[1].um_I.ena ;
 wire \top_I.branch[1].block[1].um_I.iw[10] ;
 wire \top_I.branch[1].block[1].um_I.iw[11] ;
 wire \top_I.branch[1].block[1].um_I.iw[12] ;
 wire \top_I.branch[1].block[1].um_I.iw[13] ;
 wire \top_I.branch[1].block[1].um_I.iw[14] ;
 wire \top_I.branch[1].block[1].um_I.iw[15] ;
 wire \top_I.branch[1].block[1].um_I.iw[16] ;
 wire \top_I.branch[1].block[1].um_I.iw[17] ;
 wire \top_I.branch[1].block[1].um_I.iw[1] ;
 wire \top_I.branch[1].block[1].um_I.iw[2] ;
 wire \top_I.branch[1].block[1].um_I.iw[3] ;
 wire \top_I.branch[1].block[1].um_I.iw[4] ;
 wire \top_I.branch[1].block[1].um_I.iw[5] ;
 wire \top_I.branch[1].block[1].um_I.iw[6] ;
 wire \top_I.branch[1].block[1].um_I.iw[7] ;
 wire \top_I.branch[1].block[1].um_I.iw[8] ;
 wire \top_I.branch[1].block[1].um_I.iw[9] ;
 wire \top_I.branch[1].block[1].um_I.k_zero ;
 wire \top_I.branch[1].block[1].um_I.pg_vdd ;
 wire \top_I.branch[1].block[2].um_I.ana[0] ;
 wire \top_I.branch[1].block[2].um_I.ana[1] ;
 wire \top_I.branch[1].block[2].um_I.ana[2] ;
 wire \top_I.branch[1].block[2].um_I.ana[3] ;
 wire \top_I.branch[1].block[2].um_I.ana[4] ;
 wire \top_I.branch[1].block[2].um_I.ana[5] ;
 wire \top_I.branch[1].block[2].um_I.ana[6] ;
 wire \top_I.branch[1].block[2].um_I.ana[7] ;
 wire \top_I.branch[1].block[2].um_I.clk ;
 wire \top_I.branch[1].block[2].um_I.ena ;
 wire \top_I.branch[1].block[2].um_I.iw[10] ;
 wire \top_I.branch[1].block[2].um_I.iw[11] ;
 wire \top_I.branch[1].block[2].um_I.iw[12] ;
 wire \top_I.branch[1].block[2].um_I.iw[13] ;
 wire \top_I.branch[1].block[2].um_I.iw[14] ;
 wire \top_I.branch[1].block[2].um_I.iw[15] ;
 wire \top_I.branch[1].block[2].um_I.iw[16] ;
 wire \top_I.branch[1].block[2].um_I.iw[17] ;
 wire \top_I.branch[1].block[2].um_I.iw[1] ;
 wire \top_I.branch[1].block[2].um_I.iw[2] ;
 wire \top_I.branch[1].block[2].um_I.iw[3] ;
 wire \top_I.branch[1].block[2].um_I.iw[4] ;
 wire \top_I.branch[1].block[2].um_I.iw[5] ;
 wire \top_I.branch[1].block[2].um_I.iw[6] ;
 wire \top_I.branch[1].block[2].um_I.iw[7] ;
 wire \top_I.branch[1].block[2].um_I.iw[8] ;
 wire \top_I.branch[1].block[2].um_I.iw[9] ;
 wire \top_I.branch[1].block[2].um_I.k_zero ;
 wire \top_I.branch[1].block[2].um_I.pg_vdd ;
 wire \top_I.branch[1].block[3].um_I.ana[0] ;
 wire \top_I.branch[1].block[3].um_I.ana[1] ;
 wire \top_I.branch[1].block[3].um_I.ana[2] ;
 wire \top_I.branch[1].block[3].um_I.ana[3] ;
 wire \top_I.branch[1].block[3].um_I.ana[4] ;
 wire \top_I.branch[1].block[3].um_I.ana[5] ;
 wire \top_I.branch[1].block[3].um_I.ana[6] ;
 wire \top_I.branch[1].block[3].um_I.ana[7] ;
 wire \top_I.branch[1].block[3].um_I.clk ;
 wire \top_I.branch[1].block[3].um_I.ena ;
 wire \top_I.branch[1].block[3].um_I.iw[10] ;
 wire \top_I.branch[1].block[3].um_I.iw[11] ;
 wire \top_I.branch[1].block[3].um_I.iw[12] ;
 wire \top_I.branch[1].block[3].um_I.iw[13] ;
 wire \top_I.branch[1].block[3].um_I.iw[14] ;
 wire \top_I.branch[1].block[3].um_I.iw[15] ;
 wire \top_I.branch[1].block[3].um_I.iw[16] ;
 wire \top_I.branch[1].block[3].um_I.iw[17] ;
 wire \top_I.branch[1].block[3].um_I.iw[1] ;
 wire \top_I.branch[1].block[3].um_I.iw[2] ;
 wire \top_I.branch[1].block[3].um_I.iw[3] ;
 wire \top_I.branch[1].block[3].um_I.iw[4] ;
 wire \top_I.branch[1].block[3].um_I.iw[5] ;
 wire \top_I.branch[1].block[3].um_I.iw[6] ;
 wire \top_I.branch[1].block[3].um_I.iw[7] ;
 wire \top_I.branch[1].block[3].um_I.iw[8] ;
 wire \top_I.branch[1].block[3].um_I.iw[9] ;
 wire \top_I.branch[1].block[3].um_I.k_zero ;
 wire \top_I.branch[1].block[3].um_I.pg_vdd ;
 wire \top_I.branch[1].block[4].um_I.ana[0] ;
 wire \top_I.branch[1].block[4].um_I.ana[1] ;
 wire \top_I.branch[1].block[4].um_I.ana[2] ;
 wire \top_I.branch[1].block[4].um_I.ana[3] ;
 wire \top_I.branch[1].block[4].um_I.ana[4] ;
 wire \top_I.branch[1].block[4].um_I.ana[5] ;
 wire \top_I.branch[1].block[4].um_I.ana[6] ;
 wire \top_I.branch[1].block[4].um_I.ana[7] ;
 wire \top_I.branch[1].block[4].um_I.clk ;
 wire \top_I.branch[1].block[4].um_I.ena ;
 wire \top_I.branch[1].block[4].um_I.iw[10] ;
 wire \top_I.branch[1].block[4].um_I.iw[11] ;
 wire \top_I.branch[1].block[4].um_I.iw[12] ;
 wire \top_I.branch[1].block[4].um_I.iw[13] ;
 wire \top_I.branch[1].block[4].um_I.iw[14] ;
 wire \top_I.branch[1].block[4].um_I.iw[15] ;
 wire \top_I.branch[1].block[4].um_I.iw[16] ;
 wire \top_I.branch[1].block[4].um_I.iw[17] ;
 wire \top_I.branch[1].block[4].um_I.iw[1] ;
 wire \top_I.branch[1].block[4].um_I.iw[2] ;
 wire \top_I.branch[1].block[4].um_I.iw[3] ;
 wire \top_I.branch[1].block[4].um_I.iw[4] ;
 wire \top_I.branch[1].block[4].um_I.iw[5] ;
 wire \top_I.branch[1].block[4].um_I.iw[6] ;
 wire \top_I.branch[1].block[4].um_I.iw[7] ;
 wire \top_I.branch[1].block[4].um_I.iw[8] ;
 wire \top_I.branch[1].block[4].um_I.iw[9] ;
 wire \top_I.branch[1].block[4].um_I.k_zero ;
 wire \top_I.branch[1].block[4].um_I.pg_vdd ;
 wire \top_I.branch[1].block[5].um_I.ana[0] ;
 wire \top_I.branch[1].block[5].um_I.ana[1] ;
 wire \top_I.branch[1].block[5].um_I.ana[2] ;
 wire \top_I.branch[1].block[5].um_I.ana[3] ;
 wire \top_I.branch[1].block[5].um_I.ana[4] ;
 wire \top_I.branch[1].block[5].um_I.ana[5] ;
 wire \top_I.branch[1].block[5].um_I.ana[6] ;
 wire \top_I.branch[1].block[5].um_I.ana[7] ;
 wire \top_I.branch[1].block[5].um_I.clk ;
 wire \top_I.branch[1].block[5].um_I.ena ;
 wire \top_I.branch[1].block[5].um_I.iw[10] ;
 wire \top_I.branch[1].block[5].um_I.iw[11] ;
 wire \top_I.branch[1].block[5].um_I.iw[12] ;
 wire \top_I.branch[1].block[5].um_I.iw[13] ;
 wire \top_I.branch[1].block[5].um_I.iw[14] ;
 wire \top_I.branch[1].block[5].um_I.iw[15] ;
 wire \top_I.branch[1].block[5].um_I.iw[16] ;
 wire \top_I.branch[1].block[5].um_I.iw[17] ;
 wire \top_I.branch[1].block[5].um_I.iw[1] ;
 wire \top_I.branch[1].block[5].um_I.iw[2] ;
 wire \top_I.branch[1].block[5].um_I.iw[3] ;
 wire \top_I.branch[1].block[5].um_I.iw[4] ;
 wire \top_I.branch[1].block[5].um_I.iw[5] ;
 wire \top_I.branch[1].block[5].um_I.iw[6] ;
 wire \top_I.branch[1].block[5].um_I.iw[7] ;
 wire \top_I.branch[1].block[5].um_I.iw[8] ;
 wire \top_I.branch[1].block[5].um_I.iw[9] ;
 wire \top_I.branch[1].block[5].um_I.k_zero ;
 wire \top_I.branch[1].block[5].um_I.pg_vdd ;
 wire \top_I.branch[1].block[6].um_I.ana[0] ;
 wire \top_I.branch[1].block[6].um_I.ana[1] ;
 wire \top_I.branch[1].block[6].um_I.ana[2] ;
 wire \top_I.branch[1].block[6].um_I.ana[3] ;
 wire \top_I.branch[1].block[6].um_I.ana[4] ;
 wire \top_I.branch[1].block[6].um_I.ana[5] ;
 wire \top_I.branch[1].block[6].um_I.ana[6] ;
 wire \top_I.branch[1].block[6].um_I.ana[7] ;
 wire \top_I.branch[1].block[6].um_I.clk ;
 wire \top_I.branch[1].block[6].um_I.ena ;
 wire \top_I.branch[1].block[6].um_I.iw[10] ;
 wire \top_I.branch[1].block[6].um_I.iw[11] ;
 wire \top_I.branch[1].block[6].um_I.iw[12] ;
 wire \top_I.branch[1].block[6].um_I.iw[13] ;
 wire \top_I.branch[1].block[6].um_I.iw[14] ;
 wire \top_I.branch[1].block[6].um_I.iw[15] ;
 wire \top_I.branch[1].block[6].um_I.iw[16] ;
 wire \top_I.branch[1].block[6].um_I.iw[17] ;
 wire \top_I.branch[1].block[6].um_I.iw[1] ;
 wire \top_I.branch[1].block[6].um_I.iw[2] ;
 wire \top_I.branch[1].block[6].um_I.iw[3] ;
 wire \top_I.branch[1].block[6].um_I.iw[4] ;
 wire \top_I.branch[1].block[6].um_I.iw[5] ;
 wire \top_I.branch[1].block[6].um_I.iw[6] ;
 wire \top_I.branch[1].block[6].um_I.iw[7] ;
 wire \top_I.branch[1].block[6].um_I.iw[8] ;
 wire \top_I.branch[1].block[6].um_I.iw[9] ;
 wire \top_I.branch[1].block[6].um_I.k_zero ;
 wire \top_I.branch[1].block[6].um_I.pg_vdd ;
 wire \top_I.branch[1].block[7].um_I.ana[0] ;
 wire \top_I.branch[1].block[7].um_I.ana[1] ;
 wire \top_I.branch[1].block[7].um_I.ana[2] ;
 wire \top_I.branch[1].block[7].um_I.ana[3] ;
 wire \top_I.branch[1].block[7].um_I.ana[4] ;
 wire \top_I.branch[1].block[7].um_I.ana[5] ;
 wire \top_I.branch[1].block[7].um_I.ana[6] ;
 wire \top_I.branch[1].block[7].um_I.ana[7] ;
 wire \top_I.branch[1].block[7].um_I.clk ;
 wire \top_I.branch[1].block[7].um_I.ena ;
 wire \top_I.branch[1].block[7].um_I.iw[10] ;
 wire \top_I.branch[1].block[7].um_I.iw[11] ;
 wire \top_I.branch[1].block[7].um_I.iw[12] ;
 wire \top_I.branch[1].block[7].um_I.iw[13] ;
 wire \top_I.branch[1].block[7].um_I.iw[14] ;
 wire \top_I.branch[1].block[7].um_I.iw[15] ;
 wire \top_I.branch[1].block[7].um_I.iw[16] ;
 wire \top_I.branch[1].block[7].um_I.iw[17] ;
 wire \top_I.branch[1].block[7].um_I.iw[1] ;
 wire \top_I.branch[1].block[7].um_I.iw[2] ;
 wire \top_I.branch[1].block[7].um_I.iw[3] ;
 wire \top_I.branch[1].block[7].um_I.iw[4] ;
 wire \top_I.branch[1].block[7].um_I.iw[5] ;
 wire \top_I.branch[1].block[7].um_I.iw[6] ;
 wire \top_I.branch[1].block[7].um_I.iw[7] ;
 wire \top_I.branch[1].block[7].um_I.iw[8] ;
 wire \top_I.branch[1].block[7].um_I.iw[9] ;
 wire \top_I.branch[1].block[7].um_I.k_zero ;
 wire \top_I.branch[1].block[7].um_I.pg_vdd ;
 wire \top_I.branch[1].block[8].um_I.ana[0] ;
 wire \top_I.branch[1].block[8].um_I.ana[1] ;
 wire \top_I.branch[1].block[8].um_I.ana[2] ;
 wire \top_I.branch[1].block[8].um_I.ana[3] ;
 wire \top_I.branch[1].block[8].um_I.ana[4] ;
 wire \top_I.branch[1].block[8].um_I.ana[5] ;
 wire \top_I.branch[1].block[8].um_I.ana[6] ;
 wire \top_I.branch[1].block[8].um_I.ana[7] ;
 wire \top_I.branch[1].block[8].um_I.clk ;
 wire \top_I.branch[1].block[8].um_I.ena ;
 wire \top_I.branch[1].block[8].um_I.iw[10] ;
 wire \top_I.branch[1].block[8].um_I.iw[11] ;
 wire \top_I.branch[1].block[8].um_I.iw[12] ;
 wire \top_I.branch[1].block[8].um_I.iw[13] ;
 wire \top_I.branch[1].block[8].um_I.iw[14] ;
 wire \top_I.branch[1].block[8].um_I.iw[15] ;
 wire \top_I.branch[1].block[8].um_I.iw[16] ;
 wire \top_I.branch[1].block[8].um_I.iw[17] ;
 wire \top_I.branch[1].block[8].um_I.iw[1] ;
 wire \top_I.branch[1].block[8].um_I.iw[2] ;
 wire \top_I.branch[1].block[8].um_I.iw[3] ;
 wire \top_I.branch[1].block[8].um_I.iw[4] ;
 wire \top_I.branch[1].block[8].um_I.iw[5] ;
 wire \top_I.branch[1].block[8].um_I.iw[6] ;
 wire \top_I.branch[1].block[8].um_I.iw[7] ;
 wire \top_I.branch[1].block[8].um_I.iw[8] ;
 wire \top_I.branch[1].block[8].um_I.iw[9] ;
 wire \top_I.branch[1].block[8].um_I.k_zero ;
 wire \top_I.branch[1].block[8].um_I.pg_vdd ;
 wire \top_I.branch[1].block[9].um_I.ana[0] ;
 wire \top_I.branch[1].block[9].um_I.ana[1] ;
 wire \top_I.branch[1].block[9].um_I.ana[2] ;
 wire \top_I.branch[1].block[9].um_I.ana[3] ;
 wire \top_I.branch[1].block[9].um_I.ana[4] ;
 wire \top_I.branch[1].block[9].um_I.ana[5] ;
 wire \top_I.branch[1].block[9].um_I.ana[6] ;
 wire \top_I.branch[1].block[9].um_I.ana[7] ;
 wire \top_I.branch[1].block[9].um_I.clk ;
 wire \top_I.branch[1].block[9].um_I.ena ;
 wire \top_I.branch[1].block[9].um_I.iw[10] ;
 wire \top_I.branch[1].block[9].um_I.iw[11] ;
 wire \top_I.branch[1].block[9].um_I.iw[12] ;
 wire \top_I.branch[1].block[9].um_I.iw[13] ;
 wire \top_I.branch[1].block[9].um_I.iw[14] ;
 wire \top_I.branch[1].block[9].um_I.iw[15] ;
 wire \top_I.branch[1].block[9].um_I.iw[16] ;
 wire \top_I.branch[1].block[9].um_I.iw[17] ;
 wire \top_I.branch[1].block[9].um_I.iw[1] ;
 wire \top_I.branch[1].block[9].um_I.iw[2] ;
 wire \top_I.branch[1].block[9].um_I.iw[3] ;
 wire \top_I.branch[1].block[9].um_I.iw[4] ;
 wire \top_I.branch[1].block[9].um_I.iw[5] ;
 wire \top_I.branch[1].block[9].um_I.iw[6] ;
 wire \top_I.branch[1].block[9].um_I.iw[7] ;
 wire \top_I.branch[1].block[9].um_I.iw[8] ;
 wire \top_I.branch[1].block[9].um_I.iw[9] ;
 wire \top_I.branch[1].block[9].um_I.k_zero ;
 wire \top_I.branch[1].block[9].um_I.pg_vdd ;
 wire \top_I.branch[1].l_addr[0] ;
 wire \top_I.branch[1].l_k_one ;
 wire \top_I.branch[20].block[0].um_I.ana[0] ;
 wire \top_I.branch[20].block[0].um_I.ana[1] ;
 wire \top_I.branch[20].block[0].um_I.ana[2] ;
 wire \top_I.branch[20].block[0].um_I.ana[3] ;
 wire \top_I.branch[20].block[0].um_I.ana[4] ;
 wire \top_I.branch[20].block[0].um_I.ana[5] ;
 wire \top_I.branch[20].block[0].um_I.ana[6] ;
 wire \top_I.branch[20].block[0].um_I.ana[7] ;
 wire \top_I.branch[20].block[0].um_I.clk ;
 wire \top_I.branch[20].block[0].um_I.ena ;
 wire \top_I.branch[20].block[0].um_I.iw[10] ;
 wire \top_I.branch[20].block[0].um_I.iw[11] ;
 wire \top_I.branch[20].block[0].um_I.iw[12] ;
 wire \top_I.branch[20].block[0].um_I.iw[13] ;
 wire \top_I.branch[20].block[0].um_I.iw[14] ;
 wire \top_I.branch[20].block[0].um_I.iw[15] ;
 wire \top_I.branch[20].block[0].um_I.iw[16] ;
 wire \top_I.branch[20].block[0].um_I.iw[17] ;
 wire \top_I.branch[20].block[0].um_I.iw[1] ;
 wire \top_I.branch[20].block[0].um_I.iw[2] ;
 wire \top_I.branch[20].block[0].um_I.iw[3] ;
 wire \top_I.branch[20].block[0].um_I.iw[4] ;
 wire \top_I.branch[20].block[0].um_I.iw[5] ;
 wire \top_I.branch[20].block[0].um_I.iw[6] ;
 wire \top_I.branch[20].block[0].um_I.iw[7] ;
 wire \top_I.branch[20].block[0].um_I.iw[8] ;
 wire \top_I.branch[20].block[0].um_I.iw[9] ;
 wire \top_I.branch[20].block[0].um_I.k_zero ;
 wire \top_I.branch[20].block[0].um_I.pg_vdd ;
 wire \top_I.branch[20].block[10].um_I.ana[0] ;
 wire \top_I.branch[20].block[10].um_I.ana[1] ;
 wire \top_I.branch[20].block[10].um_I.ana[2] ;
 wire \top_I.branch[20].block[10].um_I.ana[3] ;
 wire \top_I.branch[20].block[10].um_I.ana[4] ;
 wire \top_I.branch[20].block[10].um_I.ana[5] ;
 wire \top_I.branch[20].block[10].um_I.ana[6] ;
 wire \top_I.branch[20].block[10].um_I.ana[7] ;
 wire \top_I.branch[20].block[10].um_I.clk ;
 wire \top_I.branch[20].block[10].um_I.ena ;
 wire \top_I.branch[20].block[10].um_I.iw[10] ;
 wire \top_I.branch[20].block[10].um_I.iw[11] ;
 wire \top_I.branch[20].block[10].um_I.iw[12] ;
 wire \top_I.branch[20].block[10].um_I.iw[13] ;
 wire \top_I.branch[20].block[10].um_I.iw[14] ;
 wire \top_I.branch[20].block[10].um_I.iw[15] ;
 wire \top_I.branch[20].block[10].um_I.iw[16] ;
 wire \top_I.branch[20].block[10].um_I.iw[17] ;
 wire \top_I.branch[20].block[10].um_I.iw[1] ;
 wire \top_I.branch[20].block[10].um_I.iw[2] ;
 wire \top_I.branch[20].block[10].um_I.iw[3] ;
 wire \top_I.branch[20].block[10].um_I.iw[4] ;
 wire \top_I.branch[20].block[10].um_I.iw[5] ;
 wire \top_I.branch[20].block[10].um_I.iw[6] ;
 wire \top_I.branch[20].block[10].um_I.iw[7] ;
 wire \top_I.branch[20].block[10].um_I.iw[8] ;
 wire \top_I.branch[20].block[10].um_I.iw[9] ;
 wire \top_I.branch[20].block[10].um_I.k_zero ;
 wire \top_I.branch[20].block[10].um_I.pg_vdd ;
 wire \top_I.branch[20].block[11].um_I.ana[0] ;
 wire \top_I.branch[20].block[11].um_I.ana[1] ;
 wire \top_I.branch[20].block[11].um_I.ana[2] ;
 wire \top_I.branch[20].block[11].um_I.ana[3] ;
 wire \top_I.branch[20].block[11].um_I.ana[4] ;
 wire \top_I.branch[20].block[11].um_I.ana[5] ;
 wire \top_I.branch[20].block[11].um_I.ana[6] ;
 wire \top_I.branch[20].block[11].um_I.ana[7] ;
 wire \top_I.branch[20].block[11].um_I.clk ;
 wire \top_I.branch[20].block[11].um_I.ena ;
 wire \top_I.branch[20].block[11].um_I.iw[10] ;
 wire \top_I.branch[20].block[11].um_I.iw[11] ;
 wire \top_I.branch[20].block[11].um_I.iw[12] ;
 wire \top_I.branch[20].block[11].um_I.iw[13] ;
 wire \top_I.branch[20].block[11].um_I.iw[14] ;
 wire \top_I.branch[20].block[11].um_I.iw[15] ;
 wire \top_I.branch[20].block[11].um_I.iw[16] ;
 wire \top_I.branch[20].block[11].um_I.iw[17] ;
 wire \top_I.branch[20].block[11].um_I.iw[1] ;
 wire \top_I.branch[20].block[11].um_I.iw[2] ;
 wire \top_I.branch[20].block[11].um_I.iw[3] ;
 wire \top_I.branch[20].block[11].um_I.iw[4] ;
 wire \top_I.branch[20].block[11].um_I.iw[5] ;
 wire \top_I.branch[20].block[11].um_I.iw[6] ;
 wire \top_I.branch[20].block[11].um_I.iw[7] ;
 wire \top_I.branch[20].block[11].um_I.iw[8] ;
 wire \top_I.branch[20].block[11].um_I.iw[9] ;
 wire \top_I.branch[20].block[11].um_I.k_zero ;
 wire \top_I.branch[20].block[11].um_I.pg_vdd ;
 wire \top_I.branch[20].block[12].um_I.ana[0] ;
 wire \top_I.branch[20].block[12].um_I.ana[1] ;
 wire \top_I.branch[20].block[12].um_I.ana[2] ;
 wire \top_I.branch[20].block[12].um_I.ana[3] ;
 wire \top_I.branch[20].block[12].um_I.ana[4] ;
 wire \top_I.branch[20].block[12].um_I.ana[5] ;
 wire \top_I.branch[20].block[12].um_I.ana[6] ;
 wire \top_I.branch[20].block[12].um_I.ana[7] ;
 wire \top_I.branch[20].block[12].um_I.clk ;
 wire \top_I.branch[20].block[12].um_I.ena ;
 wire \top_I.branch[20].block[12].um_I.iw[10] ;
 wire \top_I.branch[20].block[12].um_I.iw[11] ;
 wire \top_I.branch[20].block[12].um_I.iw[12] ;
 wire \top_I.branch[20].block[12].um_I.iw[13] ;
 wire \top_I.branch[20].block[12].um_I.iw[14] ;
 wire \top_I.branch[20].block[12].um_I.iw[15] ;
 wire \top_I.branch[20].block[12].um_I.iw[16] ;
 wire \top_I.branch[20].block[12].um_I.iw[17] ;
 wire \top_I.branch[20].block[12].um_I.iw[1] ;
 wire \top_I.branch[20].block[12].um_I.iw[2] ;
 wire \top_I.branch[20].block[12].um_I.iw[3] ;
 wire \top_I.branch[20].block[12].um_I.iw[4] ;
 wire \top_I.branch[20].block[12].um_I.iw[5] ;
 wire \top_I.branch[20].block[12].um_I.iw[6] ;
 wire \top_I.branch[20].block[12].um_I.iw[7] ;
 wire \top_I.branch[20].block[12].um_I.iw[8] ;
 wire \top_I.branch[20].block[12].um_I.iw[9] ;
 wire \top_I.branch[20].block[12].um_I.k_zero ;
 wire \top_I.branch[20].block[12].um_I.pg_vdd ;
 wire \top_I.branch[20].block[13].um_I.ana[0] ;
 wire \top_I.branch[20].block[13].um_I.ana[1] ;
 wire \top_I.branch[20].block[13].um_I.ana[2] ;
 wire \top_I.branch[20].block[13].um_I.ana[3] ;
 wire \top_I.branch[20].block[13].um_I.ana[4] ;
 wire \top_I.branch[20].block[13].um_I.ana[5] ;
 wire \top_I.branch[20].block[13].um_I.ana[6] ;
 wire \top_I.branch[20].block[13].um_I.ana[7] ;
 wire \top_I.branch[20].block[13].um_I.clk ;
 wire \top_I.branch[20].block[13].um_I.ena ;
 wire \top_I.branch[20].block[13].um_I.iw[10] ;
 wire \top_I.branch[20].block[13].um_I.iw[11] ;
 wire \top_I.branch[20].block[13].um_I.iw[12] ;
 wire \top_I.branch[20].block[13].um_I.iw[13] ;
 wire \top_I.branch[20].block[13].um_I.iw[14] ;
 wire \top_I.branch[20].block[13].um_I.iw[15] ;
 wire \top_I.branch[20].block[13].um_I.iw[16] ;
 wire \top_I.branch[20].block[13].um_I.iw[17] ;
 wire \top_I.branch[20].block[13].um_I.iw[1] ;
 wire \top_I.branch[20].block[13].um_I.iw[2] ;
 wire \top_I.branch[20].block[13].um_I.iw[3] ;
 wire \top_I.branch[20].block[13].um_I.iw[4] ;
 wire \top_I.branch[20].block[13].um_I.iw[5] ;
 wire \top_I.branch[20].block[13].um_I.iw[6] ;
 wire \top_I.branch[20].block[13].um_I.iw[7] ;
 wire \top_I.branch[20].block[13].um_I.iw[8] ;
 wire \top_I.branch[20].block[13].um_I.iw[9] ;
 wire \top_I.branch[20].block[13].um_I.k_zero ;
 wire \top_I.branch[20].block[13].um_I.pg_vdd ;
 wire \top_I.branch[20].block[14].um_I.ana[0] ;
 wire \top_I.branch[20].block[14].um_I.ana[1] ;
 wire \top_I.branch[20].block[14].um_I.ana[2] ;
 wire \top_I.branch[20].block[14].um_I.ana[3] ;
 wire \top_I.branch[20].block[14].um_I.ana[4] ;
 wire \top_I.branch[20].block[14].um_I.ana[5] ;
 wire \top_I.branch[20].block[14].um_I.ana[6] ;
 wire \top_I.branch[20].block[14].um_I.ana[7] ;
 wire \top_I.branch[20].block[14].um_I.clk ;
 wire \top_I.branch[20].block[14].um_I.ena ;
 wire \top_I.branch[20].block[14].um_I.iw[10] ;
 wire \top_I.branch[20].block[14].um_I.iw[11] ;
 wire \top_I.branch[20].block[14].um_I.iw[12] ;
 wire \top_I.branch[20].block[14].um_I.iw[13] ;
 wire \top_I.branch[20].block[14].um_I.iw[14] ;
 wire \top_I.branch[20].block[14].um_I.iw[15] ;
 wire \top_I.branch[20].block[14].um_I.iw[16] ;
 wire \top_I.branch[20].block[14].um_I.iw[17] ;
 wire \top_I.branch[20].block[14].um_I.iw[1] ;
 wire \top_I.branch[20].block[14].um_I.iw[2] ;
 wire \top_I.branch[20].block[14].um_I.iw[3] ;
 wire \top_I.branch[20].block[14].um_I.iw[4] ;
 wire \top_I.branch[20].block[14].um_I.iw[5] ;
 wire \top_I.branch[20].block[14].um_I.iw[6] ;
 wire \top_I.branch[20].block[14].um_I.iw[7] ;
 wire \top_I.branch[20].block[14].um_I.iw[8] ;
 wire \top_I.branch[20].block[14].um_I.iw[9] ;
 wire \top_I.branch[20].block[14].um_I.k_zero ;
 wire \top_I.branch[20].block[14].um_I.pg_vdd ;
 wire \top_I.branch[20].block[15].um_I.ana[0] ;
 wire \top_I.branch[20].block[15].um_I.ana[1] ;
 wire \top_I.branch[20].block[15].um_I.ana[2] ;
 wire \top_I.branch[20].block[15].um_I.ana[3] ;
 wire \top_I.branch[20].block[15].um_I.ana[4] ;
 wire \top_I.branch[20].block[15].um_I.ana[5] ;
 wire \top_I.branch[20].block[15].um_I.ana[6] ;
 wire \top_I.branch[20].block[15].um_I.ana[7] ;
 wire \top_I.branch[20].block[15].um_I.clk ;
 wire \top_I.branch[20].block[15].um_I.ena ;
 wire \top_I.branch[20].block[15].um_I.iw[10] ;
 wire \top_I.branch[20].block[15].um_I.iw[11] ;
 wire \top_I.branch[20].block[15].um_I.iw[12] ;
 wire \top_I.branch[20].block[15].um_I.iw[13] ;
 wire \top_I.branch[20].block[15].um_I.iw[14] ;
 wire \top_I.branch[20].block[15].um_I.iw[15] ;
 wire \top_I.branch[20].block[15].um_I.iw[16] ;
 wire \top_I.branch[20].block[15].um_I.iw[17] ;
 wire \top_I.branch[20].block[15].um_I.iw[1] ;
 wire \top_I.branch[20].block[15].um_I.iw[2] ;
 wire \top_I.branch[20].block[15].um_I.iw[3] ;
 wire \top_I.branch[20].block[15].um_I.iw[4] ;
 wire \top_I.branch[20].block[15].um_I.iw[5] ;
 wire \top_I.branch[20].block[15].um_I.iw[6] ;
 wire \top_I.branch[20].block[15].um_I.iw[7] ;
 wire \top_I.branch[20].block[15].um_I.iw[8] ;
 wire \top_I.branch[20].block[15].um_I.iw[9] ;
 wire \top_I.branch[20].block[15].um_I.k_zero ;
 wire \top_I.branch[20].block[15].um_I.pg_vdd ;
 wire \top_I.branch[20].block[1].um_I.ana[0] ;
 wire \top_I.branch[20].block[1].um_I.ana[1] ;
 wire \top_I.branch[20].block[1].um_I.ana[2] ;
 wire \top_I.branch[20].block[1].um_I.ana[3] ;
 wire \top_I.branch[20].block[1].um_I.ana[4] ;
 wire \top_I.branch[20].block[1].um_I.ana[5] ;
 wire \top_I.branch[20].block[1].um_I.ana[6] ;
 wire \top_I.branch[20].block[1].um_I.ana[7] ;
 wire \top_I.branch[20].block[1].um_I.clk ;
 wire \top_I.branch[20].block[1].um_I.ena ;
 wire \top_I.branch[20].block[1].um_I.iw[10] ;
 wire \top_I.branch[20].block[1].um_I.iw[11] ;
 wire \top_I.branch[20].block[1].um_I.iw[12] ;
 wire \top_I.branch[20].block[1].um_I.iw[13] ;
 wire \top_I.branch[20].block[1].um_I.iw[14] ;
 wire \top_I.branch[20].block[1].um_I.iw[15] ;
 wire \top_I.branch[20].block[1].um_I.iw[16] ;
 wire \top_I.branch[20].block[1].um_I.iw[17] ;
 wire \top_I.branch[20].block[1].um_I.iw[1] ;
 wire \top_I.branch[20].block[1].um_I.iw[2] ;
 wire \top_I.branch[20].block[1].um_I.iw[3] ;
 wire \top_I.branch[20].block[1].um_I.iw[4] ;
 wire \top_I.branch[20].block[1].um_I.iw[5] ;
 wire \top_I.branch[20].block[1].um_I.iw[6] ;
 wire \top_I.branch[20].block[1].um_I.iw[7] ;
 wire \top_I.branch[20].block[1].um_I.iw[8] ;
 wire \top_I.branch[20].block[1].um_I.iw[9] ;
 wire \top_I.branch[20].block[1].um_I.k_zero ;
 wire \top_I.branch[20].block[1].um_I.pg_vdd ;
 wire \top_I.branch[20].block[2].um_I.ana[0] ;
 wire \top_I.branch[20].block[2].um_I.ana[1] ;
 wire \top_I.branch[20].block[2].um_I.ana[2] ;
 wire \top_I.branch[20].block[2].um_I.ana[3] ;
 wire \top_I.branch[20].block[2].um_I.ana[4] ;
 wire \top_I.branch[20].block[2].um_I.ana[5] ;
 wire \top_I.branch[20].block[2].um_I.ana[6] ;
 wire \top_I.branch[20].block[2].um_I.ana[7] ;
 wire \top_I.branch[20].block[2].um_I.clk ;
 wire \top_I.branch[20].block[2].um_I.ena ;
 wire \top_I.branch[20].block[2].um_I.iw[10] ;
 wire \top_I.branch[20].block[2].um_I.iw[11] ;
 wire \top_I.branch[20].block[2].um_I.iw[12] ;
 wire \top_I.branch[20].block[2].um_I.iw[13] ;
 wire \top_I.branch[20].block[2].um_I.iw[14] ;
 wire \top_I.branch[20].block[2].um_I.iw[15] ;
 wire \top_I.branch[20].block[2].um_I.iw[16] ;
 wire \top_I.branch[20].block[2].um_I.iw[17] ;
 wire \top_I.branch[20].block[2].um_I.iw[1] ;
 wire \top_I.branch[20].block[2].um_I.iw[2] ;
 wire \top_I.branch[20].block[2].um_I.iw[3] ;
 wire \top_I.branch[20].block[2].um_I.iw[4] ;
 wire \top_I.branch[20].block[2].um_I.iw[5] ;
 wire \top_I.branch[20].block[2].um_I.iw[6] ;
 wire \top_I.branch[20].block[2].um_I.iw[7] ;
 wire \top_I.branch[20].block[2].um_I.iw[8] ;
 wire \top_I.branch[20].block[2].um_I.iw[9] ;
 wire \top_I.branch[20].block[2].um_I.k_zero ;
 wire \top_I.branch[20].block[2].um_I.pg_vdd ;
 wire \top_I.branch[20].block[3].um_I.ana[0] ;
 wire \top_I.branch[20].block[3].um_I.ana[1] ;
 wire \top_I.branch[20].block[3].um_I.ana[2] ;
 wire \top_I.branch[20].block[3].um_I.ana[3] ;
 wire \top_I.branch[20].block[3].um_I.ana[4] ;
 wire \top_I.branch[20].block[3].um_I.ana[5] ;
 wire \top_I.branch[20].block[3].um_I.ana[6] ;
 wire \top_I.branch[20].block[3].um_I.ana[7] ;
 wire \top_I.branch[20].block[3].um_I.clk ;
 wire \top_I.branch[20].block[3].um_I.ena ;
 wire \top_I.branch[20].block[3].um_I.iw[10] ;
 wire \top_I.branch[20].block[3].um_I.iw[11] ;
 wire \top_I.branch[20].block[3].um_I.iw[12] ;
 wire \top_I.branch[20].block[3].um_I.iw[13] ;
 wire \top_I.branch[20].block[3].um_I.iw[14] ;
 wire \top_I.branch[20].block[3].um_I.iw[15] ;
 wire \top_I.branch[20].block[3].um_I.iw[16] ;
 wire \top_I.branch[20].block[3].um_I.iw[17] ;
 wire \top_I.branch[20].block[3].um_I.iw[1] ;
 wire \top_I.branch[20].block[3].um_I.iw[2] ;
 wire \top_I.branch[20].block[3].um_I.iw[3] ;
 wire \top_I.branch[20].block[3].um_I.iw[4] ;
 wire \top_I.branch[20].block[3].um_I.iw[5] ;
 wire \top_I.branch[20].block[3].um_I.iw[6] ;
 wire \top_I.branch[20].block[3].um_I.iw[7] ;
 wire \top_I.branch[20].block[3].um_I.iw[8] ;
 wire \top_I.branch[20].block[3].um_I.iw[9] ;
 wire \top_I.branch[20].block[3].um_I.k_zero ;
 wire \top_I.branch[20].block[3].um_I.pg_vdd ;
 wire \top_I.branch[20].block[4].um_I.ana[0] ;
 wire \top_I.branch[20].block[4].um_I.ana[1] ;
 wire \top_I.branch[20].block[4].um_I.ana[2] ;
 wire \top_I.branch[20].block[4].um_I.ana[3] ;
 wire \top_I.branch[20].block[4].um_I.ana[4] ;
 wire \top_I.branch[20].block[4].um_I.ana[5] ;
 wire \top_I.branch[20].block[4].um_I.ana[6] ;
 wire \top_I.branch[20].block[4].um_I.ana[7] ;
 wire \top_I.branch[20].block[4].um_I.clk ;
 wire \top_I.branch[20].block[4].um_I.ena ;
 wire \top_I.branch[20].block[4].um_I.iw[10] ;
 wire \top_I.branch[20].block[4].um_I.iw[11] ;
 wire \top_I.branch[20].block[4].um_I.iw[12] ;
 wire \top_I.branch[20].block[4].um_I.iw[13] ;
 wire \top_I.branch[20].block[4].um_I.iw[14] ;
 wire \top_I.branch[20].block[4].um_I.iw[15] ;
 wire \top_I.branch[20].block[4].um_I.iw[16] ;
 wire \top_I.branch[20].block[4].um_I.iw[17] ;
 wire \top_I.branch[20].block[4].um_I.iw[1] ;
 wire \top_I.branch[20].block[4].um_I.iw[2] ;
 wire \top_I.branch[20].block[4].um_I.iw[3] ;
 wire \top_I.branch[20].block[4].um_I.iw[4] ;
 wire \top_I.branch[20].block[4].um_I.iw[5] ;
 wire \top_I.branch[20].block[4].um_I.iw[6] ;
 wire \top_I.branch[20].block[4].um_I.iw[7] ;
 wire \top_I.branch[20].block[4].um_I.iw[8] ;
 wire \top_I.branch[20].block[4].um_I.iw[9] ;
 wire \top_I.branch[20].block[4].um_I.k_zero ;
 wire \top_I.branch[20].block[4].um_I.pg_vdd ;
 wire \top_I.branch[20].block[5].um_I.ana[0] ;
 wire \top_I.branch[20].block[5].um_I.ana[1] ;
 wire \top_I.branch[20].block[5].um_I.ana[2] ;
 wire \top_I.branch[20].block[5].um_I.ana[3] ;
 wire \top_I.branch[20].block[5].um_I.ana[4] ;
 wire \top_I.branch[20].block[5].um_I.ana[5] ;
 wire \top_I.branch[20].block[5].um_I.ana[6] ;
 wire \top_I.branch[20].block[5].um_I.ana[7] ;
 wire \top_I.branch[20].block[5].um_I.clk ;
 wire \top_I.branch[20].block[5].um_I.ena ;
 wire \top_I.branch[20].block[5].um_I.iw[10] ;
 wire \top_I.branch[20].block[5].um_I.iw[11] ;
 wire \top_I.branch[20].block[5].um_I.iw[12] ;
 wire \top_I.branch[20].block[5].um_I.iw[13] ;
 wire \top_I.branch[20].block[5].um_I.iw[14] ;
 wire \top_I.branch[20].block[5].um_I.iw[15] ;
 wire \top_I.branch[20].block[5].um_I.iw[16] ;
 wire \top_I.branch[20].block[5].um_I.iw[17] ;
 wire \top_I.branch[20].block[5].um_I.iw[1] ;
 wire \top_I.branch[20].block[5].um_I.iw[2] ;
 wire \top_I.branch[20].block[5].um_I.iw[3] ;
 wire \top_I.branch[20].block[5].um_I.iw[4] ;
 wire \top_I.branch[20].block[5].um_I.iw[5] ;
 wire \top_I.branch[20].block[5].um_I.iw[6] ;
 wire \top_I.branch[20].block[5].um_I.iw[7] ;
 wire \top_I.branch[20].block[5].um_I.iw[8] ;
 wire \top_I.branch[20].block[5].um_I.iw[9] ;
 wire \top_I.branch[20].block[5].um_I.k_zero ;
 wire \top_I.branch[20].block[5].um_I.pg_vdd ;
 wire \top_I.branch[20].block[6].um_I.ana[0] ;
 wire \top_I.branch[20].block[6].um_I.ana[1] ;
 wire \top_I.branch[20].block[6].um_I.ana[2] ;
 wire \top_I.branch[20].block[6].um_I.ana[3] ;
 wire \top_I.branch[20].block[6].um_I.ana[4] ;
 wire \top_I.branch[20].block[6].um_I.ana[5] ;
 wire \top_I.branch[20].block[6].um_I.ana[6] ;
 wire \top_I.branch[20].block[6].um_I.ana[7] ;
 wire \top_I.branch[20].block[6].um_I.clk ;
 wire \top_I.branch[20].block[6].um_I.ena ;
 wire \top_I.branch[20].block[6].um_I.iw[10] ;
 wire \top_I.branch[20].block[6].um_I.iw[11] ;
 wire \top_I.branch[20].block[6].um_I.iw[12] ;
 wire \top_I.branch[20].block[6].um_I.iw[13] ;
 wire \top_I.branch[20].block[6].um_I.iw[14] ;
 wire \top_I.branch[20].block[6].um_I.iw[15] ;
 wire \top_I.branch[20].block[6].um_I.iw[16] ;
 wire \top_I.branch[20].block[6].um_I.iw[17] ;
 wire \top_I.branch[20].block[6].um_I.iw[1] ;
 wire \top_I.branch[20].block[6].um_I.iw[2] ;
 wire \top_I.branch[20].block[6].um_I.iw[3] ;
 wire \top_I.branch[20].block[6].um_I.iw[4] ;
 wire \top_I.branch[20].block[6].um_I.iw[5] ;
 wire \top_I.branch[20].block[6].um_I.iw[6] ;
 wire \top_I.branch[20].block[6].um_I.iw[7] ;
 wire \top_I.branch[20].block[6].um_I.iw[8] ;
 wire \top_I.branch[20].block[6].um_I.iw[9] ;
 wire \top_I.branch[20].block[6].um_I.k_zero ;
 wire \top_I.branch[20].block[6].um_I.pg_vdd ;
 wire \top_I.branch[20].block[7].um_I.ana[0] ;
 wire \top_I.branch[20].block[7].um_I.ana[1] ;
 wire \top_I.branch[20].block[7].um_I.ana[2] ;
 wire \top_I.branch[20].block[7].um_I.ana[3] ;
 wire \top_I.branch[20].block[7].um_I.ana[4] ;
 wire \top_I.branch[20].block[7].um_I.ana[5] ;
 wire \top_I.branch[20].block[7].um_I.ana[6] ;
 wire \top_I.branch[20].block[7].um_I.ana[7] ;
 wire \top_I.branch[20].block[7].um_I.clk ;
 wire \top_I.branch[20].block[7].um_I.ena ;
 wire \top_I.branch[20].block[7].um_I.iw[10] ;
 wire \top_I.branch[20].block[7].um_I.iw[11] ;
 wire \top_I.branch[20].block[7].um_I.iw[12] ;
 wire \top_I.branch[20].block[7].um_I.iw[13] ;
 wire \top_I.branch[20].block[7].um_I.iw[14] ;
 wire \top_I.branch[20].block[7].um_I.iw[15] ;
 wire \top_I.branch[20].block[7].um_I.iw[16] ;
 wire \top_I.branch[20].block[7].um_I.iw[17] ;
 wire \top_I.branch[20].block[7].um_I.iw[1] ;
 wire \top_I.branch[20].block[7].um_I.iw[2] ;
 wire \top_I.branch[20].block[7].um_I.iw[3] ;
 wire \top_I.branch[20].block[7].um_I.iw[4] ;
 wire \top_I.branch[20].block[7].um_I.iw[5] ;
 wire \top_I.branch[20].block[7].um_I.iw[6] ;
 wire \top_I.branch[20].block[7].um_I.iw[7] ;
 wire \top_I.branch[20].block[7].um_I.iw[8] ;
 wire \top_I.branch[20].block[7].um_I.iw[9] ;
 wire \top_I.branch[20].block[7].um_I.k_zero ;
 wire \top_I.branch[20].block[7].um_I.pg_vdd ;
 wire \top_I.branch[20].block[8].um_I.ana[0] ;
 wire \top_I.branch[20].block[8].um_I.ana[1] ;
 wire \top_I.branch[20].block[8].um_I.ana[2] ;
 wire \top_I.branch[20].block[8].um_I.ana[3] ;
 wire \top_I.branch[20].block[8].um_I.ana[4] ;
 wire \top_I.branch[20].block[8].um_I.ana[5] ;
 wire \top_I.branch[20].block[8].um_I.ana[6] ;
 wire \top_I.branch[20].block[8].um_I.ana[7] ;
 wire \top_I.branch[20].block[8].um_I.clk ;
 wire \top_I.branch[20].block[8].um_I.ena ;
 wire \top_I.branch[20].block[8].um_I.iw[10] ;
 wire \top_I.branch[20].block[8].um_I.iw[11] ;
 wire \top_I.branch[20].block[8].um_I.iw[12] ;
 wire \top_I.branch[20].block[8].um_I.iw[13] ;
 wire \top_I.branch[20].block[8].um_I.iw[14] ;
 wire \top_I.branch[20].block[8].um_I.iw[15] ;
 wire \top_I.branch[20].block[8].um_I.iw[16] ;
 wire \top_I.branch[20].block[8].um_I.iw[17] ;
 wire \top_I.branch[20].block[8].um_I.iw[1] ;
 wire \top_I.branch[20].block[8].um_I.iw[2] ;
 wire \top_I.branch[20].block[8].um_I.iw[3] ;
 wire \top_I.branch[20].block[8].um_I.iw[4] ;
 wire \top_I.branch[20].block[8].um_I.iw[5] ;
 wire \top_I.branch[20].block[8].um_I.iw[6] ;
 wire \top_I.branch[20].block[8].um_I.iw[7] ;
 wire \top_I.branch[20].block[8].um_I.iw[8] ;
 wire \top_I.branch[20].block[8].um_I.iw[9] ;
 wire \top_I.branch[20].block[8].um_I.k_zero ;
 wire \top_I.branch[20].block[8].um_I.pg_vdd ;
 wire \top_I.branch[20].block[9].um_I.ana[0] ;
 wire \top_I.branch[20].block[9].um_I.ana[1] ;
 wire \top_I.branch[20].block[9].um_I.ana[2] ;
 wire \top_I.branch[20].block[9].um_I.ana[3] ;
 wire \top_I.branch[20].block[9].um_I.ana[4] ;
 wire \top_I.branch[20].block[9].um_I.ana[5] ;
 wire \top_I.branch[20].block[9].um_I.ana[6] ;
 wire \top_I.branch[20].block[9].um_I.ana[7] ;
 wire \top_I.branch[20].block[9].um_I.clk ;
 wire \top_I.branch[20].block[9].um_I.ena ;
 wire \top_I.branch[20].block[9].um_I.iw[10] ;
 wire \top_I.branch[20].block[9].um_I.iw[11] ;
 wire \top_I.branch[20].block[9].um_I.iw[12] ;
 wire \top_I.branch[20].block[9].um_I.iw[13] ;
 wire \top_I.branch[20].block[9].um_I.iw[14] ;
 wire \top_I.branch[20].block[9].um_I.iw[15] ;
 wire \top_I.branch[20].block[9].um_I.iw[16] ;
 wire \top_I.branch[20].block[9].um_I.iw[17] ;
 wire \top_I.branch[20].block[9].um_I.iw[1] ;
 wire \top_I.branch[20].block[9].um_I.iw[2] ;
 wire \top_I.branch[20].block[9].um_I.iw[3] ;
 wire \top_I.branch[20].block[9].um_I.iw[4] ;
 wire \top_I.branch[20].block[9].um_I.iw[5] ;
 wire \top_I.branch[20].block[9].um_I.iw[6] ;
 wire \top_I.branch[20].block[9].um_I.iw[7] ;
 wire \top_I.branch[20].block[9].um_I.iw[8] ;
 wire \top_I.branch[20].block[9].um_I.iw[9] ;
 wire \top_I.branch[20].block[9].um_I.k_zero ;
 wire \top_I.branch[20].block[9].um_I.pg_vdd ;
 wire \top_I.branch[20].l_addr[0] ;
 wire \top_I.branch[20].l_addr[1] ;
 wire \top_I.branch[21].block[0].um_I.ana[0] ;
 wire \top_I.branch[21].block[0].um_I.ana[1] ;
 wire \top_I.branch[21].block[0].um_I.ana[2] ;
 wire \top_I.branch[21].block[0].um_I.ana[3] ;
 wire \top_I.branch[21].block[0].um_I.ana[4] ;
 wire \top_I.branch[21].block[0].um_I.ana[5] ;
 wire \top_I.branch[21].block[0].um_I.ana[6] ;
 wire \top_I.branch[21].block[0].um_I.ana[7] ;
 wire \top_I.branch[21].block[0].um_I.clk ;
 wire \top_I.branch[21].block[0].um_I.ena ;
 wire \top_I.branch[21].block[0].um_I.iw[10] ;
 wire \top_I.branch[21].block[0].um_I.iw[11] ;
 wire \top_I.branch[21].block[0].um_I.iw[12] ;
 wire \top_I.branch[21].block[0].um_I.iw[13] ;
 wire \top_I.branch[21].block[0].um_I.iw[14] ;
 wire \top_I.branch[21].block[0].um_I.iw[15] ;
 wire \top_I.branch[21].block[0].um_I.iw[16] ;
 wire \top_I.branch[21].block[0].um_I.iw[17] ;
 wire \top_I.branch[21].block[0].um_I.iw[1] ;
 wire \top_I.branch[21].block[0].um_I.iw[2] ;
 wire \top_I.branch[21].block[0].um_I.iw[3] ;
 wire \top_I.branch[21].block[0].um_I.iw[4] ;
 wire \top_I.branch[21].block[0].um_I.iw[5] ;
 wire \top_I.branch[21].block[0].um_I.iw[6] ;
 wire \top_I.branch[21].block[0].um_I.iw[7] ;
 wire \top_I.branch[21].block[0].um_I.iw[8] ;
 wire \top_I.branch[21].block[0].um_I.iw[9] ;
 wire \top_I.branch[21].block[0].um_I.k_zero ;
 wire \top_I.branch[21].block[0].um_I.pg_vdd ;
 wire \top_I.branch[21].block[10].um_I.ana[0] ;
 wire \top_I.branch[21].block[10].um_I.ana[1] ;
 wire \top_I.branch[21].block[10].um_I.ana[2] ;
 wire \top_I.branch[21].block[10].um_I.ana[3] ;
 wire \top_I.branch[21].block[10].um_I.ana[4] ;
 wire \top_I.branch[21].block[10].um_I.ana[5] ;
 wire \top_I.branch[21].block[10].um_I.ana[6] ;
 wire \top_I.branch[21].block[10].um_I.ana[7] ;
 wire \top_I.branch[21].block[10].um_I.clk ;
 wire \top_I.branch[21].block[10].um_I.ena ;
 wire \top_I.branch[21].block[10].um_I.iw[10] ;
 wire \top_I.branch[21].block[10].um_I.iw[11] ;
 wire \top_I.branch[21].block[10].um_I.iw[12] ;
 wire \top_I.branch[21].block[10].um_I.iw[13] ;
 wire \top_I.branch[21].block[10].um_I.iw[14] ;
 wire \top_I.branch[21].block[10].um_I.iw[15] ;
 wire \top_I.branch[21].block[10].um_I.iw[16] ;
 wire \top_I.branch[21].block[10].um_I.iw[17] ;
 wire \top_I.branch[21].block[10].um_I.iw[1] ;
 wire \top_I.branch[21].block[10].um_I.iw[2] ;
 wire \top_I.branch[21].block[10].um_I.iw[3] ;
 wire \top_I.branch[21].block[10].um_I.iw[4] ;
 wire \top_I.branch[21].block[10].um_I.iw[5] ;
 wire \top_I.branch[21].block[10].um_I.iw[6] ;
 wire \top_I.branch[21].block[10].um_I.iw[7] ;
 wire \top_I.branch[21].block[10].um_I.iw[8] ;
 wire \top_I.branch[21].block[10].um_I.iw[9] ;
 wire \top_I.branch[21].block[10].um_I.k_zero ;
 wire \top_I.branch[21].block[10].um_I.pg_vdd ;
 wire \top_I.branch[21].block[11].um_I.ana[0] ;
 wire \top_I.branch[21].block[11].um_I.ana[1] ;
 wire \top_I.branch[21].block[11].um_I.ana[2] ;
 wire \top_I.branch[21].block[11].um_I.ana[3] ;
 wire \top_I.branch[21].block[11].um_I.ana[4] ;
 wire \top_I.branch[21].block[11].um_I.ana[5] ;
 wire \top_I.branch[21].block[11].um_I.ana[6] ;
 wire \top_I.branch[21].block[11].um_I.ana[7] ;
 wire \top_I.branch[21].block[11].um_I.clk ;
 wire \top_I.branch[21].block[11].um_I.ena ;
 wire \top_I.branch[21].block[11].um_I.iw[10] ;
 wire \top_I.branch[21].block[11].um_I.iw[11] ;
 wire \top_I.branch[21].block[11].um_I.iw[12] ;
 wire \top_I.branch[21].block[11].um_I.iw[13] ;
 wire \top_I.branch[21].block[11].um_I.iw[14] ;
 wire \top_I.branch[21].block[11].um_I.iw[15] ;
 wire \top_I.branch[21].block[11].um_I.iw[16] ;
 wire \top_I.branch[21].block[11].um_I.iw[17] ;
 wire \top_I.branch[21].block[11].um_I.iw[1] ;
 wire \top_I.branch[21].block[11].um_I.iw[2] ;
 wire \top_I.branch[21].block[11].um_I.iw[3] ;
 wire \top_I.branch[21].block[11].um_I.iw[4] ;
 wire \top_I.branch[21].block[11].um_I.iw[5] ;
 wire \top_I.branch[21].block[11].um_I.iw[6] ;
 wire \top_I.branch[21].block[11].um_I.iw[7] ;
 wire \top_I.branch[21].block[11].um_I.iw[8] ;
 wire \top_I.branch[21].block[11].um_I.iw[9] ;
 wire \top_I.branch[21].block[11].um_I.k_zero ;
 wire \top_I.branch[21].block[11].um_I.pg_vdd ;
 wire \top_I.branch[21].block[12].um_I.ana[0] ;
 wire \top_I.branch[21].block[12].um_I.ana[1] ;
 wire \top_I.branch[21].block[12].um_I.ana[2] ;
 wire \top_I.branch[21].block[12].um_I.ana[3] ;
 wire \top_I.branch[21].block[12].um_I.ana[4] ;
 wire \top_I.branch[21].block[12].um_I.ana[5] ;
 wire \top_I.branch[21].block[12].um_I.ana[6] ;
 wire \top_I.branch[21].block[12].um_I.ana[7] ;
 wire \top_I.branch[21].block[12].um_I.clk ;
 wire \top_I.branch[21].block[12].um_I.ena ;
 wire \top_I.branch[21].block[12].um_I.iw[10] ;
 wire \top_I.branch[21].block[12].um_I.iw[11] ;
 wire \top_I.branch[21].block[12].um_I.iw[12] ;
 wire \top_I.branch[21].block[12].um_I.iw[13] ;
 wire \top_I.branch[21].block[12].um_I.iw[14] ;
 wire \top_I.branch[21].block[12].um_I.iw[15] ;
 wire \top_I.branch[21].block[12].um_I.iw[16] ;
 wire \top_I.branch[21].block[12].um_I.iw[17] ;
 wire \top_I.branch[21].block[12].um_I.iw[1] ;
 wire \top_I.branch[21].block[12].um_I.iw[2] ;
 wire \top_I.branch[21].block[12].um_I.iw[3] ;
 wire \top_I.branch[21].block[12].um_I.iw[4] ;
 wire \top_I.branch[21].block[12].um_I.iw[5] ;
 wire \top_I.branch[21].block[12].um_I.iw[6] ;
 wire \top_I.branch[21].block[12].um_I.iw[7] ;
 wire \top_I.branch[21].block[12].um_I.iw[8] ;
 wire \top_I.branch[21].block[12].um_I.iw[9] ;
 wire \top_I.branch[21].block[12].um_I.k_zero ;
 wire \top_I.branch[21].block[12].um_I.pg_vdd ;
 wire \top_I.branch[21].block[13].um_I.ana[0] ;
 wire \top_I.branch[21].block[13].um_I.ana[1] ;
 wire \top_I.branch[21].block[13].um_I.ana[2] ;
 wire \top_I.branch[21].block[13].um_I.ana[3] ;
 wire \top_I.branch[21].block[13].um_I.ana[4] ;
 wire \top_I.branch[21].block[13].um_I.ana[5] ;
 wire \top_I.branch[21].block[13].um_I.ana[6] ;
 wire \top_I.branch[21].block[13].um_I.ana[7] ;
 wire \top_I.branch[21].block[13].um_I.clk ;
 wire \top_I.branch[21].block[13].um_I.ena ;
 wire \top_I.branch[21].block[13].um_I.iw[10] ;
 wire \top_I.branch[21].block[13].um_I.iw[11] ;
 wire \top_I.branch[21].block[13].um_I.iw[12] ;
 wire \top_I.branch[21].block[13].um_I.iw[13] ;
 wire \top_I.branch[21].block[13].um_I.iw[14] ;
 wire \top_I.branch[21].block[13].um_I.iw[15] ;
 wire \top_I.branch[21].block[13].um_I.iw[16] ;
 wire \top_I.branch[21].block[13].um_I.iw[17] ;
 wire \top_I.branch[21].block[13].um_I.iw[1] ;
 wire \top_I.branch[21].block[13].um_I.iw[2] ;
 wire \top_I.branch[21].block[13].um_I.iw[3] ;
 wire \top_I.branch[21].block[13].um_I.iw[4] ;
 wire \top_I.branch[21].block[13].um_I.iw[5] ;
 wire \top_I.branch[21].block[13].um_I.iw[6] ;
 wire \top_I.branch[21].block[13].um_I.iw[7] ;
 wire \top_I.branch[21].block[13].um_I.iw[8] ;
 wire \top_I.branch[21].block[13].um_I.iw[9] ;
 wire \top_I.branch[21].block[13].um_I.k_zero ;
 wire \top_I.branch[21].block[13].um_I.pg_vdd ;
 wire \top_I.branch[21].block[14].um_I.ana[0] ;
 wire \top_I.branch[21].block[14].um_I.ana[1] ;
 wire \top_I.branch[21].block[14].um_I.ana[2] ;
 wire \top_I.branch[21].block[14].um_I.ana[3] ;
 wire \top_I.branch[21].block[14].um_I.ana[4] ;
 wire \top_I.branch[21].block[14].um_I.ana[5] ;
 wire \top_I.branch[21].block[14].um_I.ana[6] ;
 wire \top_I.branch[21].block[14].um_I.ana[7] ;
 wire \top_I.branch[21].block[14].um_I.clk ;
 wire \top_I.branch[21].block[14].um_I.ena ;
 wire \top_I.branch[21].block[14].um_I.iw[10] ;
 wire \top_I.branch[21].block[14].um_I.iw[11] ;
 wire \top_I.branch[21].block[14].um_I.iw[12] ;
 wire \top_I.branch[21].block[14].um_I.iw[13] ;
 wire \top_I.branch[21].block[14].um_I.iw[14] ;
 wire \top_I.branch[21].block[14].um_I.iw[15] ;
 wire \top_I.branch[21].block[14].um_I.iw[16] ;
 wire \top_I.branch[21].block[14].um_I.iw[17] ;
 wire \top_I.branch[21].block[14].um_I.iw[1] ;
 wire \top_I.branch[21].block[14].um_I.iw[2] ;
 wire \top_I.branch[21].block[14].um_I.iw[3] ;
 wire \top_I.branch[21].block[14].um_I.iw[4] ;
 wire \top_I.branch[21].block[14].um_I.iw[5] ;
 wire \top_I.branch[21].block[14].um_I.iw[6] ;
 wire \top_I.branch[21].block[14].um_I.iw[7] ;
 wire \top_I.branch[21].block[14].um_I.iw[8] ;
 wire \top_I.branch[21].block[14].um_I.iw[9] ;
 wire \top_I.branch[21].block[14].um_I.k_zero ;
 wire \top_I.branch[21].block[14].um_I.pg_vdd ;
 wire \top_I.branch[21].block[15].um_I.ana[0] ;
 wire \top_I.branch[21].block[15].um_I.ana[1] ;
 wire \top_I.branch[21].block[15].um_I.ana[2] ;
 wire \top_I.branch[21].block[15].um_I.ana[3] ;
 wire \top_I.branch[21].block[15].um_I.ana[4] ;
 wire \top_I.branch[21].block[15].um_I.ana[5] ;
 wire \top_I.branch[21].block[15].um_I.ana[6] ;
 wire \top_I.branch[21].block[15].um_I.ana[7] ;
 wire \top_I.branch[21].block[15].um_I.clk ;
 wire \top_I.branch[21].block[15].um_I.ena ;
 wire \top_I.branch[21].block[15].um_I.iw[10] ;
 wire \top_I.branch[21].block[15].um_I.iw[11] ;
 wire \top_I.branch[21].block[15].um_I.iw[12] ;
 wire \top_I.branch[21].block[15].um_I.iw[13] ;
 wire \top_I.branch[21].block[15].um_I.iw[14] ;
 wire \top_I.branch[21].block[15].um_I.iw[15] ;
 wire \top_I.branch[21].block[15].um_I.iw[16] ;
 wire \top_I.branch[21].block[15].um_I.iw[17] ;
 wire \top_I.branch[21].block[15].um_I.iw[1] ;
 wire \top_I.branch[21].block[15].um_I.iw[2] ;
 wire \top_I.branch[21].block[15].um_I.iw[3] ;
 wire \top_I.branch[21].block[15].um_I.iw[4] ;
 wire \top_I.branch[21].block[15].um_I.iw[5] ;
 wire \top_I.branch[21].block[15].um_I.iw[6] ;
 wire \top_I.branch[21].block[15].um_I.iw[7] ;
 wire \top_I.branch[21].block[15].um_I.iw[8] ;
 wire \top_I.branch[21].block[15].um_I.iw[9] ;
 wire \top_I.branch[21].block[15].um_I.k_zero ;
 wire \top_I.branch[21].block[15].um_I.pg_vdd ;
 wire \top_I.branch[21].block[1].um_I.ana[0] ;
 wire \top_I.branch[21].block[1].um_I.ana[1] ;
 wire \top_I.branch[21].block[1].um_I.ana[2] ;
 wire \top_I.branch[21].block[1].um_I.ana[3] ;
 wire \top_I.branch[21].block[1].um_I.ana[4] ;
 wire \top_I.branch[21].block[1].um_I.ana[5] ;
 wire \top_I.branch[21].block[1].um_I.ana[6] ;
 wire \top_I.branch[21].block[1].um_I.ana[7] ;
 wire \top_I.branch[21].block[1].um_I.clk ;
 wire \top_I.branch[21].block[1].um_I.ena ;
 wire \top_I.branch[21].block[1].um_I.iw[10] ;
 wire \top_I.branch[21].block[1].um_I.iw[11] ;
 wire \top_I.branch[21].block[1].um_I.iw[12] ;
 wire \top_I.branch[21].block[1].um_I.iw[13] ;
 wire \top_I.branch[21].block[1].um_I.iw[14] ;
 wire \top_I.branch[21].block[1].um_I.iw[15] ;
 wire \top_I.branch[21].block[1].um_I.iw[16] ;
 wire \top_I.branch[21].block[1].um_I.iw[17] ;
 wire \top_I.branch[21].block[1].um_I.iw[1] ;
 wire \top_I.branch[21].block[1].um_I.iw[2] ;
 wire \top_I.branch[21].block[1].um_I.iw[3] ;
 wire \top_I.branch[21].block[1].um_I.iw[4] ;
 wire \top_I.branch[21].block[1].um_I.iw[5] ;
 wire \top_I.branch[21].block[1].um_I.iw[6] ;
 wire \top_I.branch[21].block[1].um_I.iw[7] ;
 wire \top_I.branch[21].block[1].um_I.iw[8] ;
 wire \top_I.branch[21].block[1].um_I.iw[9] ;
 wire \top_I.branch[21].block[1].um_I.k_zero ;
 wire \top_I.branch[21].block[1].um_I.pg_vdd ;
 wire \top_I.branch[21].block[2].um_I.ana[0] ;
 wire \top_I.branch[21].block[2].um_I.ana[1] ;
 wire \top_I.branch[21].block[2].um_I.ana[2] ;
 wire \top_I.branch[21].block[2].um_I.ana[3] ;
 wire \top_I.branch[21].block[2].um_I.ana[4] ;
 wire \top_I.branch[21].block[2].um_I.ana[5] ;
 wire \top_I.branch[21].block[2].um_I.ana[6] ;
 wire \top_I.branch[21].block[2].um_I.ana[7] ;
 wire \top_I.branch[21].block[2].um_I.clk ;
 wire \top_I.branch[21].block[2].um_I.ena ;
 wire \top_I.branch[21].block[2].um_I.iw[10] ;
 wire \top_I.branch[21].block[2].um_I.iw[11] ;
 wire \top_I.branch[21].block[2].um_I.iw[12] ;
 wire \top_I.branch[21].block[2].um_I.iw[13] ;
 wire \top_I.branch[21].block[2].um_I.iw[14] ;
 wire \top_I.branch[21].block[2].um_I.iw[15] ;
 wire \top_I.branch[21].block[2].um_I.iw[16] ;
 wire \top_I.branch[21].block[2].um_I.iw[17] ;
 wire \top_I.branch[21].block[2].um_I.iw[1] ;
 wire \top_I.branch[21].block[2].um_I.iw[2] ;
 wire \top_I.branch[21].block[2].um_I.iw[3] ;
 wire \top_I.branch[21].block[2].um_I.iw[4] ;
 wire \top_I.branch[21].block[2].um_I.iw[5] ;
 wire \top_I.branch[21].block[2].um_I.iw[6] ;
 wire \top_I.branch[21].block[2].um_I.iw[7] ;
 wire \top_I.branch[21].block[2].um_I.iw[8] ;
 wire \top_I.branch[21].block[2].um_I.iw[9] ;
 wire \top_I.branch[21].block[2].um_I.k_zero ;
 wire \top_I.branch[21].block[2].um_I.pg_vdd ;
 wire \top_I.branch[21].block[3].um_I.ana[0] ;
 wire \top_I.branch[21].block[3].um_I.ana[1] ;
 wire \top_I.branch[21].block[3].um_I.ana[2] ;
 wire \top_I.branch[21].block[3].um_I.ana[3] ;
 wire \top_I.branch[21].block[3].um_I.ana[4] ;
 wire \top_I.branch[21].block[3].um_I.ana[5] ;
 wire \top_I.branch[21].block[3].um_I.ana[6] ;
 wire \top_I.branch[21].block[3].um_I.ana[7] ;
 wire \top_I.branch[21].block[3].um_I.clk ;
 wire \top_I.branch[21].block[3].um_I.ena ;
 wire \top_I.branch[21].block[3].um_I.iw[10] ;
 wire \top_I.branch[21].block[3].um_I.iw[11] ;
 wire \top_I.branch[21].block[3].um_I.iw[12] ;
 wire \top_I.branch[21].block[3].um_I.iw[13] ;
 wire \top_I.branch[21].block[3].um_I.iw[14] ;
 wire \top_I.branch[21].block[3].um_I.iw[15] ;
 wire \top_I.branch[21].block[3].um_I.iw[16] ;
 wire \top_I.branch[21].block[3].um_I.iw[17] ;
 wire \top_I.branch[21].block[3].um_I.iw[1] ;
 wire \top_I.branch[21].block[3].um_I.iw[2] ;
 wire \top_I.branch[21].block[3].um_I.iw[3] ;
 wire \top_I.branch[21].block[3].um_I.iw[4] ;
 wire \top_I.branch[21].block[3].um_I.iw[5] ;
 wire \top_I.branch[21].block[3].um_I.iw[6] ;
 wire \top_I.branch[21].block[3].um_I.iw[7] ;
 wire \top_I.branch[21].block[3].um_I.iw[8] ;
 wire \top_I.branch[21].block[3].um_I.iw[9] ;
 wire \top_I.branch[21].block[3].um_I.k_zero ;
 wire \top_I.branch[21].block[3].um_I.pg_vdd ;
 wire \top_I.branch[21].block[4].um_I.ana[0] ;
 wire \top_I.branch[21].block[4].um_I.ana[1] ;
 wire \top_I.branch[21].block[4].um_I.ana[2] ;
 wire \top_I.branch[21].block[4].um_I.ana[3] ;
 wire \top_I.branch[21].block[4].um_I.ana[4] ;
 wire \top_I.branch[21].block[4].um_I.ana[5] ;
 wire \top_I.branch[21].block[4].um_I.ana[6] ;
 wire \top_I.branch[21].block[4].um_I.ana[7] ;
 wire \top_I.branch[21].block[4].um_I.clk ;
 wire \top_I.branch[21].block[4].um_I.ena ;
 wire \top_I.branch[21].block[4].um_I.iw[10] ;
 wire \top_I.branch[21].block[4].um_I.iw[11] ;
 wire \top_I.branch[21].block[4].um_I.iw[12] ;
 wire \top_I.branch[21].block[4].um_I.iw[13] ;
 wire \top_I.branch[21].block[4].um_I.iw[14] ;
 wire \top_I.branch[21].block[4].um_I.iw[15] ;
 wire \top_I.branch[21].block[4].um_I.iw[16] ;
 wire \top_I.branch[21].block[4].um_I.iw[17] ;
 wire \top_I.branch[21].block[4].um_I.iw[1] ;
 wire \top_I.branch[21].block[4].um_I.iw[2] ;
 wire \top_I.branch[21].block[4].um_I.iw[3] ;
 wire \top_I.branch[21].block[4].um_I.iw[4] ;
 wire \top_I.branch[21].block[4].um_I.iw[5] ;
 wire \top_I.branch[21].block[4].um_I.iw[6] ;
 wire \top_I.branch[21].block[4].um_I.iw[7] ;
 wire \top_I.branch[21].block[4].um_I.iw[8] ;
 wire \top_I.branch[21].block[4].um_I.iw[9] ;
 wire \top_I.branch[21].block[4].um_I.k_zero ;
 wire \top_I.branch[21].block[4].um_I.pg_vdd ;
 wire \top_I.branch[21].block[5].um_I.ana[0] ;
 wire \top_I.branch[21].block[5].um_I.ana[1] ;
 wire \top_I.branch[21].block[5].um_I.ana[2] ;
 wire \top_I.branch[21].block[5].um_I.ana[3] ;
 wire \top_I.branch[21].block[5].um_I.ana[4] ;
 wire \top_I.branch[21].block[5].um_I.ana[5] ;
 wire \top_I.branch[21].block[5].um_I.ana[6] ;
 wire \top_I.branch[21].block[5].um_I.ana[7] ;
 wire \top_I.branch[21].block[5].um_I.clk ;
 wire \top_I.branch[21].block[5].um_I.ena ;
 wire \top_I.branch[21].block[5].um_I.iw[10] ;
 wire \top_I.branch[21].block[5].um_I.iw[11] ;
 wire \top_I.branch[21].block[5].um_I.iw[12] ;
 wire \top_I.branch[21].block[5].um_I.iw[13] ;
 wire \top_I.branch[21].block[5].um_I.iw[14] ;
 wire \top_I.branch[21].block[5].um_I.iw[15] ;
 wire \top_I.branch[21].block[5].um_I.iw[16] ;
 wire \top_I.branch[21].block[5].um_I.iw[17] ;
 wire \top_I.branch[21].block[5].um_I.iw[1] ;
 wire \top_I.branch[21].block[5].um_I.iw[2] ;
 wire \top_I.branch[21].block[5].um_I.iw[3] ;
 wire \top_I.branch[21].block[5].um_I.iw[4] ;
 wire \top_I.branch[21].block[5].um_I.iw[5] ;
 wire \top_I.branch[21].block[5].um_I.iw[6] ;
 wire \top_I.branch[21].block[5].um_I.iw[7] ;
 wire \top_I.branch[21].block[5].um_I.iw[8] ;
 wire \top_I.branch[21].block[5].um_I.iw[9] ;
 wire \top_I.branch[21].block[5].um_I.k_zero ;
 wire \top_I.branch[21].block[5].um_I.pg_vdd ;
 wire \top_I.branch[21].block[6].um_I.ana[0] ;
 wire \top_I.branch[21].block[6].um_I.ana[1] ;
 wire \top_I.branch[21].block[6].um_I.ana[2] ;
 wire \top_I.branch[21].block[6].um_I.ana[3] ;
 wire \top_I.branch[21].block[6].um_I.ana[4] ;
 wire \top_I.branch[21].block[6].um_I.ana[5] ;
 wire \top_I.branch[21].block[6].um_I.ana[6] ;
 wire \top_I.branch[21].block[6].um_I.ana[7] ;
 wire \top_I.branch[21].block[6].um_I.clk ;
 wire \top_I.branch[21].block[6].um_I.ena ;
 wire \top_I.branch[21].block[6].um_I.iw[10] ;
 wire \top_I.branch[21].block[6].um_I.iw[11] ;
 wire \top_I.branch[21].block[6].um_I.iw[12] ;
 wire \top_I.branch[21].block[6].um_I.iw[13] ;
 wire \top_I.branch[21].block[6].um_I.iw[14] ;
 wire \top_I.branch[21].block[6].um_I.iw[15] ;
 wire \top_I.branch[21].block[6].um_I.iw[16] ;
 wire \top_I.branch[21].block[6].um_I.iw[17] ;
 wire \top_I.branch[21].block[6].um_I.iw[1] ;
 wire \top_I.branch[21].block[6].um_I.iw[2] ;
 wire \top_I.branch[21].block[6].um_I.iw[3] ;
 wire \top_I.branch[21].block[6].um_I.iw[4] ;
 wire \top_I.branch[21].block[6].um_I.iw[5] ;
 wire \top_I.branch[21].block[6].um_I.iw[6] ;
 wire \top_I.branch[21].block[6].um_I.iw[7] ;
 wire \top_I.branch[21].block[6].um_I.iw[8] ;
 wire \top_I.branch[21].block[6].um_I.iw[9] ;
 wire \top_I.branch[21].block[6].um_I.k_zero ;
 wire \top_I.branch[21].block[6].um_I.pg_vdd ;
 wire \top_I.branch[21].block[7].um_I.ana[0] ;
 wire \top_I.branch[21].block[7].um_I.ana[1] ;
 wire \top_I.branch[21].block[7].um_I.ana[2] ;
 wire \top_I.branch[21].block[7].um_I.ana[3] ;
 wire \top_I.branch[21].block[7].um_I.ana[4] ;
 wire \top_I.branch[21].block[7].um_I.ana[5] ;
 wire \top_I.branch[21].block[7].um_I.ana[6] ;
 wire \top_I.branch[21].block[7].um_I.ana[7] ;
 wire \top_I.branch[21].block[7].um_I.clk ;
 wire \top_I.branch[21].block[7].um_I.ena ;
 wire \top_I.branch[21].block[7].um_I.iw[10] ;
 wire \top_I.branch[21].block[7].um_I.iw[11] ;
 wire \top_I.branch[21].block[7].um_I.iw[12] ;
 wire \top_I.branch[21].block[7].um_I.iw[13] ;
 wire \top_I.branch[21].block[7].um_I.iw[14] ;
 wire \top_I.branch[21].block[7].um_I.iw[15] ;
 wire \top_I.branch[21].block[7].um_I.iw[16] ;
 wire \top_I.branch[21].block[7].um_I.iw[17] ;
 wire \top_I.branch[21].block[7].um_I.iw[1] ;
 wire \top_I.branch[21].block[7].um_I.iw[2] ;
 wire \top_I.branch[21].block[7].um_I.iw[3] ;
 wire \top_I.branch[21].block[7].um_I.iw[4] ;
 wire \top_I.branch[21].block[7].um_I.iw[5] ;
 wire \top_I.branch[21].block[7].um_I.iw[6] ;
 wire \top_I.branch[21].block[7].um_I.iw[7] ;
 wire \top_I.branch[21].block[7].um_I.iw[8] ;
 wire \top_I.branch[21].block[7].um_I.iw[9] ;
 wire \top_I.branch[21].block[7].um_I.k_zero ;
 wire \top_I.branch[21].block[7].um_I.pg_vdd ;
 wire \top_I.branch[21].block[8].um_I.ana[0] ;
 wire \top_I.branch[21].block[8].um_I.ana[1] ;
 wire \top_I.branch[21].block[8].um_I.ana[2] ;
 wire \top_I.branch[21].block[8].um_I.ana[3] ;
 wire \top_I.branch[21].block[8].um_I.ana[4] ;
 wire \top_I.branch[21].block[8].um_I.ana[5] ;
 wire \top_I.branch[21].block[8].um_I.ana[6] ;
 wire \top_I.branch[21].block[8].um_I.ana[7] ;
 wire \top_I.branch[21].block[8].um_I.clk ;
 wire \top_I.branch[21].block[8].um_I.ena ;
 wire \top_I.branch[21].block[8].um_I.iw[10] ;
 wire \top_I.branch[21].block[8].um_I.iw[11] ;
 wire \top_I.branch[21].block[8].um_I.iw[12] ;
 wire \top_I.branch[21].block[8].um_I.iw[13] ;
 wire \top_I.branch[21].block[8].um_I.iw[14] ;
 wire \top_I.branch[21].block[8].um_I.iw[15] ;
 wire \top_I.branch[21].block[8].um_I.iw[16] ;
 wire \top_I.branch[21].block[8].um_I.iw[17] ;
 wire \top_I.branch[21].block[8].um_I.iw[1] ;
 wire \top_I.branch[21].block[8].um_I.iw[2] ;
 wire \top_I.branch[21].block[8].um_I.iw[3] ;
 wire \top_I.branch[21].block[8].um_I.iw[4] ;
 wire \top_I.branch[21].block[8].um_I.iw[5] ;
 wire \top_I.branch[21].block[8].um_I.iw[6] ;
 wire \top_I.branch[21].block[8].um_I.iw[7] ;
 wire \top_I.branch[21].block[8].um_I.iw[8] ;
 wire \top_I.branch[21].block[8].um_I.iw[9] ;
 wire \top_I.branch[21].block[8].um_I.k_zero ;
 wire \top_I.branch[21].block[8].um_I.pg_vdd ;
 wire \top_I.branch[21].block[9].um_I.ana[0] ;
 wire \top_I.branch[21].block[9].um_I.ana[1] ;
 wire \top_I.branch[21].block[9].um_I.ana[2] ;
 wire \top_I.branch[21].block[9].um_I.ana[3] ;
 wire \top_I.branch[21].block[9].um_I.ana[4] ;
 wire \top_I.branch[21].block[9].um_I.ana[5] ;
 wire \top_I.branch[21].block[9].um_I.ana[6] ;
 wire \top_I.branch[21].block[9].um_I.ana[7] ;
 wire \top_I.branch[21].block[9].um_I.clk ;
 wire \top_I.branch[21].block[9].um_I.ena ;
 wire \top_I.branch[21].block[9].um_I.iw[10] ;
 wire \top_I.branch[21].block[9].um_I.iw[11] ;
 wire \top_I.branch[21].block[9].um_I.iw[12] ;
 wire \top_I.branch[21].block[9].um_I.iw[13] ;
 wire \top_I.branch[21].block[9].um_I.iw[14] ;
 wire \top_I.branch[21].block[9].um_I.iw[15] ;
 wire \top_I.branch[21].block[9].um_I.iw[16] ;
 wire \top_I.branch[21].block[9].um_I.iw[17] ;
 wire \top_I.branch[21].block[9].um_I.iw[1] ;
 wire \top_I.branch[21].block[9].um_I.iw[2] ;
 wire \top_I.branch[21].block[9].um_I.iw[3] ;
 wire \top_I.branch[21].block[9].um_I.iw[4] ;
 wire \top_I.branch[21].block[9].um_I.iw[5] ;
 wire \top_I.branch[21].block[9].um_I.iw[6] ;
 wire \top_I.branch[21].block[9].um_I.iw[7] ;
 wire \top_I.branch[21].block[9].um_I.iw[8] ;
 wire \top_I.branch[21].block[9].um_I.iw[9] ;
 wire \top_I.branch[21].block[9].um_I.k_zero ;
 wire \top_I.branch[21].block[9].um_I.pg_vdd ;
 wire \top_I.branch[21].l_addr[0] ;
 wire \top_I.branch[21].l_addr[1] ;
 wire \top_I.branch[22].block[0].um_I.ana[0] ;
 wire \top_I.branch[22].block[0].um_I.ana[1] ;
 wire \top_I.branch[22].block[0].um_I.ana[2] ;
 wire \top_I.branch[22].block[0].um_I.ana[3] ;
 wire \top_I.branch[22].block[0].um_I.ana[4] ;
 wire \top_I.branch[22].block[0].um_I.ana[5] ;
 wire \top_I.branch[22].block[0].um_I.ana[6] ;
 wire \top_I.branch[22].block[0].um_I.ana[7] ;
 wire \top_I.branch[22].block[0].um_I.clk ;
 wire \top_I.branch[22].block[0].um_I.ena ;
 wire \top_I.branch[22].block[0].um_I.iw[10] ;
 wire \top_I.branch[22].block[0].um_I.iw[11] ;
 wire \top_I.branch[22].block[0].um_I.iw[12] ;
 wire \top_I.branch[22].block[0].um_I.iw[13] ;
 wire \top_I.branch[22].block[0].um_I.iw[14] ;
 wire \top_I.branch[22].block[0].um_I.iw[15] ;
 wire \top_I.branch[22].block[0].um_I.iw[16] ;
 wire \top_I.branch[22].block[0].um_I.iw[17] ;
 wire \top_I.branch[22].block[0].um_I.iw[1] ;
 wire \top_I.branch[22].block[0].um_I.iw[2] ;
 wire \top_I.branch[22].block[0].um_I.iw[3] ;
 wire \top_I.branch[22].block[0].um_I.iw[4] ;
 wire \top_I.branch[22].block[0].um_I.iw[5] ;
 wire \top_I.branch[22].block[0].um_I.iw[6] ;
 wire \top_I.branch[22].block[0].um_I.iw[7] ;
 wire \top_I.branch[22].block[0].um_I.iw[8] ;
 wire \top_I.branch[22].block[0].um_I.iw[9] ;
 wire \top_I.branch[22].block[0].um_I.k_zero ;
 wire \top_I.branch[22].block[0].um_I.pg_vdd ;
 wire \top_I.branch[22].block[10].um_I.ana[0] ;
 wire \top_I.branch[22].block[10].um_I.ana[1] ;
 wire \top_I.branch[22].block[10].um_I.ana[2] ;
 wire \top_I.branch[22].block[10].um_I.ana[3] ;
 wire \top_I.branch[22].block[10].um_I.ana[4] ;
 wire \top_I.branch[22].block[10].um_I.ana[5] ;
 wire \top_I.branch[22].block[10].um_I.ana[6] ;
 wire \top_I.branch[22].block[10].um_I.ana[7] ;
 wire \top_I.branch[22].block[10].um_I.clk ;
 wire \top_I.branch[22].block[10].um_I.ena ;
 wire \top_I.branch[22].block[10].um_I.iw[10] ;
 wire \top_I.branch[22].block[10].um_I.iw[11] ;
 wire \top_I.branch[22].block[10].um_I.iw[12] ;
 wire \top_I.branch[22].block[10].um_I.iw[13] ;
 wire \top_I.branch[22].block[10].um_I.iw[14] ;
 wire \top_I.branch[22].block[10].um_I.iw[15] ;
 wire \top_I.branch[22].block[10].um_I.iw[16] ;
 wire \top_I.branch[22].block[10].um_I.iw[17] ;
 wire \top_I.branch[22].block[10].um_I.iw[1] ;
 wire \top_I.branch[22].block[10].um_I.iw[2] ;
 wire \top_I.branch[22].block[10].um_I.iw[3] ;
 wire \top_I.branch[22].block[10].um_I.iw[4] ;
 wire \top_I.branch[22].block[10].um_I.iw[5] ;
 wire \top_I.branch[22].block[10].um_I.iw[6] ;
 wire \top_I.branch[22].block[10].um_I.iw[7] ;
 wire \top_I.branch[22].block[10].um_I.iw[8] ;
 wire \top_I.branch[22].block[10].um_I.iw[9] ;
 wire \top_I.branch[22].block[10].um_I.k_zero ;
 wire \top_I.branch[22].block[10].um_I.pg_vdd ;
 wire \top_I.branch[22].block[11].um_I.ana[0] ;
 wire \top_I.branch[22].block[11].um_I.ana[1] ;
 wire \top_I.branch[22].block[11].um_I.ana[2] ;
 wire \top_I.branch[22].block[11].um_I.ana[3] ;
 wire \top_I.branch[22].block[11].um_I.ana[4] ;
 wire \top_I.branch[22].block[11].um_I.ana[5] ;
 wire \top_I.branch[22].block[11].um_I.ana[6] ;
 wire \top_I.branch[22].block[11].um_I.ana[7] ;
 wire \top_I.branch[22].block[11].um_I.clk ;
 wire \top_I.branch[22].block[11].um_I.ena ;
 wire \top_I.branch[22].block[11].um_I.iw[10] ;
 wire \top_I.branch[22].block[11].um_I.iw[11] ;
 wire \top_I.branch[22].block[11].um_I.iw[12] ;
 wire \top_I.branch[22].block[11].um_I.iw[13] ;
 wire \top_I.branch[22].block[11].um_I.iw[14] ;
 wire \top_I.branch[22].block[11].um_I.iw[15] ;
 wire \top_I.branch[22].block[11].um_I.iw[16] ;
 wire \top_I.branch[22].block[11].um_I.iw[17] ;
 wire \top_I.branch[22].block[11].um_I.iw[1] ;
 wire \top_I.branch[22].block[11].um_I.iw[2] ;
 wire \top_I.branch[22].block[11].um_I.iw[3] ;
 wire \top_I.branch[22].block[11].um_I.iw[4] ;
 wire \top_I.branch[22].block[11].um_I.iw[5] ;
 wire \top_I.branch[22].block[11].um_I.iw[6] ;
 wire \top_I.branch[22].block[11].um_I.iw[7] ;
 wire \top_I.branch[22].block[11].um_I.iw[8] ;
 wire \top_I.branch[22].block[11].um_I.iw[9] ;
 wire \top_I.branch[22].block[11].um_I.k_zero ;
 wire \top_I.branch[22].block[11].um_I.pg_vdd ;
 wire \top_I.branch[22].block[12].um_I.ana[0] ;
 wire \top_I.branch[22].block[12].um_I.ana[1] ;
 wire \top_I.branch[22].block[12].um_I.ana[2] ;
 wire \top_I.branch[22].block[12].um_I.ana[3] ;
 wire \top_I.branch[22].block[12].um_I.ana[4] ;
 wire \top_I.branch[22].block[12].um_I.ana[5] ;
 wire \top_I.branch[22].block[12].um_I.ana[6] ;
 wire \top_I.branch[22].block[12].um_I.ana[7] ;
 wire \top_I.branch[22].block[12].um_I.clk ;
 wire \top_I.branch[22].block[12].um_I.ena ;
 wire \top_I.branch[22].block[12].um_I.iw[10] ;
 wire \top_I.branch[22].block[12].um_I.iw[11] ;
 wire \top_I.branch[22].block[12].um_I.iw[12] ;
 wire \top_I.branch[22].block[12].um_I.iw[13] ;
 wire \top_I.branch[22].block[12].um_I.iw[14] ;
 wire \top_I.branch[22].block[12].um_I.iw[15] ;
 wire \top_I.branch[22].block[12].um_I.iw[16] ;
 wire \top_I.branch[22].block[12].um_I.iw[17] ;
 wire \top_I.branch[22].block[12].um_I.iw[1] ;
 wire \top_I.branch[22].block[12].um_I.iw[2] ;
 wire \top_I.branch[22].block[12].um_I.iw[3] ;
 wire \top_I.branch[22].block[12].um_I.iw[4] ;
 wire \top_I.branch[22].block[12].um_I.iw[5] ;
 wire \top_I.branch[22].block[12].um_I.iw[6] ;
 wire \top_I.branch[22].block[12].um_I.iw[7] ;
 wire \top_I.branch[22].block[12].um_I.iw[8] ;
 wire \top_I.branch[22].block[12].um_I.iw[9] ;
 wire \top_I.branch[22].block[12].um_I.k_zero ;
 wire \top_I.branch[22].block[12].um_I.pg_vdd ;
 wire \top_I.branch[22].block[13].um_I.ana[0] ;
 wire \top_I.branch[22].block[13].um_I.ana[1] ;
 wire \top_I.branch[22].block[13].um_I.ana[2] ;
 wire \top_I.branch[22].block[13].um_I.ana[3] ;
 wire \top_I.branch[22].block[13].um_I.ana[4] ;
 wire \top_I.branch[22].block[13].um_I.ana[5] ;
 wire \top_I.branch[22].block[13].um_I.ana[6] ;
 wire \top_I.branch[22].block[13].um_I.ana[7] ;
 wire \top_I.branch[22].block[13].um_I.clk ;
 wire \top_I.branch[22].block[13].um_I.ena ;
 wire \top_I.branch[22].block[13].um_I.iw[10] ;
 wire \top_I.branch[22].block[13].um_I.iw[11] ;
 wire \top_I.branch[22].block[13].um_I.iw[12] ;
 wire \top_I.branch[22].block[13].um_I.iw[13] ;
 wire \top_I.branch[22].block[13].um_I.iw[14] ;
 wire \top_I.branch[22].block[13].um_I.iw[15] ;
 wire \top_I.branch[22].block[13].um_I.iw[16] ;
 wire \top_I.branch[22].block[13].um_I.iw[17] ;
 wire \top_I.branch[22].block[13].um_I.iw[1] ;
 wire \top_I.branch[22].block[13].um_I.iw[2] ;
 wire \top_I.branch[22].block[13].um_I.iw[3] ;
 wire \top_I.branch[22].block[13].um_I.iw[4] ;
 wire \top_I.branch[22].block[13].um_I.iw[5] ;
 wire \top_I.branch[22].block[13].um_I.iw[6] ;
 wire \top_I.branch[22].block[13].um_I.iw[7] ;
 wire \top_I.branch[22].block[13].um_I.iw[8] ;
 wire \top_I.branch[22].block[13].um_I.iw[9] ;
 wire \top_I.branch[22].block[13].um_I.k_zero ;
 wire \top_I.branch[22].block[13].um_I.pg_vdd ;
 wire \top_I.branch[22].block[14].um_I.ana[0] ;
 wire \top_I.branch[22].block[14].um_I.ana[1] ;
 wire \top_I.branch[22].block[14].um_I.ana[2] ;
 wire \top_I.branch[22].block[14].um_I.ana[3] ;
 wire \top_I.branch[22].block[14].um_I.ana[4] ;
 wire \top_I.branch[22].block[14].um_I.ana[5] ;
 wire \top_I.branch[22].block[14].um_I.ana[6] ;
 wire \top_I.branch[22].block[14].um_I.ana[7] ;
 wire \top_I.branch[22].block[14].um_I.clk ;
 wire \top_I.branch[22].block[14].um_I.ena ;
 wire \top_I.branch[22].block[14].um_I.iw[10] ;
 wire \top_I.branch[22].block[14].um_I.iw[11] ;
 wire \top_I.branch[22].block[14].um_I.iw[12] ;
 wire \top_I.branch[22].block[14].um_I.iw[13] ;
 wire \top_I.branch[22].block[14].um_I.iw[14] ;
 wire \top_I.branch[22].block[14].um_I.iw[15] ;
 wire \top_I.branch[22].block[14].um_I.iw[16] ;
 wire \top_I.branch[22].block[14].um_I.iw[17] ;
 wire \top_I.branch[22].block[14].um_I.iw[1] ;
 wire \top_I.branch[22].block[14].um_I.iw[2] ;
 wire \top_I.branch[22].block[14].um_I.iw[3] ;
 wire \top_I.branch[22].block[14].um_I.iw[4] ;
 wire \top_I.branch[22].block[14].um_I.iw[5] ;
 wire \top_I.branch[22].block[14].um_I.iw[6] ;
 wire \top_I.branch[22].block[14].um_I.iw[7] ;
 wire \top_I.branch[22].block[14].um_I.iw[8] ;
 wire \top_I.branch[22].block[14].um_I.iw[9] ;
 wire \top_I.branch[22].block[14].um_I.k_zero ;
 wire \top_I.branch[22].block[14].um_I.pg_vdd ;
 wire \top_I.branch[22].block[15].um_I.ana[0] ;
 wire \top_I.branch[22].block[15].um_I.ana[1] ;
 wire \top_I.branch[22].block[15].um_I.ana[2] ;
 wire \top_I.branch[22].block[15].um_I.ana[3] ;
 wire \top_I.branch[22].block[15].um_I.ana[4] ;
 wire \top_I.branch[22].block[15].um_I.ana[5] ;
 wire \top_I.branch[22].block[15].um_I.ana[6] ;
 wire \top_I.branch[22].block[15].um_I.ana[7] ;
 wire \top_I.branch[22].block[15].um_I.clk ;
 wire \top_I.branch[22].block[15].um_I.ena ;
 wire \top_I.branch[22].block[15].um_I.iw[10] ;
 wire \top_I.branch[22].block[15].um_I.iw[11] ;
 wire \top_I.branch[22].block[15].um_I.iw[12] ;
 wire \top_I.branch[22].block[15].um_I.iw[13] ;
 wire \top_I.branch[22].block[15].um_I.iw[14] ;
 wire \top_I.branch[22].block[15].um_I.iw[15] ;
 wire \top_I.branch[22].block[15].um_I.iw[16] ;
 wire \top_I.branch[22].block[15].um_I.iw[17] ;
 wire \top_I.branch[22].block[15].um_I.iw[1] ;
 wire \top_I.branch[22].block[15].um_I.iw[2] ;
 wire \top_I.branch[22].block[15].um_I.iw[3] ;
 wire \top_I.branch[22].block[15].um_I.iw[4] ;
 wire \top_I.branch[22].block[15].um_I.iw[5] ;
 wire \top_I.branch[22].block[15].um_I.iw[6] ;
 wire \top_I.branch[22].block[15].um_I.iw[7] ;
 wire \top_I.branch[22].block[15].um_I.iw[8] ;
 wire \top_I.branch[22].block[15].um_I.iw[9] ;
 wire \top_I.branch[22].block[15].um_I.k_zero ;
 wire \top_I.branch[22].block[15].um_I.pg_vdd ;
 wire \top_I.branch[22].block[1].um_I.ana[0] ;
 wire \top_I.branch[22].block[1].um_I.ana[1] ;
 wire \top_I.branch[22].block[1].um_I.ana[2] ;
 wire \top_I.branch[22].block[1].um_I.ana[3] ;
 wire \top_I.branch[22].block[1].um_I.ana[4] ;
 wire \top_I.branch[22].block[1].um_I.ana[5] ;
 wire \top_I.branch[22].block[1].um_I.ana[6] ;
 wire \top_I.branch[22].block[1].um_I.ana[7] ;
 wire \top_I.branch[22].block[1].um_I.clk ;
 wire \top_I.branch[22].block[1].um_I.ena ;
 wire \top_I.branch[22].block[1].um_I.iw[10] ;
 wire \top_I.branch[22].block[1].um_I.iw[11] ;
 wire \top_I.branch[22].block[1].um_I.iw[12] ;
 wire \top_I.branch[22].block[1].um_I.iw[13] ;
 wire \top_I.branch[22].block[1].um_I.iw[14] ;
 wire \top_I.branch[22].block[1].um_I.iw[15] ;
 wire \top_I.branch[22].block[1].um_I.iw[16] ;
 wire \top_I.branch[22].block[1].um_I.iw[17] ;
 wire \top_I.branch[22].block[1].um_I.iw[1] ;
 wire \top_I.branch[22].block[1].um_I.iw[2] ;
 wire \top_I.branch[22].block[1].um_I.iw[3] ;
 wire \top_I.branch[22].block[1].um_I.iw[4] ;
 wire \top_I.branch[22].block[1].um_I.iw[5] ;
 wire \top_I.branch[22].block[1].um_I.iw[6] ;
 wire \top_I.branch[22].block[1].um_I.iw[7] ;
 wire \top_I.branch[22].block[1].um_I.iw[8] ;
 wire \top_I.branch[22].block[1].um_I.iw[9] ;
 wire \top_I.branch[22].block[1].um_I.k_zero ;
 wire \top_I.branch[22].block[1].um_I.pg_vdd ;
 wire \top_I.branch[22].block[2].um_I.ana[0] ;
 wire \top_I.branch[22].block[2].um_I.ana[1] ;
 wire \top_I.branch[22].block[2].um_I.ana[2] ;
 wire \top_I.branch[22].block[2].um_I.ana[3] ;
 wire \top_I.branch[22].block[2].um_I.ana[4] ;
 wire \top_I.branch[22].block[2].um_I.ana[5] ;
 wire \top_I.branch[22].block[2].um_I.ana[6] ;
 wire \top_I.branch[22].block[2].um_I.ana[7] ;
 wire \top_I.branch[22].block[2].um_I.clk ;
 wire \top_I.branch[22].block[2].um_I.ena ;
 wire \top_I.branch[22].block[2].um_I.iw[10] ;
 wire \top_I.branch[22].block[2].um_I.iw[11] ;
 wire \top_I.branch[22].block[2].um_I.iw[12] ;
 wire \top_I.branch[22].block[2].um_I.iw[13] ;
 wire \top_I.branch[22].block[2].um_I.iw[14] ;
 wire \top_I.branch[22].block[2].um_I.iw[15] ;
 wire \top_I.branch[22].block[2].um_I.iw[16] ;
 wire \top_I.branch[22].block[2].um_I.iw[17] ;
 wire \top_I.branch[22].block[2].um_I.iw[1] ;
 wire \top_I.branch[22].block[2].um_I.iw[2] ;
 wire \top_I.branch[22].block[2].um_I.iw[3] ;
 wire \top_I.branch[22].block[2].um_I.iw[4] ;
 wire \top_I.branch[22].block[2].um_I.iw[5] ;
 wire \top_I.branch[22].block[2].um_I.iw[6] ;
 wire \top_I.branch[22].block[2].um_I.iw[7] ;
 wire \top_I.branch[22].block[2].um_I.iw[8] ;
 wire \top_I.branch[22].block[2].um_I.iw[9] ;
 wire \top_I.branch[22].block[2].um_I.k_zero ;
 wire \top_I.branch[22].block[2].um_I.pg_vdd ;
 wire \top_I.branch[22].block[3].um_I.ana[0] ;
 wire \top_I.branch[22].block[3].um_I.ana[1] ;
 wire \top_I.branch[22].block[3].um_I.ana[2] ;
 wire \top_I.branch[22].block[3].um_I.ana[3] ;
 wire \top_I.branch[22].block[3].um_I.ana[4] ;
 wire \top_I.branch[22].block[3].um_I.ana[5] ;
 wire \top_I.branch[22].block[3].um_I.ana[6] ;
 wire \top_I.branch[22].block[3].um_I.ana[7] ;
 wire \top_I.branch[22].block[3].um_I.clk ;
 wire \top_I.branch[22].block[3].um_I.ena ;
 wire \top_I.branch[22].block[3].um_I.iw[10] ;
 wire \top_I.branch[22].block[3].um_I.iw[11] ;
 wire \top_I.branch[22].block[3].um_I.iw[12] ;
 wire \top_I.branch[22].block[3].um_I.iw[13] ;
 wire \top_I.branch[22].block[3].um_I.iw[14] ;
 wire \top_I.branch[22].block[3].um_I.iw[15] ;
 wire \top_I.branch[22].block[3].um_I.iw[16] ;
 wire \top_I.branch[22].block[3].um_I.iw[17] ;
 wire \top_I.branch[22].block[3].um_I.iw[1] ;
 wire \top_I.branch[22].block[3].um_I.iw[2] ;
 wire \top_I.branch[22].block[3].um_I.iw[3] ;
 wire \top_I.branch[22].block[3].um_I.iw[4] ;
 wire \top_I.branch[22].block[3].um_I.iw[5] ;
 wire \top_I.branch[22].block[3].um_I.iw[6] ;
 wire \top_I.branch[22].block[3].um_I.iw[7] ;
 wire \top_I.branch[22].block[3].um_I.iw[8] ;
 wire \top_I.branch[22].block[3].um_I.iw[9] ;
 wire \top_I.branch[22].block[3].um_I.k_zero ;
 wire \top_I.branch[22].block[3].um_I.pg_vdd ;
 wire \top_I.branch[22].block[4].um_I.ana[0] ;
 wire \top_I.branch[22].block[4].um_I.ana[1] ;
 wire \top_I.branch[22].block[4].um_I.ana[2] ;
 wire \top_I.branch[22].block[4].um_I.ana[3] ;
 wire \top_I.branch[22].block[4].um_I.ana[4] ;
 wire \top_I.branch[22].block[4].um_I.ana[5] ;
 wire \top_I.branch[22].block[4].um_I.ana[6] ;
 wire \top_I.branch[22].block[4].um_I.ana[7] ;
 wire \top_I.branch[22].block[4].um_I.clk ;
 wire \top_I.branch[22].block[4].um_I.ena ;
 wire \top_I.branch[22].block[4].um_I.iw[10] ;
 wire \top_I.branch[22].block[4].um_I.iw[11] ;
 wire \top_I.branch[22].block[4].um_I.iw[12] ;
 wire \top_I.branch[22].block[4].um_I.iw[13] ;
 wire \top_I.branch[22].block[4].um_I.iw[14] ;
 wire \top_I.branch[22].block[4].um_I.iw[15] ;
 wire \top_I.branch[22].block[4].um_I.iw[16] ;
 wire \top_I.branch[22].block[4].um_I.iw[17] ;
 wire \top_I.branch[22].block[4].um_I.iw[1] ;
 wire \top_I.branch[22].block[4].um_I.iw[2] ;
 wire \top_I.branch[22].block[4].um_I.iw[3] ;
 wire \top_I.branch[22].block[4].um_I.iw[4] ;
 wire \top_I.branch[22].block[4].um_I.iw[5] ;
 wire \top_I.branch[22].block[4].um_I.iw[6] ;
 wire \top_I.branch[22].block[4].um_I.iw[7] ;
 wire \top_I.branch[22].block[4].um_I.iw[8] ;
 wire \top_I.branch[22].block[4].um_I.iw[9] ;
 wire \top_I.branch[22].block[4].um_I.k_zero ;
 wire \top_I.branch[22].block[4].um_I.pg_vdd ;
 wire \top_I.branch[22].block[5].um_I.ana[0] ;
 wire \top_I.branch[22].block[5].um_I.ana[1] ;
 wire \top_I.branch[22].block[5].um_I.ana[2] ;
 wire \top_I.branch[22].block[5].um_I.ana[3] ;
 wire \top_I.branch[22].block[5].um_I.ana[4] ;
 wire \top_I.branch[22].block[5].um_I.ana[5] ;
 wire \top_I.branch[22].block[5].um_I.ana[6] ;
 wire \top_I.branch[22].block[5].um_I.ana[7] ;
 wire \top_I.branch[22].block[5].um_I.clk ;
 wire \top_I.branch[22].block[5].um_I.ena ;
 wire \top_I.branch[22].block[5].um_I.iw[10] ;
 wire \top_I.branch[22].block[5].um_I.iw[11] ;
 wire \top_I.branch[22].block[5].um_I.iw[12] ;
 wire \top_I.branch[22].block[5].um_I.iw[13] ;
 wire \top_I.branch[22].block[5].um_I.iw[14] ;
 wire \top_I.branch[22].block[5].um_I.iw[15] ;
 wire \top_I.branch[22].block[5].um_I.iw[16] ;
 wire \top_I.branch[22].block[5].um_I.iw[17] ;
 wire \top_I.branch[22].block[5].um_I.iw[1] ;
 wire \top_I.branch[22].block[5].um_I.iw[2] ;
 wire \top_I.branch[22].block[5].um_I.iw[3] ;
 wire \top_I.branch[22].block[5].um_I.iw[4] ;
 wire \top_I.branch[22].block[5].um_I.iw[5] ;
 wire \top_I.branch[22].block[5].um_I.iw[6] ;
 wire \top_I.branch[22].block[5].um_I.iw[7] ;
 wire \top_I.branch[22].block[5].um_I.iw[8] ;
 wire \top_I.branch[22].block[5].um_I.iw[9] ;
 wire \top_I.branch[22].block[5].um_I.k_zero ;
 wire \top_I.branch[22].block[5].um_I.pg_vdd ;
 wire \top_I.branch[22].block[6].um_I.ana[0] ;
 wire \top_I.branch[22].block[6].um_I.ana[1] ;
 wire \top_I.branch[22].block[6].um_I.ana[2] ;
 wire \top_I.branch[22].block[6].um_I.ana[3] ;
 wire \top_I.branch[22].block[6].um_I.ana[4] ;
 wire \top_I.branch[22].block[6].um_I.ana[5] ;
 wire \top_I.branch[22].block[6].um_I.ana[6] ;
 wire \top_I.branch[22].block[6].um_I.ana[7] ;
 wire \top_I.branch[22].block[6].um_I.clk ;
 wire \top_I.branch[22].block[6].um_I.ena ;
 wire \top_I.branch[22].block[6].um_I.iw[10] ;
 wire \top_I.branch[22].block[6].um_I.iw[11] ;
 wire \top_I.branch[22].block[6].um_I.iw[12] ;
 wire \top_I.branch[22].block[6].um_I.iw[13] ;
 wire \top_I.branch[22].block[6].um_I.iw[14] ;
 wire \top_I.branch[22].block[6].um_I.iw[15] ;
 wire \top_I.branch[22].block[6].um_I.iw[16] ;
 wire \top_I.branch[22].block[6].um_I.iw[17] ;
 wire \top_I.branch[22].block[6].um_I.iw[1] ;
 wire \top_I.branch[22].block[6].um_I.iw[2] ;
 wire \top_I.branch[22].block[6].um_I.iw[3] ;
 wire \top_I.branch[22].block[6].um_I.iw[4] ;
 wire \top_I.branch[22].block[6].um_I.iw[5] ;
 wire \top_I.branch[22].block[6].um_I.iw[6] ;
 wire \top_I.branch[22].block[6].um_I.iw[7] ;
 wire \top_I.branch[22].block[6].um_I.iw[8] ;
 wire \top_I.branch[22].block[6].um_I.iw[9] ;
 wire \top_I.branch[22].block[6].um_I.k_zero ;
 wire \top_I.branch[22].block[6].um_I.pg_vdd ;
 wire \top_I.branch[22].block[7].um_I.ana[0] ;
 wire \top_I.branch[22].block[7].um_I.ana[1] ;
 wire \top_I.branch[22].block[7].um_I.ana[2] ;
 wire \top_I.branch[22].block[7].um_I.ana[3] ;
 wire \top_I.branch[22].block[7].um_I.ana[4] ;
 wire \top_I.branch[22].block[7].um_I.ana[5] ;
 wire \top_I.branch[22].block[7].um_I.ana[6] ;
 wire \top_I.branch[22].block[7].um_I.ana[7] ;
 wire \top_I.branch[22].block[7].um_I.clk ;
 wire \top_I.branch[22].block[7].um_I.ena ;
 wire \top_I.branch[22].block[7].um_I.iw[10] ;
 wire \top_I.branch[22].block[7].um_I.iw[11] ;
 wire \top_I.branch[22].block[7].um_I.iw[12] ;
 wire \top_I.branch[22].block[7].um_I.iw[13] ;
 wire \top_I.branch[22].block[7].um_I.iw[14] ;
 wire \top_I.branch[22].block[7].um_I.iw[15] ;
 wire \top_I.branch[22].block[7].um_I.iw[16] ;
 wire \top_I.branch[22].block[7].um_I.iw[17] ;
 wire \top_I.branch[22].block[7].um_I.iw[1] ;
 wire \top_I.branch[22].block[7].um_I.iw[2] ;
 wire \top_I.branch[22].block[7].um_I.iw[3] ;
 wire \top_I.branch[22].block[7].um_I.iw[4] ;
 wire \top_I.branch[22].block[7].um_I.iw[5] ;
 wire \top_I.branch[22].block[7].um_I.iw[6] ;
 wire \top_I.branch[22].block[7].um_I.iw[7] ;
 wire \top_I.branch[22].block[7].um_I.iw[8] ;
 wire \top_I.branch[22].block[7].um_I.iw[9] ;
 wire \top_I.branch[22].block[7].um_I.k_zero ;
 wire \top_I.branch[22].block[7].um_I.pg_vdd ;
 wire \top_I.branch[22].block[8].um_I.ana[0] ;
 wire \top_I.branch[22].block[8].um_I.ana[1] ;
 wire \top_I.branch[22].block[8].um_I.ana[2] ;
 wire \top_I.branch[22].block[8].um_I.ana[3] ;
 wire \top_I.branch[22].block[8].um_I.ana[4] ;
 wire \top_I.branch[22].block[8].um_I.ana[5] ;
 wire \top_I.branch[22].block[8].um_I.ana[6] ;
 wire \top_I.branch[22].block[8].um_I.ana[7] ;
 wire \top_I.branch[22].block[8].um_I.clk ;
 wire \top_I.branch[22].block[8].um_I.ena ;
 wire \top_I.branch[22].block[8].um_I.iw[10] ;
 wire \top_I.branch[22].block[8].um_I.iw[11] ;
 wire \top_I.branch[22].block[8].um_I.iw[12] ;
 wire \top_I.branch[22].block[8].um_I.iw[13] ;
 wire \top_I.branch[22].block[8].um_I.iw[14] ;
 wire \top_I.branch[22].block[8].um_I.iw[15] ;
 wire \top_I.branch[22].block[8].um_I.iw[16] ;
 wire \top_I.branch[22].block[8].um_I.iw[17] ;
 wire \top_I.branch[22].block[8].um_I.iw[1] ;
 wire \top_I.branch[22].block[8].um_I.iw[2] ;
 wire \top_I.branch[22].block[8].um_I.iw[3] ;
 wire \top_I.branch[22].block[8].um_I.iw[4] ;
 wire \top_I.branch[22].block[8].um_I.iw[5] ;
 wire \top_I.branch[22].block[8].um_I.iw[6] ;
 wire \top_I.branch[22].block[8].um_I.iw[7] ;
 wire \top_I.branch[22].block[8].um_I.iw[8] ;
 wire \top_I.branch[22].block[8].um_I.iw[9] ;
 wire \top_I.branch[22].block[8].um_I.k_zero ;
 wire \top_I.branch[22].block[8].um_I.pg_vdd ;
 wire \top_I.branch[22].block[9].um_I.ana[0] ;
 wire \top_I.branch[22].block[9].um_I.ana[1] ;
 wire \top_I.branch[22].block[9].um_I.ana[2] ;
 wire \top_I.branch[22].block[9].um_I.ana[3] ;
 wire \top_I.branch[22].block[9].um_I.ana[4] ;
 wire \top_I.branch[22].block[9].um_I.ana[5] ;
 wire \top_I.branch[22].block[9].um_I.ana[6] ;
 wire \top_I.branch[22].block[9].um_I.ana[7] ;
 wire \top_I.branch[22].block[9].um_I.clk ;
 wire \top_I.branch[22].block[9].um_I.ena ;
 wire \top_I.branch[22].block[9].um_I.iw[10] ;
 wire \top_I.branch[22].block[9].um_I.iw[11] ;
 wire \top_I.branch[22].block[9].um_I.iw[12] ;
 wire \top_I.branch[22].block[9].um_I.iw[13] ;
 wire \top_I.branch[22].block[9].um_I.iw[14] ;
 wire \top_I.branch[22].block[9].um_I.iw[15] ;
 wire \top_I.branch[22].block[9].um_I.iw[16] ;
 wire \top_I.branch[22].block[9].um_I.iw[17] ;
 wire \top_I.branch[22].block[9].um_I.iw[1] ;
 wire \top_I.branch[22].block[9].um_I.iw[2] ;
 wire \top_I.branch[22].block[9].um_I.iw[3] ;
 wire \top_I.branch[22].block[9].um_I.iw[4] ;
 wire \top_I.branch[22].block[9].um_I.iw[5] ;
 wire \top_I.branch[22].block[9].um_I.iw[6] ;
 wire \top_I.branch[22].block[9].um_I.iw[7] ;
 wire \top_I.branch[22].block[9].um_I.iw[8] ;
 wire \top_I.branch[22].block[9].um_I.iw[9] ;
 wire \top_I.branch[22].block[9].um_I.k_zero ;
 wire \top_I.branch[22].block[9].um_I.pg_vdd ;
 wire \top_I.branch[22].l_addr[0] ;
 wire \top_I.branch[22].l_addr[2] ;
 wire \top_I.branch[23].block[0].um_I.ana[0] ;
 wire \top_I.branch[23].block[0].um_I.ana[1] ;
 wire \top_I.branch[23].block[0].um_I.ana[2] ;
 wire \top_I.branch[23].block[0].um_I.ana[3] ;
 wire \top_I.branch[23].block[0].um_I.ana[4] ;
 wire \top_I.branch[23].block[0].um_I.ana[5] ;
 wire \top_I.branch[23].block[0].um_I.ana[6] ;
 wire \top_I.branch[23].block[0].um_I.ana[7] ;
 wire \top_I.branch[23].block[0].um_I.clk ;
 wire \top_I.branch[23].block[0].um_I.ena ;
 wire \top_I.branch[23].block[0].um_I.iw[10] ;
 wire \top_I.branch[23].block[0].um_I.iw[11] ;
 wire \top_I.branch[23].block[0].um_I.iw[12] ;
 wire \top_I.branch[23].block[0].um_I.iw[13] ;
 wire \top_I.branch[23].block[0].um_I.iw[14] ;
 wire \top_I.branch[23].block[0].um_I.iw[15] ;
 wire \top_I.branch[23].block[0].um_I.iw[16] ;
 wire \top_I.branch[23].block[0].um_I.iw[17] ;
 wire \top_I.branch[23].block[0].um_I.iw[1] ;
 wire \top_I.branch[23].block[0].um_I.iw[2] ;
 wire \top_I.branch[23].block[0].um_I.iw[3] ;
 wire \top_I.branch[23].block[0].um_I.iw[4] ;
 wire \top_I.branch[23].block[0].um_I.iw[5] ;
 wire \top_I.branch[23].block[0].um_I.iw[6] ;
 wire \top_I.branch[23].block[0].um_I.iw[7] ;
 wire \top_I.branch[23].block[0].um_I.iw[8] ;
 wire \top_I.branch[23].block[0].um_I.iw[9] ;
 wire \top_I.branch[23].block[0].um_I.k_zero ;
 wire \top_I.branch[23].block[0].um_I.pg_vdd ;
 wire \top_I.branch[23].block[10].um_I.ana[0] ;
 wire \top_I.branch[23].block[10].um_I.ana[1] ;
 wire \top_I.branch[23].block[10].um_I.ana[2] ;
 wire \top_I.branch[23].block[10].um_I.ana[3] ;
 wire \top_I.branch[23].block[10].um_I.ana[4] ;
 wire \top_I.branch[23].block[10].um_I.ana[5] ;
 wire \top_I.branch[23].block[10].um_I.ana[6] ;
 wire \top_I.branch[23].block[10].um_I.ana[7] ;
 wire \top_I.branch[23].block[10].um_I.clk ;
 wire \top_I.branch[23].block[10].um_I.ena ;
 wire \top_I.branch[23].block[10].um_I.iw[10] ;
 wire \top_I.branch[23].block[10].um_I.iw[11] ;
 wire \top_I.branch[23].block[10].um_I.iw[12] ;
 wire \top_I.branch[23].block[10].um_I.iw[13] ;
 wire \top_I.branch[23].block[10].um_I.iw[14] ;
 wire \top_I.branch[23].block[10].um_I.iw[15] ;
 wire \top_I.branch[23].block[10].um_I.iw[16] ;
 wire \top_I.branch[23].block[10].um_I.iw[17] ;
 wire \top_I.branch[23].block[10].um_I.iw[1] ;
 wire \top_I.branch[23].block[10].um_I.iw[2] ;
 wire \top_I.branch[23].block[10].um_I.iw[3] ;
 wire \top_I.branch[23].block[10].um_I.iw[4] ;
 wire \top_I.branch[23].block[10].um_I.iw[5] ;
 wire \top_I.branch[23].block[10].um_I.iw[6] ;
 wire \top_I.branch[23].block[10].um_I.iw[7] ;
 wire \top_I.branch[23].block[10].um_I.iw[8] ;
 wire \top_I.branch[23].block[10].um_I.iw[9] ;
 wire \top_I.branch[23].block[10].um_I.k_zero ;
 wire \top_I.branch[23].block[10].um_I.pg_vdd ;
 wire \top_I.branch[23].block[11].um_I.ana[0] ;
 wire \top_I.branch[23].block[11].um_I.ana[1] ;
 wire \top_I.branch[23].block[11].um_I.ana[2] ;
 wire \top_I.branch[23].block[11].um_I.ana[3] ;
 wire \top_I.branch[23].block[11].um_I.ana[4] ;
 wire \top_I.branch[23].block[11].um_I.ana[5] ;
 wire \top_I.branch[23].block[11].um_I.ana[6] ;
 wire \top_I.branch[23].block[11].um_I.ana[7] ;
 wire \top_I.branch[23].block[11].um_I.clk ;
 wire \top_I.branch[23].block[11].um_I.ena ;
 wire \top_I.branch[23].block[11].um_I.iw[10] ;
 wire \top_I.branch[23].block[11].um_I.iw[11] ;
 wire \top_I.branch[23].block[11].um_I.iw[12] ;
 wire \top_I.branch[23].block[11].um_I.iw[13] ;
 wire \top_I.branch[23].block[11].um_I.iw[14] ;
 wire \top_I.branch[23].block[11].um_I.iw[15] ;
 wire \top_I.branch[23].block[11].um_I.iw[16] ;
 wire \top_I.branch[23].block[11].um_I.iw[17] ;
 wire \top_I.branch[23].block[11].um_I.iw[1] ;
 wire \top_I.branch[23].block[11].um_I.iw[2] ;
 wire \top_I.branch[23].block[11].um_I.iw[3] ;
 wire \top_I.branch[23].block[11].um_I.iw[4] ;
 wire \top_I.branch[23].block[11].um_I.iw[5] ;
 wire \top_I.branch[23].block[11].um_I.iw[6] ;
 wire \top_I.branch[23].block[11].um_I.iw[7] ;
 wire \top_I.branch[23].block[11].um_I.iw[8] ;
 wire \top_I.branch[23].block[11].um_I.iw[9] ;
 wire \top_I.branch[23].block[11].um_I.k_zero ;
 wire \top_I.branch[23].block[11].um_I.pg_vdd ;
 wire \top_I.branch[23].block[12].um_I.ana[0] ;
 wire \top_I.branch[23].block[12].um_I.ana[1] ;
 wire \top_I.branch[23].block[12].um_I.ana[2] ;
 wire \top_I.branch[23].block[12].um_I.ana[3] ;
 wire \top_I.branch[23].block[12].um_I.ana[4] ;
 wire \top_I.branch[23].block[12].um_I.ana[5] ;
 wire \top_I.branch[23].block[12].um_I.ana[6] ;
 wire \top_I.branch[23].block[12].um_I.ana[7] ;
 wire \top_I.branch[23].block[12].um_I.clk ;
 wire \top_I.branch[23].block[12].um_I.ena ;
 wire \top_I.branch[23].block[12].um_I.iw[10] ;
 wire \top_I.branch[23].block[12].um_I.iw[11] ;
 wire \top_I.branch[23].block[12].um_I.iw[12] ;
 wire \top_I.branch[23].block[12].um_I.iw[13] ;
 wire \top_I.branch[23].block[12].um_I.iw[14] ;
 wire \top_I.branch[23].block[12].um_I.iw[15] ;
 wire \top_I.branch[23].block[12].um_I.iw[16] ;
 wire \top_I.branch[23].block[12].um_I.iw[17] ;
 wire \top_I.branch[23].block[12].um_I.iw[1] ;
 wire \top_I.branch[23].block[12].um_I.iw[2] ;
 wire \top_I.branch[23].block[12].um_I.iw[3] ;
 wire \top_I.branch[23].block[12].um_I.iw[4] ;
 wire \top_I.branch[23].block[12].um_I.iw[5] ;
 wire \top_I.branch[23].block[12].um_I.iw[6] ;
 wire \top_I.branch[23].block[12].um_I.iw[7] ;
 wire \top_I.branch[23].block[12].um_I.iw[8] ;
 wire \top_I.branch[23].block[12].um_I.iw[9] ;
 wire \top_I.branch[23].block[12].um_I.k_zero ;
 wire \top_I.branch[23].block[12].um_I.pg_vdd ;
 wire \top_I.branch[23].block[13].um_I.ana[0] ;
 wire \top_I.branch[23].block[13].um_I.ana[1] ;
 wire \top_I.branch[23].block[13].um_I.ana[2] ;
 wire \top_I.branch[23].block[13].um_I.ana[3] ;
 wire \top_I.branch[23].block[13].um_I.ana[4] ;
 wire \top_I.branch[23].block[13].um_I.ana[5] ;
 wire \top_I.branch[23].block[13].um_I.ana[6] ;
 wire \top_I.branch[23].block[13].um_I.ana[7] ;
 wire \top_I.branch[23].block[13].um_I.clk ;
 wire \top_I.branch[23].block[13].um_I.ena ;
 wire \top_I.branch[23].block[13].um_I.iw[10] ;
 wire \top_I.branch[23].block[13].um_I.iw[11] ;
 wire \top_I.branch[23].block[13].um_I.iw[12] ;
 wire \top_I.branch[23].block[13].um_I.iw[13] ;
 wire \top_I.branch[23].block[13].um_I.iw[14] ;
 wire \top_I.branch[23].block[13].um_I.iw[15] ;
 wire \top_I.branch[23].block[13].um_I.iw[16] ;
 wire \top_I.branch[23].block[13].um_I.iw[17] ;
 wire \top_I.branch[23].block[13].um_I.iw[1] ;
 wire \top_I.branch[23].block[13].um_I.iw[2] ;
 wire \top_I.branch[23].block[13].um_I.iw[3] ;
 wire \top_I.branch[23].block[13].um_I.iw[4] ;
 wire \top_I.branch[23].block[13].um_I.iw[5] ;
 wire \top_I.branch[23].block[13].um_I.iw[6] ;
 wire \top_I.branch[23].block[13].um_I.iw[7] ;
 wire \top_I.branch[23].block[13].um_I.iw[8] ;
 wire \top_I.branch[23].block[13].um_I.iw[9] ;
 wire \top_I.branch[23].block[13].um_I.k_zero ;
 wire \top_I.branch[23].block[13].um_I.pg_vdd ;
 wire \top_I.branch[23].block[14].um_I.ana[0] ;
 wire \top_I.branch[23].block[14].um_I.ana[1] ;
 wire \top_I.branch[23].block[14].um_I.ana[2] ;
 wire \top_I.branch[23].block[14].um_I.ana[3] ;
 wire \top_I.branch[23].block[14].um_I.ana[4] ;
 wire \top_I.branch[23].block[14].um_I.ana[5] ;
 wire \top_I.branch[23].block[14].um_I.ana[6] ;
 wire \top_I.branch[23].block[14].um_I.ana[7] ;
 wire \top_I.branch[23].block[14].um_I.clk ;
 wire \top_I.branch[23].block[14].um_I.ena ;
 wire \top_I.branch[23].block[14].um_I.iw[10] ;
 wire \top_I.branch[23].block[14].um_I.iw[11] ;
 wire \top_I.branch[23].block[14].um_I.iw[12] ;
 wire \top_I.branch[23].block[14].um_I.iw[13] ;
 wire \top_I.branch[23].block[14].um_I.iw[14] ;
 wire \top_I.branch[23].block[14].um_I.iw[15] ;
 wire \top_I.branch[23].block[14].um_I.iw[16] ;
 wire \top_I.branch[23].block[14].um_I.iw[17] ;
 wire \top_I.branch[23].block[14].um_I.iw[1] ;
 wire \top_I.branch[23].block[14].um_I.iw[2] ;
 wire \top_I.branch[23].block[14].um_I.iw[3] ;
 wire \top_I.branch[23].block[14].um_I.iw[4] ;
 wire \top_I.branch[23].block[14].um_I.iw[5] ;
 wire \top_I.branch[23].block[14].um_I.iw[6] ;
 wire \top_I.branch[23].block[14].um_I.iw[7] ;
 wire \top_I.branch[23].block[14].um_I.iw[8] ;
 wire \top_I.branch[23].block[14].um_I.iw[9] ;
 wire \top_I.branch[23].block[14].um_I.k_zero ;
 wire \top_I.branch[23].block[14].um_I.pg_vdd ;
 wire \top_I.branch[23].block[15].um_I.ana[0] ;
 wire \top_I.branch[23].block[15].um_I.ana[1] ;
 wire \top_I.branch[23].block[15].um_I.ana[2] ;
 wire \top_I.branch[23].block[15].um_I.ana[3] ;
 wire \top_I.branch[23].block[15].um_I.ana[4] ;
 wire \top_I.branch[23].block[15].um_I.ana[5] ;
 wire \top_I.branch[23].block[15].um_I.ana[6] ;
 wire \top_I.branch[23].block[15].um_I.ana[7] ;
 wire \top_I.branch[23].block[15].um_I.clk ;
 wire \top_I.branch[23].block[15].um_I.ena ;
 wire \top_I.branch[23].block[15].um_I.iw[10] ;
 wire \top_I.branch[23].block[15].um_I.iw[11] ;
 wire \top_I.branch[23].block[15].um_I.iw[12] ;
 wire \top_I.branch[23].block[15].um_I.iw[13] ;
 wire \top_I.branch[23].block[15].um_I.iw[14] ;
 wire \top_I.branch[23].block[15].um_I.iw[15] ;
 wire \top_I.branch[23].block[15].um_I.iw[16] ;
 wire \top_I.branch[23].block[15].um_I.iw[17] ;
 wire \top_I.branch[23].block[15].um_I.iw[1] ;
 wire \top_I.branch[23].block[15].um_I.iw[2] ;
 wire \top_I.branch[23].block[15].um_I.iw[3] ;
 wire \top_I.branch[23].block[15].um_I.iw[4] ;
 wire \top_I.branch[23].block[15].um_I.iw[5] ;
 wire \top_I.branch[23].block[15].um_I.iw[6] ;
 wire \top_I.branch[23].block[15].um_I.iw[7] ;
 wire \top_I.branch[23].block[15].um_I.iw[8] ;
 wire \top_I.branch[23].block[15].um_I.iw[9] ;
 wire \top_I.branch[23].block[15].um_I.k_zero ;
 wire \top_I.branch[23].block[15].um_I.pg_vdd ;
 wire \top_I.branch[23].block[1].um_I.ana[0] ;
 wire \top_I.branch[23].block[1].um_I.ana[1] ;
 wire \top_I.branch[23].block[1].um_I.ana[2] ;
 wire \top_I.branch[23].block[1].um_I.ana[3] ;
 wire \top_I.branch[23].block[1].um_I.ana[4] ;
 wire \top_I.branch[23].block[1].um_I.ana[5] ;
 wire \top_I.branch[23].block[1].um_I.ana[6] ;
 wire \top_I.branch[23].block[1].um_I.ana[7] ;
 wire \top_I.branch[23].block[1].um_I.clk ;
 wire \top_I.branch[23].block[1].um_I.ena ;
 wire \top_I.branch[23].block[1].um_I.iw[10] ;
 wire \top_I.branch[23].block[1].um_I.iw[11] ;
 wire \top_I.branch[23].block[1].um_I.iw[12] ;
 wire \top_I.branch[23].block[1].um_I.iw[13] ;
 wire \top_I.branch[23].block[1].um_I.iw[14] ;
 wire \top_I.branch[23].block[1].um_I.iw[15] ;
 wire \top_I.branch[23].block[1].um_I.iw[16] ;
 wire \top_I.branch[23].block[1].um_I.iw[17] ;
 wire \top_I.branch[23].block[1].um_I.iw[1] ;
 wire \top_I.branch[23].block[1].um_I.iw[2] ;
 wire \top_I.branch[23].block[1].um_I.iw[3] ;
 wire \top_I.branch[23].block[1].um_I.iw[4] ;
 wire \top_I.branch[23].block[1].um_I.iw[5] ;
 wire \top_I.branch[23].block[1].um_I.iw[6] ;
 wire \top_I.branch[23].block[1].um_I.iw[7] ;
 wire \top_I.branch[23].block[1].um_I.iw[8] ;
 wire \top_I.branch[23].block[1].um_I.iw[9] ;
 wire \top_I.branch[23].block[1].um_I.k_zero ;
 wire \top_I.branch[23].block[1].um_I.pg_vdd ;
 wire \top_I.branch[23].block[2].um_I.ana[0] ;
 wire \top_I.branch[23].block[2].um_I.ana[1] ;
 wire \top_I.branch[23].block[2].um_I.ana[2] ;
 wire \top_I.branch[23].block[2].um_I.ana[3] ;
 wire \top_I.branch[23].block[2].um_I.ana[4] ;
 wire \top_I.branch[23].block[2].um_I.ana[5] ;
 wire \top_I.branch[23].block[2].um_I.ana[6] ;
 wire \top_I.branch[23].block[2].um_I.ana[7] ;
 wire \top_I.branch[23].block[2].um_I.clk ;
 wire \top_I.branch[23].block[2].um_I.ena ;
 wire \top_I.branch[23].block[2].um_I.iw[10] ;
 wire \top_I.branch[23].block[2].um_I.iw[11] ;
 wire \top_I.branch[23].block[2].um_I.iw[12] ;
 wire \top_I.branch[23].block[2].um_I.iw[13] ;
 wire \top_I.branch[23].block[2].um_I.iw[14] ;
 wire \top_I.branch[23].block[2].um_I.iw[15] ;
 wire \top_I.branch[23].block[2].um_I.iw[16] ;
 wire \top_I.branch[23].block[2].um_I.iw[17] ;
 wire \top_I.branch[23].block[2].um_I.iw[1] ;
 wire \top_I.branch[23].block[2].um_I.iw[2] ;
 wire \top_I.branch[23].block[2].um_I.iw[3] ;
 wire \top_I.branch[23].block[2].um_I.iw[4] ;
 wire \top_I.branch[23].block[2].um_I.iw[5] ;
 wire \top_I.branch[23].block[2].um_I.iw[6] ;
 wire \top_I.branch[23].block[2].um_I.iw[7] ;
 wire \top_I.branch[23].block[2].um_I.iw[8] ;
 wire \top_I.branch[23].block[2].um_I.iw[9] ;
 wire \top_I.branch[23].block[2].um_I.k_zero ;
 wire \top_I.branch[23].block[2].um_I.pg_vdd ;
 wire \top_I.branch[23].block[3].um_I.ana[0] ;
 wire \top_I.branch[23].block[3].um_I.ana[1] ;
 wire \top_I.branch[23].block[3].um_I.ana[2] ;
 wire \top_I.branch[23].block[3].um_I.ana[3] ;
 wire \top_I.branch[23].block[3].um_I.ana[4] ;
 wire \top_I.branch[23].block[3].um_I.ana[5] ;
 wire \top_I.branch[23].block[3].um_I.ana[6] ;
 wire \top_I.branch[23].block[3].um_I.ana[7] ;
 wire \top_I.branch[23].block[3].um_I.clk ;
 wire \top_I.branch[23].block[3].um_I.ena ;
 wire \top_I.branch[23].block[3].um_I.iw[10] ;
 wire \top_I.branch[23].block[3].um_I.iw[11] ;
 wire \top_I.branch[23].block[3].um_I.iw[12] ;
 wire \top_I.branch[23].block[3].um_I.iw[13] ;
 wire \top_I.branch[23].block[3].um_I.iw[14] ;
 wire \top_I.branch[23].block[3].um_I.iw[15] ;
 wire \top_I.branch[23].block[3].um_I.iw[16] ;
 wire \top_I.branch[23].block[3].um_I.iw[17] ;
 wire \top_I.branch[23].block[3].um_I.iw[1] ;
 wire \top_I.branch[23].block[3].um_I.iw[2] ;
 wire \top_I.branch[23].block[3].um_I.iw[3] ;
 wire \top_I.branch[23].block[3].um_I.iw[4] ;
 wire \top_I.branch[23].block[3].um_I.iw[5] ;
 wire \top_I.branch[23].block[3].um_I.iw[6] ;
 wire \top_I.branch[23].block[3].um_I.iw[7] ;
 wire \top_I.branch[23].block[3].um_I.iw[8] ;
 wire \top_I.branch[23].block[3].um_I.iw[9] ;
 wire \top_I.branch[23].block[3].um_I.k_zero ;
 wire \top_I.branch[23].block[3].um_I.pg_vdd ;
 wire \top_I.branch[23].block[4].um_I.ana[0] ;
 wire \top_I.branch[23].block[4].um_I.ana[1] ;
 wire \top_I.branch[23].block[4].um_I.ana[2] ;
 wire \top_I.branch[23].block[4].um_I.ana[3] ;
 wire \top_I.branch[23].block[4].um_I.ana[4] ;
 wire \top_I.branch[23].block[4].um_I.ana[5] ;
 wire \top_I.branch[23].block[4].um_I.ana[6] ;
 wire \top_I.branch[23].block[4].um_I.ana[7] ;
 wire \top_I.branch[23].block[4].um_I.clk ;
 wire \top_I.branch[23].block[4].um_I.ena ;
 wire \top_I.branch[23].block[4].um_I.iw[10] ;
 wire \top_I.branch[23].block[4].um_I.iw[11] ;
 wire \top_I.branch[23].block[4].um_I.iw[12] ;
 wire \top_I.branch[23].block[4].um_I.iw[13] ;
 wire \top_I.branch[23].block[4].um_I.iw[14] ;
 wire \top_I.branch[23].block[4].um_I.iw[15] ;
 wire \top_I.branch[23].block[4].um_I.iw[16] ;
 wire \top_I.branch[23].block[4].um_I.iw[17] ;
 wire \top_I.branch[23].block[4].um_I.iw[1] ;
 wire \top_I.branch[23].block[4].um_I.iw[2] ;
 wire \top_I.branch[23].block[4].um_I.iw[3] ;
 wire \top_I.branch[23].block[4].um_I.iw[4] ;
 wire \top_I.branch[23].block[4].um_I.iw[5] ;
 wire \top_I.branch[23].block[4].um_I.iw[6] ;
 wire \top_I.branch[23].block[4].um_I.iw[7] ;
 wire \top_I.branch[23].block[4].um_I.iw[8] ;
 wire \top_I.branch[23].block[4].um_I.iw[9] ;
 wire \top_I.branch[23].block[4].um_I.k_zero ;
 wire \top_I.branch[23].block[4].um_I.pg_vdd ;
 wire \top_I.branch[23].block[5].um_I.ana[0] ;
 wire \top_I.branch[23].block[5].um_I.ana[1] ;
 wire \top_I.branch[23].block[5].um_I.ana[2] ;
 wire \top_I.branch[23].block[5].um_I.ana[3] ;
 wire \top_I.branch[23].block[5].um_I.ana[4] ;
 wire \top_I.branch[23].block[5].um_I.ana[5] ;
 wire \top_I.branch[23].block[5].um_I.ana[6] ;
 wire \top_I.branch[23].block[5].um_I.ana[7] ;
 wire \top_I.branch[23].block[5].um_I.clk ;
 wire \top_I.branch[23].block[5].um_I.ena ;
 wire \top_I.branch[23].block[5].um_I.iw[10] ;
 wire \top_I.branch[23].block[5].um_I.iw[11] ;
 wire \top_I.branch[23].block[5].um_I.iw[12] ;
 wire \top_I.branch[23].block[5].um_I.iw[13] ;
 wire \top_I.branch[23].block[5].um_I.iw[14] ;
 wire \top_I.branch[23].block[5].um_I.iw[15] ;
 wire \top_I.branch[23].block[5].um_I.iw[16] ;
 wire \top_I.branch[23].block[5].um_I.iw[17] ;
 wire \top_I.branch[23].block[5].um_I.iw[1] ;
 wire \top_I.branch[23].block[5].um_I.iw[2] ;
 wire \top_I.branch[23].block[5].um_I.iw[3] ;
 wire \top_I.branch[23].block[5].um_I.iw[4] ;
 wire \top_I.branch[23].block[5].um_I.iw[5] ;
 wire \top_I.branch[23].block[5].um_I.iw[6] ;
 wire \top_I.branch[23].block[5].um_I.iw[7] ;
 wire \top_I.branch[23].block[5].um_I.iw[8] ;
 wire \top_I.branch[23].block[5].um_I.iw[9] ;
 wire \top_I.branch[23].block[5].um_I.k_zero ;
 wire \top_I.branch[23].block[5].um_I.pg_vdd ;
 wire \top_I.branch[23].block[6].um_I.ana[0] ;
 wire \top_I.branch[23].block[6].um_I.ana[1] ;
 wire \top_I.branch[23].block[6].um_I.ana[2] ;
 wire \top_I.branch[23].block[6].um_I.ana[3] ;
 wire \top_I.branch[23].block[6].um_I.ana[4] ;
 wire \top_I.branch[23].block[6].um_I.ana[5] ;
 wire \top_I.branch[23].block[6].um_I.ana[6] ;
 wire \top_I.branch[23].block[6].um_I.ana[7] ;
 wire \top_I.branch[23].block[6].um_I.clk ;
 wire \top_I.branch[23].block[6].um_I.ena ;
 wire \top_I.branch[23].block[6].um_I.iw[10] ;
 wire \top_I.branch[23].block[6].um_I.iw[11] ;
 wire \top_I.branch[23].block[6].um_I.iw[12] ;
 wire \top_I.branch[23].block[6].um_I.iw[13] ;
 wire \top_I.branch[23].block[6].um_I.iw[14] ;
 wire \top_I.branch[23].block[6].um_I.iw[15] ;
 wire \top_I.branch[23].block[6].um_I.iw[16] ;
 wire \top_I.branch[23].block[6].um_I.iw[17] ;
 wire \top_I.branch[23].block[6].um_I.iw[1] ;
 wire \top_I.branch[23].block[6].um_I.iw[2] ;
 wire \top_I.branch[23].block[6].um_I.iw[3] ;
 wire \top_I.branch[23].block[6].um_I.iw[4] ;
 wire \top_I.branch[23].block[6].um_I.iw[5] ;
 wire \top_I.branch[23].block[6].um_I.iw[6] ;
 wire \top_I.branch[23].block[6].um_I.iw[7] ;
 wire \top_I.branch[23].block[6].um_I.iw[8] ;
 wire \top_I.branch[23].block[6].um_I.iw[9] ;
 wire \top_I.branch[23].block[6].um_I.k_zero ;
 wire \top_I.branch[23].block[6].um_I.pg_vdd ;
 wire \top_I.branch[23].block[7].um_I.ana[0] ;
 wire \top_I.branch[23].block[7].um_I.ana[1] ;
 wire \top_I.branch[23].block[7].um_I.ana[2] ;
 wire \top_I.branch[23].block[7].um_I.ana[3] ;
 wire \top_I.branch[23].block[7].um_I.ana[4] ;
 wire \top_I.branch[23].block[7].um_I.ana[5] ;
 wire \top_I.branch[23].block[7].um_I.ana[6] ;
 wire \top_I.branch[23].block[7].um_I.ana[7] ;
 wire \top_I.branch[23].block[7].um_I.clk ;
 wire \top_I.branch[23].block[7].um_I.ena ;
 wire \top_I.branch[23].block[7].um_I.iw[10] ;
 wire \top_I.branch[23].block[7].um_I.iw[11] ;
 wire \top_I.branch[23].block[7].um_I.iw[12] ;
 wire \top_I.branch[23].block[7].um_I.iw[13] ;
 wire \top_I.branch[23].block[7].um_I.iw[14] ;
 wire \top_I.branch[23].block[7].um_I.iw[15] ;
 wire \top_I.branch[23].block[7].um_I.iw[16] ;
 wire \top_I.branch[23].block[7].um_I.iw[17] ;
 wire \top_I.branch[23].block[7].um_I.iw[1] ;
 wire \top_I.branch[23].block[7].um_I.iw[2] ;
 wire \top_I.branch[23].block[7].um_I.iw[3] ;
 wire \top_I.branch[23].block[7].um_I.iw[4] ;
 wire \top_I.branch[23].block[7].um_I.iw[5] ;
 wire \top_I.branch[23].block[7].um_I.iw[6] ;
 wire \top_I.branch[23].block[7].um_I.iw[7] ;
 wire \top_I.branch[23].block[7].um_I.iw[8] ;
 wire \top_I.branch[23].block[7].um_I.iw[9] ;
 wire \top_I.branch[23].block[7].um_I.k_zero ;
 wire \top_I.branch[23].block[7].um_I.pg_vdd ;
 wire \top_I.branch[23].block[8].um_I.ana[0] ;
 wire \top_I.branch[23].block[8].um_I.ana[1] ;
 wire \top_I.branch[23].block[8].um_I.ana[2] ;
 wire \top_I.branch[23].block[8].um_I.ana[3] ;
 wire \top_I.branch[23].block[8].um_I.ana[4] ;
 wire \top_I.branch[23].block[8].um_I.ana[5] ;
 wire \top_I.branch[23].block[8].um_I.ana[6] ;
 wire \top_I.branch[23].block[8].um_I.ana[7] ;
 wire \top_I.branch[23].block[8].um_I.clk ;
 wire \top_I.branch[23].block[8].um_I.ena ;
 wire \top_I.branch[23].block[8].um_I.iw[10] ;
 wire \top_I.branch[23].block[8].um_I.iw[11] ;
 wire \top_I.branch[23].block[8].um_I.iw[12] ;
 wire \top_I.branch[23].block[8].um_I.iw[13] ;
 wire \top_I.branch[23].block[8].um_I.iw[14] ;
 wire \top_I.branch[23].block[8].um_I.iw[15] ;
 wire \top_I.branch[23].block[8].um_I.iw[16] ;
 wire \top_I.branch[23].block[8].um_I.iw[17] ;
 wire \top_I.branch[23].block[8].um_I.iw[1] ;
 wire \top_I.branch[23].block[8].um_I.iw[2] ;
 wire \top_I.branch[23].block[8].um_I.iw[3] ;
 wire \top_I.branch[23].block[8].um_I.iw[4] ;
 wire \top_I.branch[23].block[8].um_I.iw[5] ;
 wire \top_I.branch[23].block[8].um_I.iw[6] ;
 wire \top_I.branch[23].block[8].um_I.iw[7] ;
 wire \top_I.branch[23].block[8].um_I.iw[8] ;
 wire \top_I.branch[23].block[8].um_I.iw[9] ;
 wire \top_I.branch[23].block[8].um_I.k_zero ;
 wire \top_I.branch[23].block[8].um_I.pg_vdd ;
 wire \top_I.branch[23].block[9].um_I.ana[0] ;
 wire \top_I.branch[23].block[9].um_I.ana[1] ;
 wire \top_I.branch[23].block[9].um_I.ana[2] ;
 wire \top_I.branch[23].block[9].um_I.ana[3] ;
 wire \top_I.branch[23].block[9].um_I.ana[4] ;
 wire \top_I.branch[23].block[9].um_I.ana[5] ;
 wire \top_I.branch[23].block[9].um_I.ana[6] ;
 wire \top_I.branch[23].block[9].um_I.ana[7] ;
 wire \top_I.branch[23].block[9].um_I.clk ;
 wire \top_I.branch[23].block[9].um_I.ena ;
 wire \top_I.branch[23].block[9].um_I.iw[10] ;
 wire \top_I.branch[23].block[9].um_I.iw[11] ;
 wire \top_I.branch[23].block[9].um_I.iw[12] ;
 wire \top_I.branch[23].block[9].um_I.iw[13] ;
 wire \top_I.branch[23].block[9].um_I.iw[14] ;
 wire \top_I.branch[23].block[9].um_I.iw[15] ;
 wire \top_I.branch[23].block[9].um_I.iw[16] ;
 wire \top_I.branch[23].block[9].um_I.iw[17] ;
 wire \top_I.branch[23].block[9].um_I.iw[1] ;
 wire \top_I.branch[23].block[9].um_I.iw[2] ;
 wire \top_I.branch[23].block[9].um_I.iw[3] ;
 wire \top_I.branch[23].block[9].um_I.iw[4] ;
 wire \top_I.branch[23].block[9].um_I.iw[5] ;
 wire \top_I.branch[23].block[9].um_I.iw[6] ;
 wire \top_I.branch[23].block[9].um_I.iw[7] ;
 wire \top_I.branch[23].block[9].um_I.iw[8] ;
 wire \top_I.branch[23].block[9].um_I.iw[9] ;
 wire \top_I.branch[23].block[9].um_I.k_zero ;
 wire \top_I.branch[23].block[9].um_I.pg_vdd ;
 wire \top_I.branch[23].l_addr[0] ;
 wire \top_I.branch[23].l_addr[2] ;
 wire \top_I.branch[24].block[0].um_I.ana[0] ;
 wire \top_I.branch[24].block[0].um_I.ana[1] ;
 wire \top_I.branch[24].block[0].um_I.ana[2] ;
 wire \top_I.branch[24].block[0].um_I.ana[3] ;
 wire \top_I.branch[24].block[0].um_I.ana[4] ;
 wire \top_I.branch[24].block[0].um_I.ana[5] ;
 wire \top_I.branch[24].block[0].um_I.ana[6] ;
 wire \top_I.branch[24].block[0].um_I.ana[7] ;
 wire \top_I.branch[24].block[0].um_I.clk ;
 wire \top_I.branch[24].block[0].um_I.ena ;
 wire \top_I.branch[24].block[0].um_I.iw[10] ;
 wire \top_I.branch[24].block[0].um_I.iw[11] ;
 wire \top_I.branch[24].block[0].um_I.iw[12] ;
 wire \top_I.branch[24].block[0].um_I.iw[13] ;
 wire \top_I.branch[24].block[0].um_I.iw[14] ;
 wire \top_I.branch[24].block[0].um_I.iw[15] ;
 wire \top_I.branch[24].block[0].um_I.iw[16] ;
 wire \top_I.branch[24].block[0].um_I.iw[17] ;
 wire \top_I.branch[24].block[0].um_I.iw[1] ;
 wire \top_I.branch[24].block[0].um_I.iw[2] ;
 wire \top_I.branch[24].block[0].um_I.iw[3] ;
 wire \top_I.branch[24].block[0].um_I.iw[4] ;
 wire \top_I.branch[24].block[0].um_I.iw[5] ;
 wire \top_I.branch[24].block[0].um_I.iw[6] ;
 wire \top_I.branch[24].block[0].um_I.iw[7] ;
 wire \top_I.branch[24].block[0].um_I.iw[8] ;
 wire \top_I.branch[24].block[0].um_I.iw[9] ;
 wire \top_I.branch[24].block[0].um_I.k_zero ;
 wire \top_I.branch[24].block[0].um_I.pg_vdd ;
 wire \top_I.branch[24].block[10].um_I.ana[0] ;
 wire \top_I.branch[24].block[10].um_I.ana[1] ;
 wire \top_I.branch[24].block[10].um_I.ana[2] ;
 wire \top_I.branch[24].block[10].um_I.ana[3] ;
 wire \top_I.branch[24].block[10].um_I.ana[4] ;
 wire \top_I.branch[24].block[10].um_I.ana[5] ;
 wire \top_I.branch[24].block[10].um_I.ana[6] ;
 wire \top_I.branch[24].block[10].um_I.ana[7] ;
 wire \top_I.branch[24].block[10].um_I.clk ;
 wire \top_I.branch[24].block[10].um_I.ena ;
 wire \top_I.branch[24].block[10].um_I.iw[10] ;
 wire \top_I.branch[24].block[10].um_I.iw[11] ;
 wire \top_I.branch[24].block[10].um_I.iw[12] ;
 wire \top_I.branch[24].block[10].um_I.iw[13] ;
 wire \top_I.branch[24].block[10].um_I.iw[14] ;
 wire \top_I.branch[24].block[10].um_I.iw[15] ;
 wire \top_I.branch[24].block[10].um_I.iw[16] ;
 wire \top_I.branch[24].block[10].um_I.iw[17] ;
 wire \top_I.branch[24].block[10].um_I.iw[1] ;
 wire \top_I.branch[24].block[10].um_I.iw[2] ;
 wire \top_I.branch[24].block[10].um_I.iw[3] ;
 wire \top_I.branch[24].block[10].um_I.iw[4] ;
 wire \top_I.branch[24].block[10].um_I.iw[5] ;
 wire \top_I.branch[24].block[10].um_I.iw[6] ;
 wire \top_I.branch[24].block[10].um_I.iw[7] ;
 wire \top_I.branch[24].block[10].um_I.iw[8] ;
 wire \top_I.branch[24].block[10].um_I.iw[9] ;
 wire \top_I.branch[24].block[10].um_I.k_zero ;
 wire \top_I.branch[24].block[10].um_I.pg_vdd ;
 wire \top_I.branch[24].block[11].um_I.ana[0] ;
 wire \top_I.branch[24].block[11].um_I.ana[1] ;
 wire \top_I.branch[24].block[11].um_I.ana[2] ;
 wire \top_I.branch[24].block[11].um_I.ana[3] ;
 wire \top_I.branch[24].block[11].um_I.ana[4] ;
 wire \top_I.branch[24].block[11].um_I.ana[5] ;
 wire \top_I.branch[24].block[11].um_I.ana[6] ;
 wire \top_I.branch[24].block[11].um_I.ana[7] ;
 wire \top_I.branch[24].block[11].um_I.clk ;
 wire \top_I.branch[24].block[11].um_I.ena ;
 wire \top_I.branch[24].block[11].um_I.iw[10] ;
 wire \top_I.branch[24].block[11].um_I.iw[11] ;
 wire \top_I.branch[24].block[11].um_I.iw[12] ;
 wire \top_I.branch[24].block[11].um_I.iw[13] ;
 wire \top_I.branch[24].block[11].um_I.iw[14] ;
 wire \top_I.branch[24].block[11].um_I.iw[15] ;
 wire \top_I.branch[24].block[11].um_I.iw[16] ;
 wire \top_I.branch[24].block[11].um_I.iw[17] ;
 wire \top_I.branch[24].block[11].um_I.iw[1] ;
 wire \top_I.branch[24].block[11].um_I.iw[2] ;
 wire \top_I.branch[24].block[11].um_I.iw[3] ;
 wire \top_I.branch[24].block[11].um_I.iw[4] ;
 wire \top_I.branch[24].block[11].um_I.iw[5] ;
 wire \top_I.branch[24].block[11].um_I.iw[6] ;
 wire \top_I.branch[24].block[11].um_I.iw[7] ;
 wire \top_I.branch[24].block[11].um_I.iw[8] ;
 wire \top_I.branch[24].block[11].um_I.iw[9] ;
 wire \top_I.branch[24].block[11].um_I.k_zero ;
 wire \top_I.branch[24].block[11].um_I.pg_vdd ;
 wire \top_I.branch[24].block[12].um_I.ana[0] ;
 wire \top_I.branch[24].block[12].um_I.ana[1] ;
 wire \top_I.branch[24].block[12].um_I.ana[2] ;
 wire \top_I.branch[24].block[12].um_I.ana[3] ;
 wire \top_I.branch[24].block[12].um_I.ana[4] ;
 wire \top_I.branch[24].block[12].um_I.ana[5] ;
 wire \top_I.branch[24].block[12].um_I.ana[6] ;
 wire \top_I.branch[24].block[12].um_I.ana[7] ;
 wire \top_I.branch[24].block[12].um_I.clk ;
 wire \top_I.branch[24].block[12].um_I.ena ;
 wire \top_I.branch[24].block[12].um_I.iw[10] ;
 wire \top_I.branch[24].block[12].um_I.iw[11] ;
 wire \top_I.branch[24].block[12].um_I.iw[12] ;
 wire \top_I.branch[24].block[12].um_I.iw[13] ;
 wire \top_I.branch[24].block[12].um_I.iw[14] ;
 wire \top_I.branch[24].block[12].um_I.iw[15] ;
 wire \top_I.branch[24].block[12].um_I.iw[16] ;
 wire \top_I.branch[24].block[12].um_I.iw[17] ;
 wire \top_I.branch[24].block[12].um_I.iw[1] ;
 wire \top_I.branch[24].block[12].um_I.iw[2] ;
 wire \top_I.branch[24].block[12].um_I.iw[3] ;
 wire \top_I.branch[24].block[12].um_I.iw[4] ;
 wire \top_I.branch[24].block[12].um_I.iw[5] ;
 wire \top_I.branch[24].block[12].um_I.iw[6] ;
 wire \top_I.branch[24].block[12].um_I.iw[7] ;
 wire \top_I.branch[24].block[12].um_I.iw[8] ;
 wire \top_I.branch[24].block[12].um_I.iw[9] ;
 wire \top_I.branch[24].block[12].um_I.k_zero ;
 wire \top_I.branch[24].block[12].um_I.pg_vdd ;
 wire \top_I.branch[24].block[13].um_I.ana[0] ;
 wire \top_I.branch[24].block[13].um_I.ana[1] ;
 wire \top_I.branch[24].block[13].um_I.ana[2] ;
 wire \top_I.branch[24].block[13].um_I.ana[3] ;
 wire \top_I.branch[24].block[13].um_I.ana[4] ;
 wire \top_I.branch[24].block[13].um_I.ana[5] ;
 wire \top_I.branch[24].block[13].um_I.ana[6] ;
 wire \top_I.branch[24].block[13].um_I.ana[7] ;
 wire \top_I.branch[24].block[13].um_I.clk ;
 wire \top_I.branch[24].block[13].um_I.ena ;
 wire \top_I.branch[24].block[13].um_I.iw[10] ;
 wire \top_I.branch[24].block[13].um_I.iw[11] ;
 wire \top_I.branch[24].block[13].um_I.iw[12] ;
 wire \top_I.branch[24].block[13].um_I.iw[13] ;
 wire \top_I.branch[24].block[13].um_I.iw[14] ;
 wire \top_I.branch[24].block[13].um_I.iw[15] ;
 wire \top_I.branch[24].block[13].um_I.iw[16] ;
 wire \top_I.branch[24].block[13].um_I.iw[17] ;
 wire \top_I.branch[24].block[13].um_I.iw[1] ;
 wire \top_I.branch[24].block[13].um_I.iw[2] ;
 wire \top_I.branch[24].block[13].um_I.iw[3] ;
 wire \top_I.branch[24].block[13].um_I.iw[4] ;
 wire \top_I.branch[24].block[13].um_I.iw[5] ;
 wire \top_I.branch[24].block[13].um_I.iw[6] ;
 wire \top_I.branch[24].block[13].um_I.iw[7] ;
 wire \top_I.branch[24].block[13].um_I.iw[8] ;
 wire \top_I.branch[24].block[13].um_I.iw[9] ;
 wire \top_I.branch[24].block[13].um_I.k_zero ;
 wire \top_I.branch[24].block[13].um_I.pg_vdd ;
 wire \top_I.branch[24].block[14].um_I.ana[0] ;
 wire \top_I.branch[24].block[14].um_I.ana[1] ;
 wire \top_I.branch[24].block[14].um_I.ana[2] ;
 wire \top_I.branch[24].block[14].um_I.ana[3] ;
 wire \top_I.branch[24].block[14].um_I.ana[4] ;
 wire \top_I.branch[24].block[14].um_I.ana[5] ;
 wire \top_I.branch[24].block[14].um_I.ana[6] ;
 wire \top_I.branch[24].block[14].um_I.ana[7] ;
 wire \top_I.branch[24].block[14].um_I.clk ;
 wire \top_I.branch[24].block[14].um_I.ena ;
 wire \top_I.branch[24].block[14].um_I.iw[10] ;
 wire \top_I.branch[24].block[14].um_I.iw[11] ;
 wire \top_I.branch[24].block[14].um_I.iw[12] ;
 wire \top_I.branch[24].block[14].um_I.iw[13] ;
 wire \top_I.branch[24].block[14].um_I.iw[14] ;
 wire \top_I.branch[24].block[14].um_I.iw[15] ;
 wire \top_I.branch[24].block[14].um_I.iw[16] ;
 wire \top_I.branch[24].block[14].um_I.iw[17] ;
 wire \top_I.branch[24].block[14].um_I.iw[1] ;
 wire \top_I.branch[24].block[14].um_I.iw[2] ;
 wire \top_I.branch[24].block[14].um_I.iw[3] ;
 wire \top_I.branch[24].block[14].um_I.iw[4] ;
 wire \top_I.branch[24].block[14].um_I.iw[5] ;
 wire \top_I.branch[24].block[14].um_I.iw[6] ;
 wire \top_I.branch[24].block[14].um_I.iw[7] ;
 wire \top_I.branch[24].block[14].um_I.iw[8] ;
 wire \top_I.branch[24].block[14].um_I.iw[9] ;
 wire \top_I.branch[24].block[14].um_I.k_zero ;
 wire \top_I.branch[24].block[14].um_I.pg_vdd ;
 wire \top_I.branch[24].block[15].um_I.ana[0] ;
 wire \top_I.branch[24].block[15].um_I.ana[1] ;
 wire \top_I.branch[24].block[15].um_I.ana[2] ;
 wire \top_I.branch[24].block[15].um_I.ana[3] ;
 wire \top_I.branch[24].block[15].um_I.ana[4] ;
 wire \top_I.branch[24].block[15].um_I.ana[5] ;
 wire \top_I.branch[24].block[15].um_I.ana[6] ;
 wire \top_I.branch[24].block[15].um_I.ana[7] ;
 wire \top_I.branch[24].block[15].um_I.clk ;
 wire \top_I.branch[24].block[15].um_I.ena ;
 wire \top_I.branch[24].block[15].um_I.iw[10] ;
 wire \top_I.branch[24].block[15].um_I.iw[11] ;
 wire \top_I.branch[24].block[15].um_I.iw[12] ;
 wire \top_I.branch[24].block[15].um_I.iw[13] ;
 wire \top_I.branch[24].block[15].um_I.iw[14] ;
 wire \top_I.branch[24].block[15].um_I.iw[15] ;
 wire \top_I.branch[24].block[15].um_I.iw[16] ;
 wire \top_I.branch[24].block[15].um_I.iw[17] ;
 wire \top_I.branch[24].block[15].um_I.iw[1] ;
 wire \top_I.branch[24].block[15].um_I.iw[2] ;
 wire \top_I.branch[24].block[15].um_I.iw[3] ;
 wire \top_I.branch[24].block[15].um_I.iw[4] ;
 wire \top_I.branch[24].block[15].um_I.iw[5] ;
 wire \top_I.branch[24].block[15].um_I.iw[6] ;
 wire \top_I.branch[24].block[15].um_I.iw[7] ;
 wire \top_I.branch[24].block[15].um_I.iw[8] ;
 wire \top_I.branch[24].block[15].um_I.iw[9] ;
 wire \top_I.branch[24].block[15].um_I.k_zero ;
 wire \top_I.branch[24].block[15].um_I.pg_vdd ;
 wire \top_I.branch[24].block[1].um_I.ana[0] ;
 wire \top_I.branch[24].block[1].um_I.ana[1] ;
 wire \top_I.branch[24].block[1].um_I.ana[2] ;
 wire \top_I.branch[24].block[1].um_I.ana[3] ;
 wire \top_I.branch[24].block[1].um_I.ana[4] ;
 wire \top_I.branch[24].block[1].um_I.ana[5] ;
 wire \top_I.branch[24].block[1].um_I.ana[6] ;
 wire \top_I.branch[24].block[1].um_I.ana[7] ;
 wire \top_I.branch[24].block[1].um_I.clk ;
 wire \top_I.branch[24].block[1].um_I.ena ;
 wire \top_I.branch[24].block[1].um_I.iw[10] ;
 wire \top_I.branch[24].block[1].um_I.iw[11] ;
 wire \top_I.branch[24].block[1].um_I.iw[12] ;
 wire \top_I.branch[24].block[1].um_I.iw[13] ;
 wire \top_I.branch[24].block[1].um_I.iw[14] ;
 wire \top_I.branch[24].block[1].um_I.iw[15] ;
 wire \top_I.branch[24].block[1].um_I.iw[16] ;
 wire \top_I.branch[24].block[1].um_I.iw[17] ;
 wire \top_I.branch[24].block[1].um_I.iw[1] ;
 wire \top_I.branch[24].block[1].um_I.iw[2] ;
 wire \top_I.branch[24].block[1].um_I.iw[3] ;
 wire \top_I.branch[24].block[1].um_I.iw[4] ;
 wire \top_I.branch[24].block[1].um_I.iw[5] ;
 wire \top_I.branch[24].block[1].um_I.iw[6] ;
 wire \top_I.branch[24].block[1].um_I.iw[7] ;
 wire \top_I.branch[24].block[1].um_I.iw[8] ;
 wire \top_I.branch[24].block[1].um_I.iw[9] ;
 wire \top_I.branch[24].block[1].um_I.k_zero ;
 wire \top_I.branch[24].block[1].um_I.pg_vdd ;
 wire \top_I.branch[24].block[2].um_I.ana[0] ;
 wire \top_I.branch[24].block[2].um_I.ana[1] ;
 wire \top_I.branch[24].block[2].um_I.ana[2] ;
 wire \top_I.branch[24].block[2].um_I.ana[3] ;
 wire \top_I.branch[24].block[2].um_I.ana[4] ;
 wire \top_I.branch[24].block[2].um_I.ana[5] ;
 wire \top_I.branch[24].block[2].um_I.ana[6] ;
 wire \top_I.branch[24].block[2].um_I.ana[7] ;
 wire \top_I.branch[24].block[2].um_I.clk ;
 wire \top_I.branch[24].block[2].um_I.ena ;
 wire \top_I.branch[24].block[2].um_I.iw[10] ;
 wire \top_I.branch[24].block[2].um_I.iw[11] ;
 wire \top_I.branch[24].block[2].um_I.iw[12] ;
 wire \top_I.branch[24].block[2].um_I.iw[13] ;
 wire \top_I.branch[24].block[2].um_I.iw[14] ;
 wire \top_I.branch[24].block[2].um_I.iw[15] ;
 wire \top_I.branch[24].block[2].um_I.iw[16] ;
 wire \top_I.branch[24].block[2].um_I.iw[17] ;
 wire \top_I.branch[24].block[2].um_I.iw[1] ;
 wire \top_I.branch[24].block[2].um_I.iw[2] ;
 wire \top_I.branch[24].block[2].um_I.iw[3] ;
 wire \top_I.branch[24].block[2].um_I.iw[4] ;
 wire \top_I.branch[24].block[2].um_I.iw[5] ;
 wire \top_I.branch[24].block[2].um_I.iw[6] ;
 wire \top_I.branch[24].block[2].um_I.iw[7] ;
 wire \top_I.branch[24].block[2].um_I.iw[8] ;
 wire \top_I.branch[24].block[2].um_I.iw[9] ;
 wire \top_I.branch[24].block[2].um_I.k_zero ;
 wire \top_I.branch[24].block[2].um_I.pg_vdd ;
 wire \top_I.branch[24].block[3].um_I.ana[0] ;
 wire \top_I.branch[24].block[3].um_I.ana[1] ;
 wire \top_I.branch[24].block[3].um_I.ana[2] ;
 wire \top_I.branch[24].block[3].um_I.ana[3] ;
 wire \top_I.branch[24].block[3].um_I.ana[4] ;
 wire \top_I.branch[24].block[3].um_I.ana[5] ;
 wire \top_I.branch[24].block[3].um_I.ana[6] ;
 wire \top_I.branch[24].block[3].um_I.ana[7] ;
 wire \top_I.branch[24].block[3].um_I.clk ;
 wire \top_I.branch[24].block[3].um_I.ena ;
 wire \top_I.branch[24].block[3].um_I.iw[10] ;
 wire \top_I.branch[24].block[3].um_I.iw[11] ;
 wire \top_I.branch[24].block[3].um_I.iw[12] ;
 wire \top_I.branch[24].block[3].um_I.iw[13] ;
 wire \top_I.branch[24].block[3].um_I.iw[14] ;
 wire \top_I.branch[24].block[3].um_I.iw[15] ;
 wire \top_I.branch[24].block[3].um_I.iw[16] ;
 wire \top_I.branch[24].block[3].um_I.iw[17] ;
 wire \top_I.branch[24].block[3].um_I.iw[1] ;
 wire \top_I.branch[24].block[3].um_I.iw[2] ;
 wire \top_I.branch[24].block[3].um_I.iw[3] ;
 wire \top_I.branch[24].block[3].um_I.iw[4] ;
 wire \top_I.branch[24].block[3].um_I.iw[5] ;
 wire \top_I.branch[24].block[3].um_I.iw[6] ;
 wire \top_I.branch[24].block[3].um_I.iw[7] ;
 wire \top_I.branch[24].block[3].um_I.iw[8] ;
 wire \top_I.branch[24].block[3].um_I.iw[9] ;
 wire \top_I.branch[24].block[3].um_I.k_zero ;
 wire \top_I.branch[24].block[3].um_I.pg_vdd ;
 wire \top_I.branch[24].block[4].um_I.ana[0] ;
 wire \top_I.branch[24].block[4].um_I.ana[1] ;
 wire \top_I.branch[24].block[4].um_I.ana[2] ;
 wire \top_I.branch[24].block[4].um_I.ana[3] ;
 wire \top_I.branch[24].block[4].um_I.ana[4] ;
 wire \top_I.branch[24].block[4].um_I.ana[5] ;
 wire \top_I.branch[24].block[4].um_I.ana[6] ;
 wire \top_I.branch[24].block[4].um_I.ana[7] ;
 wire \top_I.branch[24].block[4].um_I.clk ;
 wire \top_I.branch[24].block[4].um_I.ena ;
 wire \top_I.branch[24].block[4].um_I.iw[10] ;
 wire \top_I.branch[24].block[4].um_I.iw[11] ;
 wire \top_I.branch[24].block[4].um_I.iw[12] ;
 wire \top_I.branch[24].block[4].um_I.iw[13] ;
 wire \top_I.branch[24].block[4].um_I.iw[14] ;
 wire \top_I.branch[24].block[4].um_I.iw[15] ;
 wire \top_I.branch[24].block[4].um_I.iw[16] ;
 wire \top_I.branch[24].block[4].um_I.iw[17] ;
 wire \top_I.branch[24].block[4].um_I.iw[1] ;
 wire \top_I.branch[24].block[4].um_I.iw[2] ;
 wire \top_I.branch[24].block[4].um_I.iw[3] ;
 wire \top_I.branch[24].block[4].um_I.iw[4] ;
 wire \top_I.branch[24].block[4].um_I.iw[5] ;
 wire \top_I.branch[24].block[4].um_I.iw[6] ;
 wire \top_I.branch[24].block[4].um_I.iw[7] ;
 wire \top_I.branch[24].block[4].um_I.iw[8] ;
 wire \top_I.branch[24].block[4].um_I.iw[9] ;
 wire \top_I.branch[24].block[4].um_I.k_zero ;
 wire \top_I.branch[24].block[4].um_I.pg_vdd ;
 wire \top_I.branch[24].block[5].um_I.ana[0] ;
 wire \top_I.branch[24].block[5].um_I.ana[1] ;
 wire \top_I.branch[24].block[5].um_I.ana[2] ;
 wire \top_I.branch[24].block[5].um_I.ana[3] ;
 wire \top_I.branch[24].block[5].um_I.ana[4] ;
 wire \top_I.branch[24].block[5].um_I.ana[5] ;
 wire \top_I.branch[24].block[5].um_I.ana[6] ;
 wire \top_I.branch[24].block[5].um_I.ana[7] ;
 wire \top_I.branch[24].block[5].um_I.clk ;
 wire \top_I.branch[24].block[5].um_I.ena ;
 wire \top_I.branch[24].block[5].um_I.iw[10] ;
 wire \top_I.branch[24].block[5].um_I.iw[11] ;
 wire \top_I.branch[24].block[5].um_I.iw[12] ;
 wire \top_I.branch[24].block[5].um_I.iw[13] ;
 wire \top_I.branch[24].block[5].um_I.iw[14] ;
 wire \top_I.branch[24].block[5].um_I.iw[15] ;
 wire \top_I.branch[24].block[5].um_I.iw[16] ;
 wire \top_I.branch[24].block[5].um_I.iw[17] ;
 wire \top_I.branch[24].block[5].um_I.iw[1] ;
 wire \top_I.branch[24].block[5].um_I.iw[2] ;
 wire \top_I.branch[24].block[5].um_I.iw[3] ;
 wire \top_I.branch[24].block[5].um_I.iw[4] ;
 wire \top_I.branch[24].block[5].um_I.iw[5] ;
 wire \top_I.branch[24].block[5].um_I.iw[6] ;
 wire \top_I.branch[24].block[5].um_I.iw[7] ;
 wire \top_I.branch[24].block[5].um_I.iw[8] ;
 wire \top_I.branch[24].block[5].um_I.iw[9] ;
 wire \top_I.branch[24].block[5].um_I.k_zero ;
 wire \top_I.branch[24].block[5].um_I.pg_vdd ;
 wire \top_I.branch[24].block[6].um_I.ana[0] ;
 wire \top_I.branch[24].block[6].um_I.ana[1] ;
 wire \top_I.branch[24].block[6].um_I.ana[2] ;
 wire \top_I.branch[24].block[6].um_I.ana[3] ;
 wire \top_I.branch[24].block[6].um_I.ana[4] ;
 wire \top_I.branch[24].block[6].um_I.ana[5] ;
 wire \top_I.branch[24].block[6].um_I.ana[6] ;
 wire \top_I.branch[24].block[6].um_I.ana[7] ;
 wire \top_I.branch[24].block[6].um_I.clk ;
 wire \top_I.branch[24].block[6].um_I.ena ;
 wire \top_I.branch[24].block[6].um_I.iw[10] ;
 wire \top_I.branch[24].block[6].um_I.iw[11] ;
 wire \top_I.branch[24].block[6].um_I.iw[12] ;
 wire \top_I.branch[24].block[6].um_I.iw[13] ;
 wire \top_I.branch[24].block[6].um_I.iw[14] ;
 wire \top_I.branch[24].block[6].um_I.iw[15] ;
 wire \top_I.branch[24].block[6].um_I.iw[16] ;
 wire \top_I.branch[24].block[6].um_I.iw[17] ;
 wire \top_I.branch[24].block[6].um_I.iw[1] ;
 wire \top_I.branch[24].block[6].um_I.iw[2] ;
 wire \top_I.branch[24].block[6].um_I.iw[3] ;
 wire \top_I.branch[24].block[6].um_I.iw[4] ;
 wire \top_I.branch[24].block[6].um_I.iw[5] ;
 wire \top_I.branch[24].block[6].um_I.iw[6] ;
 wire \top_I.branch[24].block[6].um_I.iw[7] ;
 wire \top_I.branch[24].block[6].um_I.iw[8] ;
 wire \top_I.branch[24].block[6].um_I.iw[9] ;
 wire \top_I.branch[24].block[6].um_I.k_zero ;
 wire \top_I.branch[24].block[6].um_I.pg_vdd ;
 wire \top_I.branch[24].block[7].um_I.ana[0] ;
 wire \top_I.branch[24].block[7].um_I.ana[1] ;
 wire \top_I.branch[24].block[7].um_I.ana[2] ;
 wire \top_I.branch[24].block[7].um_I.ana[3] ;
 wire \top_I.branch[24].block[7].um_I.ana[4] ;
 wire \top_I.branch[24].block[7].um_I.ana[5] ;
 wire \top_I.branch[24].block[7].um_I.ana[6] ;
 wire \top_I.branch[24].block[7].um_I.ana[7] ;
 wire \top_I.branch[24].block[7].um_I.clk ;
 wire \top_I.branch[24].block[7].um_I.ena ;
 wire \top_I.branch[24].block[7].um_I.iw[10] ;
 wire \top_I.branch[24].block[7].um_I.iw[11] ;
 wire \top_I.branch[24].block[7].um_I.iw[12] ;
 wire \top_I.branch[24].block[7].um_I.iw[13] ;
 wire \top_I.branch[24].block[7].um_I.iw[14] ;
 wire \top_I.branch[24].block[7].um_I.iw[15] ;
 wire \top_I.branch[24].block[7].um_I.iw[16] ;
 wire \top_I.branch[24].block[7].um_I.iw[17] ;
 wire \top_I.branch[24].block[7].um_I.iw[1] ;
 wire \top_I.branch[24].block[7].um_I.iw[2] ;
 wire \top_I.branch[24].block[7].um_I.iw[3] ;
 wire \top_I.branch[24].block[7].um_I.iw[4] ;
 wire \top_I.branch[24].block[7].um_I.iw[5] ;
 wire \top_I.branch[24].block[7].um_I.iw[6] ;
 wire \top_I.branch[24].block[7].um_I.iw[7] ;
 wire \top_I.branch[24].block[7].um_I.iw[8] ;
 wire \top_I.branch[24].block[7].um_I.iw[9] ;
 wire \top_I.branch[24].block[7].um_I.k_zero ;
 wire \top_I.branch[24].block[7].um_I.pg_vdd ;
 wire \top_I.branch[24].block[8].um_I.ana[0] ;
 wire \top_I.branch[24].block[8].um_I.ana[1] ;
 wire \top_I.branch[24].block[8].um_I.ana[2] ;
 wire \top_I.branch[24].block[8].um_I.ana[3] ;
 wire \top_I.branch[24].block[8].um_I.ana[4] ;
 wire \top_I.branch[24].block[8].um_I.ana[5] ;
 wire \top_I.branch[24].block[8].um_I.ana[6] ;
 wire \top_I.branch[24].block[8].um_I.ana[7] ;
 wire \top_I.branch[24].block[8].um_I.clk ;
 wire \top_I.branch[24].block[8].um_I.ena ;
 wire \top_I.branch[24].block[8].um_I.iw[10] ;
 wire \top_I.branch[24].block[8].um_I.iw[11] ;
 wire \top_I.branch[24].block[8].um_I.iw[12] ;
 wire \top_I.branch[24].block[8].um_I.iw[13] ;
 wire \top_I.branch[24].block[8].um_I.iw[14] ;
 wire \top_I.branch[24].block[8].um_I.iw[15] ;
 wire \top_I.branch[24].block[8].um_I.iw[16] ;
 wire \top_I.branch[24].block[8].um_I.iw[17] ;
 wire \top_I.branch[24].block[8].um_I.iw[1] ;
 wire \top_I.branch[24].block[8].um_I.iw[2] ;
 wire \top_I.branch[24].block[8].um_I.iw[3] ;
 wire \top_I.branch[24].block[8].um_I.iw[4] ;
 wire \top_I.branch[24].block[8].um_I.iw[5] ;
 wire \top_I.branch[24].block[8].um_I.iw[6] ;
 wire \top_I.branch[24].block[8].um_I.iw[7] ;
 wire \top_I.branch[24].block[8].um_I.iw[8] ;
 wire \top_I.branch[24].block[8].um_I.iw[9] ;
 wire \top_I.branch[24].block[8].um_I.k_zero ;
 wire \top_I.branch[24].block[8].um_I.pg_vdd ;
 wire \top_I.branch[24].block[9].um_I.ana[0] ;
 wire \top_I.branch[24].block[9].um_I.ana[1] ;
 wire \top_I.branch[24].block[9].um_I.ana[2] ;
 wire \top_I.branch[24].block[9].um_I.ana[3] ;
 wire \top_I.branch[24].block[9].um_I.ana[4] ;
 wire \top_I.branch[24].block[9].um_I.ana[5] ;
 wire \top_I.branch[24].block[9].um_I.ana[6] ;
 wire \top_I.branch[24].block[9].um_I.ana[7] ;
 wire \top_I.branch[24].block[9].um_I.clk ;
 wire \top_I.branch[24].block[9].um_I.ena ;
 wire \top_I.branch[24].block[9].um_I.iw[10] ;
 wire \top_I.branch[24].block[9].um_I.iw[11] ;
 wire \top_I.branch[24].block[9].um_I.iw[12] ;
 wire \top_I.branch[24].block[9].um_I.iw[13] ;
 wire \top_I.branch[24].block[9].um_I.iw[14] ;
 wire \top_I.branch[24].block[9].um_I.iw[15] ;
 wire \top_I.branch[24].block[9].um_I.iw[16] ;
 wire \top_I.branch[24].block[9].um_I.iw[17] ;
 wire \top_I.branch[24].block[9].um_I.iw[1] ;
 wire \top_I.branch[24].block[9].um_I.iw[2] ;
 wire \top_I.branch[24].block[9].um_I.iw[3] ;
 wire \top_I.branch[24].block[9].um_I.iw[4] ;
 wire \top_I.branch[24].block[9].um_I.iw[5] ;
 wire \top_I.branch[24].block[9].um_I.iw[6] ;
 wire \top_I.branch[24].block[9].um_I.iw[7] ;
 wire \top_I.branch[24].block[9].um_I.iw[8] ;
 wire \top_I.branch[24].block[9].um_I.iw[9] ;
 wire \top_I.branch[24].block[9].um_I.k_zero ;
 wire \top_I.branch[24].block[9].um_I.pg_vdd ;
 wire \top_I.branch[24].l_addr[0] ;
 wire \top_I.branch[24].l_addr[2] ;
 wire \top_I.branch[25].block[0].um_I.ana[0] ;
 wire \top_I.branch[25].block[0].um_I.ana[1] ;
 wire \top_I.branch[25].block[0].um_I.ana[2] ;
 wire \top_I.branch[25].block[0].um_I.ana[3] ;
 wire \top_I.branch[25].block[0].um_I.ana[4] ;
 wire \top_I.branch[25].block[0].um_I.ana[5] ;
 wire \top_I.branch[25].block[0].um_I.ana[6] ;
 wire \top_I.branch[25].block[0].um_I.ana[7] ;
 wire \top_I.branch[25].block[0].um_I.clk ;
 wire \top_I.branch[25].block[0].um_I.ena ;
 wire \top_I.branch[25].block[0].um_I.iw[10] ;
 wire \top_I.branch[25].block[0].um_I.iw[11] ;
 wire \top_I.branch[25].block[0].um_I.iw[12] ;
 wire \top_I.branch[25].block[0].um_I.iw[13] ;
 wire \top_I.branch[25].block[0].um_I.iw[14] ;
 wire \top_I.branch[25].block[0].um_I.iw[15] ;
 wire \top_I.branch[25].block[0].um_I.iw[16] ;
 wire \top_I.branch[25].block[0].um_I.iw[17] ;
 wire \top_I.branch[25].block[0].um_I.iw[1] ;
 wire \top_I.branch[25].block[0].um_I.iw[2] ;
 wire \top_I.branch[25].block[0].um_I.iw[3] ;
 wire \top_I.branch[25].block[0].um_I.iw[4] ;
 wire \top_I.branch[25].block[0].um_I.iw[5] ;
 wire \top_I.branch[25].block[0].um_I.iw[6] ;
 wire \top_I.branch[25].block[0].um_I.iw[7] ;
 wire \top_I.branch[25].block[0].um_I.iw[8] ;
 wire \top_I.branch[25].block[0].um_I.iw[9] ;
 wire \top_I.branch[25].block[0].um_I.k_zero ;
 wire \top_I.branch[25].block[0].um_I.pg_vdd ;
 wire \top_I.branch[25].block[10].um_I.ana[0] ;
 wire \top_I.branch[25].block[10].um_I.ana[1] ;
 wire \top_I.branch[25].block[10].um_I.ana[2] ;
 wire \top_I.branch[25].block[10].um_I.ana[3] ;
 wire \top_I.branch[25].block[10].um_I.ana[4] ;
 wire \top_I.branch[25].block[10].um_I.ana[5] ;
 wire \top_I.branch[25].block[10].um_I.ana[6] ;
 wire \top_I.branch[25].block[10].um_I.ana[7] ;
 wire \top_I.branch[25].block[10].um_I.clk ;
 wire \top_I.branch[25].block[10].um_I.ena ;
 wire \top_I.branch[25].block[10].um_I.iw[10] ;
 wire \top_I.branch[25].block[10].um_I.iw[11] ;
 wire \top_I.branch[25].block[10].um_I.iw[12] ;
 wire \top_I.branch[25].block[10].um_I.iw[13] ;
 wire \top_I.branch[25].block[10].um_I.iw[14] ;
 wire \top_I.branch[25].block[10].um_I.iw[15] ;
 wire \top_I.branch[25].block[10].um_I.iw[16] ;
 wire \top_I.branch[25].block[10].um_I.iw[17] ;
 wire \top_I.branch[25].block[10].um_I.iw[1] ;
 wire \top_I.branch[25].block[10].um_I.iw[2] ;
 wire \top_I.branch[25].block[10].um_I.iw[3] ;
 wire \top_I.branch[25].block[10].um_I.iw[4] ;
 wire \top_I.branch[25].block[10].um_I.iw[5] ;
 wire \top_I.branch[25].block[10].um_I.iw[6] ;
 wire \top_I.branch[25].block[10].um_I.iw[7] ;
 wire \top_I.branch[25].block[10].um_I.iw[8] ;
 wire \top_I.branch[25].block[10].um_I.iw[9] ;
 wire \top_I.branch[25].block[10].um_I.k_zero ;
 wire \top_I.branch[25].block[10].um_I.pg_vdd ;
 wire \top_I.branch[25].block[11].um_I.ana[0] ;
 wire \top_I.branch[25].block[11].um_I.ana[1] ;
 wire \top_I.branch[25].block[11].um_I.ana[2] ;
 wire \top_I.branch[25].block[11].um_I.ana[3] ;
 wire \top_I.branch[25].block[11].um_I.ana[4] ;
 wire \top_I.branch[25].block[11].um_I.ana[5] ;
 wire \top_I.branch[25].block[11].um_I.ana[6] ;
 wire \top_I.branch[25].block[11].um_I.ana[7] ;
 wire \top_I.branch[25].block[11].um_I.clk ;
 wire \top_I.branch[25].block[11].um_I.ena ;
 wire \top_I.branch[25].block[11].um_I.iw[10] ;
 wire \top_I.branch[25].block[11].um_I.iw[11] ;
 wire \top_I.branch[25].block[11].um_I.iw[12] ;
 wire \top_I.branch[25].block[11].um_I.iw[13] ;
 wire \top_I.branch[25].block[11].um_I.iw[14] ;
 wire \top_I.branch[25].block[11].um_I.iw[15] ;
 wire \top_I.branch[25].block[11].um_I.iw[16] ;
 wire \top_I.branch[25].block[11].um_I.iw[17] ;
 wire \top_I.branch[25].block[11].um_I.iw[1] ;
 wire \top_I.branch[25].block[11].um_I.iw[2] ;
 wire \top_I.branch[25].block[11].um_I.iw[3] ;
 wire \top_I.branch[25].block[11].um_I.iw[4] ;
 wire \top_I.branch[25].block[11].um_I.iw[5] ;
 wire \top_I.branch[25].block[11].um_I.iw[6] ;
 wire \top_I.branch[25].block[11].um_I.iw[7] ;
 wire \top_I.branch[25].block[11].um_I.iw[8] ;
 wire \top_I.branch[25].block[11].um_I.iw[9] ;
 wire \top_I.branch[25].block[11].um_I.k_zero ;
 wire \top_I.branch[25].block[11].um_I.pg_vdd ;
 wire \top_I.branch[25].block[12].um_I.ana[0] ;
 wire \top_I.branch[25].block[12].um_I.ana[1] ;
 wire \top_I.branch[25].block[12].um_I.ana[2] ;
 wire \top_I.branch[25].block[12].um_I.ana[3] ;
 wire \top_I.branch[25].block[12].um_I.ana[4] ;
 wire \top_I.branch[25].block[12].um_I.ana[5] ;
 wire \top_I.branch[25].block[12].um_I.ana[6] ;
 wire \top_I.branch[25].block[12].um_I.ana[7] ;
 wire \top_I.branch[25].block[12].um_I.clk ;
 wire \top_I.branch[25].block[12].um_I.ena ;
 wire \top_I.branch[25].block[12].um_I.iw[10] ;
 wire \top_I.branch[25].block[12].um_I.iw[11] ;
 wire \top_I.branch[25].block[12].um_I.iw[12] ;
 wire \top_I.branch[25].block[12].um_I.iw[13] ;
 wire \top_I.branch[25].block[12].um_I.iw[14] ;
 wire \top_I.branch[25].block[12].um_I.iw[15] ;
 wire \top_I.branch[25].block[12].um_I.iw[16] ;
 wire \top_I.branch[25].block[12].um_I.iw[17] ;
 wire \top_I.branch[25].block[12].um_I.iw[1] ;
 wire \top_I.branch[25].block[12].um_I.iw[2] ;
 wire \top_I.branch[25].block[12].um_I.iw[3] ;
 wire \top_I.branch[25].block[12].um_I.iw[4] ;
 wire \top_I.branch[25].block[12].um_I.iw[5] ;
 wire \top_I.branch[25].block[12].um_I.iw[6] ;
 wire \top_I.branch[25].block[12].um_I.iw[7] ;
 wire \top_I.branch[25].block[12].um_I.iw[8] ;
 wire \top_I.branch[25].block[12].um_I.iw[9] ;
 wire \top_I.branch[25].block[12].um_I.k_zero ;
 wire \top_I.branch[25].block[12].um_I.pg_vdd ;
 wire \top_I.branch[25].block[13].um_I.ana[0] ;
 wire \top_I.branch[25].block[13].um_I.ana[1] ;
 wire \top_I.branch[25].block[13].um_I.ana[2] ;
 wire \top_I.branch[25].block[13].um_I.ana[3] ;
 wire \top_I.branch[25].block[13].um_I.ana[4] ;
 wire \top_I.branch[25].block[13].um_I.ana[5] ;
 wire \top_I.branch[25].block[13].um_I.ana[6] ;
 wire \top_I.branch[25].block[13].um_I.ana[7] ;
 wire \top_I.branch[25].block[13].um_I.clk ;
 wire \top_I.branch[25].block[13].um_I.ena ;
 wire \top_I.branch[25].block[13].um_I.iw[10] ;
 wire \top_I.branch[25].block[13].um_I.iw[11] ;
 wire \top_I.branch[25].block[13].um_I.iw[12] ;
 wire \top_I.branch[25].block[13].um_I.iw[13] ;
 wire \top_I.branch[25].block[13].um_I.iw[14] ;
 wire \top_I.branch[25].block[13].um_I.iw[15] ;
 wire \top_I.branch[25].block[13].um_I.iw[16] ;
 wire \top_I.branch[25].block[13].um_I.iw[17] ;
 wire \top_I.branch[25].block[13].um_I.iw[1] ;
 wire \top_I.branch[25].block[13].um_I.iw[2] ;
 wire \top_I.branch[25].block[13].um_I.iw[3] ;
 wire \top_I.branch[25].block[13].um_I.iw[4] ;
 wire \top_I.branch[25].block[13].um_I.iw[5] ;
 wire \top_I.branch[25].block[13].um_I.iw[6] ;
 wire \top_I.branch[25].block[13].um_I.iw[7] ;
 wire \top_I.branch[25].block[13].um_I.iw[8] ;
 wire \top_I.branch[25].block[13].um_I.iw[9] ;
 wire \top_I.branch[25].block[13].um_I.k_zero ;
 wire \top_I.branch[25].block[13].um_I.pg_vdd ;
 wire \top_I.branch[25].block[14].um_I.ana[0] ;
 wire \top_I.branch[25].block[14].um_I.ana[1] ;
 wire \top_I.branch[25].block[14].um_I.ana[2] ;
 wire \top_I.branch[25].block[14].um_I.ana[3] ;
 wire \top_I.branch[25].block[14].um_I.ana[4] ;
 wire \top_I.branch[25].block[14].um_I.ana[5] ;
 wire \top_I.branch[25].block[14].um_I.ana[6] ;
 wire \top_I.branch[25].block[14].um_I.ana[7] ;
 wire \top_I.branch[25].block[14].um_I.clk ;
 wire \top_I.branch[25].block[14].um_I.ena ;
 wire \top_I.branch[25].block[14].um_I.iw[10] ;
 wire \top_I.branch[25].block[14].um_I.iw[11] ;
 wire \top_I.branch[25].block[14].um_I.iw[12] ;
 wire \top_I.branch[25].block[14].um_I.iw[13] ;
 wire \top_I.branch[25].block[14].um_I.iw[14] ;
 wire \top_I.branch[25].block[14].um_I.iw[15] ;
 wire \top_I.branch[25].block[14].um_I.iw[16] ;
 wire \top_I.branch[25].block[14].um_I.iw[17] ;
 wire \top_I.branch[25].block[14].um_I.iw[1] ;
 wire \top_I.branch[25].block[14].um_I.iw[2] ;
 wire \top_I.branch[25].block[14].um_I.iw[3] ;
 wire \top_I.branch[25].block[14].um_I.iw[4] ;
 wire \top_I.branch[25].block[14].um_I.iw[5] ;
 wire \top_I.branch[25].block[14].um_I.iw[6] ;
 wire \top_I.branch[25].block[14].um_I.iw[7] ;
 wire \top_I.branch[25].block[14].um_I.iw[8] ;
 wire \top_I.branch[25].block[14].um_I.iw[9] ;
 wire \top_I.branch[25].block[14].um_I.k_zero ;
 wire \top_I.branch[25].block[14].um_I.pg_vdd ;
 wire \top_I.branch[25].block[15].um_I.ana[0] ;
 wire \top_I.branch[25].block[15].um_I.ana[1] ;
 wire \top_I.branch[25].block[15].um_I.ana[2] ;
 wire \top_I.branch[25].block[15].um_I.ana[3] ;
 wire \top_I.branch[25].block[15].um_I.ana[4] ;
 wire \top_I.branch[25].block[15].um_I.ana[5] ;
 wire \top_I.branch[25].block[15].um_I.ana[6] ;
 wire \top_I.branch[25].block[15].um_I.ana[7] ;
 wire \top_I.branch[25].block[15].um_I.clk ;
 wire \top_I.branch[25].block[15].um_I.ena ;
 wire \top_I.branch[25].block[15].um_I.iw[10] ;
 wire \top_I.branch[25].block[15].um_I.iw[11] ;
 wire \top_I.branch[25].block[15].um_I.iw[12] ;
 wire \top_I.branch[25].block[15].um_I.iw[13] ;
 wire \top_I.branch[25].block[15].um_I.iw[14] ;
 wire \top_I.branch[25].block[15].um_I.iw[15] ;
 wire \top_I.branch[25].block[15].um_I.iw[16] ;
 wire \top_I.branch[25].block[15].um_I.iw[17] ;
 wire \top_I.branch[25].block[15].um_I.iw[1] ;
 wire \top_I.branch[25].block[15].um_I.iw[2] ;
 wire \top_I.branch[25].block[15].um_I.iw[3] ;
 wire \top_I.branch[25].block[15].um_I.iw[4] ;
 wire \top_I.branch[25].block[15].um_I.iw[5] ;
 wire \top_I.branch[25].block[15].um_I.iw[6] ;
 wire \top_I.branch[25].block[15].um_I.iw[7] ;
 wire \top_I.branch[25].block[15].um_I.iw[8] ;
 wire \top_I.branch[25].block[15].um_I.iw[9] ;
 wire \top_I.branch[25].block[15].um_I.k_zero ;
 wire \top_I.branch[25].block[15].um_I.pg_vdd ;
 wire \top_I.branch[25].block[1].um_I.ana[0] ;
 wire \top_I.branch[25].block[1].um_I.ana[1] ;
 wire \top_I.branch[25].block[1].um_I.ana[2] ;
 wire \top_I.branch[25].block[1].um_I.ana[3] ;
 wire \top_I.branch[25].block[1].um_I.ana[4] ;
 wire \top_I.branch[25].block[1].um_I.ana[5] ;
 wire \top_I.branch[25].block[1].um_I.ana[6] ;
 wire \top_I.branch[25].block[1].um_I.ana[7] ;
 wire \top_I.branch[25].block[1].um_I.clk ;
 wire \top_I.branch[25].block[1].um_I.ena ;
 wire \top_I.branch[25].block[1].um_I.iw[10] ;
 wire \top_I.branch[25].block[1].um_I.iw[11] ;
 wire \top_I.branch[25].block[1].um_I.iw[12] ;
 wire \top_I.branch[25].block[1].um_I.iw[13] ;
 wire \top_I.branch[25].block[1].um_I.iw[14] ;
 wire \top_I.branch[25].block[1].um_I.iw[15] ;
 wire \top_I.branch[25].block[1].um_I.iw[16] ;
 wire \top_I.branch[25].block[1].um_I.iw[17] ;
 wire \top_I.branch[25].block[1].um_I.iw[1] ;
 wire \top_I.branch[25].block[1].um_I.iw[2] ;
 wire \top_I.branch[25].block[1].um_I.iw[3] ;
 wire \top_I.branch[25].block[1].um_I.iw[4] ;
 wire \top_I.branch[25].block[1].um_I.iw[5] ;
 wire \top_I.branch[25].block[1].um_I.iw[6] ;
 wire \top_I.branch[25].block[1].um_I.iw[7] ;
 wire \top_I.branch[25].block[1].um_I.iw[8] ;
 wire \top_I.branch[25].block[1].um_I.iw[9] ;
 wire \top_I.branch[25].block[1].um_I.k_zero ;
 wire \top_I.branch[25].block[1].um_I.pg_vdd ;
 wire \top_I.branch[25].block[2].um_I.ana[0] ;
 wire \top_I.branch[25].block[2].um_I.ana[1] ;
 wire \top_I.branch[25].block[2].um_I.ana[2] ;
 wire \top_I.branch[25].block[2].um_I.ana[3] ;
 wire \top_I.branch[25].block[2].um_I.ana[4] ;
 wire \top_I.branch[25].block[2].um_I.ana[5] ;
 wire \top_I.branch[25].block[2].um_I.ana[6] ;
 wire \top_I.branch[25].block[2].um_I.ana[7] ;
 wire \top_I.branch[25].block[2].um_I.clk ;
 wire \top_I.branch[25].block[2].um_I.ena ;
 wire \top_I.branch[25].block[2].um_I.iw[10] ;
 wire \top_I.branch[25].block[2].um_I.iw[11] ;
 wire \top_I.branch[25].block[2].um_I.iw[12] ;
 wire \top_I.branch[25].block[2].um_I.iw[13] ;
 wire \top_I.branch[25].block[2].um_I.iw[14] ;
 wire \top_I.branch[25].block[2].um_I.iw[15] ;
 wire \top_I.branch[25].block[2].um_I.iw[16] ;
 wire \top_I.branch[25].block[2].um_I.iw[17] ;
 wire \top_I.branch[25].block[2].um_I.iw[1] ;
 wire \top_I.branch[25].block[2].um_I.iw[2] ;
 wire \top_I.branch[25].block[2].um_I.iw[3] ;
 wire \top_I.branch[25].block[2].um_I.iw[4] ;
 wire \top_I.branch[25].block[2].um_I.iw[5] ;
 wire \top_I.branch[25].block[2].um_I.iw[6] ;
 wire \top_I.branch[25].block[2].um_I.iw[7] ;
 wire \top_I.branch[25].block[2].um_I.iw[8] ;
 wire \top_I.branch[25].block[2].um_I.iw[9] ;
 wire \top_I.branch[25].block[2].um_I.k_zero ;
 wire \top_I.branch[25].block[2].um_I.pg_vdd ;
 wire \top_I.branch[25].block[3].um_I.ana[0] ;
 wire \top_I.branch[25].block[3].um_I.ana[1] ;
 wire \top_I.branch[25].block[3].um_I.ana[2] ;
 wire \top_I.branch[25].block[3].um_I.ana[3] ;
 wire \top_I.branch[25].block[3].um_I.ana[4] ;
 wire \top_I.branch[25].block[3].um_I.ana[5] ;
 wire \top_I.branch[25].block[3].um_I.ana[6] ;
 wire \top_I.branch[25].block[3].um_I.ana[7] ;
 wire \top_I.branch[25].block[3].um_I.clk ;
 wire \top_I.branch[25].block[3].um_I.ena ;
 wire \top_I.branch[25].block[3].um_I.iw[10] ;
 wire \top_I.branch[25].block[3].um_I.iw[11] ;
 wire \top_I.branch[25].block[3].um_I.iw[12] ;
 wire \top_I.branch[25].block[3].um_I.iw[13] ;
 wire \top_I.branch[25].block[3].um_I.iw[14] ;
 wire \top_I.branch[25].block[3].um_I.iw[15] ;
 wire \top_I.branch[25].block[3].um_I.iw[16] ;
 wire \top_I.branch[25].block[3].um_I.iw[17] ;
 wire \top_I.branch[25].block[3].um_I.iw[1] ;
 wire \top_I.branch[25].block[3].um_I.iw[2] ;
 wire \top_I.branch[25].block[3].um_I.iw[3] ;
 wire \top_I.branch[25].block[3].um_I.iw[4] ;
 wire \top_I.branch[25].block[3].um_I.iw[5] ;
 wire \top_I.branch[25].block[3].um_I.iw[6] ;
 wire \top_I.branch[25].block[3].um_I.iw[7] ;
 wire \top_I.branch[25].block[3].um_I.iw[8] ;
 wire \top_I.branch[25].block[3].um_I.iw[9] ;
 wire \top_I.branch[25].block[3].um_I.k_zero ;
 wire \top_I.branch[25].block[3].um_I.pg_vdd ;
 wire \top_I.branch[25].block[4].um_I.ana[0] ;
 wire \top_I.branch[25].block[4].um_I.ana[1] ;
 wire \top_I.branch[25].block[4].um_I.ana[2] ;
 wire \top_I.branch[25].block[4].um_I.ana[3] ;
 wire \top_I.branch[25].block[4].um_I.ana[4] ;
 wire \top_I.branch[25].block[4].um_I.ana[5] ;
 wire \top_I.branch[25].block[4].um_I.ana[6] ;
 wire \top_I.branch[25].block[4].um_I.ana[7] ;
 wire \top_I.branch[25].block[4].um_I.clk ;
 wire \top_I.branch[25].block[4].um_I.ena ;
 wire \top_I.branch[25].block[4].um_I.iw[10] ;
 wire \top_I.branch[25].block[4].um_I.iw[11] ;
 wire \top_I.branch[25].block[4].um_I.iw[12] ;
 wire \top_I.branch[25].block[4].um_I.iw[13] ;
 wire \top_I.branch[25].block[4].um_I.iw[14] ;
 wire \top_I.branch[25].block[4].um_I.iw[15] ;
 wire \top_I.branch[25].block[4].um_I.iw[16] ;
 wire \top_I.branch[25].block[4].um_I.iw[17] ;
 wire \top_I.branch[25].block[4].um_I.iw[1] ;
 wire \top_I.branch[25].block[4].um_I.iw[2] ;
 wire \top_I.branch[25].block[4].um_I.iw[3] ;
 wire \top_I.branch[25].block[4].um_I.iw[4] ;
 wire \top_I.branch[25].block[4].um_I.iw[5] ;
 wire \top_I.branch[25].block[4].um_I.iw[6] ;
 wire \top_I.branch[25].block[4].um_I.iw[7] ;
 wire \top_I.branch[25].block[4].um_I.iw[8] ;
 wire \top_I.branch[25].block[4].um_I.iw[9] ;
 wire \top_I.branch[25].block[4].um_I.k_zero ;
 wire \top_I.branch[25].block[4].um_I.pg_vdd ;
 wire \top_I.branch[25].block[5].um_I.ana[0] ;
 wire \top_I.branch[25].block[5].um_I.ana[1] ;
 wire \top_I.branch[25].block[5].um_I.ana[2] ;
 wire \top_I.branch[25].block[5].um_I.ana[3] ;
 wire \top_I.branch[25].block[5].um_I.ana[4] ;
 wire \top_I.branch[25].block[5].um_I.ana[5] ;
 wire \top_I.branch[25].block[5].um_I.ana[6] ;
 wire \top_I.branch[25].block[5].um_I.ana[7] ;
 wire \top_I.branch[25].block[5].um_I.clk ;
 wire \top_I.branch[25].block[5].um_I.ena ;
 wire \top_I.branch[25].block[5].um_I.iw[10] ;
 wire \top_I.branch[25].block[5].um_I.iw[11] ;
 wire \top_I.branch[25].block[5].um_I.iw[12] ;
 wire \top_I.branch[25].block[5].um_I.iw[13] ;
 wire \top_I.branch[25].block[5].um_I.iw[14] ;
 wire \top_I.branch[25].block[5].um_I.iw[15] ;
 wire \top_I.branch[25].block[5].um_I.iw[16] ;
 wire \top_I.branch[25].block[5].um_I.iw[17] ;
 wire \top_I.branch[25].block[5].um_I.iw[1] ;
 wire \top_I.branch[25].block[5].um_I.iw[2] ;
 wire \top_I.branch[25].block[5].um_I.iw[3] ;
 wire \top_I.branch[25].block[5].um_I.iw[4] ;
 wire \top_I.branch[25].block[5].um_I.iw[5] ;
 wire \top_I.branch[25].block[5].um_I.iw[6] ;
 wire \top_I.branch[25].block[5].um_I.iw[7] ;
 wire \top_I.branch[25].block[5].um_I.iw[8] ;
 wire \top_I.branch[25].block[5].um_I.iw[9] ;
 wire \top_I.branch[25].block[5].um_I.k_zero ;
 wire \top_I.branch[25].block[5].um_I.pg_vdd ;
 wire \top_I.branch[25].block[6].um_I.ana[0] ;
 wire \top_I.branch[25].block[6].um_I.ana[1] ;
 wire \top_I.branch[25].block[6].um_I.ana[2] ;
 wire \top_I.branch[25].block[6].um_I.ana[3] ;
 wire \top_I.branch[25].block[6].um_I.ana[4] ;
 wire \top_I.branch[25].block[6].um_I.ana[5] ;
 wire \top_I.branch[25].block[6].um_I.ana[6] ;
 wire \top_I.branch[25].block[6].um_I.ana[7] ;
 wire \top_I.branch[25].block[6].um_I.clk ;
 wire \top_I.branch[25].block[6].um_I.ena ;
 wire \top_I.branch[25].block[6].um_I.iw[10] ;
 wire \top_I.branch[25].block[6].um_I.iw[11] ;
 wire \top_I.branch[25].block[6].um_I.iw[12] ;
 wire \top_I.branch[25].block[6].um_I.iw[13] ;
 wire \top_I.branch[25].block[6].um_I.iw[14] ;
 wire \top_I.branch[25].block[6].um_I.iw[15] ;
 wire \top_I.branch[25].block[6].um_I.iw[16] ;
 wire \top_I.branch[25].block[6].um_I.iw[17] ;
 wire \top_I.branch[25].block[6].um_I.iw[1] ;
 wire \top_I.branch[25].block[6].um_I.iw[2] ;
 wire \top_I.branch[25].block[6].um_I.iw[3] ;
 wire \top_I.branch[25].block[6].um_I.iw[4] ;
 wire \top_I.branch[25].block[6].um_I.iw[5] ;
 wire \top_I.branch[25].block[6].um_I.iw[6] ;
 wire \top_I.branch[25].block[6].um_I.iw[7] ;
 wire \top_I.branch[25].block[6].um_I.iw[8] ;
 wire \top_I.branch[25].block[6].um_I.iw[9] ;
 wire \top_I.branch[25].block[6].um_I.k_zero ;
 wire \top_I.branch[25].block[6].um_I.pg_vdd ;
 wire \top_I.branch[25].block[7].um_I.ana[0] ;
 wire \top_I.branch[25].block[7].um_I.ana[1] ;
 wire \top_I.branch[25].block[7].um_I.ana[2] ;
 wire \top_I.branch[25].block[7].um_I.ana[3] ;
 wire \top_I.branch[25].block[7].um_I.ana[4] ;
 wire \top_I.branch[25].block[7].um_I.ana[5] ;
 wire \top_I.branch[25].block[7].um_I.ana[6] ;
 wire \top_I.branch[25].block[7].um_I.ana[7] ;
 wire \top_I.branch[25].block[7].um_I.clk ;
 wire \top_I.branch[25].block[7].um_I.ena ;
 wire \top_I.branch[25].block[7].um_I.iw[10] ;
 wire \top_I.branch[25].block[7].um_I.iw[11] ;
 wire \top_I.branch[25].block[7].um_I.iw[12] ;
 wire \top_I.branch[25].block[7].um_I.iw[13] ;
 wire \top_I.branch[25].block[7].um_I.iw[14] ;
 wire \top_I.branch[25].block[7].um_I.iw[15] ;
 wire \top_I.branch[25].block[7].um_I.iw[16] ;
 wire \top_I.branch[25].block[7].um_I.iw[17] ;
 wire \top_I.branch[25].block[7].um_I.iw[1] ;
 wire \top_I.branch[25].block[7].um_I.iw[2] ;
 wire \top_I.branch[25].block[7].um_I.iw[3] ;
 wire \top_I.branch[25].block[7].um_I.iw[4] ;
 wire \top_I.branch[25].block[7].um_I.iw[5] ;
 wire \top_I.branch[25].block[7].um_I.iw[6] ;
 wire \top_I.branch[25].block[7].um_I.iw[7] ;
 wire \top_I.branch[25].block[7].um_I.iw[8] ;
 wire \top_I.branch[25].block[7].um_I.iw[9] ;
 wire \top_I.branch[25].block[7].um_I.k_zero ;
 wire \top_I.branch[25].block[7].um_I.pg_vdd ;
 wire \top_I.branch[25].block[8].um_I.ana[0] ;
 wire \top_I.branch[25].block[8].um_I.ana[1] ;
 wire \top_I.branch[25].block[8].um_I.ana[2] ;
 wire \top_I.branch[25].block[8].um_I.ana[3] ;
 wire \top_I.branch[25].block[8].um_I.ana[4] ;
 wire \top_I.branch[25].block[8].um_I.ana[5] ;
 wire \top_I.branch[25].block[8].um_I.ana[6] ;
 wire \top_I.branch[25].block[8].um_I.ana[7] ;
 wire \top_I.branch[25].block[8].um_I.clk ;
 wire \top_I.branch[25].block[8].um_I.ena ;
 wire \top_I.branch[25].block[8].um_I.iw[10] ;
 wire \top_I.branch[25].block[8].um_I.iw[11] ;
 wire \top_I.branch[25].block[8].um_I.iw[12] ;
 wire \top_I.branch[25].block[8].um_I.iw[13] ;
 wire \top_I.branch[25].block[8].um_I.iw[14] ;
 wire \top_I.branch[25].block[8].um_I.iw[15] ;
 wire \top_I.branch[25].block[8].um_I.iw[16] ;
 wire \top_I.branch[25].block[8].um_I.iw[17] ;
 wire \top_I.branch[25].block[8].um_I.iw[1] ;
 wire \top_I.branch[25].block[8].um_I.iw[2] ;
 wire \top_I.branch[25].block[8].um_I.iw[3] ;
 wire \top_I.branch[25].block[8].um_I.iw[4] ;
 wire \top_I.branch[25].block[8].um_I.iw[5] ;
 wire \top_I.branch[25].block[8].um_I.iw[6] ;
 wire \top_I.branch[25].block[8].um_I.iw[7] ;
 wire \top_I.branch[25].block[8].um_I.iw[8] ;
 wire \top_I.branch[25].block[8].um_I.iw[9] ;
 wire \top_I.branch[25].block[8].um_I.k_zero ;
 wire \top_I.branch[25].block[8].um_I.pg_vdd ;
 wire \top_I.branch[25].block[9].um_I.ana[0] ;
 wire \top_I.branch[25].block[9].um_I.ana[1] ;
 wire \top_I.branch[25].block[9].um_I.ana[2] ;
 wire \top_I.branch[25].block[9].um_I.ana[3] ;
 wire \top_I.branch[25].block[9].um_I.ana[4] ;
 wire \top_I.branch[25].block[9].um_I.ana[5] ;
 wire \top_I.branch[25].block[9].um_I.ana[6] ;
 wire \top_I.branch[25].block[9].um_I.ana[7] ;
 wire \top_I.branch[25].block[9].um_I.clk ;
 wire \top_I.branch[25].block[9].um_I.ena ;
 wire \top_I.branch[25].block[9].um_I.iw[10] ;
 wire \top_I.branch[25].block[9].um_I.iw[11] ;
 wire \top_I.branch[25].block[9].um_I.iw[12] ;
 wire \top_I.branch[25].block[9].um_I.iw[13] ;
 wire \top_I.branch[25].block[9].um_I.iw[14] ;
 wire \top_I.branch[25].block[9].um_I.iw[15] ;
 wire \top_I.branch[25].block[9].um_I.iw[16] ;
 wire \top_I.branch[25].block[9].um_I.iw[17] ;
 wire \top_I.branch[25].block[9].um_I.iw[1] ;
 wire \top_I.branch[25].block[9].um_I.iw[2] ;
 wire \top_I.branch[25].block[9].um_I.iw[3] ;
 wire \top_I.branch[25].block[9].um_I.iw[4] ;
 wire \top_I.branch[25].block[9].um_I.iw[5] ;
 wire \top_I.branch[25].block[9].um_I.iw[6] ;
 wire \top_I.branch[25].block[9].um_I.iw[7] ;
 wire \top_I.branch[25].block[9].um_I.iw[8] ;
 wire \top_I.branch[25].block[9].um_I.iw[9] ;
 wire \top_I.branch[25].block[9].um_I.k_zero ;
 wire \top_I.branch[25].block[9].um_I.pg_vdd ;
 wire \top_I.branch[25].l_addr[0] ;
 wire \top_I.branch[25].l_addr[2] ;
 wire \top_I.branch[26].block[0].um_I.ana[0] ;
 wire \top_I.branch[26].block[0].um_I.ana[1] ;
 wire \top_I.branch[26].block[0].um_I.ana[2] ;
 wire \top_I.branch[26].block[0].um_I.ana[3] ;
 wire \top_I.branch[26].block[0].um_I.ana[4] ;
 wire \top_I.branch[26].block[0].um_I.ana[5] ;
 wire \top_I.branch[26].block[0].um_I.ana[6] ;
 wire \top_I.branch[26].block[0].um_I.ana[7] ;
 wire \top_I.branch[26].block[0].um_I.clk ;
 wire \top_I.branch[26].block[0].um_I.ena ;
 wire \top_I.branch[26].block[0].um_I.iw[10] ;
 wire \top_I.branch[26].block[0].um_I.iw[11] ;
 wire \top_I.branch[26].block[0].um_I.iw[12] ;
 wire \top_I.branch[26].block[0].um_I.iw[13] ;
 wire \top_I.branch[26].block[0].um_I.iw[14] ;
 wire \top_I.branch[26].block[0].um_I.iw[15] ;
 wire \top_I.branch[26].block[0].um_I.iw[16] ;
 wire \top_I.branch[26].block[0].um_I.iw[17] ;
 wire \top_I.branch[26].block[0].um_I.iw[1] ;
 wire \top_I.branch[26].block[0].um_I.iw[2] ;
 wire \top_I.branch[26].block[0].um_I.iw[3] ;
 wire \top_I.branch[26].block[0].um_I.iw[4] ;
 wire \top_I.branch[26].block[0].um_I.iw[5] ;
 wire \top_I.branch[26].block[0].um_I.iw[6] ;
 wire \top_I.branch[26].block[0].um_I.iw[7] ;
 wire \top_I.branch[26].block[0].um_I.iw[8] ;
 wire \top_I.branch[26].block[0].um_I.iw[9] ;
 wire \top_I.branch[26].block[0].um_I.k_zero ;
 wire \top_I.branch[26].block[0].um_I.pg_vdd ;
 wire \top_I.branch[26].block[10].um_I.ana[0] ;
 wire \top_I.branch[26].block[10].um_I.ana[1] ;
 wire \top_I.branch[26].block[10].um_I.ana[2] ;
 wire \top_I.branch[26].block[10].um_I.ana[3] ;
 wire \top_I.branch[26].block[10].um_I.ana[4] ;
 wire \top_I.branch[26].block[10].um_I.ana[5] ;
 wire \top_I.branch[26].block[10].um_I.ana[6] ;
 wire \top_I.branch[26].block[10].um_I.ana[7] ;
 wire \top_I.branch[26].block[10].um_I.clk ;
 wire \top_I.branch[26].block[10].um_I.ena ;
 wire \top_I.branch[26].block[10].um_I.iw[10] ;
 wire \top_I.branch[26].block[10].um_I.iw[11] ;
 wire \top_I.branch[26].block[10].um_I.iw[12] ;
 wire \top_I.branch[26].block[10].um_I.iw[13] ;
 wire \top_I.branch[26].block[10].um_I.iw[14] ;
 wire \top_I.branch[26].block[10].um_I.iw[15] ;
 wire \top_I.branch[26].block[10].um_I.iw[16] ;
 wire \top_I.branch[26].block[10].um_I.iw[17] ;
 wire \top_I.branch[26].block[10].um_I.iw[1] ;
 wire \top_I.branch[26].block[10].um_I.iw[2] ;
 wire \top_I.branch[26].block[10].um_I.iw[3] ;
 wire \top_I.branch[26].block[10].um_I.iw[4] ;
 wire \top_I.branch[26].block[10].um_I.iw[5] ;
 wire \top_I.branch[26].block[10].um_I.iw[6] ;
 wire \top_I.branch[26].block[10].um_I.iw[7] ;
 wire \top_I.branch[26].block[10].um_I.iw[8] ;
 wire \top_I.branch[26].block[10].um_I.iw[9] ;
 wire \top_I.branch[26].block[10].um_I.k_zero ;
 wire \top_I.branch[26].block[10].um_I.pg_vdd ;
 wire \top_I.branch[26].block[11].um_I.ana[0] ;
 wire \top_I.branch[26].block[11].um_I.ana[1] ;
 wire \top_I.branch[26].block[11].um_I.ana[2] ;
 wire \top_I.branch[26].block[11].um_I.ana[3] ;
 wire \top_I.branch[26].block[11].um_I.ana[4] ;
 wire \top_I.branch[26].block[11].um_I.ana[5] ;
 wire \top_I.branch[26].block[11].um_I.ana[6] ;
 wire \top_I.branch[26].block[11].um_I.ana[7] ;
 wire \top_I.branch[26].block[11].um_I.clk ;
 wire \top_I.branch[26].block[11].um_I.ena ;
 wire \top_I.branch[26].block[11].um_I.iw[10] ;
 wire \top_I.branch[26].block[11].um_I.iw[11] ;
 wire \top_I.branch[26].block[11].um_I.iw[12] ;
 wire \top_I.branch[26].block[11].um_I.iw[13] ;
 wire \top_I.branch[26].block[11].um_I.iw[14] ;
 wire \top_I.branch[26].block[11].um_I.iw[15] ;
 wire \top_I.branch[26].block[11].um_I.iw[16] ;
 wire \top_I.branch[26].block[11].um_I.iw[17] ;
 wire \top_I.branch[26].block[11].um_I.iw[1] ;
 wire \top_I.branch[26].block[11].um_I.iw[2] ;
 wire \top_I.branch[26].block[11].um_I.iw[3] ;
 wire \top_I.branch[26].block[11].um_I.iw[4] ;
 wire \top_I.branch[26].block[11].um_I.iw[5] ;
 wire \top_I.branch[26].block[11].um_I.iw[6] ;
 wire \top_I.branch[26].block[11].um_I.iw[7] ;
 wire \top_I.branch[26].block[11].um_I.iw[8] ;
 wire \top_I.branch[26].block[11].um_I.iw[9] ;
 wire \top_I.branch[26].block[11].um_I.k_zero ;
 wire \top_I.branch[26].block[11].um_I.pg_vdd ;
 wire \top_I.branch[26].block[12].um_I.ana[0] ;
 wire \top_I.branch[26].block[12].um_I.ana[1] ;
 wire \top_I.branch[26].block[12].um_I.ana[2] ;
 wire \top_I.branch[26].block[12].um_I.ana[3] ;
 wire \top_I.branch[26].block[12].um_I.ana[4] ;
 wire \top_I.branch[26].block[12].um_I.ana[5] ;
 wire \top_I.branch[26].block[12].um_I.ana[6] ;
 wire \top_I.branch[26].block[12].um_I.ana[7] ;
 wire \top_I.branch[26].block[12].um_I.clk ;
 wire \top_I.branch[26].block[12].um_I.ena ;
 wire \top_I.branch[26].block[12].um_I.iw[10] ;
 wire \top_I.branch[26].block[12].um_I.iw[11] ;
 wire \top_I.branch[26].block[12].um_I.iw[12] ;
 wire \top_I.branch[26].block[12].um_I.iw[13] ;
 wire \top_I.branch[26].block[12].um_I.iw[14] ;
 wire \top_I.branch[26].block[12].um_I.iw[15] ;
 wire \top_I.branch[26].block[12].um_I.iw[16] ;
 wire \top_I.branch[26].block[12].um_I.iw[17] ;
 wire \top_I.branch[26].block[12].um_I.iw[1] ;
 wire \top_I.branch[26].block[12].um_I.iw[2] ;
 wire \top_I.branch[26].block[12].um_I.iw[3] ;
 wire \top_I.branch[26].block[12].um_I.iw[4] ;
 wire \top_I.branch[26].block[12].um_I.iw[5] ;
 wire \top_I.branch[26].block[12].um_I.iw[6] ;
 wire \top_I.branch[26].block[12].um_I.iw[7] ;
 wire \top_I.branch[26].block[12].um_I.iw[8] ;
 wire \top_I.branch[26].block[12].um_I.iw[9] ;
 wire \top_I.branch[26].block[12].um_I.k_zero ;
 wire \top_I.branch[26].block[12].um_I.pg_vdd ;
 wire \top_I.branch[26].block[13].um_I.ana[0] ;
 wire \top_I.branch[26].block[13].um_I.ana[1] ;
 wire \top_I.branch[26].block[13].um_I.ana[2] ;
 wire \top_I.branch[26].block[13].um_I.ana[3] ;
 wire \top_I.branch[26].block[13].um_I.ana[4] ;
 wire \top_I.branch[26].block[13].um_I.ana[5] ;
 wire \top_I.branch[26].block[13].um_I.ana[6] ;
 wire \top_I.branch[26].block[13].um_I.ana[7] ;
 wire \top_I.branch[26].block[13].um_I.clk ;
 wire \top_I.branch[26].block[13].um_I.ena ;
 wire \top_I.branch[26].block[13].um_I.iw[10] ;
 wire \top_I.branch[26].block[13].um_I.iw[11] ;
 wire \top_I.branch[26].block[13].um_I.iw[12] ;
 wire \top_I.branch[26].block[13].um_I.iw[13] ;
 wire \top_I.branch[26].block[13].um_I.iw[14] ;
 wire \top_I.branch[26].block[13].um_I.iw[15] ;
 wire \top_I.branch[26].block[13].um_I.iw[16] ;
 wire \top_I.branch[26].block[13].um_I.iw[17] ;
 wire \top_I.branch[26].block[13].um_I.iw[1] ;
 wire \top_I.branch[26].block[13].um_I.iw[2] ;
 wire \top_I.branch[26].block[13].um_I.iw[3] ;
 wire \top_I.branch[26].block[13].um_I.iw[4] ;
 wire \top_I.branch[26].block[13].um_I.iw[5] ;
 wire \top_I.branch[26].block[13].um_I.iw[6] ;
 wire \top_I.branch[26].block[13].um_I.iw[7] ;
 wire \top_I.branch[26].block[13].um_I.iw[8] ;
 wire \top_I.branch[26].block[13].um_I.iw[9] ;
 wire \top_I.branch[26].block[13].um_I.k_zero ;
 wire \top_I.branch[26].block[13].um_I.pg_vdd ;
 wire \top_I.branch[26].block[14].um_I.ana[0] ;
 wire \top_I.branch[26].block[14].um_I.ana[1] ;
 wire \top_I.branch[26].block[14].um_I.ana[2] ;
 wire \top_I.branch[26].block[14].um_I.ana[3] ;
 wire \top_I.branch[26].block[14].um_I.ana[4] ;
 wire \top_I.branch[26].block[14].um_I.ana[5] ;
 wire \top_I.branch[26].block[14].um_I.ana[6] ;
 wire \top_I.branch[26].block[14].um_I.ana[7] ;
 wire \top_I.branch[26].block[14].um_I.clk ;
 wire \top_I.branch[26].block[14].um_I.ena ;
 wire \top_I.branch[26].block[14].um_I.iw[10] ;
 wire \top_I.branch[26].block[14].um_I.iw[11] ;
 wire \top_I.branch[26].block[14].um_I.iw[12] ;
 wire \top_I.branch[26].block[14].um_I.iw[13] ;
 wire \top_I.branch[26].block[14].um_I.iw[14] ;
 wire \top_I.branch[26].block[14].um_I.iw[15] ;
 wire \top_I.branch[26].block[14].um_I.iw[16] ;
 wire \top_I.branch[26].block[14].um_I.iw[17] ;
 wire \top_I.branch[26].block[14].um_I.iw[1] ;
 wire \top_I.branch[26].block[14].um_I.iw[2] ;
 wire \top_I.branch[26].block[14].um_I.iw[3] ;
 wire \top_I.branch[26].block[14].um_I.iw[4] ;
 wire \top_I.branch[26].block[14].um_I.iw[5] ;
 wire \top_I.branch[26].block[14].um_I.iw[6] ;
 wire \top_I.branch[26].block[14].um_I.iw[7] ;
 wire \top_I.branch[26].block[14].um_I.iw[8] ;
 wire \top_I.branch[26].block[14].um_I.iw[9] ;
 wire \top_I.branch[26].block[14].um_I.k_zero ;
 wire \top_I.branch[26].block[14].um_I.pg_vdd ;
 wire \top_I.branch[26].block[15].um_I.ana[0] ;
 wire \top_I.branch[26].block[15].um_I.ana[1] ;
 wire \top_I.branch[26].block[15].um_I.ana[2] ;
 wire \top_I.branch[26].block[15].um_I.ana[3] ;
 wire \top_I.branch[26].block[15].um_I.ana[4] ;
 wire \top_I.branch[26].block[15].um_I.ana[5] ;
 wire \top_I.branch[26].block[15].um_I.ana[6] ;
 wire \top_I.branch[26].block[15].um_I.ana[7] ;
 wire \top_I.branch[26].block[15].um_I.clk ;
 wire \top_I.branch[26].block[15].um_I.ena ;
 wire \top_I.branch[26].block[15].um_I.iw[10] ;
 wire \top_I.branch[26].block[15].um_I.iw[11] ;
 wire \top_I.branch[26].block[15].um_I.iw[12] ;
 wire \top_I.branch[26].block[15].um_I.iw[13] ;
 wire \top_I.branch[26].block[15].um_I.iw[14] ;
 wire \top_I.branch[26].block[15].um_I.iw[15] ;
 wire \top_I.branch[26].block[15].um_I.iw[16] ;
 wire \top_I.branch[26].block[15].um_I.iw[17] ;
 wire \top_I.branch[26].block[15].um_I.iw[1] ;
 wire \top_I.branch[26].block[15].um_I.iw[2] ;
 wire \top_I.branch[26].block[15].um_I.iw[3] ;
 wire \top_I.branch[26].block[15].um_I.iw[4] ;
 wire \top_I.branch[26].block[15].um_I.iw[5] ;
 wire \top_I.branch[26].block[15].um_I.iw[6] ;
 wire \top_I.branch[26].block[15].um_I.iw[7] ;
 wire \top_I.branch[26].block[15].um_I.iw[8] ;
 wire \top_I.branch[26].block[15].um_I.iw[9] ;
 wire \top_I.branch[26].block[15].um_I.k_zero ;
 wire \top_I.branch[26].block[15].um_I.pg_vdd ;
 wire \top_I.branch[26].block[1].um_I.ana[0] ;
 wire \top_I.branch[26].block[1].um_I.ana[1] ;
 wire \top_I.branch[26].block[1].um_I.ana[2] ;
 wire \top_I.branch[26].block[1].um_I.ana[3] ;
 wire \top_I.branch[26].block[1].um_I.ana[4] ;
 wire \top_I.branch[26].block[1].um_I.ana[5] ;
 wire \top_I.branch[26].block[1].um_I.ana[6] ;
 wire \top_I.branch[26].block[1].um_I.ana[7] ;
 wire \top_I.branch[26].block[1].um_I.clk ;
 wire \top_I.branch[26].block[1].um_I.ena ;
 wire \top_I.branch[26].block[1].um_I.iw[10] ;
 wire \top_I.branch[26].block[1].um_I.iw[11] ;
 wire \top_I.branch[26].block[1].um_I.iw[12] ;
 wire \top_I.branch[26].block[1].um_I.iw[13] ;
 wire \top_I.branch[26].block[1].um_I.iw[14] ;
 wire \top_I.branch[26].block[1].um_I.iw[15] ;
 wire \top_I.branch[26].block[1].um_I.iw[16] ;
 wire \top_I.branch[26].block[1].um_I.iw[17] ;
 wire \top_I.branch[26].block[1].um_I.iw[1] ;
 wire \top_I.branch[26].block[1].um_I.iw[2] ;
 wire \top_I.branch[26].block[1].um_I.iw[3] ;
 wire \top_I.branch[26].block[1].um_I.iw[4] ;
 wire \top_I.branch[26].block[1].um_I.iw[5] ;
 wire \top_I.branch[26].block[1].um_I.iw[6] ;
 wire \top_I.branch[26].block[1].um_I.iw[7] ;
 wire \top_I.branch[26].block[1].um_I.iw[8] ;
 wire \top_I.branch[26].block[1].um_I.iw[9] ;
 wire \top_I.branch[26].block[1].um_I.k_zero ;
 wire \top_I.branch[26].block[1].um_I.pg_vdd ;
 wire \top_I.branch[26].block[2].um_I.ana[0] ;
 wire \top_I.branch[26].block[2].um_I.ana[1] ;
 wire \top_I.branch[26].block[2].um_I.ana[2] ;
 wire \top_I.branch[26].block[2].um_I.ana[3] ;
 wire \top_I.branch[26].block[2].um_I.ana[4] ;
 wire \top_I.branch[26].block[2].um_I.ana[5] ;
 wire \top_I.branch[26].block[2].um_I.ana[6] ;
 wire \top_I.branch[26].block[2].um_I.ana[7] ;
 wire \top_I.branch[26].block[2].um_I.clk ;
 wire \top_I.branch[26].block[2].um_I.ena ;
 wire \top_I.branch[26].block[2].um_I.iw[10] ;
 wire \top_I.branch[26].block[2].um_I.iw[11] ;
 wire \top_I.branch[26].block[2].um_I.iw[12] ;
 wire \top_I.branch[26].block[2].um_I.iw[13] ;
 wire \top_I.branch[26].block[2].um_I.iw[14] ;
 wire \top_I.branch[26].block[2].um_I.iw[15] ;
 wire \top_I.branch[26].block[2].um_I.iw[16] ;
 wire \top_I.branch[26].block[2].um_I.iw[17] ;
 wire \top_I.branch[26].block[2].um_I.iw[1] ;
 wire \top_I.branch[26].block[2].um_I.iw[2] ;
 wire \top_I.branch[26].block[2].um_I.iw[3] ;
 wire \top_I.branch[26].block[2].um_I.iw[4] ;
 wire \top_I.branch[26].block[2].um_I.iw[5] ;
 wire \top_I.branch[26].block[2].um_I.iw[6] ;
 wire \top_I.branch[26].block[2].um_I.iw[7] ;
 wire \top_I.branch[26].block[2].um_I.iw[8] ;
 wire \top_I.branch[26].block[2].um_I.iw[9] ;
 wire \top_I.branch[26].block[2].um_I.k_zero ;
 wire \top_I.branch[26].block[2].um_I.pg_vdd ;
 wire \top_I.branch[26].block[3].um_I.ana[0] ;
 wire \top_I.branch[26].block[3].um_I.ana[1] ;
 wire \top_I.branch[26].block[3].um_I.ana[2] ;
 wire \top_I.branch[26].block[3].um_I.ana[3] ;
 wire \top_I.branch[26].block[3].um_I.ana[4] ;
 wire \top_I.branch[26].block[3].um_I.ana[5] ;
 wire \top_I.branch[26].block[3].um_I.ana[6] ;
 wire \top_I.branch[26].block[3].um_I.ana[7] ;
 wire \top_I.branch[26].block[3].um_I.clk ;
 wire \top_I.branch[26].block[3].um_I.ena ;
 wire \top_I.branch[26].block[3].um_I.iw[10] ;
 wire \top_I.branch[26].block[3].um_I.iw[11] ;
 wire \top_I.branch[26].block[3].um_I.iw[12] ;
 wire \top_I.branch[26].block[3].um_I.iw[13] ;
 wire \top_I.branch[26].block[3].um_I.iw[14] ;
 wire \top_I.branch[26].block[3].um_I.iw[15] ;
 wire \top_I.branch[26].block[3].um_I.iw[16] ;
 wire \top_I.branch[26].block[3].um_I.iw[17] ;
 wire \top_I.branch[26].block[3].um_I.iw[1] ;
 wire \top_I.branch[26].block[3].um_I.iw[2] ;
 wire \top_I.branch[26].block[3].um_I.iw[3] ;
 wire \top_I.branch[26].block[3].um_I.iw[4] ;
 wire \top_I.branch[26].block[3].um_I.iw[5] ;
 wire \top_I.branch[26].block[3].um_I.iw[6] ;
 wire \top_I.branch[26].block[3].um_I.iw[7] ;
 wire \top_I.branch[26].block[3].um_I.iw[8] ;
 wire \top_I.branch[26].block[3].um_I.iw[9] ;
 wire \top_I.branch[26].block[3].um_I.k_zero ;
 wire \top_I.branch[26].block[3].um_I.pg_vdd ;
 wire \top_I.branch[26].block[4].um_I.ana[0] ;
 wire \top_I.branch[26].block[4].um_I.ana[1] ;
 wire \top_I.branch[26].block[4].um_I.ana[2] ;
 wire \top_I.branch[26].block[4].um_I.ana[3] ;
 wire \top_I.branch[26].block[4].um_I.ana[4] ;
 wire \top_I.branch[26].block[4].um_I.ana[5] ;
 wire \top_I.branch[26].block[4].um_I.ana[6] ;
 wire \top_I.branch[26].block[4].um_I.ana[7] ;
 wire \top_I.branch[26].block[4].um_I.clk ;
 wire \top_I.branch[26].block[4].um_I.ena ;
 wire \top_I.branch[26].block[4].um_I.iw[10] ;
 wire \top_I.branch[26].block[4].um_I.iw[11] ;
 wire \top_I.branch[26].block[4].um_I.iw[12] ;
 wire \top_I.branch[26].block[4].um_I.iw[13] ;
 wire \top_I.branch[26].block[4].um_I.iw[14] ;
 wire \top_I.branch[26].block[4].um_I.iw[15] ;
 wire \top_I.branch[26].block[4].um_I.iw[16] ;
 wire \top_I.branch[26].block[4].um_I.iw[17] ;
 wire \top_I.branch[26].block[4].um_I.iw[1] ;
 wire \top_I.branch[26].block[4].um_I.iw[2] ;
 wire \top_I.branch[26].block[4].um_I.iw[3] ;
 wire \top_I.branch[26].block[4].um_I.iw[4] ;
 wire \top_I.branch[26].block[4].um_I.iw[5] ;
 wire \top_I.branch[26].block[4].um_I.iw[6] ;
 wire \top_I.branch[26].block[4].um_I.iw[7] ;
 wire \top_I.branch[26].block[4].um_I.iw[8] ;
 wire \top_I.branch[26].block[4].um_I.iw[9] ;
 wire \top_I.branch[26].block[4].um_I.k_zero ;
 wire \top_I.branch[26].block[4].um_I.pg_vdd ;
 wire \top_I.branch[26].block[5].um_I.ana[0] ;
 wire \top_I.branch[26].block[5].um_I.ana[1] ;
 wire \top_I.branch[26].block[5].um_I.ana[2] ;
 wire \top_I.branch[26].block[5].um_I.ana[3] ;
 wire \top_I.branch[26].block[5].um_I.ana[4] ;
 wire \top_I.branch[26].block[5].um_I.ana[5] ;
 wire \top_I.branch[26].block[5].um_I.ana[6] ;
 wire \top_I.branch[26].block[5].um_I.ana[7] ;
 wire \top_I.branch[26].block[5].um_I.clk ;
 wire \top_I.branch[26].block[5].um_I.ena ;
 wire \top_I.branch[26].block[5].um_I.iw[10] ;
 wire \top_I.branch[26].block[5].um_I.iw[11] ;
 wire \top_I.branch[26].block[5].um_I.iw[12] ;
 wire \top_I.branch[26].block[5].um_I.iw[13] ;
 wire \top_I.branch[26].block[5].um_I.iw[14] ;
 wire \top_I.branch[26].block[5].um_I.iw[15] ;
 wire \top_I.branch[26].block[5].um_I.iw[16] ;
 wire \top_I.branch[26].block[5].um_I.iw[17] ;
 wire \top_I.branch[26].block[5].um_I.iw[1] ;
 wire \top_I.branch[26].block[5].um_I.iw[2] ;
 wire \top_I.branch[26].block[5].um_I.iw[3] ;
 wire \top_I.branch[26].block[5].um_I.iw[4] ;
 wire \top_I.branch[26].block[5].um_I.iw[5] ;
 wire \top_I.branch[26].block[5].um_I.iw[6] ;
 wire \top_I.branch[26].block[5].um_I.iw[7] ;
 wire \top_I.branch[26].block[5].um_I.iw[8] ;
 wire \top_I.branch[26].block[5].um_I.iw[9] ;
 wire \top_I.branch[26].block[5].um_I.k_zero ;
 wire \top_I.branch[26].block[5].um_I.pg_vdd ;
 wire \top_I.branch[26].block[6].um_I.ana[0] ;
 wire \top_I.branch[26].block[6].um_I.ana[1] ;
 wire \top_I.branch[26].block[6].um_I.ana[2] ;
 wire \top_I.branch[26].block[6].um_I.ana[3] ;
 wire \top_I.branch[26].block[6].um_I.ana[4] ;
 wire \top_I.branch[26].block[6].um_I.ana[5] ;
 wire \top_I.branch[26].block[6].um_I.ana[6] ;
 wire \top_I.branch[26].block[6].um_I.ana[7] ;
 wire \top_I.branch[26].block[6].um_I.clk ;
 wire \top_I.branch[26].block[6].um_I.ena ;
 wire \top_I.branch[26].block[6].um_I.iw[10] ;
 wire \top_I.branch[26].block[6].um_I.iw[11] ;
 wire \top_I.branch[26].block[6].um_I.iw[12] ;
 wire \top_I.branch[26].block[6].um_I.iw[13] ;
 wire \top_I.branch[26].block[6].um_I.iw[14] ;
 wire \top_I.branch[26].block[6].um_I.iw[15] ;
 wire \top_I.branch[26].block[6].um_I.iw[16] ;
 wire \top_I.branch[26].block[6].um_I.iw[17] ;
 wire \top_I.branch[26].block[6].um_I.iw[1] ;
 wire \top_I.branch[26].block[6].um_I.iw[2] ;
 wire \top_I.branch[26].block[6].um_I.iw[3] ;
 wire \top_I.branch[26].block[6].um_I.iw[4] ;
 wire \top_I.branch[26].block[6].um_I.iw[5] ;
 wire \top_I.branch[26].block[6].um_I.iw[6] ;
 wire \top_I.branch[26].block[6].um_I.iw[7] ;
 wire \top_I.branch[26].block[6].um_I.iw[8] ;
 wire \top_I.branch[26].block[6].um_I.iw[9] ;
 wire \top_I.branch[26].block[6].um_I.k_zero ;
 wire \top_I.branch[26].block[6].um_I.pg_vdd ;
 wire \top_I.branch[26].block[7].um_I.ana[0] ;
 wire \top_I.branch[26].block[7].um_I.ana[1] ;
 wire \top_I.branch[26].block[7].um_I.ana[2] ;
 wire \top_I.branch[26].block[7].um_I.ana[3] ;
 wire \top_I.branch[26].block[7].um_I.ana[4] ;
 wire \top_I.branch[26].block[7].um_I.ana[5] ;
 wire \top_I.branch[26].block[7].um_I.ana[6] ;
 wire \top_I.branch[26].block[7].um_I.ana[7] ;
 wire \top_I.branch[26].block[7].um_I.clk ;
 wire \top_I.branch[26].block[7].um_I.ena ;
 wire \top_I.branch[26].block[7].um_I.iw[10] ;
 wire \top_I.branch[26].block[7].um_I.iw[11] ;
 wire \top_I.branch[26].block[7].um_I.iw[12] ;
 wire \top_I.branch[26].block[7].um_I.iw[13] ;
 wire \top_I.branch[26].block[7].um_I.iw[14] ;
 wire \top_I.branch[26].block[7].um_I.iw[15] ;
 wire \top_I.branch[26].block[7].um_I.iw[16] ;
 wire \top_I.branch[26].block[7].um_I.iw[17] ;
 wire \top_I.branch[26].block[7].um_I.iw[1] ;
 wire \top_I.branch[26].block[7].um_I.iw[2] ;
 wire \top_I.branch[26].block[7].um_I.iw[3] ;
 wire \top_I.branch[26].block[7].um_I.iw[4] ;
 wire \top_I.branch[26].block[7].um_I.iw[5] ;
 wire \top_I.branch[26].block[7].um_I.iw[6] ;
 wire \top_I.branch[26].block[7].um_I.iw[7] ;
 wire \top_I.branch[26].block[7].um_I.iw[8] ;
 wire \top_I.branch[26].block[7].um_I.iw[9] ;
 wire \top_I.branch[26].block[7].um_I.k_zero ;
 wire \top_I.branch[26].block[7].um_I.pg_vdd ;
 wire \top_I.branch[26].block[8].um_I.ana[0] ;
 wire \top_I.branch[26].block[8].um_I.ana[1] ;
 wire \top_I.branch[26].block[8].um_I.ana[2] ;
 wire \top_I.branch[26].block[8].um_I.ana[3] ;
 wire \top_I.branch[26].block[8].um_I.ana[4] ;
 wire \top_I.branch[26].block[8].um_I.ana[5] ;
 wire \top_I.branch[26].block[8].um_I.ana[6] ;
 wire \top_I.branch[26].block[8].um_I.ana[7] ;
 wire \top_I.branch[26].block[8].um_I.clk ;
 wire \top_I.branch[26].block[8].um_I.ena ;
 wire \top_I.branch[26].block[8].um_I.iw[10] ;
 wire \top_I.branch[26].block[8].um_I.iw[11] ;
 wire \top_I.branch[26].block[8].um_I.iw[12] ;
 wire \top_I.branch[26].block[8].um_I.iw[13] ;
 wire \top_I.branch[26].block[8].um_I.iw[14] ;
 wire \top_I.branch[26].block[8].um_I.iw[15] ;
 wire \top_I.branch[26].block[8].um_I.iw[16] ;
 wire \top_I.branch[26].block[8].um_I.iw[17] ;
 wire \top_I.branch[26].block[8].um_I.iw[1] ;
 wire \top_I.branch[26].block[8].um_I.iw[2] ;
 wire \top_I.branch[26].block[8].um_I.iw[3] ;
 wire \top_I.branch[26].block[8].um_I.iw[4] ;
 wire \top_I.branch[26].block[8].um_I.iw[5] ;
 wire \top_I.branch[26].block[8].um_I.iw[6] ;
 wire \top_I.branch[26].block[8].um_I.iw[7] ;
 wire \top_I.branch[26].block[8].um_I.iw[8] ;
 wire \top_I.branch[26].block[8].um_I.iw[9] ;
 wire \top_I.branch[26].block[8].um_I.k_zero ;
 wire \top_I.branch[26].block[8].um_I.pg_vdd ;
 wire \top_I.branch[26].block[9].um_I.ana[0] ;
 wire \top_I.branch[26].block[9].um_I.ana[1] ;
 wire \top_I.branch[26].block[9].um_I.ana[2] ;
 wire \top_I.branch[26].block[9].um_I.ana[3] ;
 wire \top_I.branch[26].block[9].um_I.ana[4] ;
 wire \top_I.branch[26].block[9].um_I.ana[5] ;
 wire \top_I.branch[26].block[9].um_I.ana[6] ;
 wire \top_I.branch[26].block[9].um_I.ana[7] ;
 wire \top_I.branch[26].block[9].um_I.clk ;
 wire \top_I.branch[26].block[9].um_I.ena ;
 wire \top_I.branch[26].block[9].um_I.iw[10] ;
 wire \top_I.branch[26].block[9].um_I.iw[11] ;
 wire \top_I.branch[26].block[9].um_I.iw[12] ;
 wire \top_I.branch[26].block[9].um_I.iw[13] ;
 wire \top_I.branch[26].block[9].um_I.iw[14] ;
 wire \top_I.branch[26].block[9].um_I.iw[15] ;
 wire \top_I.branch[26].block[9].um_I.iw[16] ;
 wire \top_I.branch[26].block[9].um_I.iw[17] ;
 wire \top_I.branch[26].block[9].um_I.iw[1] ;
 wire \top_I.branch[26].block[9].um_I.iw[2] ;
 wire \top_I.branch[26].block[9].um_I.iw[3] ;
 wire \top_I.branch[26].block[9].um_I.iw[4] ;
 wire \top_I.branch[26].block[9].um_I.iw[5] ;
 wire \top_I.branch[26].block[9].um_I.iw[6] ;
 wire \top_I.branch[26].block[9].um_I.iw[7] ;
 wire \top_I.branch[26].block[9].um_I.iw[8] ;
 wire \top_I.branch[26].block[9].um_I.iw[9] ;
 wire \top_I.branch[26].block[9].um_I.k_zero ;
 wire \top_I.branch[26].block[9].um_I.pg_vdd ;
 wire \top_I.branch[26].l_addr[0] ;
 wire \top_I.branch[26].l_addr[1] ;
 wire \top_I.branch[27].block[0].um_I.ana[0] ;
 wire \top_I.branch[27].block[0].um_I.ana[1] ;
 wire \top_I.branch[27].block[0].um_I.ana[2] ;
 wire \top_I.branch[27].block[0].um_I.ana[3] ;
 wire \top_I.branch[27].block[0].um_I.ana[4] ;
 wire \top_I.branch[27].block[0].um_I.ana[5] ;
 wire \top_I.branch[27].block[0].um_I.ana[6] ;
 wire \top_I.branch[27].block[0].um_I.ana[7] ;
 wire \top_I.branch[27].block[0].um_I.clk ;
 wire \top_I.branch[27].block[0].um_I.ena ;
 wire \top_I.branch[27].block[0].um_I.iw[10] ;
 wire \top_I.branch[27].block[0].um_I.iw[11] ;
 wire \top_I.branch[27].block[0].um_I.iw[12] ;
 wire \top_I.branch[27].block[0].um_I.iw[13] ;
 wire \top_I.branch[27].block[0].um_I.iw[14] ;
 wire \top_I.branch[27].block[0].um_I.iw[15] ;
 wire \top_I.branch[27].block[0].um_I.iw[16] ;
 wire \top_I.branch[27].block[0].um_I.iw[17] ;
 wire \top_I.branch[27].block[0].um_I.iw[1] ;
 wire \top_I.branch[27].block[0].um_I.iw[2] ;
 wire \top_I.branch[27].block[0].um_I.iw[3] ;
 wire \top_I.branch[27].block[0].um_I.iw[4] ;
 wire \top_I.branch[27].block[0].um_I.iw[5] ;
 wire \top_I.branch[27].block[0].um_I.iw[6] ;
 wire \top_I.branch[27].block[0].um_I.iw[7] ;
 wire \top_I.branch[27].block[0].um_I.iw[8] ;
 wire \top_I.branch[27].block[0].um_I.iw[9] ;
 wire \top_I.branch[27].block[0].um_I.k_zero ;
 wire \top_I.branch[27].block[0].um_I.pg_vdd ;
 wire \top_I.branch[27].block[10].um_I.ana[0] ;
 wire \top_I.branch[27].block[10].um_I.ana[1] ;
 wire \top_I.branch[27].block[10].um_I.ana[2] ;
 wire \top_I.branch[27].block[10].um_I.ana[3] ;
 wire \top_I.branch[27].block[10].um_I.ana[4] ;
 wire \top_I.branch[27].block[10].um_I.ana[5] ;
 wire \top_I.branch[27].block[10].um_I.ana[6] ;
 wire \top_I.branch[27].block[10].um_I.ana[7] ;
 wire \top_I.branch[27].block[10].um_I.clk ;
 wire \top_I.branch[27].block[10].um_I.ena ;
 wire \top_I.branch[27].block[10].um_I.iw[10] ;
 wire \top_I.branch[27].block[10].um_I.iw[11] ;
 wire \top_I.branch[27].block[10].um_I.iw[12] ;
 wire \top_I.branch[27].block[10].um_I.iw[13] ;
 wire \top_I.branch[27].block[10].um_I.iw[14] ;
 wire \top_I.branch[27].block[10].um_I.iw[15] ;
 wire \top_I.branch[27].block[10].um_I.iw[16] ;
 wire \top_I.branch[27].block[10].um_I.iw[17] ;
 wire \top_I.branch[27].block[10].um_I.iw[1] ;
 wire \top_I.branch[27].block[10].um_I.iw[2] ;
 wire \top_I.branch[27].block[10].um_I.iw[3] ;
 wire \top_I.branch[27].block[10].um_I.iw[4] ;
 wire \top_I.branch[27].block[10].um_I.iw[5] ;
 wire \top_I.branch[27].block[10].um_I.iw[6] ;
 wire \top_I.branch[27].block[10].um_I.iw[7] ;
 wire \top_I.branch[27].block[10].um_I.iw[8] ;
 wire \top_I.branch[27].block[10].um_I.iw[9] ;
 wire \top_I.branch[27].block[10].um_I.k_zero ;
 wire \top_I.branch[27].block[10].um_I.pg_vdd ;
 wire \top_I.branch[27].block[11].um_I.ana[0] ;
 wire \top_I.branch[27].block[11].um_I.ana[1] ;
 wire \top_I.branch[27].block[11].um_I.ana[2] ;
 wire \top_I.branch[27].block[11].um_I.ana[3] ;
 wire \top_I.branch[27].block[11].um_I.ana[4] ;
 wire \top_I.branch[27].block[11].um_I.ana[5] ;
 wire \top_I.branch[27].block[11].um_I.ana[6] ;
 wire \top_I.branch[27].block[11].um_I.ana[7] ;
 wire \top_I.branch[27].block[11].um_I.clk ;
 wire \top_I.branch[27].block[11].um_I.ena ;
 wire \top_I.branch[27].block[11].um_I.iw[10] ;
 wire \top_I.branch[27].block[11].um_I.iw[11] ;
 wire \top_I.branch[27].block[11].um_I.iw[12] ;
 wire \top_I.branch[27].block[11].um_I.iw[13] ;
 wire \top_I.branch[27].block[11].um_I.iw[14] ;
 wire \top_I.branch[27].block[11].um_I.iw[15] ;
 wire \top_I.branch[27].block[11].um_I.iw[16] ;
 wire \top_I.branch[27].block[11].um_I.iw[17] ;
 wire \top_I.branch[27].block[11].um_I.iw[1] ;
 wire \top_I.branch[27].block[11].um_I.iw[2] ;
 wire \top_I.branch[27].block[11].um_I.iw[3] ;
 wire \top_I.branch[27].block[11].um_I.iw[4] ;
 wire \top_I.branch[27].block[11].um_I.iw[5] ;
 wire \top_I.branch[27].block[11].um_I.iw[6] ;
 wire \top_I.branch[27].block[11].um_I.iw[7] ;
 wire \top_I.branch[27].block[11].um_I.iw[8] ;
 wire \top_I.branch[27].block[11].um_I.iw[9] ;
 wire \top_I.branch[27].block[11].um_I.k_zero ;
 wire \top_I.branch[27].block[11].um_I.pg_vdd ;
 wire \top_I.branch[27].block[12].um_I.ana[0] ;
 wire \top_I.branch[27].block[12].um_I.ana[1] ;
 wire \top_I.branch[27].block[12].um_I.ana[2] ;
 wire \top_I.branch[27].block[12].um_I.ana[3] ;
 wire \top_I.branch[27].block[12].um_I.ana[4] ;
 wire \top_I.branch[27].block[12].um_I.ana[5] ;
 wire \top_I.branch[27].block[12].um_I.ana[6] ;
 wire \top_I.branch[27].block[12].um_I.ana[7] ;
 wire \top_I.branch[27].block[12].um_I.clk ;
 wire \top_I.branch[27].block[12].um_I.ena ;
 wire \top_I.branch[27].block[12].um_I.iw[10] ;
 wire \top_I.branch[27].block[12].um_I.iw[11] ;
 wire \top_I.branch[27].block[12].um_I.iw[12] ;
 wire \top_I.branch[27].block[12].um_I.iw[13] ;
 wire \top_I.branch[27].block[12].um_I.iw[14] ;
 wire \top_I.branch[27].block[12].um_I.iw[15] ;
 wire \top_I.branch[27].block[12].um_I.iw[16] ;
 wire \top_I.branch[27].block[12].um_I.iw[17] ;
 wire \top_I.branch[27].block[12].um_I.iw[1] ;
 wire \top_I.branch[27].block[12].um_I.iw[2] ;
 wire \top_I.branch[27].block[12].um_I.iw[3] ;
 wire \top_I.branch[27].block[12].um_I.iw[4] ;
 wire \top_I.branch[27].block[12].um_I.iw[5] ;
 wire \top_I.branch[27].block[12].um_I.iw[6] ;
 wire \top_I.branch[27].block[12].um_I.iw[7] ;
 wire \top_I.branch[27].block[12].um_I.iw[8] ;
 wire \top_I.branch[27].block[12].um_I.iw[9] ;
 wire \top_I.branch[27].block[12].um_I.k_zero ;
 wire \top_I.branch[27].block[12].um_I.pg_vdd ;
 wire \top_I.branch[27].block[13].um_I.ana[0] ;
 wire \top_I.branch[27].block[13].um_I.ana[1] ;
 wire \top_I.branch[27].block[13].um_I.ana[2] ;
 wire \top_I.branch[27].block[13].um_I.ana[3] ;
 wire \top_I.branch[27].block[13].um_I.ana[4] ;
 wire \top_I.branch[27].block[13].um_I.ana[5] ;
 wire \top_I.branch[27].block[13].um_I.ana[6] ;
 wire \top_I.branch[27].block[13].um_I.ana[7] ;
 wire \top_I.branch[27].block[13].um_I.clk ;
 wire \top_I.branch[27].block[13].um_I.ena ;
 wire \top_I.branch[27].block[13].um_I.iw[10] ;
 wire \top_I.branch[27].block[13].um_I.iw[11] ;
 wire \top_I.branch[27].block[13].um_I.iw[12] ;
 wire \top_I.branch[27].block[13].um_I.iw[13] ;
 wire \top_I.branch[27].block[13].um_I.iw[14] ;
 wire \top_I.branch[27].block[13].um_I.iw[15] ;
 wire \top_I.branch[27].block[13].um_I.iw[16] ;
 wire \top_I.branch[27].block[13].um_I.iw[17] ;
 wire \top_I.branch[27].block[13].um_I.iw[1] ;
 wire \top_I.branch[27].block[13].um_I.iw[2] ;
 wire \top_I.branch[27].block[13].um_I.iw[3] ;
 wire \top_I.branch[27].block[13].um_I.iw[4] ;
 wire \top_I.branch[27].block[13].um_I.iw[5] ;
 wire \top_I.branch[27].block[13].um_I.iw[6] ;
 wire \top_I.branch[27].block[13].um_I.iw[7] ;
 wire \top_I.branch[27].block[13].um_I.iw[8] ;
 wire \top_I.branch[27].block[13].um_I.iw[9] ;
 wire \top_I.branch[27].block[13].um_I.k_zero ;
 wire \top_I.branch[27].block[13].um_I.pg_vdd ;
 wire \top_I.branch[27].block[14].um_I.ana[0] ;
 wire \top_I.branch[27].block[14].um_I.ana[1] ;
 wire \top_I.branch[27].block[14].um_I.ana[2] ;
 wire \top_I.branch[27].block[14].um_I.ana[3] ;
 wire \top_I.branch[27].block[14].um_I.ana[4] ;
 wire \top_I.branch[27].block[14].um_I.ana[5] ;
 wire \top_I.branch[27].block[14].um_I.ana[6] ;
 wire \top_I.branch[27].block[14].um_I.ana[7] ;
 wire \top_I.branch[27].block[14].um_I.clk ;
 wire \top_I.branch[27].block[14].um_I.ena ;
 wire \top_I.branch[27].block[14].um_I.iw[10] ;
 wire \top_I.branch[27].block[14].um_I.iw[11] ;
 wire \top_I.branch[27].block[14].um_I.iw[12] ;
 wire \top_I.branch[27].block[14].um_I.iw[13] ;
 wire \top_I.branch[27].block[14].um_I.iw[14] ;
 wire \top_I.branch[27].block[14].um_I.iw[15] ;
 wire \top_I.branch[27].block[14].um_I.iw[16] ;
 wire \top_I.branch[27].block[14].um_I.iw[17] ;
 wire \top_I.branch[27].block[14].um_I.iw[1] ;
 wire \top_I.branch[27].block[14].um_I.iw[2] ;
 wire \top_I.branch[27].block[14].um_I.iw[3] ;
 wire \top_I.branch[27].block[14].um_I.iw[4] ;
 wire \top_I.branch[27].block[14].um_I.iw[5] ;
 wire \top_I.branch[27].block[14].um_I.iw[6] ;
 wire \top_I.branch[27].block[14].um_I.iw[7] ;
 wire \top_I.branch[27].block[14].um_I.iw[8] ;
 wire \top_I.branch[27].block[14].um_I.iw[9] ;
 wire \top_I.branch[27].block[14].um_I.k_zero ;
 wire \top_I.branch[27].block[14].um_I.pg_vdd ;
 wire \top_I.branch[27].block[15].um_I.ana[0] ;
 wire \top_I.branch[27].block[15].um_I.ana[1] ;
 wire \top_I.branch[27].block[15].um_I.ana[2] ;
 wire \top_I.branch[27].block[15].um_I.ana[3] ;
 wire \top_I.branch[27].block[15].um_I.ana[4] ;
 wire \top_I.branch[27].block[15].um_I.ana[5] ;
 wire \top_I.branch[27].block[15].um_I.ana[6] ;
 wire \top_I.branch[27].block[15].um_I.ana[7] ;
 wire \top_I.branch[27].block[15].um_I.clk ;
 wire \top_I.branch[27].block[15].um_I.ena ;
 wire \top_I.branch[27].block[15].um_I.iw[10] ;
 wire \top_I.branch[27].block[15].um_I.iw[11] ;
 wire \top_I.branch[27].block[15].um_I.iw[12] ;
 wire \top_I.branch[27].block[15].um_I.iw[13] ;
 wire \top_I.branch[27].block[15].um_I.iw[14] ;
 wire \top_I.branch[27].block[15].um_I.iw[15] ;
 wire \top_I.branch[27].block[15].um_I.iw[16] ;
 wire \top_I.branch[27].block[15].um_I.iw[17] ;
 wire \top_I.branch[27].block[15].um_I.iw[1] ;
 wire \top_I.branch[27].block[15].um_I.iw[2] ;
 wire \top_I.branch[27].block[15].um_I.iw[3] ;
 wire \top_I.branch[27].block[15].um_I.iw[4] ;
 wire \top_I.branch[27].block[15].um_I.iw[5] ;
 wire \top_I.branch[27].block[15].um_I.iw[6] ;
 wire \top_I.branch[27].block[15].um_I.iw[7] ;
 wire \top_I.branch[27].block[15].um_I.iw[8] ;
 wire \top_I.branch[27].block[15].um_I.iw[9] ;
 wire \top_I.branch[27].block[15].um_I.k_zero ;
 wire \top_I.branch[27].block[15].um_I.pg_vdd ;
 wire \top_I.branch[27].block[1].um_I.ana[0] ;
 wire \top_I.branch[27].block[1].um_I.ana[1] ;
 wire \top_I.branch[27].block[1].um_I.ana[2] ;
 wire \top_I.branch[27].block[1].um_I.ana[3] ;
 wire \top_I.branch[27].block[1].um_I.ana[4] ;
 wire \top_I.branch[27].block[1].um_I.ana[5] ;
 wire \top_I.branch[27].block[1].um_I.ana[6] ;
 wire \top_I.branch[27].block[1].um_I.ana[7] ;
 wire \top_I.branch[27].block[1].um_I.clk ;
 wire \top_I.branch[27].block[1].um_I.ena ;
 wire \top_I.branch[27].block[1].um_I.iw[10] ;
 wire \top_I.branch[27].block[1].um_I.iw[11] ;
 wire \top_I.branch[27].block[1].um_I.iw[12] ;
 wire \top_I.branch[27].block[1].um_I.iw[13] ;
 wire \top_I.branch[27].block[1].um_I.iw[14] ;
 wire \top_I.branch[27].block[1].um_I.iw[15] ;
 wire \top_I.branch[27].block[1].um_I.iw[16] ;
 wire \top_I.branch[27].block[1].um_I.iw[17] ;
 wire \top_I.branch[27].block[1].um_I.iw[1] ;
 wire \top_I.branch[27].block[1].um_I.iw[2] ;
 wire \top_I.branch[27].block[1].um_I.iw[3] ;
 wire \top_I.branch[27].block[1].um_I.iw[4] ;
 wire \top_I.branch[27].block[1].um_I.iw[5] ;
 wire \top_I.branch[27].block[1].um_I.iw[6] ;
 wire \top_I.branch[27].block[1].um_I.iw[7] ;
 wire \top_I.branch[27].block[1].um_I.iw[8] ;
 wire \top_I.branch[27].block[1].um_I.iw[9] ;
 wire \top_I.branch[27].block[1].um_I.k_zero ;
 wire \top_I.branch[27].block[1].um_I.pg_vdd ;
 wire \top_I.branch[27].block[2].um_I.ana[0] ;
 wire \top_I.branch[27].block[2].um_I.ana[1] ;
 wire \top_I.branch[27].block[2].um_I.ana[2] ;
 wire \top_I.branch[27].block[2].um_I.ana[3] ;
 wire \top_I.branch[27].block[2].um_I.ana[4] ;
 wire \top_I.branch[27].block[2].um_I.ana[5] ;
 wire \top_I.branch[27].block[2].um_I.ana[6] ;
 wire \top_I.branch[27].block[2].um_I.ana[7] ;
 wire \top_I.branch[27].block[2].um_I.clk ;
 wire \top_I.branch[27].block[2].um_I.ena ;
 wire \top_I.branch[27].block[2].um_I.iw[10] ;
 wire \top_I.branch[27].block[2].um_I.iw[11] ;
 wire \top_I.branch[27].block[2].um_I.iw[12] ;
 wire \top_I.branch[27].block[2].um_I.iw[13] ;
 wire \top_I.branch[27].block[2].um_I.iw[14] ;
 wire \top_I.branch[27].block[2].um_I.iw[15] ;
 wire \top_I.branch[27].block[2].um_I.iw[16] ;
 wire \top_I.branch[27].block[2].um_I.iw[17] ;
 wire \top_I.branch[27].block[2].um_I.iw[1] ;
 wire \top_I.branch[27].block[2].um_I.iw[2] ;
 wire \top_I.branch[27].block[2].um_I.iw[3] ;
 wire \top_I.branch[27].block[2].um_I.iw[4] ;
 wire \top_I.branch[27].block[2].um_I.iw[5] ;
 wire \top_I.branch[27].block[2].um_I.iw[6] ;
 wire \top_I.branch[27].block[2].um_I.iw[7] ;
 wire \top_I.branch[27].block[2].um_I.iw[8] ;
 wire \top_I.branch[27].block[2].um_I.iw[9] ;
 wire \top_I.branch[27].block[2].um_I.k_zero ;
 wire \top_I.branch[27].block[2].um_I.pg_vdd ;
 wire \top_I.branch[27].block[3].um_I.ana[0] ;
 wire \top_I.branch[27].block[3].um_I.ana[1] ;
 wire \top_I.branch[27].block[3].um_I.ana[2] ;
 wire \top_I.branch[27].block[3].um_I.ana[3] ;
 wire \top_I.branch[27].block[3].um_I.ana[4] ;
 wire \top_I.branch[27].block[3].um_I.ana[5] ;
 wire \top_I.branch[27].block[3].um_I.ana[6] ;
 wire \top_I.branch[27].block[3].um_I.ana[7] ;
 wire \top_I.branch[27].block[3].um_I.clk ;
 wire \top_I.branch[27].block[3].um_I.ena ;
 wire \top_I.branch[27].block[3].um_I.iw[10] ;
 wire \top_I.branch[27].block[3].um_I.iw[11] ;
 wire \top_I.branch[27].block[3].um_I.iw[12] ;
 wire \top_I.branch[27].block[3].um_I.iw[13] ;
 wire \top_I.branch[27].block[3].um_I.iw[14] ;
 wire \top_I.branch[27].block[3].um_I.iw[15] ;
 wire \top_I.branch[27].block[3].um_I.iw[16] ;
 wire \top_I.branch[27].block[3].um_I.iw[17] ;
 wire \top_I.branch[27].block[3].um_I.iw[1] ;
 wire \top_I.branch[27].block[3].um_I.iw[2] ;
 wire \top_I.branch[27].block[3].um_I.iw[3] ;
 wire \top_I.branch[27].block[3].um_I.iw[4] ;
 wire \top_I.branch[27].block[3].um_I.iw[5] ;
 wire \top_I.branch[27].block[3].um_I.iw[6] ;
 wire \top_I.branch[27].block[3].um_I.iw[7] ;
 wire \top_I.branch[27].block[3].um_I.iw[8] ;
 wire \top_I.branch[27].block[3].um_I.iw[9] ;
 wire \top_I.branch[27].block[3].um_I.k_zero ;
 wire \top_I.branch[27].block[3].um_I.pg_vdd ;
 wire \top_I.branch[27].block[4].um_I.ana[0] ;
 wire \top_I.branch[27].block[4].um_I.ana[1] ;
 wire \top_I.branch[27].block[4].um_I.ana[2] ;
 wire \top_I.branch[27].block[4].um_I.ana[3] ;
 wire \top_I.branch[27].block[4].um_I.ana[4] ;
 wire \top_I.branch[27].block[4].um_I.ana[5] ;
 wire \top_I.branch[27].block[4].um_I.ana[6] ;
 wire \top_I.branch[27].block[4].um_I.ana[7] ;
 wire \top_I.branch[27].block[4].um_I.clk ;
 wire \top_I.branch[27].block[4].um_I.ena ;
 wire \top_I.branch[27].block[4].um_I.iw[10] ;
 wire \top_I.branch[27].block[4].um_I.iw[11] ;
 wire \top_I.branch[27].block[4].um_I.iw[12] ;
 wire \top_I.branch[27].block[4].um_I.iw[13] ;
 wire \top_I.branch[27].block[4].um_I.iw[14] ;
 wire \top_I.branch[27].block[4].um_I.iw[15] ;
 wire \top_I.branch[27].block[4].um_I.iw[16] ;
 wire \top_I.branch[27].block[4].um_I.iw[17] ;
 wire \top_I.branch[27].block[4].um_I.iw[1] ;
 wire \top_I.branch[27].block[4].um_I.iw[2] ;
 wire \top_I.branch[27].block[4].um_I.iw[3] ;
 wire \top_I.branch[27].block[4].um_I.iw[4] ;
 wire \top_I.branch[27].block[4].um_I.iw[5] ;
 wire \top_I.branch[27].block[4].um_I.iw[6] ;
 wire \top_I.branch[27].block[4].um_I.iw[7] ;
 wire \top_I.branch[27].block[4].um_I.iw[8] ;
 wire \top_I.branch[27].block[4].um_I.iw[9] ;
 wire \top_I.branch[27].block[4].um_I.k_zero ;
 wire \top_I.branch[27].block[4].um_I.pg_vdd ;
 wire \top_I.branch[27].block[5].um_I.ana[0] ;
 wire \top_I.branch[27].block[5].um_I.ana[1] ;
 wire \top_I.branch[27].block[5].um_I.ana[2] ;
 wire \top_I.branch[27].block[5].um_I.ana[3] ;
 wire \top_I.branch[27].block[5].um_I.ana[4] ;
 wire \top_I.branch[27].block[5].um_I.ana[5] ;
 wire \top_I.branch[27].block[5].um_I.ana[6] ;
 wire \top_I.branch[27].block[5].um_I.ana[7] ;
 wire \top_I.branch[27].block[5].um_I.clk ;
 wire \top_I.branch[27].block[5].um_I.ena ;
 wire \top_I.branch[27].block[5].um_I.iw[10] ;
 wire \top_I.branch[27].block[5].um_I.iw[11] ;
 wire \top_I.branch[27].block[5].um_I.iw[12] ;
 wire \top_I.branch[27].block[5].um_I.iw[13] ;
 wire \top_I.branch[27].block[5].um_I.iw[14] ;
 wire \top_I.branch[27].block[5].um_I.iw[15] ;
 wire \top_I.branch[27].block[5].um_I.iw[16] ;
 wire \top_I.branch[27].block[5].um_I.iw[17] ;
 wire \top_I.branch[27].block[5].um_I.iw[1] ;
 wire \top_I.branch[27].block[5].um_I.iw[2] ;
 wire \top_I.branch[27].block[5].um_I.iw[3] ;
 wire \top_I.branch[27].block[5].um_I.iw[4] ;
 wire \top_I.branch[27].block[5].um_I.iw[5] ;
 wire \top_I.branch[27].block[5].um_I.iw[6] ;
 wire \top_I.branch[27].block[5].um_I.iw[7] ;
 wire \top_I.branch[27].block[5].um_I.iw[8] ;
 wire \top_I.branch[27].block[5].um_I.iw[9] ;
 wire \top_I.branch[27].block[5].um_I.k_zero ;
 wire \top_I.branch[27].block[5].um_I.pg_vdd ;
 wire \top_I.branch[27].block[6].um_I.ana[0] ;
 wire \top_I.branch[27].block[6].um_I.ana[1] ;
 wire \top_I.branch[27].block[6].um_I.ana[2] ;
 wire \top_I.branch[27].block[6].um_I.ana[3] ;
 wire \top_I.branch[27].block[6].um_I.ana[4] ;
 wire \top_I.branch[27].block[6].um_I.ana[5] ;
 wire \top_I.branch[27].block[6].um_I.ana[6] ;
 wire \top_I.branch[27].block[6].um_I.ana[7] ;
 wire \top_I.branch[27].block[6].um_I.clk ;
 wire \top_I.branch[27].block[6].um_I.ena ;
 wire \top_I.branch[27].block[6].um_I.iw[10] ;
 wire \top_I.branch[27].block[6].um_I.iw[11] ;
 wire \top_I.branch[27].block[6].um_I.iw[12] ;
 wire \top_I.branch[27].block[6].um_I.iw[13] ;
 wire \top_I.branch[27].block[6].um_I.iw[14] ;
 wire \top_I.branch[27].block[6].um_I.iw[15] ;
 wire \top_I.branch[27].block[6].um_I.iw[16] ;
 wire \top_I.branch[27].block[6].um_I.iw[17] ;
 wire \top_I.branch[27].block[6].um_I.iw[1] ;
 wire \top_I.branch[27].block[6].um_I.iw[2] ;
 wire \top_I.branch[27].block[6].um_I.iw[3] ;
 wire \top_I.branch[27].block[6].um_I.iw[4] ;
 wire \top_I.branch[27].block[6].um_I.iw[5] ;
 wire \top_I.branch[27].block[6].um_I.iw[6] ;
 wire \top_I.branch[27].block[6].um_I.iw[7] ;
 wire \top_I.branch[27].block[6].um_I.iw[8] ;
 wire \top_I.branch[27].block[6].um_I.iw[9] ;
 wire \top_I.branch[27].block[6].um_I.k_zero ;
 wire \top_I.branch[27].block[6].um_I.pg_vdd ;
 wire \top_I.branch[27].block[7].um_I.ana[0] ;
 wire \top_I.branch[27].block[7].um_I.ana[1] ;
 wire \top_I.branch[27].block[7].um_I.ana[2] ;
 wire \top_I.branch[27].block[7].um_I.ana[3] ;
 wire \top_I.branch[27].block[7].um_I.ana[4] ;
 wire \top_I.branch[27].block[7].um_I.ana[5] ;
 wire \top_I.branch[27].block[7].um_I.ana[6] ;
 wire \top_I.branch[27].block[7].um_I.ana[7] ;
 wire \top_I.branch[27].block[7].um_I.clk ;
 wire \top_I.branch[27].block[7].um_I.ena ;
 wire \top_I.branch[27].block[7].um_I.iw[10] ;
 wire \top_I.branch[27].block[7].um_I.iw[11] ;
 wire \top_I.branch[27].block[7].um_I.iw[12] ;
 wire \top_I.branch[27].block[7].um_I.iw[13] ;
 wire \top_I.branch[27].block[7].um_I.iw[14] ;
 wire \top_I.branch[27].block[7].um_I.iw[15] ;
 wire \top_I.branch[27].block[7].um_I.iw[16] ;
 wire \top_I.branch[27].block[7].um_I.iw[17] ;
 wire \top_I.branch[27].block[7].um_I.iw[1] ;
 wire \top_I.branch[27].block[7].um_I.iw[2] ;
 wire \top_I.branch[27].block[7].um_I.iw[3] ;
 wire \top_I.branch[27].block[7].um_I.iw[4] ;
 wire \top_I.branch[27].block[7].um_I.iw[5] ;
 wire \top_I.branch[27].block[7].um_I.iw[6] ;
 wire \top_I.branch[27].block[7].um_I.iw[7] ;
 wire \top_I.branch[27].block[7].um_I.iw[8] ;
 wire \top_I.branch[27].block[7].um_I.iw[9] ;
 wire \top_I.branch[27].block[7].um_I.k_zero ;
 wire \top_I.branch[27].block[7].um_I.pg_vdd ;
 wire \top_I.branch[27].block[8].um_I.ana[0] ;
 wire \top_I.branch[27].block[8].um_I.ana[1] ;
 wire \top_I.branch[27].block[8].um_I.ana[2] ;
 wire \top_I.branch[27].block[8].um_I.ana[3] ;
 wire \top_I.branch[27].block[8].um_I.ana[4] ;
 wire \top_I.branch[27].block[8].um_I.ana[5] ;
 wire \top_I.branch[27].block[8].um_I.ana[6] ;
 wire \top_I.branch[27].block[8].um_I.ana[7] ;
 wire \top_I.branch[27].block[8].um_I.clk ;
 wire \top_I.branch[27].block[8].um_I.ena ;
 wire \top_I.branch[27].block[8].um_I.iw[10] ;
 wire \top_I.branch[27].block[8].um_I.iw[11] ;
 wire \top_I.branch[27].block[8].um_I.iw[12] ;
 wire \top_I.branch[27].block[8].um_I.iw[13] ;
 wire \top_I.branch[27].block[8].um_I.iw[14] ;
 wire \top_I.branch[27].block[8].um_I.iw[15] ;
 wire \top_I.branch[27].block[8].um_I.iw[16] ;
 wire \top_I.branch[27].block[8].um_I.iw[17] ;
 wire \top_I.branch[27].block[8].um_I.iw[1] ;
 wire \top_I.branch[27].block[8].um_I.iw[2] ;
 wire \top_I.branch[27].block[8].um_I.iw[3] ;
 wire \top_I.branch[27].block[8].um_I.iw[4] ;
 wire \top_I.branch[27].block[8].um_I.iw[5] ;
 wire \top_I.branch[27].block[8].um_I.iw[6] ;
 wire \top_I.branch[27].block[8].um_I.iw[7] ;
 wire \top_I.branch[27].block[8].um_I.iw[8] ;
 wire \top_I.branch[27].block[8].um_I.iw[9] ;
 wire \top_I.branch[27].block[8].um_I.k_zero ;
 wire \top_I.branch[27].block[8].um_I.pg_vdd ;
 wire \top_I.branch[27].block[9].um_I.ana[0] ;
 wire \top_I.branch[27].block[9].um_I.ana[1] ;
 wire \top_I.branch[27].block[9].um_I.ana[2] ;
 wire \top_I.branch[27].block[9].um_I.ana[3] ;
 wire \top_I.branch[27].block[9].um_I.ana[4] ;
 wire \top_I.branch[27].block[9].um_I.ana[5] ;
 wire \top_I.branch[27].block[9].um_I.ana[6] ;
 wire \top_I.branch[27].block[9].um_I.ana[7] ;
 wire \top_I.branch[27].block[9].um_I.clk ;
 wire \top_I.branch[27].block[9].um_I.ena ;
 wire \top_I.branch[27].block[9].um_I.iw[10] ;
 wire \top_I.branch[27].block[9].um_I.iw[11] ;
 wire \top_I.branch[27].block[9].um_I.iw[12] ;
 wire \top_I.branch[27].block[9].um_I.iw[13] ;
 wire \top_I.branch[27].block[9].um_I.iw[14] ;
 wire \top_I.branch[27].block[9].um_I.iw[15] ;
 wire \top_I.branch[27].block[9].um_I.iw[16] ;
 wire \top_I.branch[27].block[9].um_I.iw[17] ;
 wire \top_I.branch[27].block[9].um_I.iw[1] ;
 wire \top_I.branch[27].block[9].um_I.iw[2] ;
 wire \top_I.branch[27].block[9].um_I.iw[3] ;
 wire \top_I.branch[27].block[9].um_I.iw[4] ;
 wire \top_I.branch[27].block[9].um_I.iw[5] ;
 wire \top_I.branch[27].block[9].um_I.iw[6] ;
 wire \top_I.branch[27].block[9].um_I.iw[7] ;
 wire \top_I.branch[27].block[9].um_I.iw[8] ;
 wire \top_I.branch[27].block[9].um_I.iw[9] ;
 wire \top_I.branch[27].block[9].um_I.k_zero ;
 wire \top_I.branch[27].block[9].um_I.pg_vdd ;
 wire \top_I.branch[27].l_addr[0] ;
 wire \top_I.branch[27].l_addr[1] ;
 wire \top_I.branch[28].block[0].um_I.ana[0] ;
 wire \top_I.branch[28].block[0].um_I.ana[1] ;
 wire \top_I.branch[28].block[0].um_I.ana[2] ;
 wire \top_I.branch[28].block[0].um_I.ana[3] ;
 wire \top_I.branch[28].block[0].um_I.ana[4] ;
 wire \top_I.branch[28].block[0].um_I.ana[5] ;
 wire \top_I.branch[28].block[0].um_I.ana[6] ;
 wire \top_I.branch[28].block[0].um_I.ana[7] ;
 wire \top_I.branch[28].block[0].um_I.clk ;
 wire \top_I.branch[28].block[0].um_I.ena ;
 wire \top_I.branch[28].block[0].um_I.iw[10] ;
 wire \top_I.branch[28].block[0].um_I.iw[11] ;
 wire \top_I.branch[28].block[0].um_I.iw[12] ;
 wire \top_I.branch[28].block[0].um_I.iw[13] ;
 wire \top_I.branch[28].block[0].um_I.iw[14] ;
 wire \top_I.branch[28].block[0].um_I.iw[15] ;
 wire \top_I.branch[28].block[0].um_I.iw[16] ;
 wire \top_I.branch[28].block[0].um_I.iw[17] ;
 wire \top_I.branch[28].block[0].um_I.iw[1] ;
 wire \top_I.branch[28].block[0].um_I.iw[2] ;
 wire \top_I.branch[28].block[0].um_I.iw[3] ;
 wire \top_I.branch[28].block[0].um_I.iw[4] ;
 wire \top_I.branch[28].block[0].um_I.iw[5] ;
 wire \top_I.branch[28].block[0].um_I.iw[6] ;
 wire \top_I.branch[28].block[0].um_I.iw[7] ;
 wire \top_I.branch[28].block[0].um_I.iw[8] ;
 wire \top_I.branch[28].block[0].um_I.iw[9] ;
 wire \top_I.branch[28].block[0].um_I.k_zero ;
 wire \top_I.branch[28].block[0].um_I.ow[0] ;
 wire \top_I.branch[28].block[0].um_I.ow[10] ;
 wire \top_I.branch[28].block[0].um_I.ow[11] ;
 wire \top_I.branch[28].block[0].um_I.ow[12] ;
 wire \top_I.branch[28].block[0].um_I.ow[13] ;
 wire \top_I.branch[28].block[0].um_I.ow[14] ;
 wire \top_I.branch[28].block[0].um_I.ow[15] ;
 wire \top_I.branch[28].block[0].um_I.ow[16] ;
 wire \top_I.branch[28].block[0].um_I.ow[17] ;
 wire \top_I.branch[28].block[0].um_I.ow[18] ;
 wire \top_I.branch[28].block[0].um_I.ow[19] ;
 wire \top_I.branch[28].block[0].um_I.ow[1] ;
 wire \top_I.branch[28].block[0].um_I.ow[20] ;
 wire \top_I.branch[28].block[0].um_I.ow[21] ;
 wire \top_I.branch[28].block[0].um_I.ow[22] ;
 wire \top_I.branch[28].block[0].um_I.ow[23] ;
 wire \top_I.branch[28].block[0].um_I.ow[2] ;
 wire \top_I.branch[28].block[0].um_I.ow[3] ;
 wire \top_I.branch[28].block[0].um_I.ow[4] ;
 wire \top_I.branch[28].block[0].um_I.ow[5] ;
 wire \top_I.branch[28].block[0].um_I.ow[6] ;
 wire \top_I.branch[28].block[0].um_I.ow[7] ;
 wire \top_I.branch[28].block[0].um_I.ow[8] ;
 wire \top_I.branch[28].block[0].um_I.ow[9] ;
 wire \top_I.branch[28].block[0].um_I.pg_vdd ;
 wire \top_I.branch[28].block[10].um_I.ana[0] ;
 wire \top_I.branch[28].block[10].um_I.ana[1] ;
 wire \top_I.branch[28].block[10].um_I.ana[2] ;
 wire \top_I.branch[28].block[10].um_I.ana[3] ;
 wire \top_I.branch[28].block[10].um_I.ana[4] ;
 wire \top_I.branch[28].block[10].um_I.ana[5] ;
 wire \top_I.branch[28].block[10].um_I.ana[6] ;
 wire \top_I.branch[28].block[10].um_I.ana[7] ;
 wire \top_I.branch[28].block[10].um_I.clk ;
 wire \top_I.branch[28].block[10].um_I.ena ;
 wire \top_I.branch[28].block[10].um_I.iw[10] ;
 wire \top_I.branch[28].block[10].um_I.iw[11] ;
 wire \top_I.branch[28].block[10].um_I.iw[12] ;
 wire \top_I.branch[28].block[10].um_I.iw[13] ;
 wire \top_I.branch[28].block[10].um_I.iw[14] ;
 wire \top_I.branch[28].block[10].um_I.iw[15] ;
 wire \top_I.branch[28].block[10].um_I.iw[16] ;
 wire \top_I.branch[28].block[10].um_I.iw[17] ;
 wire \top_I.branch[28].block[10].um_I.iw[1] ;
 wire \top_I.branch[28].block[10].um_I.iw[2] ;
 wire \top_I.branch[28].block[10].um_I.iw[3] ;
 wire \top_I.branch[28].block[10].um_I.iw[4] ;
 wire \top_I.branch[28].block[10].um_I.iw[5] ;
 wire \top_I.branch[28].block[10].um_I.iw[6] ;
 wire \top_I.branch[28].block[10].um_I.iw[7] ;
 wire \top_I.branch[28].block[10].um_I.iw[8] ;
 wire \top_I.branch[28].block[10].um_I.iw[9] ;
 wire \top_I.branch[28].block[10].um_I.k_zero ;
 wire \top_I.branch[28].block[10].um_I.ow[0] ;
 wire \top_I.branch[28].block[10].um_I.ow[10] ;
 wire \top_I.branch[28].block[10].um_I.ow[11] ;
 wire \top_I.branch[28].block[10].um_I.ow[12] ;
 wire \top_I.branch[28].block[10].um_I.ow[13] ;
 wire \top_I.branch[28].block[10].um_I.ow[14] ;
 wire \top_I.branch[28].block[10].um_I.ow[15] ;
 wire \top_I.branch[28].block[10].um_I.ow[16] ;
 wire \top_I.branch[28].block[10].um_I.ow[17] ;
 wire \top_I.branch[28].block[10].um_I.ow[18] ;
 wire \top_I.branch[28].block[10].um_I.ow[19] ;
 wire \top_I.branch[28].block[10].um_I.ow[1] ;
 wire \top_I.branch[28].block[10].um_I.ow[20] ;
 wire \top_I.branch[28].block[10].um_I.ow[21] ;
 wire \top_I.branch[28].block[10].um_I.ow[22] ;
 wire \top_I.branch[28].block[10].um_I.ow[23] ;
 wire \top_I.branch[28].block[10].um_I.ow[2] ;
 wire \top_I.branch[28].block[10].um_I.ow[3] ;
 wire \top_I.branch[28].block[10].um_I.ow[4] ;
 wire \top_I.branch[28].block[10].um_I.ow[5] ;
 wire \top_I.branch[28].block[10].um_I.ow[6] ;
 wire \top_I.branch[28].block[10].um_I.ow[7] ;
 wire \top_I.branch[28].block[10].um_I.ow[8] ;
 wire \top_I.branch[28].block[10].um_I.ow[9] ;
 wire \top_I.branch[28].block[10].um_I.pg_vdd ;
 wire \top_I.branch[28].block[11].um_I.ana[0] ;
 wire \top_I.branch[28].block[11].um_I.ana[1] ;
 wire \top_I.branch[28].block[11].um_I.ana[2] ;
 wire \top_I.branch[28].block[11].um_I.ana[3] ;
 wire \top_I.branch[28].block[11].um_I.ana[4] ;
 wire \top_I.branch[28].block[11].um_I.ana[5] ;
 wire \top_I.branch[28].block[11].um_I.ana[6] ;
 wire \top_I.branch[28].block[11].um_I.ana[7] ;
 wire \top_I.branch[28].block[11].um_I.clk ;
 wire \top_I.branch[28].block[11].um_I.ena ;
 wire \top_I.branch[28].block[11].um_I.iw[10] ;
 wire \top_I.branch[28].block[11].um_I.iw[11] ;
 wire \top_I.branch[28].block[11].um_I.iw[12] ;
 wire \top_I.branch[28].block[11].um_I.iw[13] ;
 wire \top_I.branch[28].block[11].um_I.iw[14] ;
 wire \top_I.branch[28].block[11].um_I.iw[15] ;
 wire \top_I.branch[28].block[11].um_I.iw[16] ;
 wire \top_I.branch[28].block[11].um_I.iw[17] ;
 wire \top_I.branch[28].block[11].um_I.iw[1] ;
 wire \top_I.branch[28].block[11].um_I.iw[2] ;
 wire \top_I.branch[28].block[11].um_I.iw[3] ;
 wire \top_I.branch[28].block[11].um_I.iw[4] ;
 wire \top_I.branch[28].block[11].um_I.iw[5] ;
 wire \top_I.branch[28].block[11].um_I.iw[6] ;
 wire \top_I.branch[28].block[11].um_I.iw[7] ;
 wire \top_I.branch[28].block[11].um_I.iw[8] ;
 wire \top_I.branch[28].block[11].um_I.iw[9] ;
 wire \top_I.branch[28].block[11].um_I.k_zero ;
 wire \top_I.branch[28].block[11].um_I.ow[0] ;
 wire \top_I.branch[28].block[11].um_I.ow[10] ;
 wire \top_I.branch[28].block[11].um_I.ow[11] ;
 wire \top_I.branch[28].block[11].um_I.ow[12] ;
 wire \top_I.branch[28].block[11].um_I.ow[13] ;
 wire \top_I.branch[28].block[11].um_I.ow[14] ;
 wire \top_I.branch[28].block[11].um_I.ow[15] ;
 wire \top_I.branch[28].block[11].um_I.ow[16] ;
 wire \top_I.branch[28].block[11].um_I.ow[17] ;
 wire \top_I.branch[28].block[11].um_I.ow[18] ;
 wire \top_I.branch[28].block[11].um_I.ow[19] ;
 wire \top_I.branch[28].block[11].um_I.ow[1] ;
 wire \top_I.branch[28].block[11].um_I.ow[20] ;
 wire \top_I.branch[28].block[11].um_I.ow[21] ;
 wire \top_I.branch[28].block[11].um_I.ow[22] ;
 wire \top_I.branch[28].block[11].um_I.ow[23] ;
 wire \top_I.branch[28].block[11].um_I.ow[2] ;
 wire \top_I.branch[28].block[11].um_I.ow[3] ;
 wire \top_I.branch[28].block[11].um_I.ow[4] ;
 wire \top_I.branch[28].block[11].um_I.ow[5] ;
 wire \top_I.branch[28].block[11].um_I.ow[6] ;
 wire \top_I.branch[28].block[11].um_I.ow[7] ;
 wire \top_I.branch[28].block[11].um_I.ow[8] ;
 wire \top_I.branch[28].block[11].um_I.ow[9] ;
 wire \top_I.branch[28].block[11].um_I.pg_vdd ;
 wire \top_I.branch[28].block[12].um_I.ana[0] ;
 wire \top_I.branch[28].block[12].um_I.ana[1] ;
 wire \top_I.branch[28].block[12].um_I.ana[2] ;
 wire \top_I.branch[28].block[12].um_I.ana[3] ;
 wire \top_I.branch[28].block[12].um_I.ana[4] ;
 wire \top_I.branch[28].block[12].um_I.ana[5] ;
 wire \top_I.branch[28].block[12].um_I.ana[6] ;
 wire \top_I.branch[28].block[12].um_I.ana[7] ;
 wire \top_I.branch[28].block[12].um_I.clk ;
 wire \top_I.branch[28].block[12].um_I.ena ;
 wire \top_I.branch[28].block[12].um_I.iw[10] ;
 wire \top_I.branch[28].block[12].um_I.iw[11] ;
 wire \top_I.branch[28].block[12].um_I.iw[12] ;
 wire \top_I.branch[28].block[12].um_I.iw[13] ;
 wire \top_I.branch[28].block[12].um_I.iw[14] ;
 wire \top_I.branch[28].block[12].um_I.iw[15] ;
 wire \top_I.branch[28].block[12].um_I.iw[16] ;
 wire \top_I.branch[28].block[12].um_I.iw[17] ;
 wire \top_I.branch[28].block[12].um_I.iw[1] ;
 wire \top_I.branch[28].block[12].um_I.iw[2] ;
 wire \top_I.branch[28].block[12].um_I.iw[3] ;
 wire \top_I.branch[28].block[12].um_I.iw[4] ;
 wire \top_I.branch[28].block[12].um_I.iw[5] ;
 wire \top_I.branch[28].block[12].um_I.iw[6] ;
 wire \top_I.branch[28].block[12].um_I.iw[7] ;
 wire \top_I.branch[28].block[12].um_I.iw[8] ;
 wire \top_I.branch[28].block[12].um_I.iw[9] ;
 wire \top_I.branch[28].block[12].um_I.k_zero ;
 wire \top_I.branch[28].block[12].um_I.pg_vdd ;
 wire \top_I.branch[28].block[13].um_I.ana[0] ;
 wire \top_I.branch[28].block[13].um_I.ana[1] ;
 wire \top_I.branch[28].block[13].um_I.ana[2] ;
 wire \top_I.branch[28].block[13].um_I.ana[3] ;
 wire \top_I.branch[28].block[13].um_I.ana[4] ;
 wire \top_I.branch[28].block[13].um_I.ana[5] ;
 wire \top_I.branch[28].block[13].um_I.ana[6] ;
 wire \top_I.branch[28].block[13].um_I.ana[7] ;
 wire \top_I.branch[28].block[13].um_I.clk ;
 wire \top_I.branch[28].block[13].um_I.ena ;
 wire \top_I.branch[28].block[13].um_I.iw[10] ;
 wire \top_I.branch[28].block[13].um_I.iw[11] ;
 wire \top_I.branch[28].block[13].um_I.iw[12] ;
 wire \top_I.branch[28].block[13].um_I.iw[13] ;
 wire \top_I.branch[28].block[13].um_I.iw[14] ;
 wire \top_I.branch[28].block[13].um_I.iw[15] ;
 wire \top_I.branch[28].block[13].um_I.iw[16] ;
 wire \top_I.branch[28].block[13].um_I.iw[17] ;
 wire \top_I.branch[28].block[13].um_I.iw[1] ;
 wire \top_I.branch[28].block[13].um_I.iw[2] ;
 wire \top_I.branch[28].block[13].um_I.iw[3] ;
 wire \top_I.branch[28].block[13].um_I.iw[4] ;
 wire \top_I.branch[28].block[13].um_I.iw[5] ;
 wire \top_I.branch[28].block[13].um_I.iw[6] ;
 wire \top_I.branch[28].block[13].um_I.iw[7] ;
 wire \top_I.branch[28].block[13].um_I.iw[8] ;
 wire \top_I.branch[28].block[13].um_I.iw[9] ;
 wire \top_I.branch[28].block[13].um_I.k_zero ;
 wire \top_I.branch[28].block[13].um_I.ow[0] ;
 wire \top_I.branch[28].block[13].um_I.ow[10] ;
 wire \top_I.branch[28].block[13].um_I.ow[11] ;
 wire \top_I.branch[28].block[13].um_I.ow[12] ;
 wire \top_I.branch[28].block[13].um_I.ow[13] ;
 wire \top_I.branch[28].block[13].um_I.ow[14] ;
 wire \top_I.branch[28].block[13].um_I.ow[15] ;
 wire \top_I.branch[28].block[13].um_I.ow[16] ;
 wire \top_I.branch[28].block[13].um_I.ow[17] ;
 wire \top_I.branch[28].block[13].um_I.ow[18] ;
 wire \top_I.branch[28].block[13].um_I.ow[19] ;
 wire \top_I.branch[28].block[13].um_I.ow[1] ;
 wire \top_I.branch[28].block[13].um_I.ow[20] ;
 wire \top_I.branch[28].block[13].um_I.ow[21] ;
 wire \top_I.branch[28].block[13].um_I.ow[22] ;
 wire \top_I.branch[28].block[13].um_I.ow[23] ;
 wire \top_I.branch[28].block[13].um_I.ow[2] ;
 wire \top_I.branch[28].block[13].um_I.ow[3] ;
 wire \top_I.branch[28].block[13].um_I.ow[4] ;
 wire \top_I.branch[28].block[13].um_I.ow[5] ;
 wire \top_I.branch[28].block[13].um_I.ow[6] ;
 wire \top_I.branch[28].block[13].um_I.ow[7] ;
 wire \top_I.branch[28].block[13].um_I.ow[8] ;
 wire \top_I.branch[28].block[13].um_I.ow[9] ;
 wire \top_I.branch[28].block[13].um_I.pg_vdd ;
 wire \top_I.branch[28].block[14].um_I.ana[0] ;
 wire \top_I.branch[28].block[14].um_I.ana[1] ;
 wire \top_I.branch[28].block[14].um_I.ana[2] ;
 wire \top_I.branch[28].block[14].um_I.ana[3] ;
 wire \top_I.branch[28].block[14].um_I.ana[4] ;
 wire \top_I.branch[28].block[14].um_I.ana[5] ;
 wire \top_I.branch[28].block[14].um_I.ana[6] ;
 wire \top_I.branch[28].block[14].um_I.ana[7] ;
 wire \top_I.branch[28].block[14].um_I.clk ;
 wire \top_I.branch[28].block[14].um_I.ena ;
 wire \top_I.branch[28].block[14].um_I.iw[10] ;
 wire \top_I.branch[28].block[14].um_I.iw[11] ;
 wire \top_I.branch[28].block[14].um_I.iw[12] ;
 wire \top_I.branch[28].block[14].um_I.iw[13] ;
 wire \top_I.branch[28].block[14].um_I.iw[14] ;
 wire \top_I.branch[28].block[14].um_I.iw[15] ;
 wire \top_I.branch[28].block[14].um_I.iw[16] ;
 wire \top_I.branch[28].block[14].um_I.iw[17] ;
 wire \top_I.branch[28].block[14].um_I.iw[1] ;
 wire \top_I.branch[28].block[14].um_I.iw[2] ;
 wire \top_I.branch[28].block[14].um_I.iw[3] ;
 wire \top_I.branch[28].block[14].um_I.iw[4] ;
 wire \top_I.branch[28].block[14].um_I.iw[5] ;
 wire \top_I.branch[28].block[14].um_I.iw[6] ;
 wire \top_I.branch[28].block[14].um_I.iw[7] ;
 wire \top_I.branch[28].block[14].um_I.iw[8] ;
 wire \top_I.branch[28].block[14].um_I.iw[9] ;
 wire \top_I.branch[28].block[14].um_I.k_zero ;
 wire \top_I.branch[28].block[14].um_I.ow[0] ;
 wire \top_I.branch[28].block[14].um_I.ow[10] ;
 wire \top_I.branch[28].block[14].um_I.ow[11] ;
 wire \top_I.branch[28].block[14].um_I.ow[12] ;
 wire \top_I.branch[28].block[14].um_I.ow[13] ;
 wire \top_I.branch[28].block[14].um_I.ow[14] ;
 wire \top_I.branch[28].block[14].um_I.ow[15] ;
 wire \top_I.branch[28].block[14].um_I.ow[16] ;
 wire \top_I.branch[28].block[14].um_I.ow[17] ;
 wire \top_I.branch[28].block[14].um_I.ow[18] ;
 wire \top_I.branch[28].block[14].um_I.ow[19] ;
 wire \top_I.branch[28].block[14].um_I.ow[1] ;
 wire \top_I.branch[28].block[14].um_I.ow[20] ;
 wire \top_I.branch[28].block[14].um_I.ow[21] ;
 wire \top_I.branch[28].block[14].um_I.ow[22] ;
 wire \top_I.branch[28].block[14].um_I.ow[23] ;
 wire \top_I.branch[28].block[14].um_I.ow[2] ;
 wire \top_I.branch[28].block[14].um_I.ow[3] ;
 wire \top_I.branch[28].block[14].um_I.ow[4] ;
 wire \top_I.branch[28].block[14].um_I.ow[5] ;
 wire \top_I.branch[28].block[14].um_I.ow[6] ;
 wire \top_I.branch[28].block[14].um_I.ow[7] ;
 wire \top_I.branch[28].block[14].um_I.ow[8] ;
 wire \top_I.branch[28].block[14].um_I.ow[9] ;
 wire \top_I.branch[28].block[14].um_I.pg_vdd ;
 wire \top_I.branch[28].block[15].um_I.ana[0] ;
 wire \top_I.branch[28].block[15].um_I.ana[1] ;
 wire \top_I.branch[28].block[15].um_I.ana[2] ;
 wire \top_I.branch[28].block[15].um_I.ana[3] ;
 wire \top_I.branch[28].block[15].um_I.ana[4] ;
 wire \top_I.branch[28].block[15].um_I.ana[5] ;
 wire \top_I.branch[28].block[15].um_I.ana[6] ;
 wire \top_I.branch[28].block[15].um_I.ana[7] ;
 wire \top_I.branch[28].block[15].um_I.clk ;
 wire \top_I.branch[28].block[15].um_I.ena ;
 wire \top_I.branch[28].block[15].um_I.iw[10] ;
 wire \top_I.branch[28].block[15].um_I.iw[11] ;
 wire \top_I.branch[28].block[15].um_I.iw[12] ;
 wire \top_I.branch[28].block[15].um_I.iw[13] ;
 wire \top_I.branch[28].block[15].um_I.iw[14] ;
 wire \top_I.branch[28].block[15].um_I.iw[15] ;
 wire \top_I.branch[28].block[15].um_I.iw[16] ;
 wire \top_I.branch[28].block[15].um_I.iw[17] ;
 wire \top_I.branch[28].block[15].um_I.iw[1] ;
 wire \top_I.branch[28].block[15].um_I.iw[2] ;
 wire \top_I.branch[28].block[15].um_I.iw[3] ;
 wire \top_I.branch[28].block[15].um_I.iw[4] ;
 wire \top_I.branch[28].block[15].um_I.iw[5] ;
 wire \top_I.branch[28].block[15].um_I.iw[6] ;
 wire \top_I.branch[28].block[15].um_I.iw[7] ;
 wire \top_I.branch[28].block[15].um_I.iw[8] ;
 wire \top_I.branch[28].block[15].um_I.iw[9] ;
 wire \top_I.branch[28].block[15].um_I.k_zero ;
 wire \top_I.branch[28].block[15].um_I.ow[0] ;
 wire \top_I.branch[28].block[15].um_I.ow[10] ;
 wire \top_I.branch[28].block[15].um_I.ow[11] ;
 wire \top_I.branch[28].block[15].um_I.ow[12] ;
 wire \top_I.branch[28].block[15].um_I.ow[13] ;
 wire \top_I.branch[28].block[15].um_I.ow[14] ;
 wire \top_I.branch[28].block[15].um_I.ow[15] ;
 wire \top_I.branch[28].block[15].um_I.ow[16] ;
 wire \top_I.branch[28].block[15].um_I.ow[17] ;
 wire \top_I.branch[28].block[15].um_I.ow[18] ;
 wire \top_I.branch[28].block[15].um_I.ow[19] ;
 wire \top_I.branch[28].block[15].um_I.ow[1] ;
 wire \top_I.branch[28].block[15].um_I.ow[20] ;
 wire \top_I.branch[28].block[15].um_I.ow[21] ;
 wire \top_I.branch[28].block[15].um_I.ow[22] ;
 wire \top_I.branch[28].block[15].um_I.ow[23] ;
 wire \top_I.branch[28].block[15].um_I.ow[2] ;
 wire \top_I.branch[28].block[15].um_I.ow[3] ;
 wire \top_I.branch[28].block[15].um_I.ow[4] ;
 wire \top_I.branch[28].block[15].um_I.ow[5] ;
 wire \top_I.branch[28].block[15].um_I.ow[6] ;
 wire \top_I.branch[28].block[15].um_I.ow[7] ;
 wire \top_I.branch[28].block[15].um_I.ow[8] ;
 wire \top_I.branch[28].block[15].um_I.ow[9] ;
 wire \top_I.branch[28].block[15].um_I.pg_vdd ;
 wire \top_I.branch[28].block[1].um_I.ana[0] ;
 wire \top_I.branch[28].block[1].um_I.ana[1] ;
 wire \top_I.branch[28].block[1].um_I.ana[2] ;
 wire \top_I.branch[28].block[1].um_I.ana[3] ;
 wire \top_I.branch[28].block[1].um_I.ana[4] ;
 wire \top_I.branch[28].block[1].um_I.ana[5] ;
 wire \top_I.branch[28].block[1].um_I.ana[6] ;
 wire \top_I.branch[28].block[1].um_I.ana[7] ;
 wire \top_I.branch[28].block[1].um_I.clk ;
 wire \top_I.branch[28].block[1].um_I.ena ;
 wire \top_I.branch[28].block[1].um_I.iw[10] ;
 wire \top_I.branch[28].block[1].um_I.iw[11] ;
 wire \top_I.branch[28].block[1].um_I.iw[12] ;
 wire \top_I.branch[28].block[1].um_I.iw[13] ;
 wire \top_I.branch[28].block[1].um_I.iw[14] ;
 wire \top_I.branch[28].block[1].um_I.iw[15] ;
 wire \top_I.branch[28].block[1].um_I.iw[16] ;
 wire \top_I.branch[28].block[1].um_I.iw[17] ;
 wire \top_I.branch[28].block[1].um_I.iw[1] ;
 wire \top_I.branch[28].block[1].um_I.iw[2] ;
 wire \top_I.branch[28].block[1].um_I.iw[3] ;
 wire \top_I.branch[28].block[1].um_I.iw[4] ;
 wire \top_I.branch[28].block[1].um_I.iw[5] ;
 wire \top_I.branch[28].block[1].um_I.iw[6] ;
 wire \top_I.branch[28].block[1].um_I.iw[7] ;
 wire \top_I.branch[28].block[1].um_I.iw[8] ;
 wire \top_I.branch[28].block[1].um_I.iw[9] ;
 wire \top_I.branch[28].block[1].um_I.k_zero ;
 wire \top_I.branch[28].block[1].um_I.ow[0] ;
 wire \top_I.branch[28].block[1].um_I.ow[10] ;
 wire \top_I.branch[28].block[1].um_I.ow[11] ;
 wire \top_I.branch[28].block[1].um_I.ow[12] ;
 wire \top_I.branch[28].block[1].um_I.ow[13] ;
 wire \top_I.branch[28].block[1].um_I.ow[14] ;
 wire \top_I.branch[28].block[1].um_I.ow[15] ;
 wire \top_I.branch[28].block[1].um_I.ow[16] ;
 wire \top_I.branch[28].block[1].um_I.ow[17] ;
 wire \top_I.branch[28].block[1].um_I.ow[18] ;
 wire \top_I.branch[28].block[1].um_I.ow[19] ;
 wire \top_I.branch[28].block[1].um_I.ow[1] ;
 wire \top_I.branch[28].block[1].um_I.ow[20] ;
 wire \top_I.branch[28].block[1].um_I.ow[21] ;
 wire \top_I.branch[28].block[1].um_I.ow[22] ;
 wire \top_I.branch[28].block[1].um_I.ow[23] ;
 wire \top_I.branch[28].block[1].um_I.ow[2] ;
 wire \top_I.branch[28].block[1].um_I.ow[3] ;
 wire \top_I.branch[28].block[1].um_I.ow[4] ;
 wire \top_I.branch[28].block[1].um_I.ow[5] ;
 wire \top_I.branch[28].block[1].um_I.ow[6] ;
 wire \top_I.branch[28].block[1].um_I.ow[7] ;
 wire \top_I.branch[28].block[1].um_I.ow[8] ;
 wire \top_I.branch[28].block[1].um_I.ow[9] ;
 wire \top_I.branch[28].block[1].um_I.pg_vdd ;
 wire \top_I.branch[28].block[2].um_I.ana[0] ;
 wire \top_I.branch[28].block[2].um_I.ana[1] ;
 wire \top_I.branch[28].block[2].um_I.ana[2] ;
 wire \top_I.branch[28].block[2].um_I.ana[3] ;
 wire \top_I.branch[28].block[2].um_I.ana[4] ;
 wire \top_I.branch[28].block[2].um_I.ana[5] ;
 wire \top_I.branch[28].block[2].um_I.ana[6] ;
 wire \top_I.branch[28].block[2].um_I.ana[7] ;
 wire \top_I.branch[28].block[2].um_I.clk ;
 wire \top_I.branch[28].block[2].um_I.ena ;
 wire \top_I.branch[28].block[2].um_I.iw[10] ;
 wire \top_I.branch[28].block[2].um_I.iw[11] ;
 wire \top_I.branch[28].block[2].um_I.iw[12] ;
 wire \top_I.branch[28].block[2].um_I.iw[13] ;
 wire \top_I.branch[28].block[2].um_I.iw[14] ;
 wire \top_I.branch[28].block[2].um_I.iw[15] ;
 wire \top_I.branch[28].block[2].um_I.iw[16] ;
 wire \top_I.branch[28].block[2].um_I.iw[17] ;
 wire \top_I.branch[28].block[2].um_I.iw[1] ;
 wire \top_I.branch[28].block[2].um_I.iw[2] ;
 wire \top_I.branch[28].block[2].um_I.iw[3] ;
 wire \top_I.branch[28].block[2].um_I.iw[4] ;
 wire \top_I.branch[28].block[2].um_I.iw[5] ;
 wire \top_I.branch[28].block[2].um_I.iw[6] ;
 wire \top_I.branch[28].block[2].um_I.iw[7] ;
 wire \top_I.branch[28].block[2].um_I.iw[8] ;
 wire \top_I.branch[28].block[2].um_I.iw[9] ;
 wire \top_I.branch[28].block[2].um_I.k_zero ;
 wire \top_I.branch[28].block[2].um_I.ow[0] ;
 wire \top_I.branch[28].block[2].um_I.ow[10] ;
 wire \top_I.branch[28].block[2].um_I.ow[11] ;
 wire \top_I.branch[28].block[2].um_I.ow[12] ;
 wire \top_I.branch[28].block[2].um_I.ow[13] ;
 wire \top_I.branch[28].block[2].um_I.ow[14] ;
 wire \top_I.branch[28].block[2].um_I.ow[15] ;
 wire \top_I.branch[28].block[2].um_I.ow[16] ;
 wire \top_I.branch[28].block[2].um_I.ow[17] ;
 wire \top_I.branch[28].block[2].um_I.ow[18] ;
 wire \top_I.branch[28].block[2].um_I.ow[19] ;
 wire \top_I.branch[28].block[2].um_I.ow[1] ;
 wire \top_I.branch[28].block[2].um_I.ow[20] ;
 wire \top_I.branch[28].block[2].um_I.ow[21] ;
 wire \top_I.branch[28].block[2].um_I.ow[22] ;
 wire \top_I.branch[28].block[2].um_I.ow[23] ;
 wire \top_I.branch[28].block[2].um_I.ow[2] ;
 wire \top_I.branch[28].block[2].um_I.ow[3] ;
 wire \top_I.branch[28].block[2].um_I.ow[4] ;
 wire \top_I.branch[28].block[2].um_I.ow[5] ;
 wire \top_I.branch[28].block[2].um_I.ow[6] ;
 wire \top_I.branch[28].block[2].um_I.ow[7] ;
 wire \top_I.branch[28].block[2].um_I.ow[8] ;
 wire \top_I.branch[28].block[2].um_I.ow[9] ;
 wire \top_I.branch[28].block[2].um_I.pg_vdd ;
 wire \top_I.branch[28].block[3].um_I.ana[0] ;
 wire \top_I.branch[28].block[3].um_I.ana[1] ;
 wire \top_I.branch[28].block[3].um_I.ana[2] ;
 wire \top_I.branch[28].block[3].um_I.ana[3] ;
 wire \top_I.branch[28].block[3].um_I.ana[4] ;
 wire \top_I.branch[28].block[3].um_I.ana[5] ;
 wire \top_I.branch[28].block[3].um_I.ana[6] ;
 wire \top_I.branch[28].block[3].um_I.ana[7] ;
 wire \top_I.branch[28].block[3].um_I.clk ;
 wire \top_I.branch[28].block[3].um_I.ena ;
 wire \top_I.branch[28].block[3].um_I.iw[10] ;
 wire \top_I.branch[28].block[3].um_I.iw[11] ;
 wire \top_I.branch[28].block[3].um_I.iw[12] ;
 wire \top_I.branch[28].block[3].um_I.iw[13] ;
 wire \top_I.branch[28].block[3].um_I.iw[14] ;
 wire \top_I.branch[28].block[3].um_I.iw[15] ;
 wire \top_I.branch[28].block[3].um_I.iw[16] ;
 wire \top_I.branch[28].block[3].um_I.iw[17] ;
 wire \top_I.branch[28].block[3].um_I.iw[1] ;
 wire \top_I.branch[28].block[3].um_I.iw[2] ;
 wire \top_I.branch[28].block[3].um_I.iw[3] ;
 wire \top_I.branch[28].block[3].um_I.iw[4] ;
 wire \top_I.branch[28].block[3].um_I.iw[5] ;
 wire \top_I.branch[28].block[3].um_I.iw[6] ;
 wire \top_I.branch[28].block[3].um_I.iw[7] ;
 wire \top_I.branch[28].block[3].um_I.iw[8] ;
 wire \top_I.branch[28].block[3].um_I.iw[9] ;
 wire \top_I.branch[28].block[3].um_I.k_zero ;
 wire \top_I.branch[28].block[3].um_I.ow[0] ;
 wire \top_I.branch[28].block[3].um_I.ow[10] ;
 wire \top_I.branch[28].block[3].um_I.ow[11] ;
 wire \top_I.branch[28].block[3].um_I.ow[12] ;
 wire \top_I.branch[28].block[3].um_I.ow[13] ;
 wire \top_I.branch[28].block[3].um_I.ow[14] ;
 wire \top_I.branch[28].block[3].um_I.ow[15] ;
 wire \top_I.branch[28].block[3].um_I.ow[16] ;
 wire \top_I.branch[28].block[3].um_I.ow[17] ;
 wire \top_I.branch[28].block[3].um_I.ow[18] ;
 wire \top_I.branch[28].block[3].um_I.ow[19] ;
 wire \top_I.branch[28].block[3].um_I.ow[1] ;
 wire \top_I.branch[28].block[3].um_I.ow[20] ;
 wire \top_I.branch[28].block[3].um_I.ow[21] ;
 wire \top_I.branch[28].block[3].um_I.ow[22] ;
 wire \top_I.branch[28].block[3].um_I.ow[23] ;
 wire \top_I.branch[28].block[3].um_I.ow[2] ;
 wire \top_I.branch[28].block[3].um_I.ow[3] ;
 wire \top_I.branch[28].block[3].um_I.ow[4] ;
 wire \top_I.branch[28].block[3].um_I.ow[5] ;
 wire \top_I.branch[28].block[3].um_I.ow[6] ;
 wire \top_I.branch[28].block[3].um_I.ow[7] ;
 wire \top_I.branch[28].block[3].um_I.ow[8] ;
 wire \top_I.branch[28].block[3].um_I.ow[9] ;
 wire \top_I.branch[28].block[3].um_I.pg_vdd ;
 wire \top_I.branch[28].block[4].um_I.ana[0] ;
 wire \top_I.branch[28].block[4].um_I.ana[1] ;
 wire \top_I.branch[28].block[4].um_I.ana[2] ;
 wire \top_I.branch[28].block[4].um_I.ana[3] ;
 wire \top_I.branch[28].block[4].um_I.ana[4] ;
 wire \top_I.branch[28].block[4].um_I.ana[5] ;
 wire \top_I.branch[28].block[4].um_I.ana[6] ;
 wire \top_I.branch[28].block[4].um_I.ana[7] ;
 wire \top_I.branch[28].block[4].um_I.clk ;
 wire \top_I.branch[28].block[4].um_I.ena ;
 wire \top_I.branch[28].block[4].um_I.iw[10] ;
 wire \top_I.branch[28].block[4].um_I.iw[11] ;
 wire \top_I.branch[28].block[4].um_I.iw[12] ;
 wire \top_I.branch[28].block[4].um_I.iw[13] ;
 wire \top_I.branch[28].block[4].um_I.iw[14] ;
 wire \top_I.branch[28].block[4].um_I.iw[15] ;
 wire \top_I.branch[28].block[4].um_I.iw[16] ;
 wire \top_I.branch[28].block[4].um_I.iw[17] ;
 wire \top_I.branch[28].block[4].um_I.iw[1] ;
 wire \top_I.branch[28].block[4].um_I.iw[2] ;
 wire \top_I.branch[28].block[4].um_I.iw[3] ;
 wire \top_I.branch[28].block[4].um_I.iw[4] ;
 wire \top_I.branch[28].block[4].um_I.iw[5] ;
 wire \top_I.branch[28].block[4].um_I.iw[6] ;
 wire \top_I.branch[28].block[4].um_I.iw[7] ;
 wire \top_I.branch[28].block[4].um_I.iw[8] ;
 wire \top_I.branch[28].block[4].um_I.iw[9] ;
 wire \top_I.branch[28].block[4].um_I.k_zero ;
 wire \top_I.branch[28].block[4].um_I.ow[0] ;
 wire \top_I.branch[28].block[4].um_I.ow[10] ;
 wire \top_I.branch[28].block[4].um_I.ow[11] ;
 wire \top_I.branch[28].block[4].um_I.ow[12] ;
 wire \top_I.branch[28].block[4].um_I.ow[13] ;
 wire \top_I.branch[28].block[4].um_I.ow[14] ;
 wire \top_I.branch[28].block[4].um_I.ow[15] ;
 wire \top_I.branch[28].block[4].um_I.ow[16] ;
 wire \top_I.branch[28].block[4].um_I.ow[17] ;
 wire \top_I.branch[28].block[4].um_I.ow[18] ;
 wire \top_I.branch[28].block[4].um_I.ow[19] ;
 wire \top_I.branch[28].block[4].um_I.ow[1] ;
 wire \top_I.branch[28].block[4].um_I.ow[20] ;
 wire \top_I.branch[28].block[4].um_I.ow[21] ;
 wire \top_I.branch[28].block[4].um_I.ow[22] ;
 wire \top_I.branch[28].block[4].um_I.ow[23] ;
 wire \top_I.branch[28].block[4].um_I.ow[2] ;
 wire \top_I.branch[28].block[4].um_I.ow[3] ;
 wire \top_I.branch[28].block[4].um_I.ow[4] ;
 wire \top_I.branch[28].block[4].um_I.ow[5] ;
 wire \top_I.branch[28].block[4].um_I.ow[6] ;
 wire \top_I.branch[28].block[4].um_I.ow[7] ;
 wire \top_I.branch[28].block[4].um_I.ow[8] ;
 wire \top_I.branch[28].block[4].um_I.ow[9] ;
 wire \top_I.branch[28].block[4].um_I.pg_vdd ;
 wire \top_I.branch[28].block[5].um_I.ana[0] ;
 wire \top_I.branch[28].block[5].um_I.ana[1] ;
 wire \top_I.branch[28].block[5].um_I.ana[2] ;
 wire \top_I.branch[28].block[5].um_I.ana[3] ;
 wire \top_I.branch[28].block[5].um_I.ana[4] ;
 wire \top_I.branch[28].block[5].um_I.ana[5] ;
 wire \top_I.branch[28].block[5].um_I.ana[6] ;
 wire \top_I.branch[28].block[5].um_I.ana[7] ;
 wire \top_I.branch[28].block[5].um_I.clk ;
 wire \top_I.branch[28].block[5].um_I.ena ;
 wire \top_I.branch[28].block[5].um_I.iw[10] ;
 wire \top_I.branch[28].block[5].um_I.iw[11] ;
 wire \top_I.branch[28].block[5].um_I.iw[12] ;
 wire \top_I.branch[28].block[5].um_I.iw[13] ;
 wire \top_I.branch[28].block[5].um_I.iw[14] ;
 wire \top_I.branch[28].block[5].um_I.iw[15] ;
 wire \top_I.branch[28].block[5].um_I.iw[16] ;
 wire \top_I.branch[28].block[5].um_I.iw[17] ;
 wire \top_I.branch[28].block[5].um_I.iw[1] ;
 wire \top_I.branch[28].block[5].um_I.iw[2] ;
 wire \top_I.branch[28].block[5].um_I.iw[3] ;
 wire \top_I.branch[28].block[5].um_I.iw[4] ;
 wire \top_I.branch[28].block[5].um_I.iw[5] ;
 wire \top_I.branch[28].block[5].um_I.iw[6] ;
 wire \top_I.branch[28].block[5].um_I.iw[7] ;
 wire \top_I.branch[28].block[5].um_I.iw[8] ;
 wire \top_I.branch[28].block[5].um_I.iw[9] ;
 wire \top_I.branch[28].block[5].um_I.k_zero ;
 wire \top_I.branch[28].block[5].um_I.ow[0] ;
 wire \top_I.branch[28].block[5].um_I.ow[10] ;
 wire \top_I.branch[28].block[5].um_I.ow[11] ;
 wire \top_I.branch[28].block[5].um_I.ow[12] ;
 wire \top_I.branch[28].block[5].um_I.ow[13] ;
 wire \top_I.branch[28].block[5].um_I.ow[14] ;
 wire \top_I.branch[28].block[5].um_I.ow[15] ;
 wire \top_I.branch[28].block[5].um_I.ow[16] ;
 wire \top_I.branch[28].block[5].um_I.ow[17] ;
 wire \top_I.branch[28].block[5].um_I.ow[18] ;
 wire \top_I.branch[28].block[5].um_I.ow[19] ;
 wire \top_I.branch[28].block[5].um_I.ow[1] ;
 wire \top_I.branch[28].block[5].um_I.ow[20] ;
 wire \top_I.branch[28].block[5].um_I.ow[21] ;
 wire \top_I.branch[28].block[5].um_I.ow[22] ;
 wire \top_I.branch[28].block[5].um_I.ow[23] ;
 wire \top_I.branch[28].block[5].um_I.ow[2] ;
 wire \top_I.branch[28].block[5].um_I.ow[3] ;
 wire \top_I.branch[28].block[5].um_I.ow[4] ;
 wire \top_I.branch[28].block[5].um_I.ow[5] ;
 wire \top_I.branch[28].block[5].um_I.ow[6] ;
 wire \top_I.branch[28].block[5].um_I.ow[7] ;
 wire \top_I.branch[28].block[5].um_I.ow[8] ;
 wire \top_I.branch[28].block[5].um_I.ow[9] ;
 wire \top_I.branch[28].block[5].um_I.pg_vdd ;
 wire \top_I.branch[28].block[6].um_I.ana[0] ;
 wire \top_I.branch[28].block[6].um_I.ana[1] ;
 wire \top_I.branch[28].block[6].um_I.ana[2] ;
 wire \top_I.branch[28].block[6].um_I.ana[3] ;
 wire \top_I.branch[28].block[6].um_I.ana[4] ;
 wire \top_I.branch[28].block[6].um_I.ana[5] ;
 wire \top_I.branch[28].block[6].um_I.ana[6] ;
 wire \top_I.branch[28].block[6].um_I.ana[7] ;
 wire \top_I.branch[28].block[6].um_I.clk ;
 wire \top_I.branch[28].block[6].um_I.ena ;
 wire \top_I.branch[28].block[6].um_I.iw[10] ;
 wire \top_I.branch[28].block[6].um_I.iw[11] ;
 wire \top_I.branch[28].block[6].um_I.iw[12] ;
 wire \top_I.branch[28].block[6].um_I.iw[13] ;
 wire \top_I.branch[28].block[6].um_I.iw[14] ;
 wire \top_I.branch[28].block[6].um_I.iw[15] ;
 wire \top_I.branch[28].block[6].um_I.iw[16] ;
 wire \top_I.branch[28].block[6].um_I.iw[17] ;
 wire \top_I.branch[28].block[6].um_I.iw[1] ;
 wire \top_I.branch[28].block[6].um_I.iw[2] ;
 wire \top_I.branch[28].block[6].um_I.iw[3] ;
 wire \top_I.branch[28].block[6].um_I.iw[4] ;
 wire \top_I.branch[28].block[6].um_I.iw[5] ;
 wire \top_I.branch[28].block[6].um_I.iw[6] ;
 wire \top_I.branch[28].block[6].um_I.iw[7] ;
 wire \top_I.branch[28].block[6].um_I.iw[8] ;
 wire \top_I.branch[28].block[6].um_I.iw[9] ;
 wire \top_I.branch[28].block[6].um_I.k_zero ;
 wire \top_I.branch[28].block[6].um_I.ow[0] ;
 wire \top_I.branch[28].block[6].um_I.ow[10] ;
 wire \top_I.branch[28].block[6].um_I.ow[11] ;
 wire \top_I.branch[28].block[6].um_I.ow[12] ;
 wire \top_I.branch[28].block[6].um_I.ow[13] ;
 wire \top_I.branch[28].block[6].um_I.ow[14] ;
 wire \top_I.branch[28].block[6].um_I.ow[15] ;
 wire \top_I.branch[28].block[6].um_I.ow[16] ;
 wire \top_I.branch[28].block[6].um_I.ow[17] ;
 wire \top_I.branch[28].block[6].um_I.ow[18] ;
 wire \top_I.branch[28].block[6].um_I.ow[19] ;
 wire \top_I.branch[28].block[6].um_I.ow[1] ;
 wire \top_I.branch[28].block[6].um_I.ow[20] ;
 wire \top_I.branch[28].block[6].um_I.ow[21] ;
 wire \top_I.branch[28].block[6].um_I.ow[22] ;
 wire \top_I.branch[28].block[6].um_I.ow[23] ;
 wire \top_I.branch[28].block[6].um_I.ow[2] ;
 wire \top_I.branch[28].block[6].um_I.ow[3] ;
 wire \top_I.branch[28].block[6].um_I.ow[4] ;
 wire \top_I.branch[28].block[6].um_I.ow[5] ;
 wire \top_I.branch[28].block[6].um_I.ow[6] ;
 wire \top_I.branch[28].block[6].um_I.ow[7] ;
 wire \top_I.branch[28].block[6].um_I.ow[8] ;
 wire \top_I.branch[28].block[6].um_I.ow[9] ;
 wire \top_I.branch[28].block[6].um_I.pg_vdd ;
 wire \top_I.branch[28].block[7].um_I.ana[0] ;
 wire \top_I.branch[28].block[7].um_I.ana[1] ;
 wire \top_I.branch[28].block[7].um_I.ana[2] ;
 wire \top_I.branch[28].block[7].um_I.ana[3] ;
 wire \top_I.branch[28].block[7].um_I.ana[4] ;
 wire \top_I.branch[28].block[7].um_I.ana[5] ;
 wire \top_I.branch[28].block[7].um_I.ana[6] ;
 wire \top_I.branch[28].block[7].um_I.ana[7] ;
 wire \top_I.branch[28].block[7].um_I.clk ;
 wire \top_I.branch[28].block[7].um_I.ena ;
 wire \top_I.branch[28].block[7].um_I.iw[10] ;
 wire \top_I.branch[28].block[7].um_I.iw[11] ;
 wire \top_I.branch[28].block[7].um_I.iw[12] ;
 wire \top_I.branch[28].block[7].um_I.iw[13] ;
 wire \top_I.branch[28].block[7].um_I.iw[14] ;
 wire \top_I.branch[28].block[7].um_I.iw[15] ;
 wire \top_I.branch[28].block[7].um_I.iw[16] ;
 wire \top_I.branch[28].block[7].um_I.iw[17] ;
 wire \top_I.branch[28].block[7].um_I.iw[1] ;
 wire \top_I.branch[28].block[7].um_I.iw[2] ;
 wire \top_I.branch[28].block[7].um_I.iw[3] ;
 wire \top_I.branch[28].block[7].um_I.iw[4] ;
 wire \top_I.branch[28].block[7].um_I.iw[5] ;
 wire \top_I.branch[28].block[7].um_I.iw[6] ;
 wire \top_I.branch[28].block[7].um_I.iw[7] ;
 wire \top_I.branch[28].block[7].um_I.iw[8] ;
 wire \top_I.branch[28].block[7].um_I.iw[9] ;
 wire \top_I.branch[28].block[7].um_I.k_zero ;
 wire \top_I.branch[28].block[7].um_I.ow[0] ;
 wire \top_I.branch[28].block[7].um_I.ow[10] ;
 wire \top_I.branch[28].block[7].um_I.ow[11] ;
 wire \top_I.branch[28].block[7].um_I.ow[12] ;
 wire \top_I.branch[28].block[7].um_I.ow[13] ;
 wire \top_I.branch[28].block[7].um_I.ow[14] ;
 wire \top_I.branch[28].block[7].um_I.ow[15] ;
 wire \top_I.branch[28].block[7].um_I.ow[16] ;
 wire \top_I.branch[28].block[7].um_I.ow[17] ;
 wire \top_I.branch[28].block[7].um_I.ow[18] ;
 wire \top_I.branch[28].block[7].um_I.ow[19] ;
 wire \top_I.branch[28].block[7].um_I.ow[1] ;
 wire \top_I.branch[28].block[7].um_I.ow[20] ;
 wire \top_I.branch[28].block[7].um_I.ow[21] ;
 wire \top_I.branch[28].block[7].um_I.ow[22] ;
 wire \top_I.branch[28].block[7].um_I.ow[23] ;
 wire \top_I.branch[28].block[7].um_I.ow[2] ;
 wire \top_I.branch[28].block[7].um_I.ow[3] ;
 wire \top_I.branch[28].block[7].um_I.ow[4] ;
 wire \top_I.branch[28].block[7].um_I.ow[5] ;
 wire \top_I.branch[28].block[7].um_I.ow[6] ;
 wire \top_I.branch[28].block[7].um_I.ow[7] ;
 wire \top_I.branch[28].block[7].um_I.ow[8] ;
 wire \top_I.branch[28].block[7].um_I.ow[9] ;
 wire \top_I.branch[28].block[7].um_I.pg_vdd ;
 wire \top_I.branch[28].block[8].um_I.ana[0] ;
 wire \top_I.branch[28].block[8].um_I.ana[1] ;
 wire \top_I.branch[28].block[8].um_I.ana[2] ;
 wire \top_I.branch[28].block[8].um_I.ana[3] ;
 wire \top_I.branch[28].block[8].um_I.ana[4] ;
 wire \top_I.branch[28].block[8].um_I.ana[5] ;
 wire \top_I.branch[28].block[8].um_I.ana[6] ;
 wire \top_I.branch[28].block[8].um_I.ana[7] ;
 wire \top_I.branch[28].block[8].um_I.clk ;
 wire \top_I.branch[28].block[8].um_I.ena ;
 wire \top_I.branch[28].block[8].um_I.iw[10] ;
 wire \top_I.branch[28].block[8].um_I.iw[11] ;
 wire \top_I.branch[28].block[8].um_I.iw[12] ;
 wire \top_I.branch[28].block[8].um_I.iw[13] ;
 wire \top_I.branch[28].block[8].um_I.iw[14] ;
 wire \top_I.branch[28].block[8].um_I.iw[15] ;
 wire \top_I.branch[28].block[8].um_I.iw[16] ;
 wire \top_I.branch[28].block[8].um_I.iw[17] ;
 wire \top_I.branch[28].block[8].um_I.iw[1] ;
 wire \top_I.branch[28].block[8].um_I.iw[2] ;
 wire \top_I.branch[28].block[8].um_I.iw[3] ;
 wire \top_I.branch[28].block[8].um_I.iw[4] ;
 wire \top_I.branch[28].block[8].um_I.iw[5] ;
 wire \top_I.branch[28].block[8].um_I.iw[6] ;
 wire \top_I.branch[28].block[8].um_I.iw[7] ;
 wire \top_I.branch[28].block[8].um_I.iw[8] ;
 wire \top_I.branch[28].block[8].um_I.iw[9] ;
 wire \top_I.branch[28].block[8].um_I.k_zero ;
 wire \top_I.branch[28].block[8].um_I.ow[0] ;
 wire \top_I.branch[28].block[8].um_I.ow[10] ;
 wire \top_I.branch[28].block[8].um_I.ow[11] ;
 wire \top_I.branch[28].block[8].um_I.ow[12] ;
 wire \top_I.branch[28].block[8].um_I.ow[13] ;
 wire \top_I.branch[28].block[8].um_I.ow[14] ;
 wire \top_I.branch[28].block[8].um_I.ow[15] ;
 wire \top_I.branch[28].block[8].um_I.ow[16] ;
 wire \top_I.branch[28].block[8].um_I.ow[17] ;
 wire \top_I.branch[28].block[8].um_I.ow[18] ;
 wire \top_I.branch[28].block[8].um_I.ow[19] ;
 wire \top_I.branch[28].block[8].um_I.ow[1] ;
 wire \top_I.branch[28].block[8].um_I.ow[20] ;
 wire \top_I.branch[28].block[8].um_I.ow[21] ;
 wire \top_I.branch[28].block[8].um_I.ow[22] ;
 wire \top_I.branch[28].block[8].um_I.ow[23] ;
 wire \top_I.branch[28].block[8].um_I.ow[2] ;
 wire \top_I.branch[28].block[8].um_I.ow[3] ;
 wire \top_I.branch[28].block[8].um_I.ow[4] ;
 wire \top_I.branch[28].block[8].um_I.ow[5] ;
 wire \top_I.branch[28].block[8].um_I.ow[6] ;
 wire \top_I.branch[28].block[8].um_I.ow[7] ;
 wire \top_I.branch[28].block[8].um_I.ow[8] ;
 wire \top_I.branch[28].block[8].um_I.ow[9] ;
 wire \top_I.branch[28].block[8].um_I.pg_vdd ;
 wire \top_I.branch[28].block[9].um_I.ana[0] ;
 wire \top_I.branch[28].block[9].um_I.ana[1] ;
 wire \top_I.branch[28].block[9].um_I.ana[2] ;
 wire \top_I.branch[28].block[9].um_I.ana[3] ;
 wire \top_I.branch[28].block[9].um_I.ana[4] ;
 wire \top_I.branch[28].block[9].um_I.ana[5] ;
 wire \top_I.branch[28].block[9].um_I.ana[6] ;
 wire \top_I.branch[28].block[9].um_I.ana[7] ;
 wire \top_I.branch[28].block[9].um_I.clk ;
 wire \top_I.branch[28].block[9].um_I.ena ;
 wire \top_I.branch[28].block[9].um_I.iw[10] ;
 wire \top_I.branch[28].block[9].um_I.iw[11] ;
 wire \top_I.branch[28].block[9].um_I.iw[12] ;
 wire \top_I.branch[28].block[9].um_I.iw[13] ;
 wire \top_I.branch[28].block[9].um_I.iw[14] ;
 wire \top_I.branch[28].block[9].um_I.iw[15] ;
 wire \top_I.branch[28].block[9].um_I.iw[16] ;
 wire \top_I.branch[28].block[9].um_I.iw[17] ;
 wire \top_I.branch[28].block[9].um_I.iw[1] ;
 wire \top_I.branch[28].block[9].um_I.iw[2] ;
 wire \top_I.branch[28].block[9].um_I.iw[3] ;
 wire \top_I.branch[28].block[9].um_I.iw[4] ;
 wire \top_I.branch[28].block[9].um_I.iw[5] ;
 wire \top_I.branch[28].block[9].um_I.iw[6] ;
 wire \top_I.branch[28].block[9].um_I.iw[7] ;
 wire \top_I.branch[28].block[9].um_I.iw[8] ;
 wire \top_I.branch[28].block[9].um_I.iw[9] ;
 wire \top_I.branch[28].block[9].um_I.k_zero ;
 wire \top_I.branch[28].block[9].um_I.ow[0] ;
 wire \top_I.branch[28].block[9].um_I.ow[10] ;
 wire \top_I.branch[28].block[9].um_I.ow[11] ;
 wire \top_I.branch[28].block[9].um_I.ow[12] ;
 wire \top_I.branch[28].block[9].um_I.ow[13] ;
 wire \top_I.branch[28].block[9].um_I.ow[14] ;
 wire \top_I.branch[28].block[9].um_I.ow[15] ;
 wire \top_I.branch[28].block[9].um_I.ow[16] ;
 wire \top_I.branch[28].block[9].um_I.ow[17] ;
 wire \top_I.branch[28].block[9].um_I.ow[18] ;
 wire \top_I.branch[28].block[9].um_I.ow[19] ;
 wire \top_I.branch[28].block[9].um_I.ow[1] ;
 wire \top_I.branch[28].block[9].um_I.ow[20] ;
 wire \top_I.branch[28].block[9].um_I.ow[21] ;
 wire \top_I.branch[28].block[9].um_I.ow[22] ;
 wire \top_I.branch[28].block[9].um_I.ow[23] ;
 wire \top_I.branch[28].block[9].um_I.ow[2] ;
 wire \top_I.branch[28].block[9].um_I.ow[3] ;
 wire \top_I.branch[28].block[9].um_I.ow[4] ;
 wire \top_I.branch[28].block[9].um_I.ow[5] ;
 wire \top_I.branch[28].block[9].um_I.ow[6] ;
 wire \top_I.branch[28].block[9].um_I.ow[7] ;
 wire \top_I.branch[28].block[9].um_I.ow[8] ;
 wire \top_I.branch[28].block[9].um_I.ow[9] ;
 wire \top_I.branch[28].block[9].um_I.pg_vdd ;
 wire \top_I.branch[28].l_addr[0] ;
 wire \top_I.branch[28].l_addr[1] ;
 wire \top_I.branch[29].block[0].um_I.ana[0] ;
 wire \top_I.branch[29].block[0].um_I.ana[1] ;
 wire \top_I.branch[29].block[0].um_I.ana[2] ;
 wire \top_I.branch[29].block[0].um_I.ana[3] ;
 wire \top_I.branch[29].block[0].um_I.ana[4] ;
 wire \top_I.branch[29].block[0].um_I.ana[5] ;
 wire \top_I.branch[29].block[0].um_I.ana[6] ;
 wire \top_I.branch[29].block[0].um_I.ana[7] ;
 wire \top_I.branch[29].block[0].um_I.clk ;
 wire \top_I.branch[29].block[0].um_I.ena ;
 wire \top_I.branch[29].block[0].um_I.iw[10] ;
 wire \top_I.branch[29].block[0].um_I.iw[11] ;
 wire \top_I.branch[29].block[0].um_I.iw[12] ;
 wire \top_I.branch[29].block[0].um_I.iw[13] ;
 wire \top_I.branch[29].block[0].um_I.iw[14] ;
 wire \top_I.branch[29].block[0].um_I.iw[15] ;
 wire \top_I.branch[29].block[0].um_I.iw[16] ;
 wire \top_I.branch[29].block[0].um_I.iw[17] ;
 wire \top_I.branch[29].block[0].um_I.iw[1] ;
 wire \top_I.branch[29].block[0].um_I.iw[2] ;
 wire \top_I.branch[29].block[0].um_I.iw[3] ;
 wire \top_I.branch[29].block[0].um_I.iw[4] ;
 wire \top_I.branch[29].block[0].um_I.iw[5] ;
 wire \top_I.branch[29].block[0].um_I.iw[6] ;
 wire \top_I.branch[29].block[0].um_I.iw[7] ;
 wire \top_I.branch[29].block[0].um_I.iw[8] ;
 wire \top_I.branch[29].block[0].um_I.iw[9] ;
 wire \top_I.branch[29].block[0].um_I.k_zero ;
 wire \top_I.branch[29].block[0].um_I.pg_vdd ;
 wire \top_I.branch[29].block[10].um_I.ana[0] ;
 wire \top_I.branch[29].block[10].um_I.ana[1] ;
 wire \top_I.branch[29].block[10].um_I.ana[2] ;
 wire \top_I.branch[29].block[10].um_I.ana[3] ;
 wire \top_I.branch[29].block[10].um_I.ana[4] ;
 wire \top_I.branch[29].block[10].um_I.ana[5] ;
 wire \top_I.branch[29].block[10].um_I.ana[6] ;
 wire \top_I.branch[29].block[10].um_I.ana[7] ;
 wire \top_I.branch[29].block[10].um_I.clk ;
 wire \top_I.branch[29].block[10].um_I.ena ;
 wire \top_I.branch[29].block[10].um_I.iw[10] ;
 wire \top_I.branch[29].block[10].um_I.iw[11] ;
 wire \top_I.branch[29].block[10].um_I.iw[12] ;
 wire \top_I.branch[29].block[10].um_I.iw[13] ;
 wire \top_I.branch[29].block[10].um_I.iw[14] ;
 wire \top_I.branch[29].block[10].um_I.iw[15] ;
 wire \top_I.branch[29].block[10].um_I.iw[16] ;
 wire \top_I.branch[29].block[10].um_I.iw[17] ;
 wire \top_I.branch[29].block[10].um_I.iw[1] ;
 wire \top_I.branch[29].block[10].um_I.iw[2] ;
 wire \top_I.branch[29].block[10].um_I.iw[3] ;
 wire \top_I.branch[29].block[10].um_I.iw[4] ;
 wire \top_I.branch[29].block[10].um_I.iw[5] ;
 wire \top_I.branch[29].block[10].um_I.iw[6] ;
 wire \top_I.branch[29].block[10].um_I.iw[7] ;
 wire \top_I.branch[29].block[10].um_I.iw[8] ;
 wire \top_I.branch[29].block[10].um_I.iw[9] ;
 wire \top_I.branch[29].block[10].um_I.k_zero ;
 wire \top_I.branch[29].block[10].um_I.pg_vdd ;
 wire \top_I.branch[29].block[11].um_I.ana[0] ;
 wire \top_I.branch[29].block[11].um_I.ana[1] ;
 wire \top_I.branch[29].block[11].um_I.ana[2] ;
 wire \top_I.branch[29].block[11].um_I.ana[3] ;
 wire \top_I.branch[29].block[11].um_I.ana[4] ;
 wire \top_I.branch[29].block[11].um_I.ana[5] ;
 wire \top_I.branch[29].block[11].um_I.ana[6] ;
 wire \top_I.branch[29].block[11].um_I.ana[7] ;
 wire \top_I.branch[29].block[11].um_I.clk ;
 wire \top_I.branch[29].block[11].um_I.ena ;
 wire \top_I.branch[29].block[11].um_I.iw[10] ;
 wire \top_I.branch[29].block[11].um_I.iw[11] ;
 wire \top_I.branch[29].block[11].um_I.iw[12] ;
 wire \top_I.branch[29].block[11].um_I.iw[13] ;
 wire \top_I.branch[29].block[11].um_I.iw[14] ;
 wire \top_I.branch[29].block[11].um_I.iw[15] ;
 wire \top_I.branch[29].block[11].um_I.iw[16] ;
 wire \top_I.branch[29].block[11].um_I.iw[17] ;
 wire \top_I.branch[29].block[11].um_I.iw[1] ;
 wire \top_I.branch[29].block[11].um_I.iw[2] ;
 wire \top_I.branch[29].block[11].um_I.iw[3] ;
 wire \top_I.branch[29].block[11].um_I.iw[4] ;
 wire \top_I.branch[29].block[11].um_I.iw[5] ;
 wire \top_I.branch[29].block[11].um_I.iw[6] ;
 wire \top_I.branch[29].block[11].um_I.iw[7] ;
 wire \top_I.branch[29].block[11].um_I.iw[8] ;
 wire \top_I.branch[29].block[11].um_I.iw[9] ;
 wire \top_I.branch[29].block[11].um_I.k_zero ;
 wire \top_I.branch[29].block[11].um_I.pg_vdd ;
 wire \top_I.branch[29].block[12].um_I.ana[0] ;
 wire \top_I.branch[29].block[12].um_I.ana[1] ;
 wire \top_I.branch[29].block[12].um_I.ana[2] ;
 wire \top_I.branch[29].block[12].um_I.ana[3] ;
 wire \top_I.branch[29].block[12].um_I.ana[4] ;
 wire \top_I.branch[29].block[12].um_I.ana[5] ;
 wire \top_I.branch[29].block[12].um_I.ana[6] ;
 wire \top_I.branch[29].block[12].um_I.ana[7] ;
 wire \top_I.branch[29].block[12].um_I.clk ;
 wire \top_I.branch[29].block[12].um_I.ena ;
 wire \top_I.branch[29].block[12].um_I.iw[10] ;
 wire \top_I.branch[29].block[12].um_I.iw[11] ;
 wire \top_I.branch[29].block[12].um_I.iw[12] ;
 wire \top_I.branch[29].block[12].um_I.iw[13] ;
 wire \top_I.branch[29].block[12].um_I.iw[14] ;
 wire \top_I.branch[29].block[12].um_I.iw[15] ;
 wire \top_I.branch[29].block[12].um_I.iw[16] ;
 wire \top_I.branch[29].block[12].um_I.iw[17] ;
 wire \top_I.branch[29].block[12].um_I.iw[1] ;
 wire \top_I.branch[29].block[12].um_I.iw[2] ;
 wire \top_I.branch[29].block[12].um_I.iw[3] ;
 wire \top_I.branch[29].block[12].um_I.iw[4] ;
 wire \top_I.branch[29].block[12].um_I.iw[5] ;
 wire \top_I.branch[29].block[12].um_I.iw[6] ;
 wire \top_I.branch[29].block[12].um_I.iw[7] ;
 wire \top_I.branch[29].block[12].um_I.iw[8] ;
 wire \top_I.branch[29].block[12].um_I.iw[9] ;
 wire \top_I.branch[29].block[12].um_I.k_zero ;
 wire \top_I.branch[29].block[12].um_I.pg_vdd ;
 wire \top_I.branch[29].block[13].um_I.ana[0] ;
 wire \top_I.branch[29].block[13].um_I.ana[1] ;
 wire \top_I.branch[29].block[13].um_I.ana[2] ;
 wire \top_I.branch[29].block[13].um_I.ana[3] ;
 wire \top_I.branch[29].block[13].um_I.ana[4] ;
 wire \top_I.branch[29].block[13].um_I.ana[5] ;
 wire \top_I.branch[29].block[13].um_I.ana[6] ;
 wire \top_I.branch[29].block[13].um_I.ana[7] ;
 wire \top_I.branch[29].block[13].um_I.clk ;
 wire \top_I.branch[29].block[13].um_I.ena ;
 wire \top_I.branch[29].block[13].um_I.iw[10] ;
 wire \top_I.branch[29].block[13].um_I.iw[11] ;
 wire \top_I.branch[29].block[13].um_I.iw[12] ;
 wire \top_I.branch[29].block[13].um_I.iw[13] ;
 wire \top_I.branch[29].block[13].um_I.iw[14] ;
 wire \top_I.branch[29].block[13].um_I.iw[15] ;
 wire \top_I.branch[29].block[13].um_I.iw[16] ;
 wire \top_I.branch[29].block[13].um_I.iw[17] ;
 wire \top_I.branch[29].block[13].um_I.iw[1] ;
 wire \top_I.branch[29].block[13].um_I.iw[2] ;
 wire \top_I.branch[29].block[13].um_I.iw[3] ;
 wire \top_I.branch[29].block[13].um_I.iw[4] ;
 wire \top_I.branch[29].block[13].um_I.iw[5] ;
 wire \top_I.branch[29].block[13].um_I.iw[6] ;
 wire \top_I.branch[29].block[13].um_I.iw[7] ;
 wire \top_I.branch[29].block[13].um_I.iw[8] ;
 wire \top_I.branch[29].block[13].um_I.iw[9] ;
 wire \top_I.branch[29].block[13].um_I.k_zero ;
 wire \top_I.branch[29].block[13].um_I.pg_vdd ;
 wire \top_I.branch[29].block[14].um_I.ana[0] ;
 wire \top_I.branch[29].block[14].um_I.ana[1] ;
 wire \top_I.branch[29].block[14].um_I.ana[2] ;
 wire \top_I.branch[29].block[14].um_I.ana[3] ;
 wire \top_I.branch[29].block[14].um_I.ana[4] ;
 wire \top_I.branch[29].block[14].um_I.ana[5] ;
 wire \top_I.branch[29].block[14].um_I.ana[6] ;
 wire \top_I.branch[29].block[14].um_I.ana[7] ;
 wire \top_I.branch[29].block[14].um_I.clk ;
 wire \top_I.branch[29].block[14].um_I.ena ;
 wire \top_I.branch[29].block[14].um_I.iw[10] ;
 wire \top_I.branch[29].block[14].um_I.iw[11] ;
 wire \top_I.branch[29].block[14].um_I.iw[12] ;
 wire \top_I.branch[29].block[14].um_I.iw[13] ;
 wire \top_I.branch[29].block[14].um_I.iw[14] ;
 wire \top_I.branch[29].block[14].um_I.iw[15] ;
 wire \top_I.branch[29].block[14].um_I.iw[16] ;
 wire \top_I.branch[29].block[14].um_I.iw[17] ;
 wire \top_I.branch[29].block[14].um_I.iw[1] ;
 wire \top_I.branch[29].block[14].um_I.iw[2] ;
 wire \top_I.branch[29].block[14].um_I.iw[3] ;
 wire \top_I.branch[29].block[14].um_I.iw[4] ;
 wire \top_I.branch[29].block[14].um_I.iw[5] ;
 wire \top_I.branch[29].block[14].um_I.iw[6] ;
 wire \top_I.branch[29].block[14].um_I.iw[7] ;
 wire \top_I.branch[29].block[14].um_I.iw[8] ;
 wire \top_I.branch[29].block[14].um_I.iw[9] ;
 wire \top_I.branch[29].block[14].um_I.k_zero ;
 wire \top_I.branch[29].block[14].um_I.pg_vdd ;
 wire \top_I.branch[29].block[15].um_I.ana[0] ;
 wire \top_I.branch[29].block[15].um_I.ana[1] ;
 wire \top_I.branch[29].block[15].um_I.ana[2] ;
 wire \top_I.branch[29].block[15].um_I.ana[3] ;
 wire \top_I.branch[29].block[15].um_I.ana[4] ;
 wire \top_I.branch[29].block[15].um_I.ana[5] ;
 wire \top_I.branch[29].block[15].um_I.ana[6] ;
 wire \top_I.branch[29].block[15].um_I.ana[7] ;
 wire \top_I.branch[29].block[15].um_I.clk ;
 wire \top_I.branch[29].block[15].um_I.ena ;
 wire \top_I.branch[29].block[15].um_I.iw[10] ;
 wire \top_I.branch[29].block[15].um_I.iw[11] ;
 wire \top_I.branch[29].block[15].um_I.iw[12] ;
 wire \top_I.branch[29].block[15].um_I.iw[13] ;
 wire \top_I.branch[29].block[15].um_I.iw[14] ;
 wire \top_I.branch[29].block[15].um_I.iw[15] ;
 wire \top_I.branch[29].block[15].um_I.iw[16] ;
 wire \top_I.branch[29].block[15].um_I.iw[17] ;
 wire \top_I.branch[29].block[15].um_I.iw[1] ;
 wire \top_I.branch[29].block[15].um_I.iw[2] ;
 wire \top_I.branch[29].block[15].um_I.iw[3] ;
 wire \top_I.branch[29].block[15].um_I.iw[4] ;
 wire \top_I.branch[29].block[15].um_I.iw[5] ;
 wire \top_I.branch[29].block[15].um_I.iw[6] ;
 wire \top_I.branch[29].block[15].um_I.iw[7] ;
 wire \top_I.branch[29].block[15].um_I.iw[8] ;
 wire \top_I.branch[29].block[15].um_I.iw[9] ;
 wire \top_I.branch[29].block[15].um_I.k_zero ;
 wire \top_I.branch[29].block[15].um_I.pg_vdd ;
 wire \top_I.branch[29].block[1].um_I.ana[0] ;
 wire \top_I.branch[29].block[1].um_I.ana[1] ;
 wire \top_I.branch[29].block[1].um_I.ana[2] ;
 wire \top_I.branch[29].block[1].um_I.ana[3] ;
 wire \top_I.branch[29].block[1].um_I.ana[4] ;
 wire \top_I.branch[29].block[1].um_I.ana[5] ;
 wire \top_I.branch[29].block[1].um_I.ana[6] ;
 wire \top_I.branch[29].block[1].um_I.ana[7] ;
 wire \top_I.branch[29].block[1].um_I.clk ;
 wire \top_I.branch[29].block[1].um_I.ena ;
 wire \top_I.branch[29].block[1].um_I.iw[10] ;
 wire \top_I.branch[29].block[1].um_I.iw[11] ;
 wire \top_I.branch[29].block[1].um_I.iw[12] ;
 wire \top_I.branch[29].block[1].um_I.iw[13] ;
 wire \top_I.branch[29].block[1].um_I.iw[14] ;
 wire \top_I.branch[29].block[1].um_I.iw[15] ;
 wire \top_I.branch[29].block[1].um_I.iw[16] ;
 wire \top_I.branch[29].block[1].um_I.iw[17] ;
 wire \top_I.branch[29].block[1].um_I.iw[1] ;
 wire \top_I.branch[29].block[1].um_I.iw[2] ;
 wire \top_I.branch[29].block[1].um_I.iw[3] ;
 wire \top_I.branch[29].block[1].um_I.iw[4] ;
 wire \top_I.branch[29].block[1].um_I.iw[5] ;
 wire \top_I.branch[29].block[1].um_I.iw[6] ;
 wire \top_I.branch[29].block[1].um_I.iw[7] ;
 wire \top_I.branch[29].block[1].um_I.iw[8] ;
 wire \top_I.branch[29].block[1].um_I.iw[9] ;
 wire \top_I.branch[29].block[1].um_I.k_zero ;
 wire \top_I.branch[29].block[1].um_I.pg_vdd ;
 wire \top_I.branch[29].block[2].um_I.ana[0] ;
 wire \top_I.branch[29].block[2].um_I.ana[1] ;
 wire \top_I.branch[29].block[2].um_I.ana[2] ;
 wire \top_I.branch[29].block[2].um_I.ana[3] ;
 wire \top_I.branch[29].block[2].um_I.ana[4] ;
 wire \top_I.branch[29].block[2].um_I.ana[5] ;
 wire \top_I.branch[29].block[2].um_I.ana[6] ;
 wire \top_I.branch[29].block[2].um_I.ana[7] ;
 wire \top_I.branch[29].block[2].um_I.clk ;
 wire \top_I.branch[29].block[2].um_I.ena ;
 wire \top_I.branch[29].block[2].um_I.iw[10] ;
 wire \top_I.branch[29].block[2].um_I.iw[11] ;
 wire \top_I.branch[29].block[2].um_I.iw[12] ;
 wire \top_I.branch[29].block[2].um_I.iw[13] ;
 wire \top_I.branch[29].block[2].um_I.iw[14] ;
 wire \top_I.branch[29].block[2].um_I.iw[15] ;
 wire \top_I.branch[29].block[2].um_I.iw[16] ;
 wire \top_I.branch[29].block[2].um_I.iw[17] ;
 wire \top_I.branch[29].block[2].um_I.iw[1] ;
 wire \top_I.branch[29].block[2].um_I.iw[2] ;
 wire \top_I.branch[29].block[2].um_I.iw[3] ;
 wire \top_I.branch[29].block[2].um_I.iw[4] ;
 wire \top_I.branch[29].block[2].um_I.iw[5] ;
 wire \top_I.branch[29].block[2].um_I.iw[6] ;
 wire \top_I.branch[29].block[2].um_I.iw[7] ;
 wire \top_I.branch[29].block[2].um_I.iw[8] ;
 wire \top_I.branch[29].block[2].um_I.iw[9] ;
 wire \top_I.branch[29].block[2].um_I.k_zero ;
 wire \top_I.branch[29].block[2].um_I.pg_vdd ;
 wire \top_I.branch[29].block[3].um_I.ana[0] ;
 wire \top_I.branch[29].block[3].um_I.ana[1] ;
 wire \top_I.branch[29].block[3].um_I.ana[2] ;
 wire \top_I.branch[29].block[3].um_I.ana[3] ;
 wire \top_I.branch[29].block[3].um_I.ana[4] ;
 wire \top_I.branch[29].block[3].um_I.ana[5] ;
 wire \top_I.branch[29].block[3].um_I.ana[6] ;
 wire \top_I.branch[29].block[3].um_I.ana[7] ;
 wire \top_I.branch[29].block[3].um_I.clk ;
 wire \top_I.branch[29].block[3].um_I.ena ;
 wire \top_I.branch[29].block[3].um_I.iw[10] ;
 wire \top_I.branch[29].block[3].um_I.iw[11] ;
 wire \top_I.branch[29].block[3].um_I.iw[12] ;
 wire \top_I.branch[29].block[3].um_I.iw[13] ;
 wire \top_I.branch[29].block[3].um_I.iw[14] ;
 wire \top_I.branch[29].block[3].um_I.iw[15] ;
 wire \top_I.branch[29].block[3].um_I.iw[16] ;
 wire \top_I.branch[29].block[3].um_I.iw[17] ;
 wire \top_I.branch[29].block[3].um_I.iw[1] ;
 wire \top_I.branch[29].block[3].um_I.iw[2] ;
 wire \top_I.branch[29].block[3].um_I.iw[3] ;
 wire \top_I.branch[29].block[3].um_I.iw[4] ;
 wire \top_I.branch[29].block[3].um_I.iw[5] ;
 wire \top_I.branch[29].block[3].um_I.iw[6] ;
 wire \top_I.branch[29].block[3].um_I.iw[7] ;
 wire \top_I.branch[29].block[3].um_I.iw[8] ;
 wire \top_I.branch[29].block[3].um_I.iw[9] ;
 wire \top_I.branch[29].block[3].um_I.k_zero ;
 wire \top_I.branch[29].block[3].um_I.pg_vdd ;
 wire \top_I.branch[29].block[4].um_I.ana[0] ;
 wire \top_I.branch[29].block[4].um_I.ana[1] ;
 wire \top_I.branch[29].block[4].um_I.ana[2] ;
 wire \top_I.branch[29].block[4].um_I.ana[3] ;
 wire \top_I.branch[29].block[4].um_I.ana[4] ;
 wire \top_I.branch[29].block[4].um_I.ana[5] ;
 wire \top_I.branch[29].block[4].um_I.ana[6] ;
 wire \top_I.branch[29].block[4].um_I.ana[7] ;
 wire \top_I.branch[29].block[4].um_I.clk ;
 wire \top_I.branch[29].block[4].um_I.ena ;
 wire \top_I.branch[29].block[4].um_I.iw[10] ;
 wire \top_I.branch[29].block[4].um_I.iw[11] ;
 wire \top_I.branch[29].block[4].um_I.iw[12] ;
 wire \top_I.branch[29].block[4].um_I.iw[13] ;
 wire \top_I.branch[29].block[4].um_I.iw[14] ;
 wire \top_I.branch[29].block[4].um_I.iw[15] ;
 wire \top_I.branch[29].block[4].um_I.iw[16] ;
 wire \top_I.branch[29].block[4].um_I.iw[17] ;
 wire \top_I.branch[29].block[4].um_I.iw[1] ;
 wire \top_I.branch[29].block[4].um_I.iw[2] ;
 wire \top_I.branch[29].block[4].um_I.iw[3] ;
 wire \top_I.branch[29].block[4].um_I.iw[4] ;
 wire \top_I.branch[29].block[4].um_I.iw[5] ;
 wire \top_I.branch[29].block[4].um_I.iw[6] ;
 wire \top_I.branch[29].block[4].um_I.iw[7] ;
 wire \top_I.branch[29].block[4].um_I.iw[8] ;
 wire \top_I.branch[29].block[4].um_I.iw[9] ;
 wire \top_I.branch[29].block[4].um_I.k_zero ;
 wire \top_I.branch[29].block[4].um_I.pg_vdd ;
 wire \top_I.branch[29].block[5].um_I.ana[0] ;
 wire \top_I.branch[29].block[5].um_I.ana[1] ;
 wire \top_I.branch[29].block[5].um_I.ana[2] ;
 wire \top_I.branch[29].block[5].um_I.ana[3] ;
 wire \top_I.branch[29].block[5].um_I.ana[4] ;
 wire \top_I.branch[29].block[5].um_I.ana[5] ;
 wire \top_I.branch[29].block[5].um_I.ana[6] ;
 wire \top_I.branch[29].block[5].um_I.ana[7] ;
 wire \top_I.branch[29].block[5].um_I.clk ;
 wire \top_I.branch[29].block[5].um_I.ena ;
 wire \top_I.branch[29].block[5].um_I.iw[10] ;
 wire \top_I.branch[29].block[5].um_I.iw[11] ;
 wire \top_I.branch[29].block[5].um_I.iw[12] ;
 wire \top_I.branch[29].block[5].um_I.iw[13] ;
 wire \top_I.branch[29].block[5].um_I.iw[14] ;
 wire \top_I.branch[29].block[5].um_I.iw[15] ;
 wire \top_I.branch[29].block[5].um_I.iw[16] ;
 wire \top_I.branch[29].block[5].um_I.iw[17] ;
 wire \top_I.branch[29].block[5].um_I.iw[1] ;
 wire \top_I.branch[29].block[5].um_I.iw[2] ;
 wire \top_I.branch[29].block[5].um_I.iw[3] ;
 wire \top_I.branch[29].block[5].um_I.iw[4] ;
 wire \top_I.branch[29].block[5].um_I.iw[5] ;
 wire \top_I.branch[29].block[5].um_I.iw[6] ;
 wire \top_I.branch[29].block[5].um_I.iw[7] ;
 wire \top_I.branch[29].block[5].um_I.iw[8] ;
 wire \top_I.branch[29].block[5].um_I.iw[9] ;
 wire \top_I.branch[29].block[5].um_I.k_zero ;
 wire \top_I.branch[29].block[5].um_I.pg_vdd ;
 wire \top_I.branch[29].block[6].um_I.ana[0] ;
 wire \top_I.branch[29].block[6].um_I.ana[1] ;
 wire \top_I.branch[29].block[6].um_I.ana[2] ;
 wire \top_I.branch[29].block[6].um_I.ana[3] ;
 wire \top_I.branch[29].block[6].um_I.ana[4] ;
 wire \top_I.branch[29].block[6].um_I.ana[5] ;
 wire \top_I.branch[29].block[6].um_I.ana[6] ;
 wire \top_I.branch[29].block[6].um_I.ana[7] ;
 wire \top_I.branch[29].block[6].um_I.clk ;
 wire \top_I.branch[29].block[6].um_I.ena ;
 wire \top_I.branch[29].block[6].um_I.iw[10] ;
 wire \top_I.branch[29].block[6].um_I.iw[11] ;
 wire \top_I.branch[29].block[6].um_I.iw[12] ;
 wire \top_I.branch[29].block[6].um_I.iw[13] ;
 wire \top_I.branch[29].block[6].um_I.iw[14] ;
 wire \top_I.branch[29].block[6].um_I.iw[15] ;
 wire \top_I.branch[29].block[6].um_I.iw[16] ;
 wire \top_I.branch[29].block[6].um_I.iw[17] ;
 wire \top_I.branch[29].block[6].um_I.iw[1] ;
 wire \top_I.branch[29].block[6].um_I.iw[2] ;
 wire \top_I.branch[29].block[6].um_I.iw[3] ;
 wire \top_I.branch[29].block[6].um_I.iw[4] ;
 wire \top_I.branch[29].block[6].um_I.iw[5] ;
 wire \top_I.branch[29].block[6].um_I.iw[6] ;
 wire \top_I.branch[29].block[6].um_I.iw[7] ;
 wire \top_I.branch[29].block[6].um_I.iw[8] ;
 wire \top_I.branch[29].block[6].um_I.iw[9] ;
 wire \top_I.branch[29].block[6].um_I.k_zero ;
 wire \top_I.branch[29].block[6].um_I.pg_vdd ;
 wire \top_I.branch[29].block[7].um_I.ana[0] ;
 wire \top_I.branch[29].block[7].um_I.ana[1] ;
 wire \top_I.branch[29].block[7].um_I.ana[2] ;
 wire \top_I.branch[29].block[7].um_I.ana[3] ;
 wire \top_I.branch[29].block[7].um_I.ana[4] ;
 wire \top_I.branch[29].block[7].um_I.ana[5] ;
 wire \top_I.branch[29].block[7].um_I.ana[6] ;
 wire \top_I.branch[29].block[7].um_I.ana[7] ;
 wire \top_I.branch[29].block[7].um_I.clk ;
 wire \top_I.branch[29].block[7].um_I.ena ;
 wire \top_I.branch[29].block[7].um_I.iw[10] ;
 wire \top_I.branch[29].block[7].um_I.iw[11] ;
 wire \top_I.branch[29].block[7].um_I.iw[12] ;
 wire \top_I.branch[29].block[7].um_I.iw[13] ;
 wire \top_I.branch[29].block[7].um_I.iw[14] ;
 wire \top_I.branch[29].block[7].um_I.iw[15] ;
 wire \top_I.branch[29].block[7].um_I.iw[16] ;
 wire \top_I.branch[29].block[7].um_I.iw[17] ;
 wire \top_I.branch[29].block[7].um_I.iw[1] ;
 wire \top_I.branch[29].block[7].um_I.iw[2] ;
 wire \top_I.branch[29].block[7].um_I.iw[3] ;
 wire \top_I.branch[29].block[7].um_I.iw[4] ;
 wire \top_I.branch[29].block[7].um_I.iw[5] ;
 wire \top_I.branch[29].block[7].um_I.iw[6] ;
 wire \top_I.branch[29].block[7].um_I.iw[7] ;
 wire \top_I.branch[29].block[7].um_I.iw[8] ;
 wire \top_I.branch[29].block[7].um_I.iw[9] ;
 wire \top_I.branch[29].block[7].um_I.k_zero ;
 wire \top_I.branch[29].block[7].um_I.pg_vdd ;
 wire \top_I.branch[29].block[8].um_I.ana[0] ;
 wire \top_I.branch[29].block[8].um_I.ana[1] ;
 wire \top_I.branch[29].block[8].um_I.ana[2] ;
 wire \top_I.branch[29].block[8].um_I.ana[3] ;
 wire \top_I.branch[29].block[8].um_I.ana[4] ;
 wire \top_I.branch[29].block[8].um_I.ana[5] ;
 wire \top_I.branch[29].block[8].um_I.ana[6] ;
 wire \top_I.branch[29].block[8].um_I.ana[7] ;
 wire \top_I.branch[29].block[8].um_I.clk ;
 wire \top_I.branch[29].block[8].um_I.ena ;
 wire \top_I.branch[29].block[8].um_I.iw[10] ;
 wire \top_I.branch[29].block[8].um_I.iw[11] ;
 wire \top_I.branch[29].block[8].um_I.iw[12] ;
 wire \top_I.branch[29].block[8].um_I.iw[13] ;
 wire \top_I.branch[29].block[8].um_I.iw[14] ;
 wire \top_I.branch[29].block[8].um_I.iw[15] ;
 wire \top_I.branch[29].block[8].um_I.iw[16] ;
 wire \top_I.branch[29].block[8].um_I.iw[17] ;
 wire \top_I.branch[29].block[8].um_I.iw[1] ;
 wire \top_I.branch[29].block[8].um_I.iw[2] ;
 wire \top_I.branch[29].block[8].um_I.iw[3] ;
 wire \top_I.branch[29].block[8].um_I.iw[4] ;
 wire \top_I.branch[29].block[8].um_I.iw[5] ;
 wire \top_I.branch[29].block[8].um_I.iw[6] ;
 wire \top_I.branch[29].block[8].um_I.iw[7] ;
 wire \top_I.branch[29].block[8].um_I.iw[8] ;
 wire \top_I.branch[29].block[8].um_I.iw[9] ;
 wire \top_I.branch[29].block[8].um_I.k_zero ;
 wire \top_I.branch[29].block[8].um_I.pg_vdd ;
 wire \top_I.branch[29].block[9].um_I.ana[0] ;
 wire \top_I.branch[29].block[9].um_I.ana[1] ;
 wire \top_I.branch[29].block[9].um_I.ana[2] ;
 wire \top_I.branch[29].block[9].um_I.ana[3] ;
 wire \top_I.branch[29].block[9].um_I.ana[4] ;
 wire \top_I.branch[29].block[9].um_I.ana[5] ;
 wire \top_I.branch[29].block[9].um_I.ana[6] ;
 wire \top_I.branch[29].block[9].um_I.ana[7] ;
 wire \top_I.branch[29].block[9].um_I.clk ;
 wire \top_I.branch[29].block[9].um_I.ena ;
 wire \top_I.branch[29].block[9].um_I.iw[10] ;
 wire \top_I.branch[29].block[9].um_I.iw[11] ;
 wire \top_I.branch[29].block[9].um_I.iw[12] ;
 wire \top_I.branch[29].block[9].um_I.iw[13] ;
 wire \top_I.branch[29].block[9].um_I.iw[14] ;
 wire \top_I.branch[29].block[9].um_I.iw[15] ;
 wire \top_I.branch[29].block[9].um_I.iw[16] ;
 wire \top_I.branch[29].block[9].um_I.iw[17] ;
 wire \top_I.branch[29].block[9].um_I.iw[1] ;
 wire \top_I.branch[29].block[9].um_I.iw[2] ;
 wire \top_I.branch[29].block[9].um_I.iw[3] ;
 wire \top_I.branch[29].block[9].um_I.iw[4] ;
 wire \top_I.branch[29].block[9].um_I.iw[5] ;
 wire \top_I.branch[29].block[9].um_I.iw[6] ;
 wire \top_I.branch[29].block[9].um_I.iw[7] ;
 wire \top_I.branch[29].block[9].um_I.iw[8] ;
 wire \top_I.branch[29].block[9].um_I.iw[9] ;
 wire \top_I.branch[29].block[9].um_I.k_zero ;
 wire \top_I.branch[29].block[9].um_I.pg_vdd ;
 wire \top_I.branch[29].l_addr[0] ;
 wire \top_I.branch[29].l_addr[1] ;
 wire \top_I.branch[2].block[0].um_I.ana[0] ;
 wire \top_I.branch[2].block[0].um_I.ana[1] ;
 wire \top_I.branch[2].block[0].um_I.ana[2] ;
 wire \top_I.branch[2].block[0].um_I.ana[3] ;
 wire \top_I.branch[2].block[0].um_I.ana[4] ;
 wire \top_I.branch[2].block[0].um_I.ana[5] ;
 wire \top_I.branch[2].block[0].um_I.ana[6] ;
 wire \top_I.branch[2].block[0].um_I.ana[7] ;
 wire \top_I.branch[2].block[0].um_I.clk ;
 wire \top_I.branch[2].block[0].um_I.ena ;
 wire \top_I.branch[2].block[0].um_I.iw[10] ;
 wire \top_I.branch[2].block[0].um_I.iw[11] ;
 wire \top_I.branch[2].block[0].um_I.iw[12] ;
 wire \top_I.branch[2].block[0].um_I.iw[13] ;
 wire \top_I.branch[2].block[0].um_I.iw[14] ;
 wire \top_I.branch[2].block[0].um_I.iw[15] ;
 wire \top_I.branch[2].block[0].um_I.iw[16] ;
 wire \top_I.branch[2].block[0].um_I.iw[17] ;
 wire \top_I.branch[2].block[0].um_I.iw[1] ;
 wire \top_I.branch[2].block[0].um_I.iw[2] ;
 wire \top_I.branch[2].block[0].um_I.iw[3] ;
 wire \top_I.branch[2].block[0].um_I.iw[4] ;
 wire \top_I.branch[2].block[0].um_I.iw[5] ;
 wire \top_I.branch[2].block[0].um_I.iw[6] ;
 wire \top_I.branch[2].block[0].um_I.iw[7] ;
 wire \top_I.branch[2].block[0].um_I.iw[8] ;
 wire \top_I.branch[2].block[0].um_I.iw[9] ;
 wire \top_I.branch[2].block[0].um_I.k_zero ;
 wire \top_I.branch[2].block[0].um_I.pg_vdd ;
 wire \top_I.branch[2].block[10].um_I.ana[0] ;
 wire \top_I.branch[2].block[10].um_I.ana[1] ;
 wire \top_I.branch[2].block[10].um_I.ana[2] ;
 wire \top_I.branch[2].block[10].um_I.ana[3] ;
 wire \top_I.branch[2].block[10].um_I.ana[4] ;
 wire \top_I.branch[2].block[10].um_I.ana[5] ;
 wire \top_I.branch[2].block[10].um_I.ana[6] ;
 wire \top_I.branch[2].block[10].um_I.ana[7] ;
 wire \top_I.branch[2].block[10].um_I.clk ;
 wire \top_I.branch[2].block[10].um_I.ena ;
 wire \top_I.branch[2].block[10].um_I.iw[10] ;
 wire \top_I.branch[2].block[10].um_I.iw[11] ;
 wire \top_I.branch[2].block[10].um_I.iw[12] ;
 wire \top_I.branch[2].block[10].um_I.iw[13] ;
 wire \top_I.branch[2].block[10].um_I.iw[14] ;
 wire \top_I.branch[2].block[10].um_I.iw[15] ;
 wire \top_I.branch[2].block[10].um_I.iw[16] ;
 wire \top_I.branch[2].block[10].um_I.iw[17] ;
 wire \top_I.branch[2].block[10].um_I.iw[1] ;
 wire \top_I.branch[2].block[10].um_I.iw[2] ;
 wire \top_I.branch[2].block[10].um_I.iw[3] ;
 wire \top_I.branch[2].block[10].um_I.iw[4] ;
 wire \top_I.branch[2].block[10].um_I.iw[5] ;
 wire \top_I.branch[2].block[10].um_I.iw[6] ;
 wire \top_I.branch[2].block[10].um_I.iw[7] ;
 wire \top_I.branch[2].block[10].um_I.iw[8] ;
 wire \top_I.branch[2].block[10].um_I.iw[9] ;
 wire \top_I.branch[2].block[10].um_I.k_zero ;
 wire \top_I.branch[2].block[10].um_I.pg_vdd ;
 wire \top_I.branch[2].block[11].um_I.ana[0] ;
 wire \top_I.branch[2].block[11].um_I.ana[1] ;
 wire \top_I.branch[2].block[11].um_I.ana[2] ;
 wire \top_I.branch[2].block[11].um_I.ana[3] ;
 wire \top_I.branch[2].block[11].um_I.ana[4] ;
 wire \top_I.branch[2].block[11].um_I.ana[5] ;
 wire \top_I.branch[2].block[11].um_I.ana[6] ;
 wire \top_I.branch[2].block[11].um_I.ana[7] ;
 wire \top_I.branch[2].block[11].um_I.clk ;
 wire \top_I.branch[2].block[11].um_I.ena ;
 wire \top_I.branch[2].block[11].um_I.iw[10] ;
 wire \top_I.branch[2].block[11].um_I.iw[11] ;
 wire \top_I.branch[2].block[11].um_I.iw[12] ;
 wire \top_I.branch[2].block[11].um_I.iw[13] ;
 wire \top_I.branch[2].block[11].um_I.iw[14] ;
 wire \top_I.branch[2].block[11].um_I.iw[15] ;
 wire \top_I.branch[2].block[11].um_I.iw[16] ;
 wire \top_I.branch[2].block[11].um_I.iw[17] ;
 wire \top_I.branch[2].block[11].um_I.iw[1] ;
 wire \top_I.branch[2].block[11].um_I.iw[2] ;
 wire \top_I.branch[2].block[11].um_I.iw[3] ;
 wire \top_I.branch[2].block[11].um_I.iw[4] ;
 wire \top_I.branch[2].block[11].um_I.iw[5] ;
 wire \top_I.branch[2].block[11].um_I.iw[6] ;
 wire \top_I.branch[2].block[11].um_I.iw[7] ;
 wire \top_I.branch[2].block[11].um_I.iw[8] ;
 wire \top_I.branch[2].block[11].um_I.iw[9] ;
 wire \top_I.branch[2].block[11].um_I.k_zero ;
 wire \top_I.branch[2].block[11].um_I.pg_vdd ;
 wire \top_I.branch[2].block[12].um_I.ana[0] ;
 wire \top_I.branch[2].block[12].um_I.ana[1] ;
 wire \top_I.branch[2].block[12].um_I.ana[2] ;
 wire \top_I.branch[2].block[12].um_I.ana[3] ;
 wire \top_I.branch[2].block[12].um_I.ana[4] ;
 wire \top_I.branch[2].block[12].um_I.ana[5] ;
 wire \top_I.branch[2].block[12].um_I.ana[6] ;
 wire \top_I.branch[2].block[12].um_I.ana[7] ;
 wire \top_I.branch[2].block[12].um_I.clk ;
 wire \top_I.branch[2].block[12].um_I.ena ;
 wire \top_I.branch[2].block[12].um_I.iw[10] ;
 wire \top_I.branch[2].block[12].um_I.iw[11] ;
 wire \top_I.branch[2].block[12].um_I.iw[12] ;
 wire \top_I.branch[2].block[12].um_I.iw[13] ;
 wire \top_I.branch[2].block[12].um_I.iw[14] ;
 wire \top_I.branch[2].block[12].um_I.iw[15] ;
 wire \top_I.branch[2].block[12].um_I.iw[16] ;
 wire \top_I.branch[2].block[12].um_I.iw[17] ;
 wire \top_I.branch[2].block[12].um_I.iw[1] ;
 wire \top_I.branch[2].block[12].um_I.iw[2] ;
 wire \top_I.branch[2].block[12].um_I.iw[3] ;
 wire \top_I.branch[2].block[12].um_I.iw[4] ;
 wire \top_I.branch[2].block[12].um_I.iw[5] ;
 wire \top_I.branch[2].block[12].um_I.iw[6] ;
 wire \top_I.branch[2].block[12].um_I.iw[7] ;
 wire \top_I.branch[2].block[12].um_I.iw[8] ;
 wire \top_I.branch[2].block[12].um_I.iw[9] ;
 wire \top_I.branch[2].block[12].um_I.k_zero ;
 wire \top_I.branch[2].block[12].um_I.pg_vdd ;
 wire \top_I.branch[2].block[13].um_I.ana[0] ;
 wire \top_I.branch[2].block[13].um_I.ana[1] ;
 wire \top_I.branch[2].block[13].um_I.ana[2] ;
 wire \top_I.branch[2].block[13].um_I.ana[3] ;
 wire \top_I.branch[2].block[13].um_I.ana[4] ;
 wire \top_I.branch[2].block[13].um_I.ana[5] ;
 wire \top_I.branch[2].block[13].um_I.ana[6] ;
 wire \top_I.branch[2].block[13].um_I.ana[7] ;
 wire \top_I.branch[2].block[13].um_I.clk ;
 wire \top_I.branch[2].block[13].um_I.ena ;
 wire \top_I.branch[2].block[13].um_I.iw[10] ;
 wire \top_I.branch[2].block[13].um_I.iw[11] ;
 wire \top_I.branch[2].block[13].um_I.iw[12] ;
 wire \top_I.branch[2].block[13].um_I.iw[13] ;
 wire \top_I.branch[2].block[13].um_I.iw[14] ;
 wire \top_I.branch[2].block[13].um_I.iw[15] ;
 wire \top_I.branch[2].block[13].um_I.iw[16] ;
 wire \top_I.branch[2].block[13].um_I.iw[17] ;
 wire \top_I.branch[2].block[13].um_I.iw[1] ;
 wire \top_I.branch[2].block[13].um_I.iw[2] ;
 wire \top_I.branch[2].block[13].um_I.iw[3] ;
 wire \top_I.branch[2].block[13].um_I.iw[4] ;
 wire \top_I.branch[2].block[13].um_I.iw[5] ;
 wire \top_I.branch[2].block[13].um_I.iw[6] ;
 wire \top_I.branch[2].block[13].um_I.iw[7] ;
 wire \top_I.branch[2].block[13].um_I.iw[8] ;
 wire \top_I.branch[2].block[13].um_I.iw[9] ;
 wire \top_I.branch[2].block[13].um_I.k_zero ;
 wire \top_I.branch[2].block[13].um_I.pg_vdd ;
 wire \top_I.branch[2].block[14].um_I.ana[0] ;
 wire \top_I.branch[2].block[14].um_I.ana[1] ;
 wire \top_I.branch[2].block[14].um_I.ana[2] ;
 wire \top_I.branch[2].block[14].um_I.ana[3] ;
 wire \top_I.branch[2].block[14].um_I.ana[4] ;
 wire \top_I.branch[2].block[14].um_I.ana[5] ;
 wire \top_I.branch[2].block[14].um_I.ana[6] ;
 wire \top_I.branch[2].block[14].um_I.ana[7] ;
 wire \top_I.branch[2].block[14].um_I.clk ;
 wire \top_I.branch[2].block[14].um_I.ena ;
 wire \top_I.branch[2].block[14].um_I.iw[10] ;
 wire \top_I.branch[2].block[14].um_I.iw[11] ;
 wire \top_I.branch[2].block[14].um_I.iw[12] ;
 wire \top_I.branch[2].block[14].um_I.iw[13] ;
 wire \top_I.branch[2].block[14].um_I.iw[14] ;
 wire \top_I.branch[2].block[14].um_I.iw[15] ;
 wire \top_I.branch[2].block[14].um_I.iw[16] ;
 wire \top_I.branch[2].block[14].um_I.iw[17] ;
 wire \top_I.branch[2].block[14].um_I.iw[1] ;
 wire \top_I.branch[2].block[14].um_I.iw[2] ;
 wire \top_I.branch[2].block[14].um_I.iw[3] ;
 wire \top_I.branch[2].block[14].um_I.iw[4] ;
 wire \top_I.branch[2].block[14].um_I.iw[5] ;
 wire \top_I.branch[2].block[14].um_I.iw[6] ;
 wire \top_I.branch[2].block[14].um_I.iw[7] ;
 wire \top_I.branch[2].block[14].um_I.iw[8] ;
 wire \top_I.branch[2].block[14].um_I.iw[9] ;
 wire \top_I.branch[2].block[14].um_I.k_zero ;
 wire \top_I.branch[2].block[14].um_I.pg_vdd ;
 wire \top_I.branch[2].block[15].um_I.ana[0] ;
 wire \top_I.branch[2].block[15].um_I.ana[1] ;
 wire \top_I.branch[2].block[15].um_I.ana[2] ;
 wire \top_I.branch[2].block[15].um_I.ana[3] ;
 wire \top_I.branch[2].block[15].um_I.ana[4] ;
 wire \top_I.branch[2].block[15].um_I.ana[5] ;
 wire \top_I.branch[2].block[15].um_I.ana[6] ;
 wire \top_I.branch[2].block[15].um_I.ana[7] ;
 wire \top_I.branch[2].block[15].um_I.clk ;
 wire \top_I.branch[2].block[15].um_I.ena ;
 wire \top_I.branch[2].block[15].um_I.iw[10] ;
 wire \top_I.branch[2].block[15].um_I.iw[11] ;
 wire \top_I.branch[2].block[15].um_I.iw[12] ;
 wire \top_I.branch[2].block[15].um_I.iw[13] ;
 wire \top_I.branch[2].block[15].um_I.iw[14] ;
 wire \top_I.branch[2].block[15].um_I.iw[15] ;
 wire \top_I.branch[2].block[15].um_I.iw[16] ;
 wire \top_I.branch[2].block[15].um_I.iw[17] ;
 wire \top_I.branch[2].block[15].um_I.iw[1] ;
 wire \top_I.branch[2].block[15].um_I.iw[2] ;
 wire \top_I.branch[2].block[15].um_I.iw[3] ;
 wire \top_I.branch[2].block[15].um_I.iw[4] ;
 wire \top_I.branch[2].block[15].um_I.iw[5] ;
 wire \top_I.branch[2].block[15].um_I.iw[6] ;
 wire \top_I.branch[2].block[15].um_I.iw[7] ;
 wire \top_I.branch[2].block[15].um_I.iw[8] ;
 wire \top_I.branch[2].block[15].um_I.iw[9] ;
 wire \top_I.branch[2].block[15].um_I.k_zero ;
 wire \top_I.branch[2].block[15].um_I.pg_vdd ;
 wire \top_I.branch[2].block[1].um_I.ana[0] ;
 wire \top_I.branch[2].block[1].um_I.ana[1] ;
 wire \top_I.branch[2].block[1].um_I.ana[2] ;
 wire \top_I.branch[2].block[1].um_I.ana[3] ;
 wire \top_I.branch[2].block[1].um_I.ana[4] ;
 wire \top_I.branch[2].block[1].um_I.ana[5] ;
 wire \top_I.branch[2].block[1].um_I.ana[6] ;
 wire \top_I.branch[2].block[1].um_I.ana[7] ;
 wire \top_I.branch[2].block[1].um_I.clk ;
 wire \top_I.branch[2].block[1].um_I.ena ;
 wire \top_I.branch[2].block[1].um_I.iw[10] ;
 wire \top_I.branch[2].block[1].um_I.iw[11] ;
 wire \top_I.branch[2].block[1].um_I.iw[12] ;
 wire \top_I.branch[2].block[1].um_I.iw[13] ;
 wire \top_I.branch[2].block[1].um_I.iw[14] ;
 wire \top_I.branch[2].block[1].um_I.iw[15] ;
 wire \top_I.branch[2].block[1].um_I.iw[16] ;
 wire \top_I.branch[2].block[1].um_I.iw[17] ;
 wire \top_I.branch[2].block[1].um_I.iw[1] ;
 wire \top_I.branch[2].block[1].um_I.iw[2] ;
 wire \top_I.branch[2].block[1].um_I.iw[3] ;
 wire \top_I.branch[2].block[1].um_I.iw[4] ;
 wire \top_I.branch[2].block[1].um_I.iw[5] ;
 wire \top_I.branch[2].block[1].um_I.iw[6] ;
 wire \top_I.branch[2].block[1].um_I.iw[7] ;
 wire \top_I.branch[2].block[1].um_I.iw[8] ;
 wire \top_I.branch[2].block[1].um_I.iw[9] ;
 wire \top_I.branch[2].block[1].um_I.k_zero ;
 wire \top_I.branch[2].block[1].um_I.pg_vdd ;
 wire \top_I.branch[2].block[2].um_I.ana[0] ;
 wire \top_I.branch[2].block[2].um_I.ana[1] ;
 wire \top_I.branch[2].block[2].um_I.ana[2] ;
 wire \top_I.branch[2].block[2].um_I.ana[3] ;
 wire \top_I.branch[2].block[2].um_I.ana[4] ;
 wire \top_I.branch[2].block[2].um_I.ana[5] ;
 wire \top_I.branch[2].block[2].um_I.ana[6] ;
 wire \top_I.branch[2].block[2].um_I.ana[7] ;
 wire \top_I.branch[2].block[2].um_I.clk ;
 wire \top_I.branch[2].block[2].um_I.ena ;
 wire \top_I.branch[2].block[2].um_I.iw[10] ;
 wire \top_I.branch[2].block[2].um_I.iw[11] ;
 wire \top_I.branch[2].block[2].um_I.iw[12] ;
 wire \top_I.branch[2].block[2].um_I.iw[13] ;
 wire \top_I.branch[2].block[2].um_I.iw[14] ;
 wire \top_I.branch[2].block[2].um_I.iw[15] ;
 wire \top_I.branch[2].block[2].um_I.iw[16] ;
 wire \top_I.branch[2].block[2].um_I.iw[17] ;
 wire \top_I.branch[2].block[2].um_I.iw[1] ;
 wire \top_I.branch[2].block[2].um_I.iw[2] ;
 wire \top_I.branch[2].block[2].um_I.iw[3] ;
 wire \top_I.branch[2].block[2].um_I.iw[4] ;
 wire \top_I.branch[2].block[2].um_I.iw[5] ;
 wire \top_I.branch[2].block[2].um_I.iw[6] ;
 wire \top_I.branch[2].block[2].um_I.iw[7] ;
 wire \top_I.branch[2].block[2].um_I.iw[8] ;
 wire \top_I.branch[2].block[2].um_I.iw[9] ;
 wire \top_I.branch[2].block[2].um_I.k_zero ;
 wire \top_I.branch[2].block[2].um_I.pg_vdd ;
 wire \top_I.branch[2].block[3].um_I.ana[0] ;
 wire \top_I.branch[2].block[3].um_I.ana[1] ;
 wire \top_I.branch[2].block[3].um_I.ana[2] ;
 wire \top_I.branch[2].block[3].um_I.ana[3] ;
 wire \top_I.branch[2].block[3].um_I.ana[4] ;
 wire \top_I.branch[2].block[3].um_I.ana[5] ;
 wire \top_I.branch[2].block[3].um_I.ana[6] ;
 wire \top_I.branch[2].block[3].um_I.ana[7] ;
 wire \top_I.branch[2].block[3].um_I.clk ;
 wire \top_I.branch[2].block[3].um_I.ena ;
 wire \top_I.branch[2].block[3].um_I.iw[10] ;
 wire \top_I.branch[2].block[3].um_I.iw[11] ;
 wire \top_I.branch[2].block[3].um_I.iw[12] ;
 wire \top_I.branch[2].block[3].um_I.iw[13] ;
 wire \top_I.branch[2].block[3].um_I.iw[14] ;
 wire \top_I.branch[2].block[3].um_I.iw[15] ;
 wire \top_I.branch[2].block[3].um_I.iw[16] ;
 wire \top_I.branch[2].block[3].um_I.iw[17] ;
 wire \top_I.branch[2].block[3].um_I.iw[1] ;
 wire \top_I.branch[2].block[3].um_I.iw[2] ;
 wire \top_I.branch[2].block[3].um_I.iw[3] ;
 wire \top_I.branch[2].block[3].um_I.iw[4] ;
 wire \top_I.branch[2].block[3].um_I.iw[5] ;
 wire \top_I.branch[2].block[3].um_I.iw[6] ;
 wire \top_I.branch[2].block[3].um_I.iw[7] ;
 wire \top_I.branch[2].block[3].um_I.iw[8] ;
 wire \top_I.branch[2].block[3].um_I.iw[9] ;
 wire \top_I.branch[2].block[3].um_I.k_zero ;
 wire \top_I.branch[2].block[3].um_I.pg_vdd ;
 wire \top_I.branch[2].block[4].um_I.ana[0] ;
 wire \top_I.branch[2].block[4].um_I.ana[1] ;
 wire \top_I.branch[2].block[4].um_I.ana[2] ;
 wire \top_I.branch[2].block[4].um_I.ana[3] ;
 wire \top_I.branch[2].block[4].um_I.ana[4] ;
 wire \top_I.branch[2].block[4].um_I.ana[5] ;
 wire \top_I.branch[2].block[4].um_I.ana[6] ;
 wire \top_I.branch[2].block[4].um_I.ana[7] ;
 wire \top_I.branch[2].block[4].um_I.clk ;
 wire \top_I.branch[2].block[4].um_I.ena ;
 wire \top_I.branch[2].block[4].um_I.iw[10] ;
 wire \top_I.branch[2].block[4].um_I.iw[11] ;
 wire \top_I.branch[2].block[4].um_I.iw[12] ;
 wire \top_I.branch[2].block[4].um_I.iw[13] ;
 wire \top_I.branch[2].block[4].um_I.iw[14] ;
 wire \top_I.branch[2].block[4].um_I.iw[15] ;
 wire \top_I.branch[2].block[4].um_I.iw[16] ;
 wire \top_I.branch[2].block[4].um_I.iw[17] ;
 wire \top_I.branch[2].block[4].um_I.iw[1] ;
 wire \top_I.branch[2].block[4].um_I.iw[2] ;
 wire \top_I.branch[2].block[4].um_I.iw[3] ;
 wire \top_I.branch[2].block[4].um_I.iw[4] ;
 wire \top_I.branch[2].block[4].um_I.iw[5] ;
 wire \top_I.branch[2].block[4].um_I.iw[6] ;
 wire \top_I.branch[2].block[4].um_I.iw[7] ;
 wire \top_I.branch[2].block[4].um_I.iw[8] ;
 wire \top_I.branch[2].block[4].um_I.iw[9] ;
 wire \top_I.branch[2].block[4].um_I.k_zero ;
 wire \top_I.branch[2].block[4].um_I.pg_vdd ;
 wire \top_I.branch[2].block[5].um_I.ana[0] ;
 wire \top_I.branch[2].block[5].um_I.ana[1] ;
 wire \top_I.branch[2].block[5].um_I.ana[2] ;
 wire \top_I.branch[2].block[5].um_I.ana[3] ;
 wire \top_I.branch[2].block[5].um_I.ana[4] ;
 wire \top_I.branch[2].block[5].um_I.ana[5] ;
 wire \top_I.branch[2].block[5].um_I.ana[6] ;
 wire \top_I.branch[2].block[5].um_I.ana[7] ;
 wire \top_I.branch[2].block[5].um_I.clk ;
 wire \top_I.branch[2].block[5].um_I.ena ;
 wire \top_I.branch[2].block[5].um_I.iw[10] ;
 wire \top_I.branch[2].block[5].um_I.iw[11] ;
 wire \top_I.branch[2].block[5].um_I.iw[12] ;
 wire \top_I.branch[2].block[5].um_I.iw[13] ;
 wire \top_I.branch[2].block[5].um_I.iw[14] ;
 wire \top_I.branch[2].block[5].um_I.iw[15] ;
 wire \top_I.branch[2].block[5].um_I.iw[16] ;
 wire \top_I.branch[2].block[5].um_I.iw[17] ;
 wire \top_I.branch[2].block[5].um_I.iw[1] ;
 wire \top_I.branch[2].block[5].um_I.iw[2] ;
 wire \top_I.branch[2].block[5].um_I.iw[3] ;
 wire \top_I.branch[2].block[5].um_I.iw[4] ;
 wire \top_I.branch[2].block[5].um_I.iw[5] ;
 wire \top_I.branch[2].block[5].um_I.iw[6] ;
 wire \top_I.branch[2].block[5].um_I.iw[7] ;
 wire \top_I.branch[2].block[5].um_I.iw[8] ;
 wire \top_I.branch[2].block[5].um_I.iw[9] ;
 wire \top_I.branch[2].block[5].um_I.k_zero ;
 wire \top_I.branch[2].block[5].um_I.pg_vdd ;
 wire \top_I.branch[2].block[6].um_I.ana[0] ;
 wire \top_I.branch[2].block[6].um_I.ana[1] ;
 wire \top_I.branch[2].block[6].um_I.ana[2] ;
 wire \top_I.branch[2].block[6].um_I.ana[3] ;
 wire \top_I.branch[2].block[6].um_I.ana[4] ;
 wire \top_I.branch[2].block[6].um_I.ana[5] ;
 wire \top_I.branch[2].block[6].um_I.ana[6] ;
 wire \top_I.branch[2].block[6].um_I.ana[7] ;
 wire \top_I.branch[2].block[6].um_I.clk ;
 wire \top_I.branch[2].block[6].um_I.ena ;
 wire \top_I.branch[2].block[6].um_I.iw[10] ;
 wire \top_I.branch[2].block[6].um_I.iw[11] ;
 wire \top_I.branch[2].block[6].um_I.iw[12] ;
 wire \top_I.branch[2].block[6].um_I.iw[13] ;
 wire \top_I.branch[2].block[6].um_I.iw[14] ;
 wire \top_I.branch[2].block[6].um_I.iw[15] ;
 wire \top_I.branch[2].block[6].um_I.iw[16] ;
 wire \top_I.branch[2].block[6].um_I.iw[17] ;
 wire \top_I.branch[2].block[6].um_I.iw[1] ;
 wire \top_I.branch[2].block[6].um_I.iw[2] ;
 wire \top_I.branch[2].block[6].um_I.iw[3] ;
 wire \top_I.branch[2].block[6].um_I.iw[4] ;
 wire \top_I.branch[2].block[6].um_I.iw[5] ;
 wire \top_I.branch[2].block[6].um_I.iw[6] ;
 wire \top_I.branch[2].block[6].um_I.iw[7] ;
 wire \top_I.branch[2].block[6].um_I.iw[8] ;
 wire \top_I.branch[2].block[6].um_I.iw[9] ;
 wire \top_I.branch[2].block[6].um_I.k_zero ;
 wire \top_I.branch[2].block[6].um_I.pg_vdd ;
 wire \top_I.branch[2].block[7].um_I.ana[0] ;
 wire \top_I.branch[2].block[7].um_I.ana[1] ;
 wire \top_I.branch[2].block[7].um_I.ana[2] ;
 wire \top_I.branch[2].block[7].um_I.ana[3] ;
 wire \top_I.branch[2].block[7].um_I.ana[4] ;
 wire \top_I.branch[2].block[7].um_I.ana[5] ;
 wire \top_I.branch[2].block[7].um_I.ana[6] ;
 wire \top_I.branch[2].block[7].um_I.ana[7] ;
 wire \top_I.branch[2].block[7].um_I.clk ;
 wire \top_I.branch[2].block[7].um_I.ena ;
 wire \top_I.branch[2].block[7].um_I.iw[10] ;
 wire \top_I.branch[2].block[7].um_I.iw[11] ;
 wire \top_I.branch[2].block[7].um_I.iw[12] ;
 wire \top_I.branch[2].block[7].um_I.iw[13] ;
 wire \top_I.branch[2].block[7].um_I.iw[14] ;
 wire \top_I.branch[2].block[7].um_I.iw[15] ;
 wire \top_I.branch[2].block[7].um_I.iw[16] ;
 wire \top_I.branch[2].block[7].um_I.iw[17] ;
 wire \top_I.branch[2].block[7].um_I.iw[1] ;
 wire \top_I.branch[2].block[7].um_I.iw[2] ;
 wire \top_I.branch[2].block[7].um_I.iw[3] ;
 wire \top_I.branch[2].block[7].um_I.iw[4] ;
 wire \top_I.branch[2].block[7].um_I.iw[5] ;
 wire \top_I.branch[2].block[7].um_I.iw[6] ;
 wire \top_I.branch[2].block[7].um_I.iw[7] ;
 wire \top_I.branch[2].block[7].um_I.iw[8] ;
 wire \top_I.branch[2].block[7].um_I.iw[9] ;
 wire \top_I.branch[2].block[7].um_I.k_zero ;
 wire \top_I.branch[2].block[7].um_I.pg_vdd ;
 wire \top_I.branch[2].block[8].um_I.ana[0] ;
 wire \top_I.branch[2].block[8].um_I.ana[1] ;
 wire \top_I.branch[2].block[8].um_I.ana[2] ;
 wire \top_I.branch[2].block[8].um_I.ana[3] ;
 wire \top_I.branch[2].block[8].um_I.ana[4] ;
 wire \top_I.branch[2].block[8].um_I.ana[5] ;
 wire \top_I.branch[2].block[8].um_I.ana[6] ;
 wire \top_I.branch[2].block[8].um_I.ana[7] ;
 wire \top_I.branch[2].block[8].um_I.clk ;
 wire \top_I.branch[2].block[8].um_I.ena ;
 wire \top_I.branch[2].block[8].um_I.iw[10] ;
 wire \top_I.branch[2].block[8].um_I.iw[11] ;
 wire \top_I.branch[2].block[8].um_I.iw[12] ;
 wire \top_I.branch[2].block[8].um_I.iw[13] ;
 wire \top_I.branch[2].block[8].um_I.iw[14] ;
 wire \top_I.branch[2].block[8].um_I.iw[15] ;
 wire \top_I.branch[2].block[8].um_I.iw[16] ;
 wire \top_I.branch[2].block[8].um_I.iw[17] ;
 wire \top_I.branch[2].block[8].um_I.iw[1] ;
 wire \top_I.branch[2].block[8].um_I.iw[2] ;
 wire \top_I.branch[2].block[8].um_I.iw[3] ;
 wire \top_I.branch[2].block[8].um_I.iw[4] ;
 wire \top_I.branch[2].block[8].um_I.iw[5] ;
 wire \top_I.branch[2].block[8].um_I.iw[6] ;
 wire \top_I.branch[2].block[8].um_I.iw[7] ;
 wire \top_I.branch[2].block[8].um_I.iw[8] ;
 wire \top_I.branch[2].block[8].um_I.iw[9] ;
 wire \top_I.branch[2].block[8].um_I.k_zero ;
 wire \top_I.branch[2].block[8].um_I.pg_vdd ;
 wire \top_I.branch[2].block[9].um_I.ana[0] ;
 wire \top_I.branch[2].block[9].um_I.ana[1] ;
 wire \top_I.branch[2].block[9].um_I.ana[2] ;
 wire \top_I.branch[2].block[9].um_I.ana[3] ;
 wire \top_I.branch[2].block[9].um_I.ana[4] ;
 wire \top_I.branch[2].block[9].um_I.ana[5] ;
 wire \top_I.branch[2].block[9].um_I.ana[6] ;
 wire \top_I.branch[2].block[9].um_I.ana[7] ;
 wire \top_I.branch[2].block[9].um_I.clk ;
 wire \top_I.branch[2].block[9].um_I.ena ;
 wire \top_I.branch[2].block[9].um_I.iw[10] ;
 wire \top_I.branch[2].block[9].um_I.iw[11] ;
 wire \top_I.branch[2].block[9].um_I.iw[12] ;
 wire \top_I.branch[2].block[9].um_I.iw[13] ;
 wire \top_I.branch[2].block[9].um_I.iw[14] ;
 wire \top_I.branch[2].block[9].um_I.iw[15] ;
 wire \top_I.branch[2].block[9].um_I.iw[16] ;
 wire \top_I.branch[2].block[9].um_I.iw[17] ;
 wire \top_I.branch[2].block[9].um_I.iw[1] ;
 wire \top_I.branch[2].block[9].um_I.iw[2] ;
 wire \top_I.branch[2].block[9].um_I.iw[3] ;
 wire \top_I.branch[2].block[9].um_I.iw[4] ;
 wire \top_I.branch[2].block[9].um_I.iw[5] ;
 wire \top_I.branch[2].block[9].um_I.iw[6] ;
 wire \top_I.branch[2].block[9].um_I.iw[7] ;
 wire \top_I.branch[2].block[9].um_I.iw[8] ;
 wire \top_I.branch[2].block[9].um_I.iw[9] ;
 wire \top_I.branch[2].block[9].um_I.k_zero ;
 wire \top_I.branch[2].block[9].um_I.pg_vdd ;
 wire \top_I.branch[2].l_addr[0] ;
 wire \top_I.branch[2].l_addr[1] ;
 wire \top_I.branch[30].block[0].um_I.ana[0] ;
 wire \top_I.branch[30].block[0].um_I.ana[1] ;
 wire \top_I.branch[30].block[0].um_I.ana[2] ;
 wire \top_I.branch[30].block[0].um_I.ana[3] ;
 wire \top_I.branch[30].block[0].um_I.ana[4] ;
 wire \top_I.branch[30].block[0].um_I.ana[5] ;
 wire \top_I.branch[30].block[0].um_I.ana[6] ;
 wire \top_I.branch[30].block[0].um_I.ana[7] ;
 wire \top_I.branch[30].block[0].um_I.clk ;
 wire \top_I.branch[30].block[0].um_I.ena ;
 wire \top_I.branch[30].block[0].um_I.iw[10] ;
 wire \top_I.branch[30].block[0].um_I.iw[11] ;
 wire \top_I.branch[30].block[0].um_I.iw[12] ;
 wire \top_I.branch[30].block[0].um_I.iw[13] ;
 wire \top_I.branch[30].block[0].um_I.iw[14] ;
 wire \top_I.branch[30].block[0].um_I.iw[15] ;
 wire \top_I.branch[30].block[0].um_I.iw[16] ;
 wire \top_I.branch[30].block[0].um_I.iw[17] ;
 wire \top_I.branch[30].block[0].um_I.iw[1] ;
 wire \top_I.branch[30].block[0].um_I.iw[2] ;
 wire \top_I.branch[30].block[0].um_I.iw[3] ;
 wire \top_I.branch[30].block[0].um_I.iw[4] ;
 wire \top_I.branch[30].block[0].um_I.iw[5] ;
 wire \top_I.branch[30].block[0].um_I.iw[6] ;
 wire \top_I.branch[30].block[0].um_I.iw[7] ;
 wire \top_I.branch[30].block[0].um_I.iw[8] ;
 wire \top_I.branch[30].block[0].um_I.iw[9] ;
 wire \top_I.branch[30].block[0].um_I.k_zero ;
 wire \top_I.branch[30].block[0].um_I.ow[0] ;
 wire \top_I.branch[30].block[0].um_I.ow[10] ;
 wire \top_I.branch[30].block[0].um_I.ow[11] ;
 wire \top_I.branch[30].block[0].um_I.ow[12] ;
 wire \top_I.branch[30].block[0].um_I.ow[13] ;
 wire \top_I.branch[30].block[0].um_I.ow[14] ;
 wire \top_I.branch[30].block[0].um_I.ow[15] ;
 wire \top_I.branch[30].block[0].um_I.ow[16] ;
 wire \top_I.branch[30].block[0].um_I.ow[17] ;
 wire \top_I.branch[30].block[0].um_I.ow[18] ;
 wire \top_I.branch[30].block[0].um_I.ow[19] ;
 wire \top_I.branch[30].block[0].um_I.ow[1] ;
 wire \top_I.branch[30].block[0].um_I.ow[20] ;
 wire \top_I.branch[30].block[0].um_I.ow[21] ;
 wire \top_I.branch[30].block[0].um_I.ow[22] ;
 wire \top_I.branch[30].block[0].um_I.ow[23] ;
 wire \top_I.branch[30].block[0].um_I.ow[2] ;
 wire \top_I.branch[30].block[0].um_I.ow[3] ;
 wire \top_I.branch[30].block[0].um_I.ow[4] ;
 wire \top_I.branch[30].block[0].um_I.ow[5] ;
 wire \top_I.branch[30].block[0].um_I.ow[6] ;
 wire \top_I.branch[30].block[0].um_I.ow[7] ;
 wire \top_I.branch[30].block[0].um_I.ow[8] ;
 wire \top_I.branch[30].block[0].um_I.ow[9] ;
 wire \top_I.branch[30].block[0].um_I.pg_vdd ;
 wire \top_I.branch[30].block[10].um_I.ana[0] ;
 wire \top_I.branch[30].block[10].um_I.ana[1] ;
 wire \top_I.branch[30].block[10].um_I.ana[2] ;
 wire \top_I.branch[30].block[10].um_I.ana[3] ;
 wire \top_I.branch[30].block[10].um_I.ana[4] ;
 wire \top_I.branch[30].block[10].um_I.ana[5] ;
 wire \top_I.branch[30].block[10].um_I.ana[6] ;
 wire \top_I.branch[30].block[10].um_I.ana[7] ;
 wire \top_I.branch[30].block[10].um_I.clk ;
 wire \top_I.branch[30].block[10].um_I.ena ;
 wire \top_I.branch[30].block[10].um_I.iw[10] ;
 wire \top_I.branch[30].block[10].um_I.iw[11] ;
 wire \top_I.branch[30].block[10].um_I.iw[12] ;
 wire \top_I.branch[30].block[10].um_I.iw[13] ;
 wire \top_I.branch[30].block[10].um_I.iw[14] ;
 wire \top_I.branch[30].block[10].um_I.iw[15] ;
 wire \top_I.branch[30].block[10].um_I.iw[16] ;
 wire \top_I.branch[30].block[10].um_I.iw[17] ;
 wire \top_I.branch[30].block[10].um_I.iw[1] ;
 wire \top_I.branch[30].block[10].um_I.iw[2] ;
 wire \top_I.branch[30].block[10].um_I.iw[3] ;
 wire \top_I.branch[30].block[10].um_I.iw[4] ;
 wire \top_I.branch[30].block[10].um_I.iw[5] ;
 wire \top_I.branch[30].block[10].um_I.iw[6] ;
 wire \top_I.branch[30].block[10].um_I.iw[7] ;
 wire \top_I.branch[30].block[10].um_I.iw[8] ;
 wire \top_I.branch[30].block[10].um_I.iw[9] ;
 wire \top_I.branch[30].block[10].um_I.k_zero ;
 wire \top_I.branch[30].block[10].um_I.pg_vdd ;
 wire \top_I.branch[30].block[11].um_I.ana[0] ;
 wire \top_I.branch[30].block[11].um_I.ana[1] ;
 wire \top_I.branch[30].block[11].um_I.ana[2] ;
 wire \top_I.branch[30].block[11].um_I.ana[3] ;
 wire \top_I.branch[30].block[11].um_I.ana[4] ;
 wire \top_I.branch[30].block[11].um_I.ana[5] ;
 wire \top_I.branch[30].block[11].um_I.ana[6] ;
 wire \top_I.branch[30].block[11].um_I.ana[7] ;
 wire \top_I.branch[30].block[11].um_I.clk ;
 wire \top_I.branch[30].block[11].um_I.ena ;
 wire \top_I.branch[30].block[11].um_I.iw[10] ;
 wire \top_I.branch[30].block[11].um_I.iw[11] ;
 wire \top_I.branch[30].block[11].um_I.iw[12] ;
 wire \top_I.branch[30].block[11].um_I.iw[13] ;
 wire \top_I.branch[30].block[11].um_I.iw[14] ;
 wire \top_I.branch[30].block[11].um_I.iw[15] ;
 wire \top_I.branch[30].block[11].um_I.iw[16] ;
 wire \top_I.branch[30].block[11].um_I.iw[17] ;
 wire \top_I.branch[30].block[11].um_I.iw[1] ;
 wire \top_I.branch[30].block[11].um_I.iw[2] ;
 wire \top_I.branch[30].block[11].um_I.iw[3] ;
 wire \top_I.branch[30].block[11].um_I.iw[4] ;
 wire \top_I.branch[30].block[11].um_I.iw[5] ;
 wire \top_I.branch[30].block[11].um_I.iw[6] ;
 wire \top_I.branch[30].block[11].um_I.iw[7] ;
 wire \top_I.branch[30].block[11].um_I.iw[8] ;
 wire \top_I.branch[30].block[11].um_I.iw[9] ;
 wire \top_I.branch[30].block[11].um_I.k_zero ;
 wire \top_I.branch[30].block[11].um_I.ow[0] ;
 wire \top_I.branch[30].block[11].um_I.ow[10] ;
 wire \top_I.branch[30].block[11].um_I.ow[11] ;
 wire \top_I.branch[30].block[11].um_I.ow[12] ;
 wire \top_I.branch[30].block[11].um_I.ow[13] ;
 wire \top_I.branch[30].block[11].um_I.ow[14] ;
 wire \top_I.branch[30].block[11].um_I.ow[15] ;
 wire \top_I.branch[30].block[11].um_I.ow[16] ;
 wire \top_I.branch[30].block[11].um_I.ow[17] ;
 wire \top_I.branch[30].block[11].um_I.ow[18] ;
 wire \top_I.branch[30].block[11].um_I.ow[19] ;
 wire \top_I.branch[30].block[11].um_I.ow[1] ;
 wire \top_I.branch[30].block[11].um_I.ow[20] ;
 wire \top_I.branch[30].block[11].um_I.ow[21] ;
 wire \top_I.branch[30].block[11].um_I.ow[22] ;
 wire \top_I.branch[30].block[11].um_I.ow[23] ;
 wire \top_I.branch[30].block[11].um_I.ow[2] ;
 wire \top_I.branch[30].block[11].um_I.ow[3] ;
 wire \top_I.branch[30].block[11].um_I.ow[4] ;
 wire \top_I.branch[30].block[11].um_I.ow[5] ;
 wire \top_I.branch[30].block[11].um_I.ow[6] ;
 wire \top_I.branch[30].block[11].um_I.ow[7] ;
 wire \top_I.branch[30].block[11].um_I.ow[8] ;
 wire \top_I.branch[30].block[11].um_I.ow[9] ;
 wire \top_I.branch[30].block[11].um_I.pg_vdd ;
 wire \top_I.branch[30].block[12].um_I.ana[0] ;
 wire \top_I.branch[30].block[12].um_I.ana[1] ;
 wire \top_I.branch[30].block[12].um_I.ana[2] ;
 wire \top_I.branch[30].block[12].um_I.ana[3] ;
 wire \top_I.branch[30].block[12].um_I.ana[4] ;
 wire \top_I.branch[30].block[12].um_I.ana[5] ;
 wire \top_I.branch[30].block[12].um_I.ana[6] ;
 wire \top_I.branch[30].block[12].um_I.ana[7] ;
 wire \top_I.branch[30].block[12].um_I.clk ;
 wire \top_I.branch[30].block[12].um_I.ena ;
 wire \top_I.branch[30].block[12].um_I.iw[10] ;
 wire \top_I.branch[30].block[12].um_I.iw[11] ;
 wire \top_I.branch[30].block[12].um_I.iw[12] ;
 wire \top_I.branch[30].block[12].um_I.iw[13] ;
 wire \top_I.branch[30].block[12].um_I.iw[14] ;
 wire \top_I.branch[30].block[12].um_I.iw[15] ;
 wire \top_I.branch[30].block[12].um_I.iw[16] ;
 wire \top_I.branch[30].block[12].um_I.iw[17] ;
 wire \top_I.branch[30].block[12].um_I.iw[1] ;
 wire \top_I.branch[30].block[12].um_I.iw[2] ;
 wire \top_I.branch[30].block[12].um_I.iw[3] ;
 wire \top_I.branch[30].block[12].um_I.iw[4] ;
 wire \top_I.branch[30].block[12].um_I.iw[5] ;
 wire \top_I.branch[30].block[12].um_I.iw[6] ;
 wire \top_I.branch[30].block[12].um_I.iw[7] ;
 wire \top_I.branch[30].block[12].um_I.iw[8] ;
 wire \top_I.branch[30].block[12].um_I.iw[9] ;
 wire \top_I.branch[30].block[12].um_I.k_zero ;
 wire \top_I.branch[30].block[12].um_I.pg_vdd ;
 wire \top_I.branch[30].block[13].um_I.ana[0] ;
 wire \top_I.branch[30].block[13].um_I.ana[1] ;
 wire \top_I.branch[30].block[13].um_I.ana[2] ;
 wire \top_I.branch[30].block[13].um_I.ana[3] ;
 wire \top_I.branch[30].block[13].um_I.ana[4] ;
 wire \top_I.branch[30].block[13].um_I.ana[5] ;
 wire \top_I.branch[30].block[13].um_I.ana[6] ;
 wire \top_I.branch[30].block[13].um_I.ana[7] ;
 wire \top_I.branch[30].block[13].um_I.clk ;
 wire \top_I.branch[30].block[13].um_I.ena ;
 wire \top_I.branch[30].block[13].um_I.iw[10] ;
 wire \top_I.branch[30].block[13].um_I.iw[11] ;
 wire \top_I.branch[30].block[13].um_I.iw[12] ;
 wire \top_I.branch[30].block[13].um_I.iw[13] ;
 wire \top_I.branch[30].block[13].um_I.iw[14] ;
 wire \top_I.branch[30].block[13].um_I.iw[15] ;
 wire \top_I.branch[30].block[13].um_I.iw[16] ;
 wire \top_I.branch[30].block[13].um_I.iw[17] ;
 wire \top_I.branch[30].block[13].um_I.iw[1] ;
 wire \top_I.branch[30].block[13].um_I.iw[2] ;
 wire \top_I.branch[30].block[13].um_I.iw[3] ;
 wire \top_I.branch[30].block[13].um_I.iw[4] ;
 wire \top_I.branch[30].block[13].um_I.iw[5] ;
 wire \top_I.branch[30].block[13].um_I.iw[6] ;
 wire \top_I.branch[30].block[13].um_I.iw[7] ;
 wire \top_I.branch[30].block[13].um_I.iw[8] ;
 wire \top_I.branch[30].block[13].um_I.iw[9] ;
 wire \top_I.branch[30].block[13].um_I.k_zero ;
 wire \top_I.branch[30].block[13].um_I.ow[0] ;
 wire \top_I.branch[30].block[13].um_I.ow[10] ;
 wire \top_I.branch[30].block[13].um_I.ow[11] ;
 wire \top_I.branch[30].block[13].um_I.ow[12] ;
 wire \top_I.branch[30].block[13].um_I.ow[13] ;
 wire \top_I.branch[30].block[13].um_I.ow[14] ;
 wire \top_I.branch[30].block[13].um_I.ow[15] ;
 wire \top_I.branch[30].block[13].um_I.ow[16] ;
 wire \top_I.branch[30].block[13].um_I.ow[17] ;
 wire \top_I.branch[30].block[13].um_I.ow[18] ;
 wire \top_I.branch[30].block[13].um_I.ow[19] ;
 wire \top_I.branch[30].block[13].um_I.ow[1] ;
 wire \top_I.branch[30].block[13].um_I.ow[20] ;
 wire \top_I.branch[30].block[13].um_I.ow[21] ;
 wire \top_I.branch[30].block[13].um_I.ow[22] ;
 wire \top_I.branch[30].block[13].um_I.ow[23] ;
 wire \top_I.branch[30].block[13].um_I.ow[2] ;
 wire \top_I.branch[30].block[13].um_I.ow[3] ;
 wire \top_I.branch[30].block[13].um_I.ow[4] ;
 wire \top_I.branch[30].block[13].um_I.ow[5] ;
 wire \top_I.branch[30].block[13].um_I.ow[6] ;
 wire \top_I.branch[30].block[13].um_I.ow[7] ;
 wire \top_I.branch[30].block[13].um_I.ow[8] ;
 wire \top_I.branch[30].block[13].um_I.ow[9] ;
 wire \top_I.branch[30].block[13].um_I.pg_vdd ;
 wire \top_I.branch[30].block[14].um_I.ana[0] ;
 wire \top_I.branch[30].block[14].um_I.ana[1] ;
 wire \top_I.branch[30].block[14].um_I.ana[2] ;
 wire \top_I.branch[30].block[14].um_I.ana[3] ;
 wire \top_I.branch[30].block[14].um_I.ana[4] ;
 wire \top_I.branch[30].block[14].um_I.ana[5] ;
 wire \top_I.branch[30].block[14].um_I.ana[6] ;
 wire \top_I.branch[30].block[14].um_I.ana[7] ;
 wire \top_I.branch[30].block[14].um_I.clk ;
 wire \top_I.branch[30].block[14].um_I.ena ;
 wire \top_I.branch[30].block[14].um_I.iw[10] ;
 wire \top_I.branch[30].block[14].um_I.iw[11] ;
 wire \top_I.branch[30].block[14].um_I.iw[12] ;
 wire \top_I.branch[30].block[14].um_I.iw[13] ;
 wire \top_I.branch[30].block[14].um_I.iw[14] ;
 wire \top_I.branch[30].block[14].um_I.iw[15] ;
 wire \top_I.branch[30].block[14].um_I.iw[16] ;
 wire \top_I.branch[30].block[14].um_I.iw[17] ;
 wire \top_I.branch[30].block[14].um_I.iw[1] ;
 wire \top_I.branch[30].block[14].um_I.iw[2] ;
 wire \top_I.branch[30].block[14].um_I.iw[3] ;
 wire \top_I.branch[30].block[14].um_I.iw[4] ;
 wire \top_I.branch[30].block[14].um_I.iw[5] ;
 wire \top_I.branch[30].block[14].um_I.iw[6] ;
 wire \top_I.branch[30].block[14].um_I.iw[7] ;
 wire \top_I.branch[30].block[14].um_I.iw[8] ;
 wire \top_I.branch[30].block[14].um_I.iw[9] ;
 wire \top_I.branch[30].block[14].um_I.k_zero ;
 wire \top_I.branch[30].block[14].um_I.pg_vdd ;
 wire \top_I.branch[30].block[15].um_I.ana[0] ;
 wire \top_I.branch[30].block[15].um_I.ana[1] ;
 wire \top_I.branch[30].block[15].um_I.ana[2] ;
 wire \top_I.branch[30].block[15].um_I.ana[3] ;
 wire \top_I.branch[30].block[15].um_I.ana[4] ;
 wire \top_I.branch[30].block[15].um_I.ana[5] ;
 wire \top_I.branch[30].block[15].um_I.ana[6] ;
 wire \top_I.branch[30].block[15].um_I.ana[7] ;
 wire \top_I.branch[30].block[15].um_I.clk ;
 wire \top_I.branch[30].block[15].um_I.ena ;
 wire \top_I.branch[30].block[15].um_I.iw[10] ;
 wire \top_I.branch[30].block[15].um_I.iw[11] ;
 wire \top_I.branch[30].block[15].um_I.iw[12] ;
 wire \top_I.branch[30].block[15].um_I.iw[13] ;
 wire \top_I.branch[30].block[15].um_I.iw[14] ;
 wire \top_I.branch[30].block[15].um_I.iw[15] ;
 wire \top_I.branch[30].block[15].um_I.iw[16] ;
 wire \top_I.branch[30].block[15].um_I.iw[17] ;
 wire \top_I.branch[30].block[15].um_I.iw[1] ;
 wire \top_I.branch[30].block[15].um_I.iw[2] ;
 wire \top_I.branch[30].block[15].um_I.iw[3] ;
 wire \top_I.branch[30].block[15].um_I.iw[4] ;
 wire \top_I.branch[30].block[15].um_I.iw[5] ;
 wire \top_I.branch[30].block[15].um_I.iw[6] ;
 wire \top_I.branch[30].block[15].um_I.iw[7] ;
 wire \top_I.branch[30].block[15].um_I.iw[8] ;
 wire \top_I.branch[30].block[15].um_I.iw[9] ;
 wire \top_I.branch[30].block[15].um_I.k_zero ;
 wire \top_I.branch[30].block[15].um_I.ow[0] ;
 wire \top_I.branch[30].block[15].um_I.ow[10] ;
 wire \top_I.branch[30].block[15].um_I.ow[11] ;
 wire \top_I.branch[30].block[15].um_I.ow[12] ;
 wire \top_I.branch[30].block[15].um_I.ow[13] ;
 wire \top_I.branch[30].block[15].um_I.ow[14] ;
 wire \top_I.branch[30].block[15].um_I.ow[15] ;
 wire \top_I.branch[30].block[15].um_I.ow[16] ;
 wire \top_I.branch[30].block[15].um_I.ow[17] ;
 wire \top_I.branch[30].block[15].um_I.ow[18] ;
 wire \top_I.branch[30].block[15].um_I.ow[19] ;
 wire \top_I.branch[30].block[15].um_I.ow[1] ;
 wire \top_I.branch[30].block[15].um_I.ow[20] ;
 wire \top_I.branch[30].block[15].um_I.ow[21] ;
 wire \top_I.branch[30].block[15].um_I.ow[22] ;
 wire \top_I.branch[30].block[15].um_I.ow[23] ;
 wire \top_I.branch[30].block[15].um_I.ow[2] ;
 wire \top_I.branch[30].block[15].um_I.ow[3] ;
 wire \top_I.branch[30].block[15].um_I.ow[4] ;
 wire \top_I.branch[30].block[15].um_I.ow[5] ;
 wire \top_I.branch[30].block[15].um_I.ow[6] ;
 wire \top_I.branch[30].block[15].um_I.ow[7] ;
 wire \top_I.branch[30].block[15].um_I.ow[8] ;
 wire \top_I.branch[30].block[15].um_I.ow[9] ;
 wire \top_I.branch[30].block[15].um_I.pg_vdd ;
 wire \top_I.branch[30].block[1].um_I.ana[0] ;
 wire \top_I.branch[30].block[1].um_I.ana[1] ;
 wire \top_I.branch[30].block[1].um_I.ana[2] ;
 wire \top_I.branch[30].block[1].um_I.ana[3] ;
 wire \top_I.branch[30].block[1].um_I.ana[4] ;
 wire \top_I.branch[30].block[1].um_I.ana[5] ;
 wire \top_I.branch[30].block[1].um_I.ana[6] ;
 wire \top_I.branch[30].block[1].um_I.ana[7] ;
 wire \top_I.branch[30].block[1].um_I.clk ;
 wire \top_I.branch[30].block[1].um_I.ena ;
 wire \top_I.branch[30].block[1].um_I.iw[10] ;
 wire \top_I.branch[30].block[1].um_I.iw[11] ;
 wire \top_I.branch[30].block[1].um_I.iw[12] ;
 wire \top_I.branch[30].block[1].um_I.iw[13] ;
 wire \top_I.branch[30].block[1].um_I.iw[14] ;
 wire \top_I.branch[30].block[1].um_I.iw[15] ;
 wire \top_I.branch[30].block[1].um_I.iw[16] ;
 wire \top_I.branch[30].block[1].um_I.iw[17] ;
 wire \top_I.branch[30].block[1].um_I.iw[1] ;
 wire \top_I.branch[30].block[1].um_I.iw[2] ;
 wire \top_I.branch[30].block[1].um_I.iw[3] ;
 wire \top_I.branch[30].block[1].um_I.iw[4] ;
 wire \top_I.branch[30].block[1].um_I.iw[5] ;
 wire \top_I.branch[30].block[1].um_I.iw[6] ;
 wire \top_I.branch[30].block[1].um_I.iw[7] ;
 wire \top_I.branch[30].block[1].um_I.iw[8] ;
 wire \top_I.branch[30].block[1].um_I.iw[9] ;
 wire \top_I.branch[30].block[1].um_I.k_zero ;
 wire \top_I.branch[30].block[1].um_I.ow[0] ;
 wire \top_I.branch[30].block[1].um_I.ow[10] ;
 wire \top_I.branch[30].block[1].um_I.ow[11] ;
 wire \top_I.branch[30].block[1].um_I.ow[12] ;
 wire \top_I.branch[30].block[1].um_I.ow[13] ;
 wire \top_I.branch[30].block[1].um_I.ow[14] ;
 wire \top_I.branch[30].block[1].um_I.ow[15] ;
 wire \top_I.branch[30].block[1].um_I.ow[16] ;
 wire \top_I.branch[30].block[1].um_I.ow[17] ;
 wire \top_I.branch[30].block[1].um_I.ow[18] ;
 wire \top_I.branch[30].block[1].um_I.ow[19] ;
 wire \top_I.branch[30].block[1].um_I.ow[1] ;
 wire \top_I.branch[30].block[1].um_I.ow[20] ;
 wire \top_I.branch[30].block[1].um_I.ow[21] ;
 wire \top_I.branch[30].block[1].um_I.ow[22] ;
 wire \top_I.branch[30].block[1].um_I.ow[23] ;
 wire \top_I.branch[30].block[1].um_I.ow[2] ;
 wire \top_I.branch[30].block[1].um_I.ow[3] ;
 wire \top_I.branch[30].block[1].um_I.ow[4] ;
 wire \top_I.branch[30].block[1].um_I.ow[5] ;
 wire \top_I.branch[30].block[1].um_I.ow[6] ;
 wire \top_I.branch[30].block[1].um_I.ow[7] ;
 wire \top_I.branch[30].block[1].um_I.ow[8] ;
 wire \top_I.branch[30].block[1].um_I.ow[9] ;
 wire \top_I.branch[30].block[1].um_I.pg_vdd ;
 wire \top_I.branch[30].block[2].um_I.ana[0] ;
 wire \top_I.branch[30].block[2].um_I.ana[1] ;
 wire \top_I.branch[30].block[2].um_I.ana[2] ;
 wire \top_I.branch[30].block[2].um_I.ana[3] ;
 wire \top_I.branch[30].block[2].um_I.ana[4] ;
 wire \top_I.branch[30].block[2].um_I.ana[5] ;
 wire \top_I.branch[30].block[2].um_I.ana[6] ;
 wire \top_I.branch[30].block[2].um_I.ana[7] ;
 wire \top_I.branch[30].block[2].um_I.clk ;
 wire \top_I.branch[30].block[2].um_I.ena ;
 wire \top_I.branch[30].block[2].um_I.iw[10] ;
 wire \top_I.branch[30].block[2].um_I.iw[11] ;
 wire \top_I.branch[30].block[2].um_I.iw[12] ;
 wire \top_I.branch[30].block[2].um_I.iw[13] ;
 wire \top_I.branch[30].block[2].um_I.iw[14] ;
 wire \top_I.branch[30].block[2].um_I.iw[15] ;
 wire \top_I.branch[30].block[2].um_I.iw[16] ;
 wire \top_I.branch[30].block[2].um_I.iw[17] ;
 wire \top_I.branch[30].block[2].um_I.iw[1] ;
 wire \top_I.branch[30].block[2].um_I.iw[2] ;
 wire \top_I.branch[30].block[2].um_I.iw[3] ;
 wire \top_I.branch[30].block[2].um_I.iw[4] ;
 wire \top_I.branch[30].block[2].um_I.iw[5] ;
 wire \top_I.branch[30].block[2].um_I.iw[6] ;
 wire \top_I.branch[30].block[2].um_I.iw[7] ;
 wire \top_I.branch[30].block[2].um_I.iw[8] ;
 wire \top_I.branch[30].block[2].um_I.iw[9] ;
 wire \top_I.branch[30].block[2].um_I.k_zero ;
 wire \top_I.branch[30].block[2].um_I.ow[0] ;
 wire \top_I.branch[30].block[2].um_I.ow[10] ;
 wire \top_I.branch[30].block[2].um_I.ow[11] ;
 wire \top_I.branch[30].block[2].um_I.ow[12] ;
 wire \top_I.branch[30].block[2].um_I.ow[13] ;
 wire \top_I.branch[30].block[2].um_I.ow[14] ;
 wire \top_I.branch[30].block[2].um_I.ow[15] ;
 wire \top_I.branch[30].block[2].um_I.ow[16] ;
 wire \top_I.branch[30].block[2].um_I.ow[17] ;
 wire \top_I.branch[30].block[2].um_I.ow[18] ;
 wire \top_I.branch[30].block[2].um_I.ow[19] ;
 wire \top_I.branch[30].block[2].um_I.ow[1] ;
 wire \top_I.branch[30].block[2].um_I.ow[20] ;
 wire \top_I.branch[30].block[2].um_I.ow[21] ;
 wire \top_I.branch[30].block[2].um_I.ow[22] ;
 wire \top_I.branch[30].block[2].um_I.ow[23] ;
 wire \top_I.branch[30].block[2].um_I.ow[2] ;
 wire \top_I.branch[30].block[2].um_I.ow[3] ;
 wire \top_I.branch[30].block[2].um_I.ow[4] ;
 wire \top_I.branch[30].block[2].um_I.ow[5] ;
 wire \top_I.branch[30].block[2].um_I.ow[6] ;
 wire \top_I.branch[30].block[2].um_I.ow[7] ;
 wire \top_I.branch[30].block[2].um_I.ow[8] ;
 wire \top_I.branch[30].block[2].um_I.ow[9] ;
 wire \top_I.branch[30].block[2].um_I.pg_vdd ;
 wire \top_I.branch[30].block[3].um_I.ana[0] ;
 wire \top_I.branch[30].block[3].um_I.ana[1] ;
 wire \top_I.branch[30].block[3].um_I.ana[2] ;
 wire \top_I.branch[30].block[3].um_I.ana[3] ;
 wire \top_I.branch[30].block[3].um_I.ana[4] ;
 wire \top_I.branch[30].block[3].um_I.ana[5] ;
 wire \top_I.branch[30].block[3].um_I.ana[6] ;
 wire \top_I.branch[30].block[3].um_I.ana[7] ;
 wire \top_I.branch[30].block[3].um_I.clk ;
 wire \top_I.branch[30].block[3].um_I.ena ;
 wire \top_I.branch[30].block[3].um_I.iw[10] ;
 wire \top_I.branch[30].block[3].um_I.iw[11] ;
 wire \top_I.branch[30].block[3].um_I.iw[12] ;
 wire \top_I.branch[30].block[3].um_I.iw[13] ;
 wire \top_I.branch[30].block[3].um_I.iw[14] ;
 wire \top_I.branch[30].block[3].um_I.iw[15] ;
 wire \top_I.branch[30].block[3].um_I.iw[16] ;
 wire \top_I.branch[30].block[3].um_I.iw[17] ;
 wire \top_I.branch[30].block[3].um_I.iw[1] ;
 wire \top_I.branch[30].block[3].um_I.iw[2] ;
 wire \top_I.branch[30].block[3].um_I.iw[3] ;
 wire \top_I.branch[30].block[3].um_I.iw[4] ;
 wire \top_I.branch[30].block[3].um_I.iw[5] ;
 wire \top_I.branch[30].block[3].um_I.iw[6] ;
 wire \top_I.branch[30].block[3].um_I.iw[7] ;
 wire \top_I.branch[30].block[3].um_I.iw[8] ;
 wire \top_I.branch[30].block[3].um_I.iw[9] ;
 wire \top_I.branch[30].block[3].um_I.k_zero ;
 wire \top_I.branch[30].block[3].um_I.ow[0] ;
 wire \top_I.branch[30].block[3].um_I.ow[10] ;
 wire \top_I.branch[30].block[3].um_I.ow[11] ;
 wire \top_I.branch[30].block[3].um_I.ow[12] ;
 wire \top_I.branch[30].block[3].um_I.ow[13] ;
 wire \top_I.branch[30].block[3].um_I.ow[14] ;
 wire \top_I.branch[30].block[3].um_I.ow[15] ;
 wire \top_I.branch[30].block[3].um_I.ow[16] ;
 wire \top_I.branch[30].block[3].um_I.ow[17] ;
 wire \top_I.branch[30].block[3].um_I.ow[18] ;
 wire \top_I.branch[30].block[3].um_I.ow[19] ;
 wire \top_I.branch[30].block[3].um_I.ow[1] ;
 wire \top_I.branch[30].block[3].um_I.ow[20] ;
 wire \top_I.branch[30].block[3].um_I.ow[21] ;
 wire \top_I.branch[30].block[3].um_I.ow[22] ;
 wire \top_I.branch[30].block[3].um_I.ow[23] ;
 wire \top_I.branch[30].block[3].um_I.ow[2] ;
 wire \top_I.branch[30].block[3].um_I.ow[3] ;
 wire \top_I.branch[30].block[3].um_I.ow[4] ;
 wire \top_I.branch[30].block[3].um_I.ow[5] ;
 wire \top_I.branch[30].block[3].um_I.ow[6] ;
 wire \top_I.branch[30].block[3].um_I.ow[7] ;
 wire \top_I.branch[30].block[3].um_I.ow[8] ;
 wire \top_I.branch[30].block[3].um_I.ow[9] ;
 wire \top_I.branch[30].block[3].um_I.pg_vdd ;
 wire \top_I.branch[30].block[4].um_I.ana[0] ;
 wire \top_I.branch[30].block[4].um_I.ana[1] ;
 wire \top_I.branch[30].block[4].um_I.ana[2] ;
 wire \top_I.branch[30].block[4].um_I.ana[3] ;
 wire \top_I.branch[30].block[4].um_I.ana[4] ;
 wire \top_I.branch[30].block[4].um_I.ana[5] ;
 wire \top_I.branch[30].block[4].um_I.ana[6] ;
 wire \top_I.branch[30].block[4].um_I.ana[7] ;
 wire \top_I.branch[30].block[4].um_I.clk ;
 wire \top_I.branch[30].block[4].um_I.ena ;
 wire \top_I.branch[30].block[4].um_I.iw[10] ;
 wire \top_I.branch[30].block[4].um_I.iw[11] ;
 wire \top_I.branch[30].block[4].um_I.iw[12] ;
 wire \top_I.branch[30].block[4].um_I.iw[13] ;
 wire \top_I.branch[30].block[4].um_I.iw[14] ;
 wire \top_I.branch[30].block[4].um_I.iw[15] ;
 wire \top_I.branch[30].block[4].um_I.iw[16] ;
 wire \top_I.branch[30].block[4].um_I.iw[17] ;
 wire \top_I.branch[30].block[4].um_I.iw[1] ;
 wire \top_I.branch[30].block[4].um_I.iw[2] ;
 wire \top_I.branch[30].block[4].um_I.iw[3] ;
 wire \top_I.branch[30].block[4].um_I.iw[4] ;
 wire \top_I.branch[30].block[4].um_I.iw[5] ;
 wire \top_I.branch[30].block[4].um_I.iw[6] ;
 wire \top_I.branch[30].block[4].um_I.iw[7] ;
 wire \top_I.branch[30].block[4].um_I.iw[8] ;
 wire \top_I.branch[30].block[4].um_I.iw[9] ;
 wire \top_I.branch[30].block[4].um_I.k_zero ;
 wire \top_I.branch[30].block[4].um_I.ow[0] ;
 wire \top_I.branch[30].block[4].um_I.ow[10] ;
 wire \top_I.branch[30].block[4].um_I.ow[11] ;
 wire \top_I.branch[30].block[4].um_I.ow[12] ;
 wire \top_I.branch[30].block[4].um_I.ow[13] ;
 wire \top_I.branch[30].block[4].um_I.ow[14] ;
 wire \top_I.branch[30].block[4].um_I.ow[15] ;
 wire \top_I.branch[30].block[4].um_I.ow[16] ;
 wire \top_I.branch[30].block[4].um_I.ow[17] ;
 wire \top_I.branch[30].block[4].um_I.ow[18] ;
 wire \top_I.branch[30].block[4].um_I.ow[19] ;
 wire \top_I.branch[30].block[4].um_I.ow[1] ;
 wire \top_I.branch[30].block[4].um_I.ow[20] ;
 wire \top_I.branch[30].block[4].um_I.ow[21] ;
 wire \top_I.branch[30].block[4].um_I.ow[22] ;
 wire \top_I.branch[30].block[4].um_I.ow[23] ;
 wire \top_I.branch[30].block[4].um_I.ow[2] ;
 wire \top_I.branch[30].block[4].um_I.ow[3] ;
 wire \top_I.branch[30].block[4].um_I.ow[4] ;
 wire \top_I.branch[30].block[4].um_I.ow[5] ;
 wire \top_I.branch[30].block[4].um_I.ow[6] ;
 wire \top_I.branch[30].block[4].um_I.ow[7] ;
 wire \top_I.branch[30].block[4].um_I.ow[8] ;
 wire \top_I.branch[30].block[4].um_I.ow[9] ;
 wire \top_I.branch[30].block[4].um_I.pg_vdd ;
 wire \top_I.branch[30].block[5].um_I.ana[0] ;
 wire \top_I.branch[30].block[5].um_I.ana[1] ;
 wire \top_I.branch[30].block[5].um_I.ana[2] ;
 wire \top_I.branch[30].block[5].um_I.ana[3] ;
 wire \top_I.branch[30].block[5].um_I.ana[4] ;
 wire \top_I.branch[30].block[5].um_I.ana[5] ;
 wire \top_I.branch[30].block[5].um_I.ana[6] ;
 wire \top_I.branch[30].block[5].um_I.ana[7] ;
 wire \top_I.branch[30].block[5].um_I.clk ;
 wire \top_I.branch[30].block[5].um_I.ena ;
 wire \top_I.branch[30].block[5].um_I.iw[10] ;
 wire \top_I.branch[30].block[5].um_I.iw[11] ;
 wire \top_I.branch[30].block[5].um_I.iw[12] ;
 wire \top_I.branch[30].block[5].um_I.iw[13] ;
 wire \top_I.branch[30].block[5].um_I.iw[14] ;
 wire \top_I.branch[30].block[5].um_I.iw[15] ;
 wire \top_I.branch[30].block[5].um_I.iw[16] ;
 wire \top_I.branch[30].block[5].um_I.iw[17] ;
 wire \top_I.branch[30].block[5].um_I.iw[1] ;
 wire \top_I.branch[30].block[5].um_I.iw[2] ;
 wire \top_I.branch[30].block[5].um_I.iw[3] ;
 wire \top_I.branch[30].block[5].um_I.iw[4] ;
 wire \top_I.branch[30].block[5].um_I.iw[5] ;
 wire \top_I.branch[30].block[5].um_I.iw[6] ;
 wire \top_I.branch[30].block[5].um_I.iw[7] ;
 wire \top_I.branch[30].block[5].um_I.iw[8] ;
 wire \top_I.branch[30].block[5].um_I.iw[9] ;
 wire \top_I.branch[30].block[5].um_I.k_zero ;
 wire \top_I.branch[30].block[5].um_I.ow[0] ;
 wire \top_I.branch[30].block[5].um_I.ow[10] ;
 wire \top_I.branch[30].block[5].um_I.ow[11] ;
 wire \top_I.branch[30].block[5].um_I.ow[12] ;
 wire \top_I.branch[30].block[5].um_I.ow[13] ;
 wire \top_I.branch[30].block[5].um_I.ow[14] ;
 wire \top_I.branch[30].block[5].um_I.ow[15] ;
 wire \top_I.branch[30].block[5].um_I.ow[16] ;
 wire \top_I.branch[30].block[5].um_I.ow[17] ;
 wire \top_I.branch[30].block[5].um_I.ow[18] ;
 wire \top_I.branch[30].block[5].um_I.ow[19] ;
 wire \top_I.branch[30].block[5].um_I.ow[1] ;
 wire \top_I.branch[30].block[5].um_I.ow[20] ;
 wire \top_I.branch[30].block[5].um_I.ow[21] ;
 wire \top_I.branch[30].block[5].um_I.ow[22] ;
 wire \top_I.branch[30].block[5].um_I.ow[23] ;
 wire \top_I.branch[30].block[5].um_I.ow[2] ;
 wire \top_I.branch[30].block[5].um_I.ow[3] ;
 wire \top_I.branch[30].block[5].um_I.ow[4] ;
 wire \top_I.branch[30].block[5].um_I.ow[5] ;
 wire \top_I.branch[30].block[5].um_I.ow[6] ;
 wire \top_I.branch[30].block[5].um_I.ow[7] ;
 wire \top_I.branch[30].block[5].um_I.ow[8] ;
 wire \top_I.branch[30].block[5].um_I.ow[9] ;
 wire \top_I.branch[30].block[5].um_I.pg_vdd ;
 wire \top_I.branch[30].block[6].um_I.ana[0] ;
 wire \top_I.branch[30].block[6].um_I.ana[1] ;
 wire \top_I.branch[30].block[6].um_I.ana[2] ;
 wire \top_I.branch[30].block[6].um_I.ana[3] ;
 wire \top_I.branch[30].block[6].um_I.ana[4] ;
 wire \top_I.branch[30].block[6].um_I.ana[5] ;
 wire \top_I.branch[30].block[6].um_I.ana[6] ;
 wire \top_I.branch[30].block[6].um_I.ana[7] ;
 wire \top_I.branch[30].block[6].um_I.clk ;
 wire \top_I.branch[30].block[6].um_I.ena ;
 wire \top_I.branch[30].block[6].um_I.iw[10] ;
 wire \top_I.branch[30].block[6].um_I.iw[11] ;
 wire \top_I.branch[30].block[6].um_I.iw[12] ;
 wire \top_I.branch[30].block[6].um_I.iw[13] ;
 wire \top_I.branch[30].block[6].um_I.iw[14] ;
 wire \top_I.branch[30].block[6].um_I.iw[15] ;
 wire \top_I.branch[30].block[6].um_I.iw[16] ;
 wire \top_I.branch[30].block[6].um_I.iw[17] ;
 wire \top_I.branch[30].block[6].um_I.iw[1] ;
 wire \top_I.branch[30].block[6].um_I.iw[2] ;
 wire \top_I.branch[30].block[6].um_I.iw[3] ;
 wire \top_I.branch[30].block[6].um_I.iw[4] ;
 wire \top_I.branch[30].block[6].um_I.iw[5] ;
 wire \top_I.branch[30].block[6].um_I.iw[6] ;
 wire \top_I.branch[30].block[6].um_I.iw[7] ;
 wire \top_I.branch[30].block[6].um_I.iw[8] ;
 wire \top_I.branch[30].block[6].um_I.iw[9] ;
 wire \top_I.branch[30].block[6].um_I.k_zero ;
 wire \top_I.branch[30].block[6].um_I.ow[0] ;
 wire \top_I.branch[30].block[6].um_I.ow[10] ;
 wire \top_I.branch[30].block[6].um_I.ow[11] ;
 wire \top_I.branch[30].block[6].um_I.ow[12] ;
 wire \top_I.branch[30].block[6].um_I.ow[13] ;
 wire \top_I.branch[30].block[6].um_I.ow[14] ;
 wire \top_I.branch[30].block[6].um_I.ow[15] ;
 wire \top_I.branch[30].block[6].um_I.ow[16] ;
 wire \top_I.branch[30].block[6].um_I.ow[17] ;
 wire \top_I.branch[30].block[6].um_I.ow[18] ;
 wire \top_I.branch[30].block[6].um_I.ow[19] ;
 wire \top_I.branch[30].block[6].um_I.ow[1] ;
 wire \top_I.branch[30].block[6].um_I.ow[20] ;
 wire \top_I.branch[30].block[6].um_I.ow[21] ;
 wire \top_I.branch[30].block[6].um_I.ow[22] ;
 wire \top_I.branch[30].block[6].um_I.ow[23] ;
 wire \top_I.branch[30].block[6].um_I.ow[2] ;
 wire \top_I.branch[30].block[6].um_I.ow[3] ;
 wire \top_I.branch[30].block[6].um_I.ow[4] ;
 wire \top_I.branch[30].block[6].um_I.ow[5] ;
 wire \top_I.branch[30].block[6].um_I.ow[6] ;
 wire \top_I.branch[30].block[6].um_I.ow[7] ;
 wire \top_I.branch[30].block[6].um_I.ow[8] ;
 wire \top_I.branch[30].block[6].um_I.ow[9] ;
 wire \top_I.branch[30].block[6].um_I.pg_vdd ;
 wire \top_I.branch[30].block[7].um_I.ana[0] ;
 wire \top_I.branch[30].block[7].um_I.ana[1] ;
 wire \top_I.branch[30].block[7].um_I.ana[2] ;
 wire \top_I.branch[30].block[7].um_I.ana[3] ;
 wire \top_I.branch[30].block[7].um_I.ana[4] ;
 wire \top_I.branch[30].block[7].um_I.ana[5] ;
 wire \top_I.branch[30].block[7].um_I.ana[6] ;
 wire \top_I.branch[30].block[7].um_I.ana[7] ;
 wire \top_I.branch[30].block[7].um_I.clk ;
 wire \top_I.branch[30].block[7].um_I.ena ;
 wire \top_I.branch[30].block[7].um_I.iw[10] ;
 wire \top_I.branch[30].block[7].um_I.iw[11] ;
 wire \top_I.branch[30].block[7].um_I.iw[12] ;
 wire \top_I.branch[30].block[7].um_I.iw[13] ;
 wire \top_I.branch[30].block[7].um_I.iw[14] ;
 wire \top_I.branch[30].block[7].um_I.iw[15] ;
 wire \top_I.branch[30].block[7].um_I.iw[16] ;
 wire \top_I.branch[30].block[7].um_I.iw[17] ;
 wire \top_I.branch[30].block[7].um_I.iw[1] ;
 wire \top_I.branch[30].block[7].um_I.iw[2] ;
 wire \top_I.branch[30].block[7].um_I.iw[3] ;
 wire \top_I.branch[30].block[7].um_I.iw[4] ;
 wire \top_I.branch[30].block[7].um_I.iw[5] ;
 wire \top_I.branch[30].block[7].um_I.iw[6] ;
 wire \top_I.branch[30].block[7].um_I.iw[7] ;
 wire \top_I.branch[30].block[7].um_I.iw[8] ;
 wire \top_I.branch[30].block[7].um_I.iw[9] ;
 wire \top_I.branch[30].block[7].um_I.k_zero ;
 wire \top_I.branch[30].block[7].um_I.ow[0] ;
 wire \top_I.branch[30].block[7].um_I.ow[10] ;
 wire \top_I.branch[30].block[7].um_I.ow[11] ;
 wire \top_I.branch[30].block[7].um_I.ow[12] ;
 wire \top_I.branch[30].block[7].um_I.ow[13] ;
 wire \top_I.branch[30].block[7].um_I.ow[14] ;
 wire \top_I.branch[30].block[7].um_I.ow[15] ;
 wire \top_I.branch[30].block[7].um_I.ow[16] ;
 wire \top_I.branch[30].block[7].um_I.ow[17] ;
 wire \top_I.branch[30].block[7].um_I.ow[18] ;
 wire \top_I.branch[30].block[7].um_I.ow[19] ;
 wire \top_I.branch[30].block[7].um_I.ow[1] ;
 wire \top_I.branch[30].block[7].um_I.ow[20] ;
 wire \top_I.branch[30].block[7].um_I.ow[21] ;
 wire \top_I.branch[30].block[7].um_I.ow[22] ;
 wire \top_I.branch[30].block[7].um_I.ow[23] ;
 wire \top_I.branch[30].block[7].um_I.ow[2] ;
 wire \top_I.branch[30].block[7].um_I.ow[3] ;
 wire \top_I.branch[30].block[7].um_I.ow[4] ;
 wire \top_I.branch[30].block[7].um_I.ow[5] ;
 wire \top_I.branch[30].block[7].um_I.ow[6] ;
 wire \top_I.branch[30].block[7].um_I.ow[7] ;
 wire \top_I.branch[30].block[7].um_I.ow[8] ;
 wire \top_I.branch[30].block[7].um_I.ow[9] ;
 wire \top_I.branch[30].block[7].um_I.pg_vdd ;
 wire \top_I.branch[30].block[8].um_I.ana[0] ;
 wire \top_I.branch[30].block[8].um_I.ana[1] ;
 wire \top_I.branch[30].block[8].um_I.ana[2] ;
 wire \top_I.branch[30].block[8].um_I.ana[3] ;
 wire \top_I.branch[30].block[8].um_I.ana[4] ;
 wire \top_I.branch[30].block[8].um_I.ana[5] ;
 wire \top_I.branch[30].block[8].um_I.ana[6] ;
 wire \top_I.branch[30].block[8].um_I.ana[7] ;
 wire \top_I.branch[30].block[8].um_I.clk ;
 wire \top_I.branch[30].block[8].um_I.ena ;
 wire \top_I.branch[30].block[8].um_I.iw[10] ;
 wire \top_I.branch[30].block[8].um_I.iw[11] ;
 wire \top_I.branch[30].block[8].um_I.iw[12] ;
 wire \top_I.branch[30].block[8].um_I.iw[13] ;
 wire \top_I.branch[30].block[8].um_I.iw[14] ;
 wire \top_I.branch[30].block[8].um_I.iw[15] ;
 wire \top_I.branch[30].block[8].um_I.iw[16] ;
 wire \top_I.branch[30].block[8].um_I.iw[17] ;
 wire \top_I.branch[30].block[8].um_I.iw[1] ;
 wire \top_I.branch[30].block[8].um_I.iw[2] ;
 wire \top_I.branch[30].block[8].um_I.iw[3] ;
 wire \top_I.branch[30].block[8].um_I.iw[4] ;
 wire \top_I.branch[30].block[8].um_I.iw[5] ;
 wire \top_I.branch[30].block[8].um_I.iw[6] ;
 wire \top_I.branch[30].block[8].um_I.iw[7] ;
 wire \top_I.branch[30].block[8].um_I.iw[8] ;
 wire \top_I.branch[30].block[8].um_I.iw[9] ;
 wire \top_I.branch[30].block[8].um_I.k_zero ;
 wire \top_I.branch[30].block[8].um_I.ow[0] ;
 wire \top_I.branch[30].block[8].um_I.ow[10] ;
 wire \top_I.branch[30].block[8].um_I.ow[11] ;
 wire \top_I.branch[30].block[8].um_I.ow[12] ;
 wire \top_I.branch[30].block[8].um_I.ow[13] ;
 wire \top_I.branch[30].block[8].um_I.ow[14] ;
 wire \top_I.branch[30].block[8].um_I.ow[15] ;
 wire \top_I.branch[30].block[8].um_I.ow[16] ;
 wire \top_I.branch[30].block[8].um_I.ow[17] ;
 wire \top_I.branch[30].block[8].um_I.ow[18] ;
 wire \top_I.branch[30].block[8].um_I.ow[19] ;
 wire \top_I.branch[30].block[8].um_I.ow[1] ;
 wire \top_I.branch[30].block[8].um_I.ow[20] ;
 wire \top_I.branch[30].block[8].um_I.ow[21] ;
 wire \top_I.branch[30].block[8].um_I.ow[22] ;
 wire \top_I.branch[30].block[8].um_I.ow[23] ;
 wire \top_I.branch[30].block[8].um_I.ow[2] ;
 wire \top_I.branch[30].block[8].um_I.ow[3] ;
 wire \top_I.branch[30].block[8].um_I.ow[4] ;
 wire \top_I.branch[30].block[8].um_I.ow[5] ;
 wire \top_I.branch[30].block[8].um_I.ow[6] ;
 wire \top_I.branch[30].block[8].um_I.ow[7] ;
 wire \top_I.branch[30].block[8].um_I.ow[8] ;
 wire \top_I.branch[30].block[8].um_I.ow[9] ;
 wire \top_I.branch[30].block[8].um_I.pg_vdd ;
 wire \top_I.branch[30].block[9].um_I.ana[0] ;
 wire \top_I.branch[30].block[9].um_I.ana[1] ;
 wire \top_I.branch[30].block[9].um_I.ana[2] ;
 wire \top_I.branch[30].block[9].um_I.ana[3] ;
 wire \top_I.branch[30].block[9].um_I.ana[4] ;
 wire \top_I.branch[30].block[9].um_I.ana[5] ;
 wire \top_I.branch[30].block[9].um_I.ana[6] ;
 wire \top_I.branch[30].block[9].um_I.ana[7] ;
 wire \top_I.branch[30].block[9].um_I.clk ;
 wire \top_I.branch[30].block[9].um_I.ena ;
 wire \top_I.branch[30].block[9].um_I.iw[10] ;
 wire \top_I.branch[30].block[9].um_I.iw[11] ;
 wire \top_I.branch[30].block[9].um_I.iw[12] ;
 wire \top_I.branch[30].block[9].um_I.iw[13] ;
 wire \top_I.branch[30].block[9].um_I.iw[14] ;
 wire \top_I.branch[30].block[9].um_I.iw[15] ;
 wire \top_I.branch[30].block[9].um_I.iw[16] ;
 wire \top_I.branch[30].block[9].um_I.iw[17] ;
 wire \top_I.branch[30].block[9].um_I.iw[1] ;
 wire \top_I.branch[30].block[9].um_I.iw[2] ;
 wire \top_I.branch[30].block[9].um_I.iw[3] ;
 wire \top_I.branch[30].block[9].um_I.iw[4] ;
 wire \top_I.branch[30].block[9].um_I.iw[5] ;
 wire \top_I.branch[30].block[9].um_I.iw[6] ;
 wire \top_I.branch[30].block[9].um_I.iw[7] ;
 wire \top_I.branch[30].block[9].um_I.iw[8] ;
 wire \top_I.branch[30].block[9].um_I.iw[9] ;
 wire \top_I.branch[30].block[9].um_I.k_zero ;
 wire \top_I.branch[30].block[9].um_I.ow[0] ;
 wire \top_I.branch[30].block[9].um_I.ow[10] ;
 wire \top_I.branch[30].block[9].um_I.ow[11] ;
 wire \top_I.branch[30].block[9].um_I.ow[12] ;
 wire \top_I.branch[30].block[9].um_I.ow[13] ;
 wire \top_I.branch[30].block[9].um_I.ow[14] ;
 wire \top_I.branch[30].block[9].um_I.ow[15] ;
 wire \top_I.branch[30].block[9].um_I.ow[16] ;
 wire \top_I.branch[30].block[9].um_I.ow[17] ;
 wire \top_I.branch[30].block[9].um_I.ow[18] ;
 wire \top_I.branch[30].block[9].um_I.ow[19] ;
 wire \top_I.branch[30].block[9].um_I.ow[1] ;
 wire \top_I.branch[30].block[9].um_I.ow[20] ;
 wire \top_I.branch[30].block[9].um_I.ow[21] ;
 wire \top_I.branch[30].block[9].um_I.ow[22] ;
 wire \top_I.branch[30].block[9].um_I.ow[23] ;
 wire \top_I.branch[30].block[9].um_I.ow[2] ;
 wire \top_I.branch[30].block[9].um_I.ow[3] ;
 wire \top_I.branch[30].block[9].um_I.ow[4] ;
 wire \top_I.branch[30].block[9].um_I.ow[5] ;
 wire \top_I.branch[30].block[9].um_I.ow[6] ;
 wire \top_I.branch[30].block[9].um_I.ow[7] ;
 wire \top_I.branch[30].block[9].um_I.ow[8] ;
 wire \top_I.branch[30].block[9].um_I.ow[9] ;
 wire \top_I.branch[30].block[9].um_I.pg_vdd ;
 wire \top_I.branch[30].l_addr[0] ;
 wire \top_I.branch[30].l_k_zero ;
 wire \top_I.branch[31].block[0].um_I.ana[0] ;
 wire \top_I.branch[31].block[0].um_I.ana[1] ;
 wire \top_I.branch[31].block[0].um_I.ana[2] ;
 wire \top_I.branch[31].block[0].um_I.ana[3] ;
 wire \top_I.branch[31].block[0].um_I.ana[4] ;
 wire \top_I.branch[31].block[0].um_I.ana[5] ;
 wire \top_I.branch[31].block[0].um_I.ana[6] ;
 wire \top_I.branch[31].block[0].um_I.ana[7] ;
 wire \top_I.branch[31].block[0].um_I.clk ;
 wire \top_I.branch[31].block[0].um_I.ena ;
 wire \top_I.branch[31].block[0].um_I.iw[10] ;
 wire \top_I.branch[31].block[0].um_I.iw[11] ;
 wire \top_I.branch[31].block[0].um_I.iw[12] ;
 wire \top_I.branch[31].block[0].um_I.iw[13] ;
 wire \top_I.branch[31].block[0].um_I.iw[14] ;
 wire \top_I.branch[31].block[0].um_I.iw[15] ;
 wire \top_I.branch[31].block[0].um_I.iw[16] ;
 wire \top_I.branch[31].block[0].um_I.iw[17] ;
 wire \top_I.branch[31].block[0].um_I.iw[1] ;
 wire \top_I.branch[31].block[0].um_I.iw[2] ;
 wire \top_I.branch[31].block[0].um_I.iw[3] ;
 wire \top_I.branch[31].block[0].um_I.iw[4] ;
 wire \top_I.branch[31].block[0].um_I.iw[5] ;
 wire \top_I.branch[31].block[0].um_I.iw[6] ;
 wire \top_I.branch[31].block[0].um_I.iw[7] ;
 wire \top_I.branch[31].block[0].um_I.iw[8] ;
 wire \top_I.branch[31].block[0].um_I.iw[9] ;
 wire \top_I.branch[31].block[0].um_I.k_zero ;
 wire \top_I.branch[31].block[0].um_I.pg_vdd ;
 wire \top_I.branch[31].block[10].um_I.ana[0] ;
 wire \top_I.branch[31].block[10].um_I.ana[1] ;
 wire \top_I.branch[31].block[10].um_I.ana[2] ;
 wire \top_I.branch[31].block[10].um_I.ana[3] ;
 wire \top_I.branch[31].block[10].um_I.ana[4] ;
 wire \top_I.branch[31].block[10].um_I.ana[5] ;
 wire \top_I.branch[31].block[10].um_I.ana[6] ;
 wire \top_I.branch[31].block[10].um_I.ana[7] ;
 wire \top_I.branch[31].block[10].um_I.clk ;
 wire \top_I.branch[31].block[10].um_I.ena ;
 wire \top_I.branch[31].block[10].um_I.iw[10] ;
 wire \top_I.branch[31].block[10].um_I.iw[11] ;
 wire \top_I.branch[31].block[10].um_I.iw[12] ;
 wire \top_I.branch[31].block[10].um_I.iw[13] ;
 wire \top_I.branch[31].block[10].um_I.iw[14] ;
 wire \top_I.branch[31].block[10].um_I.iw[15] ;
 wire \top_I.branch[31].block[10].um_I.iw[16] ;
 wire \top_I.branch[31].block[10].um_I.iw[17] ;
 wire \top_I.branch[31].block[10].um_I.iw[1] ;
 wire \top_I.branch[31].block[10].um_I.iw[2] ;
 wire \top_I.branch[31].block[10].um_I.iw[3] ;
 wire \top_I.branch[31].block[10].um_I.iw[4] ;
 wire \top_I.branch[31].block[10].um_I.iw[5] ;
 wire \top_I.branch[31].block[10].um_I.iw[6] ;
 wire \top_I.branch[31].block[10].um_I.iw[7] ;
 wire \top_I.branch[31].block[10].um_I.iw[8] ;
 wire \top_I.branch[31].block[10].um_I.iw[9] ;
 wire \top_I.branch[31].block[10].um_I.k_zero ;
 wire \top_I.branch[31].block[10].um_I.pg_vdd ;
 wire \top_I.branch[31].block[11].um_I.ana[0] ;
 wire \top_I.branch[31].block[11].um_I.ana[1] ;
 wire \top_I.branch[31].block[11].um_I.ana[2] ;
 wire \top_I.branch[31].block[11].um_I.ana[3] ;
 wire \top_I.branch[31].block[11].um_I.ana[4] ;
 wire \top_I.branch[31].block[11].um_I.ana[5] ;
 wire \top_I.branch[31].block[11].um_I.ana[6] ;
 wire \top_I.branch[31].block[11].um_I.ana[7] ;
 wire \top_I.branch[31].block[11].um_I.clk ;
 wire \top_I.branch[31].block[11].um_I.ena ;
 wire \top_I.branch[31].block[11].um_I.iw[10] ;
 wire \top_I.branch[31].block[11].um_I.iw[11] ;
 wire \top_I.branch[31].block[11].um_I.iw[12] ;
 wire \top_I.branch[31].block[11].um_I.iw[13] ;
 wire \top_I.branch[31].block[11].um_I.iw[14] ;
 wire \top_I.branch[31].block[11].um_I.iw[15] ;
 wire \top_I.branch[31].block[11].um_I.iw[16] ;
 wire \top_I.branch[31].block[11].um_I.iw[17] ;
 wire \top_I.branch[31].block[11].um_I.iw[1] ;
 wire \top_I.branch[31].block[11].um_I.iw[2] ;
 wire \top_I.branch[31].block[11].um_I.iw[3] ;
 wire \top_I.branch[31].block[11].um_I.iw[4] ;
 wire \top_I.branch[31].block[11].um_I.iw[5] ;
 wire \top_I.branch[31].block[11].um_I.iw[6] ;
 wire \top_I.branch[31].block[11].um_I.iw[7] ;
 wire \top_I.branch[31].block[11].um_I.iw[8] ;
 wire \top_I.branch[31].block[11].um_I.iw[9] ;
 wire \top_I.branch[31].block[11].um_I.k_zero ;
 wire \top_I.branch[31].block[11].um_I.pg_vdd ;
 wire \top_I.branch[31].block[12].um_I.ana[0] ;
 wire \top_I.branch[31].block[12].um_I.ana[1] ;
 wire \top_I.branch[31].block[12].um_I.ana[2] ;
 wire \top_I.branch[31].block[12].um_I.ana[3] ;
 wire \top_I.branch[31].block[12].um_I.ana[4] ;
 wire \top_I.branch[31].block[12].um_I.ana[5] ;
 wire \top_I.branch[31].block[12].um_I.ana[6] ;
 wire \top_I.branch[31].block[12].um_I.ana[7] ;
 wire \top_I.branch[31].block[12].um_I.clk ;
 wire \top_I.branch[31].block[12].um_I.ena ;
 wire \top_I.branch[31].block[12].um_I.iw[10] ;
 wire \top_I.branch[31].block[12].um_I.iw[11] ;
 wire \top_I.branch[31].block[12].um_I.iw[12] ;
 wire \top_I.branch[31].block[12].um_I.iw[13] ;
 wire \top_I.branch[31].block[12].um_I.iw[14] ;
 wire \top_I.branch[31].block[12].um_I.iw[15] ;
 wire \top_I.branch[31].block[12].um_I.iw[16] ;
 wire \top_I.branch[31].block[12].um_I.iw[17] ;
 wire \top_I.branch[31].block[12].um_I.iw[1] ;
 wire \top_I.branch[31].block[12].um_I.iw[2] ;
 wire \top_I.branch[31].block[12].um_I.iw[3] ;
 wire \top_I.branch[31].block[12].um_I.iw[4] ;
 wire \top_I.branch[31].block[12].um_I.iw[5] ;
 wire \top_I.branch[31].block[12].um_I.iw[6] ;
 wire \top_I.branch[31].block[12].um_I.iw[7] ;
 wire \top_I.branch[31].block[12].um_I.iw[8] ;
 wire \top_I.branch[31].block[12].um_I.iw[9] ;
 wire \top_I.branch[31].block[12].um_I.k_zero ;
 wire \top_I.branch[31].block[12].um_I.pg_vdd ;
 wire \top_I.branch[31].block[13].um_I.ana[0] ;
 wire \top_I.branch[31].block[13].um_I.ana[1] ;
 wire \top_I.branch[31].block[13].um_I.ana[2] ;
 wire \top_I.branch[31].block[13].um_I.ana[3] ;
 wire \top_I.branch[31].block[13].um_I.ana[4] ;
 wire \top_I.branch[31].block[13].um_I.ana[5] ;
 wire \top_I.branch[31].block[13].um_I.ana[6] ;
 wire \top_I.branch[31].block[13].um_I.ana[7] ;
 wire \top_I.branch[31].block[13].um_I.clk ;
 wire \top_I.branch[31].block[13].um_I.ena ;
 wire \top_I.branch[31].block[13].um_I.iw[10] ;
 wire \top_I.branch[31].block[13].um_I.iw[11] ;
 wire \top_I.branch[31].block[13].um_I.iw[12] ;
 wire \top_I.branch[31].block[13].um_I.iw[13] ;
 wire \top_I.branch[31].block[13].um_I.iw[14] ;
 wire \top_I.branch[31].block[13].um_I.iw[15] ;
 wire \top_I.branch[31].block[13].um_I.iw[16] ;
 wire \top_I.branch[31].block[13].um_I.iw[17] ;
 wire \top_I.branch[31].block[13].um_I.iw[1] ;
 wire \top_I.branch[31].block[13].um_I.iw[2] ;
 wire \top_I.branch[31].block[13].um_I.iw[3] ;
 wire \top_I.branch[31].block[13].um_I.iw[4] ;
 wire \top_I.branch[31].block[13].um_I.iw[5] ;
 wire \top_I.branch[31].block[13].um_I.iw[6] ;
 wire \top_I.branch[31].block[13].um_I.iw[7] ;
 wire \top_I.branch[31].block[13].um_I.iw[8] ;
 wire \top_I.branch[31].block[13].um_I.iw[9] ;
 wire \top_I.branch[31].block[13].um_I.k_zero ;
 wire \top_I.branch[31].block[13].um_I.pg_vdd ;
 wire \top_I.branch[31].block[14].um_I.ana[0] ;
 wire \top_I.branch[31].block[14].um_I.ana[1] ;
 wire \top_I.branch[31].block[14].um_I.ana[2] ;
 wire \top_I.branch[31].block[14].um_I.ana[3] ;
 wire \top_I.branch[31].block[14].um_I.ana[4] ;
 wire \top_I.branch[31].block[14].um_I.ana[5] ;
 wire \top_I.branch[31].block[14].um_I.ana[6] ;
 wire \top_I.branch[31].block[14].um_I.ana[7] ;
 wire \top_I.branch[31].block[14].um_I.clk ;
 wire \top_I.branch[31].block[14].um_I.ena ;
 wire \top_I.branch[31].block[14].um_I.iw[10] ;
 wire \top_I.branch[31].block[14].um_I.iw[11] ;
 wire \top_I.branch[31].block[14].um_I.iw[12] ;
 wire \top_I.branch[31].block[14].um_I.iw[13] ;
 wire \top_I.branch[31].block[14].um_I.iw[14] ;
 wire \top_I.branch[31].block[14].um_I.iw[15] ;
 wire \top_I.branch[31].block[14].um_I.iw[16] ;
 wire \top_I.branch[31].block[14].um_I.iw[17] ;
 wire \top_I.branch[31].block[14].um_I.iw[1] ;
 wire \top_I.branch[31].block[14].um_I.iw[2] ;
 wire \top_I.branch[31].block[14].um_I.iw[3] ;
 wire \top_I.branch[31].block[14].um_I.iw[4] ;
 wire \top_I.branch[31].block[14].um_I.iw[5] ;
 wire \top_I.branch[31].block[14].um_I.iw[6] ;
 wire \top_I.branch[31].block[14].um_I.iw[7] ;
 wire \top_I.branch[31].block[14].um_I.iw[8] ;
 wire \top_I.branch[31].block[14].um_I.iw[9] ;
 wire \top_I.branch[31].block[14].um_I.k_zero ;
 wire \top_I.branch[31].block[14].um_I.pg_vdd ;
 wire \top_I.branch[31].block[15].um_I.ana[0] ;
 wire \top_I.branch[31].block[15].um_I.ana[1] ;
 wire \top_I.branch[31].block[15].um_I.ana[2] ;
 wire \top_I.branch[31].block[15].um_I.ana[3] ;
 wire \top_I.branch[31].block[15].um_I.ana[4] ;
 wire \top_I.branch[31].block[15].um_I.ana[5] ;
 wire \top_I.branch[31].block[15].um_I.ana[6] ;
 wire \top_I.branch[31].block[15].um_I.ana[7] ;
 wire \top_I.branch[31].block[15].um_I.clk ;
 wire \top_I.branch[31].block[15].um_I.ena ;
 wire \top_I.branch[31].block[15].um_I.iw[10] ;
 wire \top_I.branch[31].block[15].um_I.iw[11] ;
 wire \top_I.branch[31].block[15].um_I.iw[12] ;
 wire \top_I.branch[31].block[15].um_I.iw[13] ;
 wire \top_I.branch[31].block[15].um_I.iw[14] ;
 wire \top_I.branch[31].block[15].um_I.iw[15] ;
 wire \top_I.branch[31].block[15].um_I.iw[16] ;
 wire \top_I.branch[31].block[15].um_I.iw[17] ;
 wire \top_I.branch[31].block[15].um_I.iw[1] ;
 wire \top_I.branch[31].block[15].um_I.iw[2] ;
 wire \top_I.branch[31].block[15].um_I.iw[3] ;
 wire \top_I.branch[31].block[15].um_I.iw[4] ;
 wire \top_I.branch[31].block[15].um_I.iw[5] ;
 wire \top_I.branch[31].block[15].um_I.iw[6] ;
 wire \top_I.branch[31].block[15].um_I.iw[7] ;
 wire \top_I.branch[31].block[15].um_I.iw[8] ;
 wire \top_I.branch[31].block[15].um_I.iw[9] ;
 wire \top_I.branch[31].block[15].um_I.k_zero ;
 wire \top_I.branch[31].block[15].um_I.pg_vdd ;
 wire \top_I.branch[31].block[1].um_I.ana[0] ;
 wire \top_I.branch[31].block[1].um_I.ana[1] ;
 wire \top_I.branch[31].block[1].um_I.ana[2] ;
 wire \top_I.branch[31].block[1].um_I.ana[3] ;
 wire \top_I.branch[31].block[1].um_I.ana[4] ;
 wire \top_I.branch[31].block[1].um_I.ana[5] ;
 wire \top_I.branch[31].block[1].um_I.ana[6] ;
 wire \top_I.branch[31].block[1].um_I.ana[7] ;
 wire \top_I.branch[31].block[1].um_I.clk ;
 wire \top_I.branch[31].block[1].um_I.ena ;
 wire \top_I.branch[31].block[1].um_I.iw[10] ;
 wire \top_I.branch[31].block[1].um_I.iw[11] ;
 wire \top_I.branch[31].block[1].um_I.iw[12] ;
 wire \top_I.branch[31].block[1].um_I.iw[13] ;
 wire \top_I.branch[31].block[1].um_I.iw[14] ;
 wire \top_I.branch[31].block[1].um_I.iw[15] ;
 wire \top_I.branch[31].block[1].um_I.iw[16] ;
 wire \top_I.branch[31].block[1].um_I.iw[17] ;
 wire \top_I.branch[31].block[1].um_I.iw[1] ;
 wire \top_I.branch[31].block[1].um_I.iw[2] ;
 wire \top_I.branch[31].block[1].um_I.iw[3] ;
 wire \top_I.branch[31].block[1].um_I.iw[4] ;
 wire \top_I.branch[31].block[1].um_I.iw[5] ;
 wire \top_I.branch[31].block[1].um_I.iw[6] ;
 wire \top_I.branch[31].block[1].um_I.iw[7] ;
 wire \top_I.branch[31].block[1].um_I.iw[8] ;
 wire \top_I.branch[31].block[1].um_I.iw[9] ;
 wire \top_I.branch[31].block[1].um_I.k_zero ;
 wire \top_I.branch[31].block[1].um_I.pg_vdd ;
 wire \top_I.branch[31].block[2].um_I.ana[0] ;
 wire \top_I.branch[31].block[2].um_I.ana[1] ;
 wire \top_I.branch[31].block[2].um_I.ana[2] ;
 wire \top_I.branch[31].block[2].um_I.ana[3] ;
 wire \top_I.branch[31].block[2].um_I.ana[4] ;
 wire \top_I.branch[31].block[2].um_I.ana[5] ;
 wire \top_I.branch[31].block[2].um_I.ana[6] ;
 wire \top_I.branch[31].block[2].um_I.ana[7] ;
 wire \top_I.branch[31].block[2].um_I.clk ;
 wire \top_I.branch[31].block[2].um_I.ena ;
 wire \top_I.branch[31].block[2].um_I.iw[10] ;
 wire \top_I.branch[31].block[2].um_I.iw[11] ;
 wire \top_I.branch[31].block[2].um_I.iw[12] ;
 wire \top_I.branch[31].block[2].um_I.iw[13] ;
 wire \top_I.branch[31].block[2].um_I.iw[14] ;
 wire \top_I.branch[31].block[2].um_I.iw[15] ;
 wire \top_I.branch[31].block[2].um_I.iw[16] ;
 wire \top_I.branch[31].block[2].um_I.iw[17] ;
 wire \top_I.branch[31].block[2].um_I.iw[1] ;
 wire \top_I.branch[31].block[2].um_I.iw[2] ;
 wire \top_I.branch[31].block[2].um_I.iw[3] ;
 wire \top_I.branch[31].block[2].um_I.iw[4] ;
 wire \top_I.branch[31].block[2].um_I.iw[5] ;
 wire \top_I.branch[31].block[2].um_I.iw[6] ;
 wire \top_I.branch[31].block[2].um_I.iw[7] ;
 wire \top_I.branch[31].block[2].um_I.iw[8] ;
 wire \top_I.branch[31].block[2].um_I.iw[9] ;
 wire \top_I.branch[31].block[2].um_I.k_zero ;
 wire \top_I.branch[31].block[2].um_I.pg_vdd ;
 wire \top_I.branch[31].block[3].um_I.ana[0] ;
 wire \top_I.branch[31].block[3].um_I.ana[1] ;
 wire \top_I.branch[31].block[3].um_I.ana[2] ;
 wire \top_I.branch[31].block[3].um_I.ana[3] ;
 wire \top_I.branch[31].block[3].um_I.ana[4] ;
 wire \top_I.branch[31].block[3].um_I.ana[5] ;
 wire \top_I.branch[31].block[3].um_I.ana[6] ;
 wire \top_I.branch[31].block[3].um_I.ana[7] ;
 wire \top_I.branch[31].block[3].um_I.clk ;
 wire \top_I.branch[31].block[3].um_I.ena ;
 wire \top_I.branch[31].block[3].um_I.iw[10] ;
 wire \top_I.branch[31].block[3].um_I.iw[11] ;
 wire \top_I.branch[31].block[3].um_I.iw[12] ;
 wire \top_I.branch[31].block[3].um_I.iw[13] ;
 wire \top_I.branch[31].block[3].um_I.iw[14] ;
 wire \top_I.branch[31].block[3].um_I.iw[15] ;
 wire \top_I.branch[31].block[3].um_I.iw[16] ;
 wire \top_I.branch[31].block[3].um_I.iw[17] ;
 wire \top_I.branch[31].block[3].um_I.iw[1] ;
 wire \top_I.branch[31].block[3].um_I.iw[2] ;
 wire \top_I.branch[31].block[3].um_I.iw[3] ;
 wire \top_I.branch[31].block[3].um_I.iw[4] ;
 wire \top_I.branch[31].block[3].um_I.iw[5] ;
 wire \top_I.branch[31].block[3].um_I.iw[6] ;
 wire \top_I.branch[31].block[3].um_I.iw[7] ;
 wire \top_I.branch[31].block[3].um_I.iw[8] ;
 wire \top_I.branch[31].block[3].um_I.iw[9] ;
 wire \top_I.branch[31].block[3].um_I.k_zero ;
 wire \top_I.branch[31].block[3].um_I.pg_vdd ;
 wire \top_I.branch[31].block[4].um_I.ana[0] ;
 wire \top_I.branch[31].block[4].um_I.ana[1] ;
 wire \top_I.branch[31].block[4].um_I.ana[2] ;
 wire \top_I.branch[31].block[4].um_I.ana[3] ;
 wire \top_I.branch[31].block[4].um_I.ana[4] ;
 wire \top_I.branch[31].block[4].um_I.ana[5] ;
 wire \top_I.branch[31].block[4].um_I.ana[6] ;
 wire \top_I.branch[31].block[4].um_I.ana[7] ;
 wire \top_I.branch[31].block[4].um_I.clk ;
 wire \top_I.branch[31].block[4].um_I.ena ;
 wire \top_I.branch[31].block[4].um_I.iw[10] ;
 wire \top_I.branch[31].block[4].um_I.iw[11] ;
 wire \top_I.branch[31].block[4].um_I.iw[12] ;
 wire \top_I.branch[31].block[4].um_I.iw[13] ;
 wire \top_I.branch[31].block[4].um_I.iw[14] ;
 wire \top_I.branch[31].block[4].um_I.iw[15] ;
 wire \top_I.branch[31].block[4].um_I.iw[16] ;
 wire \top_I.branch[31].block[4].um_I.iw[17] ;
 wire \top_I.branch[31].block[4].um_I.iw[1] ;
 wire \top_I.branch[31].block[4].um_I.iw[2] ;
 wire \top_I.branch[31].block[4].um_I.iw[3] ;
 wire \top_I.branch[31].block[4].um_I.iw[4] ;
 wire \top_I.branch[31].block[4].um_I.iw[5] ;
 wire \top_I.branch[31].block[4].um_I.iw[6] ;
 wire \top_I.branch[31].block[4].um_I.iw[7] ;
 wire \top_I.branch[31].block[4].um_I.iw[8] ;
 wire \top_I.branch[31].block[4].um_I.iw[9] ;
 wire \top_I.branch[31].block[4].um_I.k_zero ;
 wire \top_I.branch[31].block[4].um_I.pg_vdd ;
 wire \top_I.branch[31].block[5].um_I.ana[0] ;
 wire \top_I.branch[31].block[5].um_I.ana[1] ;
 wire \top_I.branch[31].block[5].um_I.ana[2] ;
 wire \top_I.branch[31].block[5].um_I.ana[3] ;
 wire \top_I.branch[31].block[5].um_I.ana[4] ;
 wire \top_I.branch[31].block[5].um_I.ana[5] ;
 wire \top_I.branch[31].block[5].um_I.ana[6] ;
 wire \top_I.branch[31].block[5].um_I.ana[7] ;
 wire \top_I.branch[31].block[5].um_I.clk ;
 wire \top_I.branch[31].block[5].um_I.ena ;
 wire \top_I.branch[31].block[5].um_I.iw[10] ;
 wire \top_I.branch[31].block[5].um_I.iw[11] ;
 wire \top_I.branch[31].block[5].um_I.iw[12] ;
 wire \top_I.branch[31].block[5].um_I.iw[13] ;
 wire \top_I.branch[31].block[5].um_I.iw[14] ;
 wire \top_I.branch[31].block[5].um_I.iw[15] ;
 wire \top_I.branch[31].block[5].um_I.iw[16] ;
 wire \top_I.branch[31].block[5].um_I.iw[17] ;
 wire \top_I.branch[31].block[5].um_I.iw[1] ;
 wire \top_I.branch[31].block[5].um_I.iw[2] ;
 wire \top_I.branch[31].block[5].um_I.iw[3] ;
 wire \top_I.branch[31].block[5].um_I.iw[4] ;
 wire \top_I.branch[31].block[5].um_I.iw[5] ;
 wire \top_I.branch[31].block[5].um_I.iw[6] ;
 wire \top_I.branch[31].block[5].um_I.iw[7] ;
 wire \top_I.branch[31].block[5].um_I.iw[8] ;
 wire \top_I.branch[31].block[5].um_I.iw[9] ;
 wire \top_I.branch[31].block[5].um_I.k_zero ;
 wire \top_I.branch[31].block[5].um_I.pg_vdd ;
 wire \top_I.branch[31].block[6].um_I.ana[0] ;
 wire \top_I.branch[31].block[6].um_I.ana[1] ;
 wire \top_I.branch[31].block[6].um_I.ana[2] ;
 wire \top_I.branch[31].block[6].um_I.ana[3] ;
 wire \top_I.branch[31].block[6].um_I.ana[4] ;
 wire \top_I.branch[31].block[6].um_I.ana[5] ;
 wire \top_I.branch[31].block[6].um_I.ana[6] ;
 wire \top_I.branch[31].block[6].um_I.ana[7] ;
 wire \top_I.branch[31].block[6].um_I.clk ;
 wire \top_I.branch[31].block[6].um_I.ena ;
 wire \top_I.branch[31].block[6].um_I.iw[10] ;
 wire \top_I.branch[31].block[6].um_I.iw[11] ;
 wire \top_I.branch[31].block[6].um_I.iw[12] ;
 wire \top_I.branch[31].block[6].um_I.iw[13] ;
 wire \top_I.branch[31].block[6].um_I.iw[14] ;
 wire \top_I.branch[31].block[6].um_I.iw[15] ;
 wire \top_I.branch[31].block[6].um_I.iw[16] ;
 wire \top_I.branch[31].block[6].um_I.iw[17] ;
 wire \top_I.branch[31].block[6].um_I.iw[1] ;
 wire \top_I.branch[31].block[6].um_I.iw[2] ;
 wire \top_I.branch[31].block[6].um_I.iw[3] ;
 wire \top_I.branch[31].block[6].um_I.iw[4] ;
 wire \top_I.branch[31].block[6].um_I.iw[5] ;
 wire \top_I.branch[31].block[6].um_I.iw[6] ;
 wire \top_I.branch[31].block[6].um_I.iw[7] ;
 wire \top_I.branch[31].block[6].um_I.iw[8] ;
 wire \top_I.branch[31].block[6].um_I.iw[9] ;
 wire \top_I.branch[31].block[6].um_I.k_zero ;
 wire \top_I.branch[31].block[6].um_I.pg_vdd ;
 wire \top_I.branch[31].block[7].um_I.ana[0] ;
 wire \top_I.branch[31].block[7].um_I.ana[1] ;
 wire \top_I.branch[31].block[7].um_I.ana[2] ;
 wire \top_I.branch[31].block[7].um_I.ana[3] ;
 wire \top_I.branch[31].block[7].um_I.ana[4] ;
 wire \top_I.branch[31].block[7].um_I.ana[5] ;
 wire \top_I.branch[31].block[7].um_I.ana[6] ;
 wire \top_I.branch[31].block[7].um_I.ana[7] ;
 wire \top_I.branch[31].block[7].um_I.clk ;
 wire \top_I.branch[31].block[7].um_I.ena ;
 wire \top_I.branch[31].block[7].um_I.iw[10] ;
 wire \top_I.branch[31].block[7].um_I.iw[11] ;
 wire \top_I.branch[31].block[7].um_I.iw[12] ;
 wire \top_I.branch[31].block[7].um_I.iw[13] ;
 wire \top_I.branch[31].block[7].um_I.iw[14] ;
 wire \top_I.branch[31].block[7].um_I.iw[15] ;
 wire \top_I.branch[31].block[7].um_I.iw[16] ;
 wire \top_I.branch[31].block[7].um_I.iw[17] ;
 wire \top_I.branch[31].block[7].um_I.iw[1] ;
 wire \top_I.branch[31].block[7].um_I.iw[2] ;
 wire \top_I.branch[31].block[7].um_I.iw[3] ;
 wire \top_I.branch[31].block[7].um_I.iw[4] ;
 wire \top_I.branch[31].block[7].um_I.iw[5] ;
 wire \top_I.branch[31].block[7].um_I.iw[6] ;
 wire \top_I.branch[31].block[7].um_I.iw[7] ;
 wire \top_I.branch[31].block[7].um_I.iw[8] ;
 wire \top_I.branch[31].block[7].um_I.iw[9] ;
 wire \top_I.branch[31].block[7].um_I.k_zero ;
 wire \top_I.branch[31].block[7].um_I.pg_vdd ;
 wire \top_I.branch[31].block[8].um_I.ana[0] ;
 wire \top_I.branch[31].block[8].um_I.ana[1] ;
 wire \top_I.branch[31].block[8].um_I.ana[2] ;
 wire \top_I.branch[31].block[8].um_I.ana[3] ;
 wire \top_I.branch[31].block[8].um_I.ana[4] ;
 wire \top_I.branch[31].block[8].um_I.ana[5] ;
 wire \top_I.branch[31].block[8].um_I.ana[6] ;
 wire \top_I.branch[31].block[8].um_I.ana[7] ;
 wire \top_I.branch[31].block[8].um_I.clk ;
 wire \top_I.branch[31].block[8].um_I.ena ;
 wire \top_I.branch[31].block[8].um_I.iw[10] ;
 wire \top_I.branch[31].block[8].um_I.iw[11] ;
 wire \top_I.branch[31].block[8].um_I.iw[12] ;
 wire \top_I.branch[31].block[8].um_I.iw[13] ;
 wire \top_I.branch[31].block[8].um_I.iw[14] ;
 wire \top_I.branch[31].block[8].um_I.iw[15] ;
 wire \top_I.branch[31].block[8].um_I.iw[16] ;
 wire \top_I.branch[31].block[8].um_I.iw[17] ;
 wire \top_I.branch[31].block[8].um_I.iw[1] ;
 wire \top_I.branch[31].block[8].um_I.iw[2] ;
 wire \top_I.branch[31].block[8].um_I.iw[3] ;
 wire \top_I.branch[31].block[8].um_I.iw[4] ;
 wire \top_I.branch[31].block[8].um_I.iw[5] ;
 wire \top_I.branch[31].block[8].um_I.iw[6] ;
 wire \top_I.branch[31].block[8].um_I.iw[7] ;
 wire \top_I.branch[31].block[8].um_I.iw[8] ;
 wire \top_I.branch[31].block[8].um_I.iw[9] ;
 wire \top_I.branch[31].block[8].um_I.k_zero ;
 wire \top_I.branch[31].block[8].um_I.pg_vdd ;
 wire \top_I.branch[31].block[9].um_I.ana[0] ;
 wire \top_I.branch[31].block[9].um_I.ana[1] ;
 wire \top_I.branch[31].block[9].um_I.ana[2] ;
 wire \top_I.branch[31].block[9].um_I.ana[3] ;
 wire \top_I.branch[31].block[9].um_I.ana[4] ;
 wire \top_I.branch[31].block[9].um_I.ana[5] ;
 wire \top_I.branch[31].block[9].um_I.ana[6] ;
 wire \top_I.branch[31].block[9].um_I.ana[7] ;
 wire \top_I.branch[31].block[9].um_I.clk ;
 wire \top_I.branch[31].block[9].um_I.ena ;
 wire \top_I.branch[31].block[9].um_I.iw[10] ;
 wire \top_I.branch[31].block[9].um_I.iw[11] ;
 wire \top_I.branch[31].block[9].um_I.iw[12] ;
 wire \top_I.branch[31].block[9].um_I.iw[13] ;
 wire \top_I.branch[31].block[9].um_I.iw[14] ;
 wire \top_I.branch[31].block[9].um_I.iw[15] ;
 wire \top_I.branch[31].block[9].um_I.iw[16] ;
 wire \top_I.branch[31].block[9].um_I.iw[17] ;
 wire \top_I.branch[31].block[9].um_I.iw[1] ;
 wire \top_I.branch[31].block[9].um_I.iw[2] ;
 wire \top_I.branch[31].block[9].um_I.iw[3] ;
 wire \top_I.branch[31].block[9].um_I.iw[4] ;
 wire \top_I.branch[31].block[9].um_I.iw[5] ;
 wire \top_I.branch[31].block[9].um_I.iw[6] ;
 wire \top_I.branch[31].block[9].um_I.iw[7] ;
 wire \top_I.branch[31].block[9].um_I.iw[8] ;
 wire \top_I.branch[31].block[9].um_I.iw[9] ;
 wire \top_I.branch[31].block[9].um_I.k_zero ;
 wire \top_I.branch[31].block[9].um_I.pg_vdd ;
 wire \top_I.branch[31].l_addr[0] ;
 wire \top_I.branch[31].l_k_zero ;
 wire \top_I.branch[3].block[0].um_I.ana[0] ;
 wire \top_I.branch[3].block[0].um_I.ana[1] ;
 wire \top_I.branch[3].block[0].um_I.ana[2] ;
 wire \top_I.branch[3].block[0].um_I.ana[3] ;
 wire \top_I.branch[3].block[0].um_I.ana[4] ;
 wire \top_I.branch[3].block[0].um_I.ana[5] ;
 wire \top_I.branch[3].block[0].um_I.ana[6] ;
 wire \top_I.branch[3].block[0].um_I.ana[7] ;
 wire \top_I.branch[3].block[0].um_I.clk ;
 wire \top_I.branch[3].block[0].um_I.ena ;
 wire \top_I.branch[3].block[0].um_I.iw[10] ;
 wire \top_I.branch[3].block[0].um_I.iw[11] ;
 wire \top_I.branch[3].block[0].um_I.iw[12] ;
 wire \top_I.branch[3].block[0].um_I.iw[13] ;
 wire \top_I.branch[3].block[0].um_I.iw[14] ;
 wire \top_I.branch[3].block[0].um_I.iw[15] ;
 wire \top_I.branch[3].block[0].um_I.iw[16] ;
 wire \top_I.branch[3].block[0].um_I.iw[17] ;
 wire \top_I.branch[3].block[0].um_I.iw[1] ;
 wire \top_I.branch[3].block[0].um_I.iw[2] ;
 wire \top_I.branch[3].block[0].um_I.iw[3] ;
 wire \top_I.branch[3].block[0].um_I.iw[4] ;
 wire \top_I.branch[3].block[0].um_I.iw[5] ;
 wire \top_I.branch[3].block[0].um_I.iw[6] ;
 wire \top_I.branch[3].block[0].um_I.iw[7] ;
 wire \top_I.branch[3].block[0].um_I.iw[8] ;
 wire \top_I.branch[3].block[0].um_I.iw[9] ;
 wire \top_I.branch[3].block[0].um_I.k_zero ;
 wire \top_I.branch[3].block[0].um_I.pg_vdd ;
 wire \top_I.branch[3].block[10].um_I.ana[0] ;
 wire \top_I.branch[3].block[10].um_I.ana[1] ;
 wire \top_I.branch[3].block[10].um_I.ana[2] ;
 wire \top_I.branch[3].block[10].um_I.ana[3] ;
 wire \top_I.branch[3].block[10].um_I.ana[4] ;
 wire \top_I.branch[3].block[10].um_I.ana[5] ;
 wire \top_I.branch[3].block[10].um_I.ana[6] ;
 wire \top_I.branch[3].block[10].um_I.ana[7] ;
 wire \top_I.branch[3].block[10].um_I.clk ;
 wire \top_I.branch[3].block[10].um_I.ena ;
 wire \top_I.branch[3].block[10].um_I.iw[10] ;
 wire \top_I.branch[3].block[10].um_I.iw[11] ;
 wire \top_I.branch[3].block[10].um_I.iw[12] ;
 wire \top_I.branch[3].block[10].um_I.iw[13] ;
 wire \top_I.branch[3].block[10].um_I.iw[14] ;
 wire \top_I.branch[3].block[10].um_I.iw[15] ;
 wire \top_I.branch[3].block[10].um_I.iw[16] ;
 wire \top_I.branch[3].block[10].um_I.iw[17] ;
 wire \top_I.branch[3].block[10].um_I.iw[1] ;
 wire \top_I.branch[3].block[10].um_I.iw[2] ;
 wire \top_I.branch[3].block[10].um_I.iw[3] ;
 wire \top_I.branch[3].block[10].um_I.iw[4] ;
 wire \top_I.branch[3].block[10].um_I.iw[5] ;
 wire \top_I.branch[3].block[10].um_I.iw[6] ;
 wire \top_I.branch[3].block[10].um_I.iw[7] ;
 wire \top_I.branch[3].block[10].um_I.iw[8] ;
 wire \top_I.branch[3].block[10].um_I.iw[9] ;
 wire \top_I.branch[3].block[10].um_I.k_zero ;
 wire \top_I.branch[3].block[10].um_I.pg_vdd ;
 wire \top_I.branch[3].block[11].um_I.ana[0] ;
 wire \top_I.branch[3].block[11].um_I.ana[1] ;
 wire \top_I.branch[3].block[11].um_I.ana[2] ;
 wire \top_I.branch[3].block[11].um_I.ana[3] ;
 wire \top_I.branch[3].block[11].um_I.ana[4] ;
 wire \top_I.branch[3].block[11].um_I.ana[5] ;
 wire \top_I.branch[3].block[11].um_I.ana[6] ;
 wire \top_I.branch[3].block[11].um_I.ana[7] ;
 wire \top_I.branch[3].block[11].um_I.clk ;
 wire \top_I.branch[3].block[11].um_I.ena ;
 wire \top_I.branch[3].block[11].um_I.iw[10] ;
 wire \top_I.branch[3].block[11].um_I.iw[11] ;
 wire \top_I.branch[3].block[11].um_I.iw[12] ;
 wire \top_I.branch[3].block[11].um_I.iw[13] ;
 wire \top_I.branch[3].block[11].um_I.iw[14] ;
 wire \top_I.branch[3].block[11].um_I.iw[15] ;
 wire \top_I.branch[3].block[11].um_I.iw[16] ;
 wire \top_I.branch[3].block[11].um_I.iw[17] ;
 wire \top_I.branch[3].block[11].um_I.iw[1] ;
 wire \top_I.branch[3].block[11].um_I.iw[2] ;
 wire \top_I.branch[3].block[11].um_I.iw[3] ;
 wire \top_I.branch[3].block[11].um_I.iw[4] ;
 wire \top_I.branch[3].block[11].um_I.iw[5] ;
 wire \top_I.branch[3].block[11].um_I.iw[6] ;
 wire \top_I.branch[3].block[11].um_I.iw[7] ;
 wire \top_I.branch[3].block[11].um_I.iw[8] ;
 wire \top_I.branch[3].block[11].um_I.iw[9] ;
 wire \top_I.branch[3].block[11].um_I.k_zero ;
 wire \top_I.branch[3].block[11].um_I.pg_vdd ;
 wire \top_I.branch[3].block[12].um_I.ana[0] ;
 wire \top_I.branch[3].block[12].um_I.ana[1] ;
 wire \top_I.branch[3].block[12].um_I.ana[2] ;
 wire \top_I.branch[3].block[12].um_I.ana[3] ;
 wire \top_I.branch[3].block[12].um_I.ana[4] ;
 wire \top_I.branch[3].block[12].um_I.ana[5] ;
 wire \top_I.branch[3].block[12].um_I.ana[6] ;
 wire \top_I.branch[3].block[12].um_I.ana[7] ;
 wire \top_I.branch[3].block[12].um_I.clk ;
 wire \top_I.branch[3].block[12].um_I.ena ;
 wire \top_I.branch[3].block[12].um_I.iw[10] ;
 wire \top_I.branch[3].block[12].um_I.iw[11] ;
 wire \top_I.branch[3].block[12].um_I.iw[12] ;
 wire \top_I.branch[3].block[12].um_I.iw[13] ;
 wire \top_I.branch[3].block[12].um_I.iw[14] ;
 wire \top_I.branch[3].block[12].um_I.iw[15] ;
 wire \top_I.branch[3].block[12].um_I.iw[16] ;
 wire \top_I.branch[3].block[12].um_I.iw[17] ;
 wire \top_I.branch[3].block[12].um_I.iw[1] ;
 wire \top_I.branch[3].block[12].um_I.iw[2] ;
 wire \top_I.branch[3].block[12].um_I.iw[3] ;
 wire \top_I.branch[3].block[12].um_I.iw[4] ;
 wire \top_I.branch[3].block[12].um_I.iw[5] ;
 wire \top_I.branch[3].block[12].um_I.iw[6] ;
 wire \top_I.branch[3].block[12].um_I.iw[7] ;
 wire \top_I.branch[3].block[12].um_I.iw[8] ;
 wire \top_I.branch[3].block[12].um_I.iw[9] ;
 wire \top_I.branch[3].block[12].um_I.k_zero ;
 wire \top_I.branch[3].block[12].um_I.pg_vdd ;
 wire \top_I.branch[3].block[13].um_I.ana[0] ;
 wire \top_I.branch[3].block[13].um_I.ana[1] ;
 wire \top_I.branch[3].block[13].um_I.ana[2] ;
 wire \top_I.branch[3].block[13].um_I.ana[3] ;
 wire \top_I.branch[3].block[13].um_I.ana[4] ;
 wire \top_I.branch[3].block[13].um_I.ana[5] ;
 wire \top_I.branch[3].block[13].um_I.ana[6] ;
 wire \top_I.branch[3].block[13].um_I.ana[7] ;
 wire \top_I.branch[3].block[13].um_I.clk ;
 wire \top_I.branch[3].block[13].um_I.ena ;
 wire \top_I.branch[3].block[13].um_I.iw[10] ;
 wire \top_I.branch[3].block[13].um_I.iw[11] ;
 wire \top_I.branch[3].block[13].um_I.iw[12] ;
 wire \top_I.branch[3].block[13].um_I.iw[13] ;
 wire \top_I.branch[3].block[13].um_I.iw[14] ;
 wire \top_I.branch[3].block[13].um_I.iw[15] ;
 wire \top_I.branch[3].block[13].um_I.iw[16] ;
 wire \top_I.branch[3].block[13].um_I.iw[17] ;
 wire \top_I.branch[3].block[13].um_I.iw[1] ;
 wire \top_I.branch[3].block[13].um_I.iw[2] ;
 wire \top_I.branch[3].block[13].um_I.iw[3] ;
 wire \top_I.branch[3].block[13].um_I.iw[4] ;
 wire \top_I.branch[3].block[13].um_I.iw[5] ;
 wire \top_I.branch[3].block[13].um_I.iw[6] ;
 wire \top_I.branch[3].block[13].um_I.iw[7] ;
 wire \top_I.branch[3].block[13].um_I.iw[8] ;
 wire \top_I.branch[3].block[13].um_I.iw[9] ;
 wire \top_I.branch[3].block[13].um_I.k_zero ;
 wire \top_I.branch[3].block[13].um_I.pg_vdd ;
 wire \top_I.branch[3].block[14].um_I.ana[0] ;
 wire \top_I.branch[3].block[14].um_I.ana[1] ;
 wire \top_I.branch[3].block[14].um_I.ana[2] ;
 wire \top_I.branch[3].block[14].um_I.ana[3] ;
 wire \top_I.branch[3].block[14].um_I.ana[4] ;
 wire \top_I.branch[3].block[14].um_I.ana[5] ;
 wire \top_I.branch[3].block[14].um_I.ana[6] ;
 wire \top_I.branch[3].block[14].um_I.ana[7] ;
 wire \top_I.branch[3].block[14].um_I.clk ;
 wire \top_I.branch[3].block[14].um_I.ena ;
 wire \top_I.branch[3].block[14].um_I.iw[10] ;
 wire \top_I.branch[3].block[14].um_I.iw[11] ;
 wire \top_I.branch[3].block[14].um_I.iw[12] ;
 wire \top_I.branch[3].block[14].um_I.iw[13] ;
 wire \top_I.branch[3].block[14].um_I.iw[14] ;
 wire \top_I.branch[3].block[14].um_I.iw[15] ;
 wire \top_I.branch[3].block[14].um_I.iw[16] ;
 wire \top_I.branch[3].block[14].um_I.iw[17] ;
 wire \top_I.branch[3].block[14].um_I.iw[1] ;
 wire \top_I.branch[3].block[14].um_I.iw[2] ;
 wire \top_I.branch[3].block[14].um_I.iw[3] ;
 wire \top_I.branch[3].block[14].um_I.iw[4] ;
 wire \top_I.branch[3].block[14].um_I.iw[5] ;
 wire \top_I.branch[3].block[14].um_I.iw[6] ;
 wire \top_I.branch[3].block[14].um_I.iw[7] ;
 wire \top_I.branch[3].block[14].um_I.iw[8] ;
 wire \top_I.branch[3].block[14].um_I.iw[9] ;
 wire \top_I.branch[3].block[14].um_I.k_zero ;
 wire \top_I.branch[3].block[14].um_I.pg_vdd ;
 wire \top_I.branch[3].block[15].um_I.ana[0] ;
 wire \top_I.branch[3].block[15].um_I.ana[1] ;
 wire \top_I.branch[3].block[15].um_I.ana[2] ;
 wire \top_I.branch[3].block[15].um_I.ana[3] ;
 wire \top_I.branch[3].block[15].um_I.ana[4] ;
 wire \top_I.branch[3].block[15].um_I.ana[5] ;
 wire \top_I.branch[3].block[15].um_I.ana[6] ;
 wire \top_I.branch[3].block[15].um_I.ana[7] ;
 wire \top_I.branch[3].block[15].um_I.clk ;
 wire \top_I.branch[3].block[15].um_I.ena ;
 wire \top_I.branch[3].block[15].um_I.iw[10] ;
 wire \top_I.branch[3].block[15].um_I.iw[11] ;
 wire \top_I.branch[3].block[15].um_I.iw[12] ;
 wire \top_I.branch[3].block[15].um_I.iw[13] ;
 wire \top_I.branch[3].block[15].um_I.iw[14] ;
 wire \top_I.branch[3].block[15].um_I.iw[15] ;
 wire \top_I.branch[3].block[15].um_I.iw[16] ;
 wire \top_I.branch[3].block[15].um_I.iw[17] ;
 wire \top_I.branch[3].block[15].um_I.iw[1] ;
 wire \top_I.branch[3].block[15].um_I.iw[2] ;
 wire \top_I.branch[3].block[15].um_I.iw[3] ;
 wire \top_I.branch[3].block[15].um_I.iw[4] ;
 wire \top_I.branch[3].block[15].um_I.iw[5] ;
 wire \top_I.branch[3].block[15].um_I.iw[6] ;
 wire \top_I.branch[3].block[15].um_I.iw[7] ;
 wire \top_I.branch[3].block[15].um_I.iw[8] ;
 wire \top_I.branch[3].block[15].um_I.iw[9] ;
 wire \top_I.branch[3].block[15].um_I.k_zero ;
 wire \top_I.branch[3].block[15].um_I.pg_vdd ;
 wire \top_I.branch[3].block[1].um_I.ana[0] ;
 wire \top_I.branch[3].block[1].um_I.ana[1] ;
 wire \top_I.branch[3].block[1].um_I.ana[2] ;
 wire \top_I.branch[3].block[1].um_I.ana[3] ;
 wire \top_I.branch[3].block[1].um_I.ana[4] ;
 wire \top_I.branch[3].block[1].um_I.ana[5] ;
 wire \top_I.branch[3].block[1].um_I.ana[6] ;
 wire \top_I.branch[3].block[1].um_I.ana[7] ;
 wire \top_I.branch[3].block[1].um_I.clk ;
 wire \top_I.branch[3].block[1].um_I.ena ;
 wire \top_I.branch[3].block[1].um_I.iw[10] ;
 wire \top_I.branch[3].block[1].um_I.iw[11] ;
 wire \top_I.branch[3].block[1].um_I.iw[12] ;
 wire \top_I.branch[3].block[1].um_I.iw[13] ;
 wire \top_I.branch[3].block[1].um_I.iw[14] ;
 wire \top_I.branch[3].block[1].um_I.iw[15] ;
 wire \top_I.branch[3].block[1].um_I.iw[16] ;
 wire \top_I.branch[3].block[1].um_I.iw[17] ;
 wire \top_I.branch[3].block[1].um_I.iw[1] ;
 wire \top_I.branch[3].block[1].um_I.iw[2] ;
 wire \top_I.branch[3].block[1].um_I.iw[3] ;
 wire \top_I.branch[3].block[1].um_I.iw[4] ;
 wire \top_I.branch[3].block[1].um_I.iw[5] ;
 wire \top_I.branch[3].block[1].um_I.iw[6] ;
 wire \top_I.branch[3].block[1].um_I.iw[7] ;
 wire \top_I.branch[3].block[1].um_I.iw[8] ;
 wire \top_I.branch[3].block[1].um_I.iw[9] ;
 wire \top_I.branch[3].block[1].um_I.k_zero ;
 wire \top_I.branch[3].block[1].um_I.pg_vdd ;
 wire \top_I.branch[3].block[2].um_I.ana[0] ;
 wire \top_I.branch[3].block[2].um_I.ana[1] ;
 wire \top_I.branch[3].block[2].um_I.ana[2] ;
 wire \top_I.branch[3].block[2].um_I.ana[3] ;
 wire \top_I.branch[3].block[2].um_I.ana[4] ;
 wire \top_I.branch[3].block[2].um_I.ana[5] ;
 wire \top_I.branch[3].block[2].um_I.ana[6] ;
 wire \top_I.branch[3].block[2].um_I.ana[7] ;
 wire \top_I.branch[3].block[2].um_I.clk ;
 wire \top_I.branch[3].block[2].um_I.ena ;
 wire \top_I.branch[3].block[2].um_I.iw[10] ;
 wire \top_I.branch[3].block[2].um_I.iw[11] ;
 wire \top_I.branch[3].block[2].um_I.iw[12] ;
 wire \top_I.branch[3].block[2].um_I.iw[13] ;
 wire \top_I.branch[3].block[2].um_I.iw[14] ;
 wire \top_I.branch[3].block[2].um_I.iw[15] ;
 wire \top_I.branch[3].block[2].um_I.iw[16] ;
 wire \top_I.branch[3].block[2].um_I.iw[17] ;
 wire \top_I.branch[3].block[2].um_I.iw[1] ;
 wire \top_I.branch[3].block[2].um_I.iw[2] ;
 wire \top_I.branch[3].block[2].um_I.iw[3] ;
 wire \top_I.branch[3].block[2].um_I.iw[4] ;
 wire \top_I.branch[3].block[2].um_I.iw[5] ;
 wire \top_I.branch[3].block[2].um_I.iw[6] ;
 wire \top_I.branch[3].block[2].um_I.iw[7] ;
 wire \top_I.branch[3].block[2].um_I.iw[8] ;
 wire \top_I.branch[3].block[2].um_I.iw[9] ;
 wire \top_I.branch[3].block[2].um_I.k_zero ;
 wire \top_I.branch[3].block[2].um_I.pg_vdd ;
 wire \top_I.branch[3].block[3].um_I.ana[0] ;
 wire \top_I.branch[3].block[3].um_I.ana[1] ;
 wire \top_I.branch[3].block[3].um_I.ana[2] ;
 wire \top_I.branch[3].block[3].um_I.ana[3] ;
 wire \top_I.branch[3].block[3].um_I.ana[4] ;
 wire \top_I.branch[3].block[3].um_I.ana[5] ;
 wire \top_I.branch[3].block[3].um_I.ana[6] ;
 wire \top_I.branch[3].block[3].um_I.ana[7] ;
 wire \top_I.branch[3].block[3].um_I.clk ;
 wire \top_I.branch[3].block[3].um_I.ena ;
 wire \top_I.branch[3].block[3].um_I.iw[10] ;
 wire \top_I.branch[3].block[3].um_I.iw[11] ;
 wire \top_I.branch[3].block[3].um_I.iw[12] ;
 wire \top_I.branch[3].block[3].um_I.iw[13] ;
 wire \top_I.branch[3].block[3].um_I.iw[14] ;
 wire \top_I.branch[3].block[3].um_I.iw[15] ;
 wire \top_I.branch[3].block[3].um_I.iw[16] ;
 wire \top_I.branch[3].block[3].um_I.iw[17] ;
 wire \top_I.branch[3].block[3].um_I.iw[1] ;
 wire \top_I.branch[3].block[3].um_I.iw[2] ;
 wire \top_I.branch[3].block[3].um_I.iw[3] ;
 wire \top_I.branch[3].block[3].um_I.iw[4] ;
 wire \top_I.branch[3].block[3].um_I.iw[5] ;
 wire \top_I.branch[3].block[3].um_I.iw[6] ;
 wire \top_I.branch[3].block[3].um_I.iw[7] ;
 wire \top_I.branch[3].block[3].um_I.iw[8] ;
 wire \top_I.branch[3].block[3].um_I.iw[9] ;
 wire \top_I.branch[3].block[3].um_I.k_zero ;
 wire \top_I.branch[3].block[3].um_I.pg_vdd ;
 wire \top_I.branch[3].block[4].um_I.ana[0] ;
 wire \top_I.branch[3].block[4].um_I.ana[1] ;
 wire \top_I.branch[3].block[4].um_I.ana[2] ;
 wire \top_I.branch[3].block[4].um_I.ana[3] ;
 wire \top_I.branch[3].block[4].um_I.ana[4] ;
 wire \top_I.branch[3].block[4].um_I.ana[5] ;
 wire \top_I.branch[3].block[4].um_I.ana[6] ;
 wire \top_I.branch[3].block[4].um_I.ana[7] ;
 wire \top_I.branch[3].block[4].um_I.clk ;
 wire \top_I.branch[3].block[4].um_I.ena ;
 wire \top_I.branch[3].block[4].um_I.iw[10] ;
 wire \top_I.branch[3].block[4].um_I.iw[11] ;
 wire \top_I.branch[3].block[4].um_I.iw[12] ;
 wire \top_I.branch[3].block[4].um_I.iw[13] ;
 wire \top_I.branch[3].block[4].um_I.iw[14] ;
 wire \top_I.branch[3].block[4].um_I.iw[15] ;
 wire \top_I.branch[3].block[4].um_I.iw[16] ;
 wire \top_I.branch[3].block[4].um_I.iw[17] ;
 wire \top_I.branch[3].block[4].um_I.iw[1] ;
 wire \top_I.branch[3].block[4].um_I.iw[2] ;
 wire \top_I.branch[3].block[4].um_I.iw[3] ;
 wire \top_I.branch[3].block[4].um_I.iw[4] ;
 wire \top_I.branch[3].block[4].um_I.iw[5] ;
 wire \top_I.branch[3].block[4].um_I.iw[6] ;
 wire \top_I.branch[3].block[4].um_I.iw[7] ;
 wire \top_I.branch[3].block[4].um_I.iw[8] ;
 wire \top_I.branch[3].block[4].um_I.iw[9] ;
 wire \top_I.branch[3].block[4].um_I.k_zero ;
 wire \top_I.branch[3].block[4].um_I.pg_vdd ;
 wire \top_I.branch[3].block[5].um_I.ana[0] ;
 wire \top_I.branch[3].block[5].um_I.ana[1] ;
 wire \top_I.branch[3].block[5].um_I.ana[2] ;
 wire \top_I.branch[3].block[5].um_I.ana[3] ;
 wire \top_I.branch[3].block[5].um_I.ana[4] ;
 wire \top_I.branch[3].block[5].um_I.ana[5] ;
 wire \top_I.branch[3].block[5].um_I.ana[6] ;
 wire \top_I.branch[3].block[5].um_I.ana[7] ;
 wire \top_I.branch[3].block[5].um_I.clk ;
 wire \top_I.branch[3].block[5].um_I.ena ;
 wire \top_I.branch[3].block[5].um_I.iw[10] ;
 wire \top_I.branch[3].block[5].um_I.iw[11] ;
 wire \top_I.branch[3].block[5].um_I.iw[12] ;
 wire \top_I.branch[3].block[5].um_I.iw[13] ;
 wire \top_I.branch[3].block[5].um_I.iw[14] ;
 wire \top_I.branch[3].block[5].um_I.iw[15] ;
 wire \top_I.branch[3].block[5].um_I.iw[16] ;
 wire \top_I.branch[3].block[5].um_I.iw[17] ;
 wire \top_I.branch[3].block[5].um_I.iw[1] ;
 wire \top_I.branch[3].block[5].um_I.iw[2] ;
 wire \top_I.branch[3].block[5].um_I.iw[3] ;
 wire \top_I.branch[3].block[5].um_I.iw[4] ;
 wire \top_I.branch[3].block[5].um_I.iw[5] ;
 wire \top_I.branch[3].block[5].um_I.iw[6] ;
 wire \top_I.branch[3].block[5].um_I.iw[7] ;
 wire \top_I.branch[3].block[5].um_I.iw[8] ;
 wire \top_I.branch[3].block[5].um_I.iw[9] ;
 wire \top_I.branch[3].block[5].um_I.k_zero ;
 wire \top_I.branch[3].block[5].um_I.pg_vdd ;
 wire \top_I.branch[3].block[6].um_I.ana[0] ;
 wire \top_I.branch[3].block[6].um_I.ana[1] ;
 wire \top_I.branch[3].block[6].um_I.ana[2] ;
 wire \top_I.branch[3].block[6].um_I.ana[3] ;
 wire \top_I.branch[3].block[6].um_I.ana[4] ;
 wire \top_I.branch[3].block[6].um_I.ana[5] ;
 wire \top_I.branch[3].block[6].um_I.ana[6] ;
 wire \top_I.branch[3].block[6].um_I.ana[7] ;
 wire \top_I.branch[3].block[6].um_I.clk ;
 wire \top_I.branch[3].block[6].um_I.ena ;
 wire \top_I.branch[3].block[6].um_I.iw[10] ;
 wire \top_I.branch[3].block[6].um_I.iw[11] ;
 wire \top_I.branch[3].block[6].um_I.iw[12] ;
 wire \top_I.branch[3].block[6].um_I.iw[13] ;
 wire \top_I.branch[3].block[6].um_I.iw[14] ;
 wire \top_I.branch[3].block[6].um_I.iw[15] ;
 wire \top_I.branch[3].block[6].um_I.iw[16] ;
 wire \top_I.branch[3].block[6].um_I.iw[17] ;
 wire \top_I.branch[3].block[6].um_I.iw[1] ;
 wire \top_I.branch[3].block[6].um_I.iw[2] ;
 wire \top_I.branch[3].block[6].um_I.iw[3] ;
 wire \top_I.branch[3].block[6].um_I.iw[4] ;
 wire \top_I.branch[3].block[6].um_I.iw[5] ;
 wire \top_I.branch[3].block[6].um_I.iw[6] ;
 wire \top_I.branch[3].block[6].um_I.iw[7] ;
 wire \top_I.branch[3].block[6].um_I.iw[8] ;
 wire \top_I.branch[3].block[6].um_I.iw[9] ;
 wire \top_I.branch[3].block[6].um_I.k_zero ;
 wire \top_I.branch[3].block[6].um_I.pg_vdd ;
 wire \top_I.branch[3].block[7].um_I.ana[0] ;
 wire \top_I.branch[3].block[7].um_I.ana[1] ;
 wire \top_I.branch[3].block[7].um_I.ana[2] ;
 wire \top_I.branch[3].block[7].um_I.ana[3] ;
 wire \top_I.branch[3].block[7].um_I.ana[4] ;
 wire \top_I.branch[3].block[7].um_I.ana[5] ;
 wire \top_I.branch[3].block[7].um_I.ana[6] ;
 wire \top_I.branch[3].block[7].um_I.ana[7] ;
 wire \top_I.branch[3].block[7].um_I.clk ;
 wire \top_I.branch[3].block[7].um_I.ena ;
 wire \top_I.branch[3].block[7].um_I.iw[10] ;
 wire \top_I.branch[3].block[7].um_I.iw[11] ;
 wire \top_I.branch[3].block[7].um_I.iw[12] ;
 wire \top_I.branch[3].block[7].um_I.iw[13] ;
 wire \top_I.branch[3].block[7].um_I.iw[14] ;
 wire \top_I.branch[3].block[7].um_I.iw[15] ;
 wire \top_I.branch[3].block[7].um_I.iw[16] ;
 wire \top_I.branch[3].block[7].um_I.iw[17] ;
 wire \top_I.branch[3].block[7].um_I.iw[1] ;
 wire \top_I.branch[3].block[7].um_I.iw[2] ;
 wire \top_I.branch[3].block[7].um_I.iw[3] ;
 wire \top_I.branch[3].block[7].um_I.iw[4] ;
 wire \top_I.branch[3].block[7].um_I.iw[5] ;
 wire \top_I.branch[3].block[7].um_I.iw[6] ;
 wire \top_I.branch[3].block[7].um_I.iw[7] ;
 wire \top_I.branch[3].block[7].um_I.iw[8] ;
 wire \top_I.branch[3].block[7].um_I.iw[9] ;
 wire \top_I.branch[3].block[7].um_I.k_zero ;
 wire \top_I.branch[3].block[7].um_I.pg_vdd ;
 wire \top_I.branch[3].block[8].um_I.ana[0] ;
 wire \top_I.branch[3].block[8].um_I.ana[1] ;
 wire \top_I.branch[3].block[8].um_I.ana[2] ;
 wire \top_I.branch[3].block[8].um_I.ana[3] ;
 wire \top_I.branch[3].block[8].um_I.ana[4] ;
 wire \top_I.branch[3].block[8].um_I.ana[5] ;
 wire \top_I.branch[3].block[8].um_I.ana[6] ;
 wire \top_I.branch[3].block[8].um_I.ana[7] ;
 wire \top_I.branch[3].block[8].um_I.clk ;
 wire \top_I.branch[3].block[8].um_I.ena ;
 wire \top_I.branch[3].block[8].um_I.iw[10] ;
 wire \top_I.branch[3].block[8].um_I.iw[11] ;
 wire \top_I.branch[3].block[8].um_I.iw[12] ;
 wire \top_I.branch[3].block[8].um_I.iw[13] ;
 wire \top_I.branch[3].block[8].um_I.iw[14] ;
 wire \top_I.branch[3].block[8].um_I.iw[15] ;
 wire \top_I.branch[3].block[8].um_I.iw[16] ;
 wire \top_I.branch[3].block[8].um_I.iw[17] ;
 wire \top_I.branch[3].block[8].um_I.iw[1] ;
 wire \top_I.branch[3].block[8].um_I.iw[2] ;
 wire \top_I.branch[3].block[8].um_I.iw[3] ;
 wire \top_I.branch[3].block[8].um_I.iw[4] ;
 wire \top_I.branch[3].block[8].um_I.iw[5] ;
 wire \top_I.branch[3].block[8].um_I.iw[6] ;
 wire \top_I.branch[3].block[8].um_I.iw[7] ;
 wire \top_I.branch[3].block[8].um_I.iw[8] ;
 wire \top_I.branch[3].block[8].um_I.iw[9] ;
 wire \top_I.branch[3].block[8].um_I.k_zero ;
 wire \top_I.branch[3].block[8].um_I.pg_vdd ;
 wire \top_I.branch[3].block[9].um_I.ana[0] ;
 wire \top_I.branch[3].block[9].um_I.ana[1] ;
 wire \top_I.branch[3].block[9].um_I.ana[2] ;
 wire \top_I.branch[3].block[9].um_I.ana[3] ;
 wire \top_I.branch[3].block[9].um_I.ana[4] ;
 wire \top_I.branch[3].block[9].um_I.ana[5] ;
 wire \top_I.branch[3].block[9].um_I.ana[6] ;
 wire \top_I.branch[3].block[9].um_I.ana[7] ;
 wire \top_I.branch[3].block[9].um_I.clk ;
 wire \top_I.branch[3].block[9].um_I.ena ;
 wire \top_I.branch[3].block[9].um_I.iw[10] ;
 wire \top_I.branch[3].block[9].um_I.iw[11] ;
 wire \top_I.branch[3].block[9].um_I.iw[12] ;
 wire \top_I.branch[3].block[9].um_I.iw[13] ;
 wire \top_I.branch[3].block[9].um_I.iw[14] ;
 wire \top_I.branch[3].block[9].um_I.iw[15] ;
 wire \top_I.branch[3].block[9].um_I.iw[16] ;
 wire \top_I.branch[3].block[9].um_I.iw[17] ;
 wire \top_I.branch[3].block[9].um_I.iw[1] ;
 wire \top_I.branch[3].block[9].um_I.iw[2] ;
 wire \top_I.branch[3].block[9].um_I.iw[3] ;
 wire \top_I.branch[3].block[9].um_I.iw[4] ;
 wire \top_I.branch[3].block[9].um_I.iw[5] ;
 wire \top_I.branch[3].block[9].um_I.iw[6] ;
 wire \top_I.branch[3].block[9].um_I.iw[7] ;
 wire \top_I.branch[3].block[9].um_I.iw[8] ;
 wire \top_I.branch[3].block[9].um_I.iw[9] ;
 wire \top_I.branch[3].block[9].um_I.k_zero ;
 wire \top_I.branch[3].block[9].um_I.pg_vdd ;
 wire \top_I.branch[3].l_addr[0] ;
 wire \top_I.branch[3].l_addr[1] ;
 wire \top_I.branch[4].block[0].um_I.ana[0] ;
 wire \top_I.branch[4].block[0].um_I.ana[1] ;
 wire \top_I.branch[4].block[0].um_I.ana[2] ;
 wire \top_I.branch[4].block[0].um_I.ana[3] ;
 wire \top_I.branch[4].block[0].um_I.ana[4] ;
 wire \top_I.branch[4].block[0].um_I.ana[5] ;
 wire \top_I.branch[4].block[0].um_I.ana[6] ;
 wire \top_I.branch[4].block[0].um_I.ana[7] ;
 wire \top_I.branch[4].block[0].um_I.clk ;
 wire \top_I.branch[4].block[0].um_I.ena ;
 wire \top_I.branch[4].block[0].um_I.iw[10] ;
 wire \top_I.branch[4].block[0].um_I.iw[11] ;
 wire \top_I.branch[4].block[0].um_I.iw[12] ;
 wire \top_I.branch[4].block[0].um_I.iw[13] ;
 wire \top_I.branch[4].block[0].um_I.iw[14] ;
 wire \top_I.branch[4].block[0].um_I.iw[15] ;
 wire \top_I.branch[4].block[0].um_I.iw[16] ;
 wire \top_I.branch[4].block[0].um_I.iw[17] ;
 wire \top_I.branch[4].block[0].um_I.iw[1] ;
 wire \top_I.branch[4].block[0].um_I.iw[2] ;
 wire \top_I.branch[4].block[0].um_I.iw[3] ;
 wire \top_I.branch[4].block[0].um_I.iw[4] ;
 wire \top_I.branch[4].block[0].um_I.iw[5] ;
 wire \top_I.branch[4].block[0].um_I.iw[6] ;
 wire \top_I.branch[4].block[0].um_I.iw[7] ;
 wire \top_I.branch[4].block[0].um_I.iw[8] ;
 wire \top_I.branch[4].block[0].um_I.iw[9] ;
 wire \top_I.branch[4].block[0].um_I.k_zero ;
 wire \top_I.branch[4].block[0].um_I.pg_vdd ;
 wire \top_I.branch[4].block[10].um_I.ana[0] ;
 wire \top_I.branch[4].block[10].um_I.ana[1] ;
 wire \top_I.branch[4].block[10].um_I.ana[2] ;
 wire \top_I.branch[4].block[10].um_I.ana[3] ;
 wire \top_I.branch[4].block[10].um_I.ana[4] ;
 wire \top_I.branch[4].block[10].um_I.ana[5] ;
 wire \top_I.branch[4].block[10].um_I.ana[6] ;
 wire \top_I.branch[4].block[10].um_I.ana[7] ;
 wire \top_I.branch[4].block[10].um_I.clk ;
 wire \top_I.branch[4].block[10].um_I.ena ;
 wire \top_I.branch[4].block[10].um_I.iw[10] ;
 wire \top_I.branch[4].block[10].um_I.iw[11] ;
 wire \top_I.branch[4].block[10].um_I.iw[12] ;
 wire \top_I.branch[4].block[10].um_I.iw[13] ;
 wire \top_I.branch[4].block[10].um_I.iw[14] ;
 wire \top_I.branch[4].block[10].um_I.iw[15] ;
 wire \top_I.branch[4].block[10].um_I.iw[16] ;
 wire \top_I.branch[4].block[10].um_I.iw[17] ;
 wire \top_I.branch[4].block[10].um_I.iw[1] ;
 wire \top_I.branch[4].block[10].um_I.iw[2] ;
 wire \top_I.branch[4].block[10].um_I.iw[3] ;
 wire \top_I.branch[4].block[10].um_I.iw[4] ;
 wire \top_I.branch[4].block[10].um_I.iw[5] ;
 wire \top_I.branch[4].block[10].um_I.iw[6] ;
 wire \top_I.branch[4].block[10].um_I.iw[7] ;
 wire \top_I.branch[4].block[10].um_I.iw[8] ;
 wire \top_I.branch[4].block[10].um_I.iw[9] ;
 wire \top_I.branch[4].block[10].um_I.k_zero ;
 wire \top_I.branch[4].block[10].um_I.pg_vdd ;
 wire \top_I.branch[4].block[11].um_I.ana[0] ;
 wire \top_I.branch[4].block[11].um_I.ana[1] ;
 wire \top_I.branch[4].block[11].um_I.ana[2] ;
 wire \top_I.branch[4].block[11].um_I.ana[3] ;
 wire \top_I.branch[4].block[11].um_I.ana[4] ;
 wire \top_I.branch[4].block[11].um_I.ana[5] ;
 wire \top_I.branch[4].block[11].um_I.ana[6] ;
 wire \top_I.branch[4].block[11].um_I.ana[7] ;
 wire \top_I.branch[4].block[11].um_I.clk ;
 wire \top_I.branch[4].block[11].um_I.ena ;
 wire \top_I.branch[4].block[11].um_I.iw[10] ;
 wire \top_I.branch[4].block[11].um_I.iw[11] ;
 wire \top_I.branch[4].block[11].um_I.iw[12] ;
 wire \top_I.branch[4].block[11].um_I.iw[13] ;
 wire \top_I.branch[4].block[11].um_I.iw[14] ;
 wire \top_I.branch[4].block[11].um_I.iw[15] ;
 wire \top_I.branch[4].block[11].um_I.iw[16] ;
 wire \top_I.branch[4].block[11].um_I.iw[17] ;
 wire \top_I.branch[4].block[11].um_I.iw[1] ;
 wire \top_I.branch[4].block[11].um_I.iw[2] ;
 wire \top_I.branch[4].block[11].um_I.iw[3] ;
 wire \top_I.branch[4].block[11].um_I.iw[4] ;
 wire \top_I.branch[4].block[11].um_I.iw[5] ;
 wire \top_I.branch[4].block[11].um_I.iw[6] ;
 wire \top_I.branch[4].block[11].um_I.iw[7] ;
 wire \top_I.branch[4].block[11].um_I.iw[8] ;
 wire \top_I.branch[4].block[11].um_I.iw[9] ;
 wire \top_I.branch[4].block[11].um_I.k_zero ;
 wire \top_I.branch[4].block[11].um_I.pg_vdd ;
 wire \top_I.branch[4].block[12].um_I.ana[0] ;
 wire \top_I.branch[4].block[12].um_I.ana[1] ;
 wire \top_I.branch[4].block[12].um_I.ana[2] ;
 wire \top_I.branch[4].block[12].um_I.ana[3] ;
 wire \top_I.branch[4].block[12].um_I.ana[4] ;
 wire \top_I.branch[4].block[12].um_I.ana[5] ;
 wire \top_I.branch[4].block[12].um_I.ana[6] ;
 wire \top_I.branch[4].block[12].um_I.ana[7] ;
 wire \top_I.branch[4].block[12].um_I.clk ;
 wire \top_I.branch[4].block[12].um_I.ena ;
 wire \top_I.branch[4].block[12].um_I.iw[10] ;
 wire \top_I.branch[4].block[12].um_I.iw[11] ;
 wire \top_I.branch[4].block[12].um_I.iw[12] ;
 wire \top_I.branch[4].block[12].um_I.iw[13] ;
 wire \top_I.branch[4].block[12].um_I.iw[14] ;
 wire \top_I.branch[4].block[12].um_I.iw[15] ;
 wire \top_I.branch[4].block[12].um_I.iw[16] ;
 wire \top_I.branch[4].block[12].um_I.iw[17] ;
 wire \top_I.branch[4].block[12].um_I.iw[1] ;
 wire \top_I.branch[4].block[12].um_I.iw[2] ;
 wire \top_I.branch[4].block[12].um_I.iw[3] ;
 wire \top_I.branch[4].block[12].um_I.iw[4] ;
 wire \top_I.branch[4].block[12].um_I.iw[5] ;
 wire \top_I.branch[4].block[12].um_I.iw[6] ;
 wire \top_I.branch[4].block[12].um_I.iw[7] ;
 wire \top_I.branch[4].block[12].um_I.iw[8] ;
 wire \top_I.branch[4].block[12].um_I.iw[9] ;
 wire \top_I.branch[4].block[12].um_I.k_zero ;
 wire \top_I.branch[4].block[12].um_I.pg_vdd ;
 wire \top_I.branch[4].block[13].um_I.ana[0] ;
 wire \top_I.branch[4].block[13].um_I.ana[1] ;
 wire \top_I.branch[4].block[13].um_I.ana[2] ;
 wire \top_I.branch[4].block[13].um_I.ana[3] ;
 wire \top_I.branch[4].block[13].um_I.ana[4] ;
 wire \top_I.branch[4].block[13].um_I.ana[5] ;
 wire \top_I.branch[4].block[13].um_I.ana[6] ;
 wire \top_I.branch[4].block[13].um_I.ana[7] ;
 wire \top_I.branch[4].block[13].um_I.clk ;
 wire \top_I.branch[4].block[13].um_I.ena ;
 wire \top_I.branch[4].block[13].um_I.iw[10] ;
 wire \top_I.branch[4].block[13].um_I.iw[11] ;
 wire \top_I.branch[4].block[13].um_I.iw[12] ;
 wire \top_I.branch[4].block[13].um_I.iw[13] ;
 wire \top_I.branch[4].block[13].um_I.iw[14] ;
 wire \top_I.branch[4].block[13].um_I.iw[15] ;
 wire \top_I.branch[4].block[13].um_I.iw[16] ;
 wire \top_I.branch[4].block[13].um_I.iw[17] ;
 wire \top_I.branch[4].block[13].um_I.iw[1] ;
 wire \top_I.branch[4].block[13].um_I.iw[2] ;
 wire \top_I.branch[4].block[13].um_I.iw[3] ;
 wire \top_I.branch[4].block[13].um_I.iw[4] ;
 wire \top_I.branch[4].block[13].um_I.iw[5] ;
 wire \top_I.branch[4].block[13].um_I.iw[6] ;
 wire \top_I.branch[4].block[13].um_I.iw[7] ;
 wire \top_I.branch[4].block[13].um_I.iw[8] ;
 wire \top_I.branch[4].block[13].um_I.iw[9] ;
 wire \top_I.branch[4].block[13].um_I.k_zero ;
 wire \top_I.branch[4].block[13].um_I.pg_vdd ;
 wire \top_I.branch[4].block[14].um_I.ana[0] ;
 wire \top_I.branch[4].block[14].um_I.ana[1] ;
 wire \top_I.branch[4].block[14].um_I.ana[2] ;
 wire \top_I.branch[4].block[14].um_I.ana[3] ;
 wire \top_I.branch[4].block[14].um_I.ana[4] ;
 wire \top_I.branch[4].block[14].um_I.ana[5] ;
 wire \top_I.branch[4].block[14].um_I.ana[6] ;
 wire \top_I.branch[4].block[14].um_I.ana[7] ;
 wire \top_I.branch[4].block[14].um_I.clk ;
 wire \top_I.branch[4].block[14].um_I.ena ;
 wire \top_I.branch[4].block[14].um_I.iw[10] ;
 wire \top_I.branch[4].block[14].um_I.iw[11] ;
 wire \top_I.branch[4].block[14].um_I.iw[12] ;
 wire \top_I.branch[4].block[14].um_I.iw[13] ;
 wire \top_I.branch[4].block[14].um_I.iw[14] ;
 wire \top_I.branch[4].block[14].um_I.iw[15] ;
 wire \top_I.branch[4].block[14].um_I.iw[16] ;
 wire \top_I.branch[4].block[14].um_I.iw[17] ;
 wire \top_I.branch[4].block[14].um_I.iw[1] ;
 wire \top_I.branch[4].block[14].um_I.iw[2] ;
 wire \top_I.branch[4].block[14].um_I.iw[3] ;
 wire \top_I.branch[4].block[14].um_I.iw[4] ;
 wire \top_I.branch[4].block[14].um_I.iw[5] ;
 wire \top_I.branch[4].block[14].um_I.iw[6] ;
 wire \top_I.branch[4].block[14].um_I.iw[7] ;
 wire \top_I.branch[4].block[14].um_I.iw[8] ;
 wire \top_I.branch[4].block[14].um_I.iw[9] ;
 wire \top_I.branch[4].block[14].um_I.k_zero ;
 wire \top_I.branch[4].block[14].um_I.pg_vdd ;
 wire \top_I.branch[4].block[15].um_I.ana[0] ;
 wire \top_I.branch[4].block[15].um_I.ana[1] ;
 wire \top_I.branch[4].block[15].um_I.ana[2] ;
 wire \top_I.branch[4].block[15].um_I.ana[3] ;
 wire \top_I.branch[4].block[15].um_I.ana[4] ;
 wire \top_I.branch[4].block[15].um_I.ana[5] ;
 wire \top_I.branch[4].block[15].um_I.ana[6] ;
 wire \top_I.branch[4].block[15].um_I.ana[7] ;
 wire \top_I.branch[4].block[15].um_I.clk ;
 wire \top_I.branch[4].block[15].um_I.ena ;
 wire \top_I.branch[4].block[15].um_I.iw[10] ;
 wire \top_I.branch[4].block[15].um_I.iw[11] ;
 wire \top_I.branch[4].block[15].um_I.iw[12] ;
 wire \top_I.branch[4].block[15].um_I.iw[13] ;
 wire \top_I.branch[4].block[15].um_I.iw[14] ;
 wire \top_I.branch[4].block[15].um_I.iw[15] ;
 wire \top_I.branch[4].block[15].um_I.iw[16] ;
 wire \top_I.branch[4].block[15].um_I.iw[17] ;
 wire \top_I.branch[4].block[15].um_I.iw[1] ;
 wire \top_I.branch[4].block[15].um_I.iw[2] ;
 wire \top_I.branch[4].block[15].um_I.iw[3] ;
 wire \top_I.branch[4].block[15].um_I.iw[4] ;
 wire \top_I.branch[4].block[15].um_I.iw[5] ;
 wire \top_I.branch[4].block[15].um_I.iw[6] ;
 wire \top_I.branch[4].block[15].um_I.iw[7] ;
 wire \top_I.branch[4].block[15].um_I.iw[8] ;
 wire \top_I.branch[4].block[15].um_I.iw[9] ;
 wire \top_I.branch[4].block[15].um_I.k_zero ;
 wire \top_I.branch[4].block[15].um_I.pg_vdd ;
 wire \top_I.branch[4].block[1].um_I.ana[0] ;
 wire \top_I.branch[4].block[1].um_I.ana[1] ;
 wire \top_I.branch[4].block[1].um_I.ana[2] ;
 wire \top_I.branch[4].block[1].um_I.ana[3] ;
 wire \top_I.branch[4].block[1].um_I.ana[4] ;
 wire \top_I.branch[4].block[1].um_I.ana[5] ;
 wire \top_I.branch[4].block[1].um_I.ana[6] ;
 wire \top_I.branch[4].block[1].um_I.ana[7] ;
 wire \top_I.branch[4].block[1].um_I.clk ;
 wire \top_I.branch[4].block[1].um_I.ena ;
 wire \top_I.branch[4].block[1].um_I.iw[10] ;
 wire \top_I.branch[4].block[1].um_I.iw[11] ;
 wire \top_I.branch[4].block[1].um_I.iw[12] ;
 wire \top_I.branch[4].block[1].um_I.iw[13] ;
 wire \top_I.branch[4].block[1].um_I.iw[14] ;
 wire \top_I.branch[4].block[1].um_I.iw[15] ;
 wire \top_I.branch[4].block[1].um_I.iw[16] ;
 wire \top_I.branch[4].block[1].um_I.iw[17] ;
 wire \top_I.branch[4].block[1].um_I.iw[1] ;
 wire \top_I.branch[4].block[1].um_I.iw[2] ;
 wire \top_I.branch[4].block[1].um_I.iw[3] ;
 wire \top_I.branch[4].block[1].um_I.iw[4] ;
 wire \top_I.branch[4].block[1].um_I.iw[5] ;
 wire \top_I.branch[4].block[1].um_I.iw[6] ;
 wire \top_I.branch[4].block[1].um_I.iw[7] ;
 wire \top_I.branch[4].block[1].um_I.iw[8] ;
 wire \top_I.branch[4].block[1].um_I.iw[9] ;
 wire \top_I.branch[4].block[1].um_I.k_zero ;
 wire \top_I.branch[4].block[1].um_I.pg_vdd ;
 wire \top_I.branch[4].block[2].um_I.ana[0] ;
 wire \top_I.branch[4].block[2].um_I.ana[1] ;
 wire \top_I.branch[4].block[2].um_I.ana[2] ;
 wire \top_I.branch[4].block[2].um_I.ana[3] ;
 wire \top_I.branch[4].block[2].um_I.ana[4] ;
 wire \top_I.branch[4].block[2].um_I.ana[5] ;
 wire \top_I.branch[4].block[2].um_I.ana[6] ;
 wire \top_I.branch[4].block[2].um_I.ana[7] ;
 wire \top_I.branch[4].block[2].um_I.clk ;
 wire \top_I.branch[4].block[2].um_I.ena ;
 wire \top_I.branch[4].block[2].um_I.iw[10] ;
 wire \top_I.branch[4].block[2].um_I.iw[11] ;
 wire \top_I.branch[4].block[2].um_I.iw[12] ;
 wire \top_I.branch[4].block[2].um_I.iw[13] ;
 wire \top_I.branch[4].block[2].um_I.iw[14] ;
 wire \top_I.branch[4].block[2].um_I.iw[15] ;
 wire \top_I.branch[4].block[2].um_I.iw[16] ;
 wire \top_I.branch[4].block[2].um_I.iw[17] ;
 wire \top_I.branch[4].block[2].um_I.iw[1] ;
 wire \top_I.branch[4].block[2].um_I.iw[2] ;
 wire \top_I.branch[4].block[2].um_I.iw[3] ;
 wire \top_I.branch[4].block[2].um_I.iw[4] ;
 wire \top_I.branch[4].block[2].um_I.iw[5] ;
 wire \top_I.branch[4].block[2].um_I.iw[6] ;
 wire \top_I.branch[4].block[2].um_I.iw[7] ;
 wire \top_I.branch[4].block[2].um_I.iw[8] ;
 wire \top_I.branch[4].block[2].um_I.iw[9] ;
 wire \top_I.branch[4].block[2].um_I.k_zero ;
 wire \top_I.branch[4].block[2].um_I.pg_vdd ;
 wire \top_I.branch[4].block[3].um_I.ana[0] ;
 wire \top_I.branch[4].block[3].um_I.ana[1] ;
 wire \top_I.branch[4].block[3].um_I.ana[2] ;
 wire \top_I.branch[4].block[3].um_I.ana[3] ;
 wire \top_I.branch[4].block[3].um_I.ana[4] ;
 wire \top_I.branch[4].block[3].um_I.ana[5] ;
 wire \top_I.branch[4].block[3].um_I.ana[6] ;
 wire \top_I.branch[4].block[3].um_I.ana[7] ;
 wire \top_I.branch[4].block[3].um_I.clk ;
 wire \top_I.branch[4].block[3].um_I.ena ;
 wire \top_I.branch[4].block[3].um_I.iw[10] ;
 wire \top_I.branch[4].block[3].um_I.iw[11] ;
 wire \top_I.branch[4].block[3].um_I.iw[12] ;
 wire \top_I.branch[4].block[3].um_I.iw[13] ;
 wire \top_I.branch[4].block[3].um_I.iw[14] ;
 wire \top_I.branch[4].block[3].um_I.iw[15] ;
 wire \top_I.branch[4].block[3].um_I.iw[16] ;
 wire \top_I.branch[4].block[3].um_I.iw[17] ;
 wire \top_I.branch[4].block[3].um_I.iw[1] ;
 wire \top_I.branch[4].block[3].um_I.iw[2] ;
 wire \top_I.branch[4].block[3].um_I.iw[3] ;
 wire \top_I.branch[4].block[3].um_I.iw[4] ;
 wire \top_I.branch[4].block[3].um_I.iw[5] ;
 wire \top_I.branch[4].block[3].um_I.iw[6] ;
 wire \top_I.branch[4].block[3].um_I.iw[7] ;
 wire \top_I.branch[4].block[3].um_I.iw[8] ;
 wire \top_I.branch[4].block[3].um_I.iw[9] ;
 wire \top_I.branch[4].block[3].um_I.k_zero ;
 wire \top_I.branch[4].block[3].um_I.pg_vdd ;
 wire \top_I.branch[4].block[4].um_I.ana[0] ;
 wire \top_I.branch[4].block[4].um_I.ana[1] ;
 wire \top_I.branch[4].block[4].um_I.ana[2] ;
 wire \top_I.branch[4].block[4].um_I.ana[3] ;
 wire \top_I.branch[4].block[4].um_I.ana[4] ;
 wire \top_I.branch[4].block[4].um_I.ana[5] ;
 wire \top_I.branch[4].block[4].um_I.ana[6] ;
 wire \top_I.branch[4].block[4].um_I.ana[7] ;
 wire \top_I.branch[4].block[4].um_I.clk ;
 wire \top_I.branch[4].block[4].um_I.ena ;
 wire \top_I.branch[4].block[4].um_I.iw[10] ;
 wire \top_I.branch[4].block[4].um_I.iw[11] ;
 wire \top_I.branch[4].block[4].um_I.iw[12] ;
 wire \top_I.branch[4].block[4].um_I.iw[13] ;
 wire \top_I.branch[4].block[4].um_I.iw[14] ;
 wire \top_I.branch[4].block[4].um_I.iw[15] ;
 wire \top_I.branch[4].block[4].um_I.iw[16] ;
 wire \top_I.branch[4].block[4].um_I.iw[17] ;
 wire \top_I.branch[4].block[4].um_I.iw[1] ;
 wire \top_I.branch[4].block[4].um_I.iw[2] ;
 wire \top_I.branch[4].block[4].um_I.iw[3] ;
 wire \top_I.branch[4].block[4].um_I.iw[4] ;
 wire \top_I.branch[4].block[4].um_I.iw[5] ;
 wire \top_I.branch[4].block[4].um_I.iw[6] ;
 wire \top_I.branch[4].block[4].um_I.iw[7] ;
 wire \top_I.branch[4].block[4].um_I.iw[8] ;
 wire \top_I.branch[4].block[4].um_I.iw[9] ;
 wire \top_I.branch[4].block[4].um_I.k_zero ;
 wire \top_I.branch[4].block[4].um_I.pg_vdd ;
 wire \top_I.branch[4].block[5].um_I.ana[0] ;
 wire \top_I.branch[4].block[5].um_I.ana[1] ;
 wire \top_I.branch[4].block[5].um_I.ana[2] ;
 wire \top_I.branch[4].block[5].um_I.ana[3] ;
 wire \top_I.branch[4].block[5].um_I.ana[4] ;
 wire \top_I.branch[4].block[5].um_I.ana[5] ;
 wire \top_I.branch[4].block[5].um_I.ana[6] ;
 wire \top_I.branch[4].block[5].um_I.ana[7] ;
 wire \top_I.branch[4].block[5].um_I.clk ;
 wire \top_I.branch[4].block[5].um_I.ena ;
 wire \top_I.branch[4].block[5].um_I.iw[10] ;
 wire \top_I.branch[4].block[5].um_I.iw[11] ;
 wire \top_I.branch[4].block[5].um_I.iw[12] ;
 wire \top_I.branch[4].block[5].um_I.iw[13] ;
 wire \top_I.branch[4].block[5].um_I.iw[14] ;
 wire \top_I.branch[4].block[5].um_I.iw[15] ;
 wire \top_I.branch[4].block[5].um_I.iw[16] ;
 wire \top_I.branch[4].block[5].um_I.iw[17] ;
 wire \top_I.branch[4].block[5].um_I.iw[1] ;
 wire \top_I.branch[4].block[5].um_I.iw[2] ;
 wire \top_I.branch[4].block[5].um_I.iw[3] ;
 wire \top_I.branch[4].block[5].um_I.iw[4] ;
 wire \top_I.branch[4].block[5].um_I.iw[5] ;
 wire \top_I.branch[4].block[5].um_I.iw[6] ;
 wire \top_I.branch[4].block[5].um_I.iw[7] ;
 wire \top_I.branch[4].block[5].um_I.iw[8] ;
 wire \top_I.branch[4].block[5].um_I.iw[9] ;
 wire \top_I.branch[4].block[5].um_I.k_zero ;
 wire \top_I.branch[4].block[5].um_I.pg_vdd ;
 wire \top_I.branch[4].block[6].um_I.ana[0] ;
 wire \top_I.branch[4].block[6].um_I.ana[1] ;
 wire \top_I.branch[4].block[6].um_I.ana[2] ;
 wire \top_I.branch[4].block[6].um_I.ana[3] ;
 wire \top_I.branch[4].block[6].um_I.ana[4] ;
 wire \top_I.branch[4].block[6].um_I.ana[5] ;
 wire \top_I.branch[4].block[6].um_I.ana[6] ;
 wire \top_I.branch[4].block[6].um_I.ana[7] ;
 wire \top_I.branch[4].block[6].um_I.clk ;
 wire \top_I.branch[4].block[6].um_I.ena ;
 wire \top_I.branch[4].block[6].um_I.iw[10] ;
 wire \top_I.branch[4].block[6].um_I.iw[11] ;
 wire \top_I.branch[4].block[6].um_I.iw[12] ;
 wire \top_I.branch[4].block[6].um_I.iw[13] ;
 wire \top_I.branch[4].block[6].um_I.iw[14] ;
 wire \top_I.branch[4].block[6].um_I.iw[15] ;
 wire \top_I.branch[4].block[6].um_I.iw[16] ;
 wire \top_I.branch[4].block[6].um_I.iw[17] ;
 wire \top_I.branch[4].block[6].um_I.iw[1] ;
 wire \top_I.branch[4].block[6].um_I.iw[2] ;
 wire \top_I.branch[4].block[6].um_I.iw[3] ;
 wire \top_I.branch[4].block[6].um_I.iw[4] ;
 wire \top_I.branch[4].block[6].um_I.iw[5] ;
 wire \top_I.branch[4].block[6].um_I.iw[6] ;
 wire \top_I.branch[4].block[6].um_I.iw[7] ;
 wire \top_I.branch[4].block[6].um_I.iw[8] ;
 wire \top_I.branch[4].block[6].um_I.iw[9] ;
 wire \top_I.branch[4].block[6].um_I.k_zero ;
 wire \top_I.branch[4].block[6].um_I.pg_vdd ;
 wire \top_I.branch[4].block[7].um_I.ana[0] ;
 wire \top_I.branch[4].block[7].um_I.ana[1] ;
 wire \top_I.branch[4].block[7].um_I.ana[2] ;
 wire \top_I.branch[4].block[7].um_I.ana[3] ;
 wire \top_I.branch[4].block[7].um_I.ana[4] ;
 wire \top_I.branch[4].block[7].um_I.ana[5] ;
 wire \top_I.branch[4].block[7].um_I.ana[6] ;
 wire \top_I.branch[4].block[7].um_I.ana[7] ;
 wire \top_I.branch[4].block[7].um_I.clk ;
 wire \top_I.branch[4].block[7].um_I.ena ;
 wire \top_I.branch[4].block[7].um_I.iw[10] ;
 wire \top_I.branch[4].block[7].um_I.iw[11] ;
 wire \top_I.branch[4].block[7].um_I.iw[12] ;
 wire \top_I.branch[4].block[7].um_I.iw[13] ;
 wire \top_I.branch[4].block[7].um_I.iw[14] ;
 wire \top_I.branch[4].block[7].um_I.iw[15] ;
 wire \top_I.branch[4].block[7].um_I.iw[16] ;
 wire \top_I.branch[4].block[7].um_I.iw[17] ;
 wire \top_I.branch[4].block[7].um_I.iw[1] ;
 wire \top_I.branch[4].block[7].um_I.iw[2] ;
 wire \top_I.branch[4].block[7].um_I.iw[3] ;
 wire \top_I.branch[4].block[7].um_I.iw[4] ;
 wire \top_I.branch[4].block[7].um_I.iw[5] ;
 wire \top_I.branch[4].block[7].um_I.iw[6] ;
 wire \top_I.branch[4].block[7].um_I.iw[7] ;
 wire \top_I.branch[4].block[7].um_I.iw[8] ;
 wire \top_I.branch[4].block[7].um_I.iw[9] ;
 wire \top_I.branch[4].block[7].um_I.k_zero ;
 wire \top_I.branch[4].block[7].um_I.pg_vdd ;
 wire \top_I.branch[4].block[8].um_I.ana[0] ;
 wire \top_I.branch[4].block[8].um_I.ana[1] ;
 wire \top_I.branch[4].block[8].um_I.ana[2] ;
 wire \top_I.branch[4].block[8].um_I.ana[3] ;
 wire \top_I.branch[4].block[8].um_I.ana[4] ;
 wire \top_I.branch[4].block[8].um_I.ana[5] ;
 wire \top_I.branch[4].block[8].um_I.ana[6] ;
 wire \top_I.branch[4].block[8].um_I.ana[7] ;
 wire \top_I.branch[4].block[8].um_I.clk ;
 wire \top_I.branch[4].block[8].um_I.ena ;
 wire \top_I.branch[4].block[8].um_I.iw[10] ;
 wire \top_I.branch[4].block[8].um_I.iw[11] ;
 wire \top_I.branch[4].block[8].um_I.iw[12] ;
 wire \top_I.branch[4].block[8].um_I.iw[13] ;
 wire \top_I.branch[4].block[8].um_I.iw[14] ;
 wire \top_I.branch[4].block[8].um_I.iw[15] ;
 wire \top_I.branch[4].block[8].um_I.iw[16] ;
 wire \top_I.branch[4].block[8].um_I.iw[17] ;
 wire \top_I.branch[4].block[8].um_I.iw[1] ;
 wire \top_I.branch[4].block[8].um_I.iw[2] ;
 wire \top_I.branch[4].block[8].um_I.iw[3] ;
 wire \top_I.branch[4].block[8].um_I.iw[4] ;
 wire \top_I.branch[4].block[8].um_I.iw[5] ;
 wire \top_I.branch[4].block[8].um_I.iw[6] ;
 wire \top_I.branch[4].block[8].um_I.iw[7] ;
 wire \top_I.branch[4].block[8].um_I.iw[8] ;
 wire \top_I.branch[4].block[8].um_I.iw[9] ;
 wire \top_I.branch[4].block[8].um_I.k_zero ;
 wire \top_I.branch[4].block[8].um_I.pg_vdd ;
 wire \top_I.branch[4].block[9].um_I.ana[0] ;
 wire \top_I.branch[4].block[9].um_I.ana[1] ;
 wire \top_I.branch[4].block[9].um_I.ana[2] ;
 wire \top_I.branch[4].block[9].um_I.ana[3] ;
 wire \top_I.branch[4].block[9].um_I.ana[4] ;
 wire \top_I.branch[4].block[9].um_I.ana[5] ;
 wire \top_I.branch[4].block[9].um_I.ana[6] ;
 wire \top_I.branch[4].block[9].um_I.ana[7] ;
 wire \top_I.branch[4].block[9].um_I.clk ;
 wire \top_I.branch[4].block[9].um_I.ena ;
 wire \top_I.branch[4].block[9].um_I.iw[10] ;
 wire \top_I.branch[4].block[9].um_I.iw[11] ;
 wire \top_I.branch[4].block[9].um_I.iw[12] ;
 wire \top_I.branch[4].block[9].um_I.iw[13] ;
 wire \top_I.branch[4].block[9].um_I.iw[14] ;
 wire \top_I.branch[4].block[9].um_I.iw[15] ;
 wire \top_I.branch[4].block[9].um_I.iw[16] ;
 wire \top_I.branch[4].block[9].um_I.iw[17] ;
 wire \top_I.branch[4].block[9].um_I.iw[1] ;
 wire \top_I.branch[4].block[9].um_I.iw[2] ;
 wire \top_I.branch[4].block[9].um_I.iw[3] ;
 wire \top_I.branch[4].block[9].um_I.iw[4] ;
 wire \top_I.branch[4].block[9].um_I.iw[5] ;
 wire \top_I.branch[4].block[9].um_I.iw[6] ;
 wire \top_I.branch[4].block[9].um_I.iw[7] ;
 wire \top_I.branch[4].block[9].um_I.iw[8] ;
 wire \top_I.branch[4].block[9].um_I.iw[9] ;
 wire \top_I.branch[4].block[9].um_I.k_zero ;
 wire \top_I.branch[4].block[9].um_I.pg_vdd ;
 wire \top_I.branch[4].l_addr[0] ;
 wire \top_I.branch[4].l_addr[1] ;
 wire \top_I.branch[5].block[0].um_I.ana[0] ;
 wire \top_I.branch[5].block[0].um_I.ana[1] ;
 wire \top_I.branch[5].block[0].um_I.ana[2] ;
 wire \top_I.branch[5].block[0].um_I.ana[3] ;
 wire \top_I.branch[5].block[0].um_I.ana[4] ;
 wire \top_I.branch[5].block[0].um_I.ana[5] ;
 wire \top_I.branch[5].block[0].um_I.ana[6] ;
 wire \top_I.branch[5].block[0].um_I.ana[7] ;
 wire \top_I.branch[5].block[0].um_I.clk ;
 wire \top_I.branch[5].block[0].um_I.ena ;
 wire \top_I.branch[5].block[0].um_I.iw[10] ;
 wire \top_I.branch[5].block[0].um_I.iw[11] ;
 wire \top_I.branch[5].block[0].um_I.iw[12] ;
 wire \top_I.branch[5].block[0].um_I.iw[13] ;
 wire \top_I.branch[5].block[0].um_I.iw[14] ;
 wire \top_I.branch[5].block[0].um_I.iw[15] ;
 wire \top_I.branch[5].block[0].um_I.iw[16] ;
 wire \top_I.branch[5].block[0].um_I.iw[17] ;
 wire \top_I.branch[5].block[0].um_I.iw[1] ;
 wire \top_I.branch[5].block[0].um_I.iw[2] ;
 wire \top_I.branch[5].block[0].um_I.iw[3] ;
 wire \top_I.branch[5].block[0].um_I.iw[4] ;
 wire \top_I.branch[5].block[0].um_I.iw[5] ;
 wire \top_I.branch[5].block[0].um_I.iw[6] ;
 wire \top_I.branch[5].block[0].um_I.iw[7] ;
 wire \top_I.branch[5].block[0].um_I.iw[8] ;
 wire \top_I.branch[5].block[0].um_I.iw[9] ;
 wire \top_I.branch[5].block[0].um_I.k_zero ;
 wire \top_I.branch[5].block[0].um_I.pg_vdd ;
 wire \top_I.branch[5].block[10].um_I.ana[0] ;
 wire \top_I.branch[5].block[10].um_I.ana[1] ;
 wire \top_I.branch[5].block[10].um_I.ana[2] ;
 wire \top_I.branch[5].block[10].um_I.ana[3] ;
 wire \top_I.branch[5].block[10].um_I.ana[4] ;
 wire \top_I.branch[5].block[10].um_I.ana[5] ;
 wire \top_I.branch[5].block[10].um_I.ana[6] ;
 wire \top_I.branch[5].block[10].um_I.ana[7] ;
 wire \top_I.branch[5].block[10].um_I.clk ;
 wire \top_I.branch[5].block[10].um_I.ena ;
 wire \top_I.branch[5].block[10].um_I.iw[10] ;
 wire \top_I.branch[5].block[10].um_I.iw[11] ;
 wire \top_I.branch[5].block[10].um_I.iw[12] ;
 wire \top_I.branch[5].block[10].um_I.iw[13] ;
 wire \top_I.branch[5].block[10].um_I.iw[14] ;
 wire \top_I.branch[5].block[10].um_I.iw[15] ;
 wire \top_I.branch[5].block[10].um_I.iw[16] ;
 wire \top_I.branch[5].block[10].um_I.iw[17] ;
 wire \top_I.branch[5].block[10].um_I.iw[1] ;
 wire \top_I.branch[5].block[10].um_I.iw[2] ;
 wire \top_I.branch[5].block[10].um_I.iw[3] ;
 wire \top_I.branch[5].block[10].um_I.iw[4] ;
 wire \top_I.branch[5].block[10].um_I.iw[5] ;
 wire \top_I.branch[5].block[10].um_I.iw[6] ;
 wire \top_I.branch[5].block[10].um_I.iw[7] ;
 wire \top_I.branch[5].block[10].um_I.iw[8] ;
 wire \top_I.branch[5].block[10].um_I.iw[9] ;
 wire \top_I.branch[5].block[10].um_I.k_zero ;
 wire \top_I.branch[5].block[10].um_I.pg_vdd ;
 wire \top_I.branch[5].block[11].um_I.ana[0] ;
 wire \top_I.branch[5].block[11].um_I.ana[1] ;
 wire \top_I.branch[5].block[11].um_I.ana[2] ;
 wire \top_I.branch[5].block[11].um_I.ana[3] ;
 wire \top_I.branch[5].block[11].um_I.ana[4] ;
 wire \top_I.branch[5].block[11].um_I.ana[5] ;
 wire \top_I.branch[5].block[11].um_I.ana[6] ;
 wire \top_I.branch[5].block[11].um_I.ana[7] ;
 wire \top_I.branch[5].block[11].um_I.clk ;
 wire \top_I.branch[5].block[11].um_I.ena ;
 wire \top_I.branch[5].block[11].um_I.iw[10] ;
 wire \top_I.branch[5].block[11].um_I.iw[11] ;
 wire \top_I.branch[5].block[11].um_I.iw[12] ;
 wire \top_I.branch[5].block[11].um_I.iw[13] ;
 wire \top_I.branch[5].block[11].um_I.iw[14] ;
 wire \top_I.branch[5].block[11].um_I.iw[15] ;
 wire \top_I.branch[5].block[11].um_I.iw[16] ;
 wire \top_I.branch[5].block[11].um_I.iw[17] ;
 wire \top_I.branch[5].block[11].um_I.iw[1] ;
 wire \top_I.branch[5].block[11].um_I.iw[2] ;
 wire \top_I.branch[5].block[11].um_I.iw[3] ;
 wire \top_I.branch[5].block[11].um_I.iw[4] ;
 wire \top_I.branch[5].block[11].um_I.iw[5] ;
 wire \top_I.branch[5].block[11].um_I.iw[6] ;
 wire \top_I.branch[5].block[11].um_I.iw[7] ;
 wire \top_I.branch[5].block[11].um_I.iw[8] ;
 wire \top_I.branch[5].block[11].um_I.iw[9] ;
 wire \top_I.branch[5].block[11].um_I.k_zero ;
 wire \top_I.branch[5].block[11].um_I.pg_vdd ;
 wire \top_I.branch[5].block[12].um_I.ana[0] ;
 wire \top_I.branch[5].block[12].um_I.ana[1] ;
 wire \top_I.branch[5].block[12].um_I.ana[2] ;
 wire \top_I.branch[5].block[12].um_I.ana[3] ;
 wire \top_I.branch[5].block[12].um_I.ana[4] ;
 wire \top_I.branch[5].block[12].um_I.ana[5] ;
 wire \top_I.branch[5].block[12].um_I.ana[6] ;
 wire \top_I.branch[5].block[12].um_I.ana[7] ;
 wire \top_I.branch[5].block[12].um_I.clk ;
 wire \top_I.branch[5].block[12].um_I.ena ;
 wire \top_I.branch[5].block[12].um_I.iw[10] ;
 wire \top_I.branch[5].block[12].um_I.iw[11] ;
 wire \top_I.branch[5].block[12].um_I.iw[12] ;
 wire \top_I.branch[5].block[12].um_I.iw[13] ;
 wire \top_I.branch[5].block[12].um_I.iw[14] ;
 wire \top_I.branch[5].block[12].um_I.iw[15] ;
 wire \top_I.branch[5].block[12].um_I.iw[16] ;
 wire \top_I.branch[5].block[12].um_I.iw[17] ;
 wire \top_I.branch[5].block[12].um_I.iw[1] ;
 wire \top_I.branch[5].block[12].um_I.iw[2] ;
 wire \top_I.branch[5].block[12].um_I.iw[3] ;
 wire \top_I.branch[5].block[12].um_I.iw[4] ;
 wire \top_I.branch[5].block[12].um_I.iw[5] ;
 wire \top_I.branch[5].block[12].um_I.iw[6] ;
 wire \top_I.branch[5].block[12].um_I.iw[7] ;
 wire \top_I.branch[5].block[12].um_I.iw[8] ;
 wire \top_I.branch[5].block[12].um_I.iw[9] ;
 wire \top_I.branch[5].block[12].um_I.k_zero ;
 wire \top_I.branch[5].block[12].um_I.pg_vdd ;
 wire \top_I.branch[5].block[13].um_I.ana[0] ;
 wire \top_I.branch[5].block[13].um_I.ana[1] ;
 wire \top_I.branch[5].block[13].um_I.ana[2] ;
 wire \top_I.branch[5].block[13].um_I.ana[3] ;
 wire \top_I.branch[5].block[13].um_I.ana[4] ;
 wire \top_I.branch[5].block[13].um_I.ana[5] ;
 wire \top_I.branch[5].block[13].um_I.ana[6] ;
 wire \top_I.branch[5].block[13].um_I.ana[7] ;
 wire \top_I.branch[5].block[13].um_I.clk ;
 wire \top_I.branch[5].block[13].um_I.ena ;
 wire \top_I.branch[5].block[13].um_I.iw[10] ;
 wire \top_I.branch[5].block[13].um_I.iw[11] ;
 wire \top_I.branch[5].block[13].um_I.iw[12] ;
 wire \top_I.branch[5].block[13].um_I.iw[13] ;
 wire \top_I.branch[5].block[13].um_I.iw[14] ;
 wire \top_I.branch[5].block[13].um_I.iw[15] ;
 wire \top_I.branch[5].block[13].um_I.iw[16] ;
 wire \top_I.branch[5].block[13].um_I.iw[17] ;
 wire \top_I.branch[5].block[13].um_I.iw[1] ;
 wire \top_I.branch[5].block[13].um_I.iw[2] ;
 wire \top_I.branch[5].block[13].um_I.iw[3] ;
 wire \top_I.branch[5].block[13].um_I.iw[4] ;
 wire \top_I.branch[5].block[13].um_I.iw[5] ;
 wire \top_I.branch[5].block[13].um_I.iw[6] ;
 wire \top_I.branch[5].block[13].um_I.iw[7] ;
 wire \top_I.branch[5].block[13].um_I.iw[8] ;
 wire \top_I.branch[5].block[13].um_I.iw[9] ;
 wire \top_I.branch[5].block[13].um_I.k_zero ;
 wire \top_I.branch[5].block[13].um_I.pg_vdd ;
 wire \top_I.branch[5].block[14].um_I.ana[0] ;
 wire \top_I.branch[5].block[14].um_I.ana[1] ;
 wire \top_I.branch[5].block[14].um_I.ana[2] ;
 wire \top_I.branch[5].block[14].um_I.ana[3] ;
 wire \top_I.branch[5].block[14].um_I.ana[4] ;
 wire \top_I.branch[5].block[14].um_I.ana[5] ;
 wire \top_I.branch[5].block[14].um_I.ana[6] ;
 wire \top_I.branch[5].block[14].um_I.ana[7] ;
 wire \top_I.branch[5].block[14].um_I.clk ;
 wire \top_I.branch[5].block[14].um_I.ena ;
 wire \top_I.branch[5].block[14].um_I.iw[10] ;
 wire \top_I.branch[5].block[14].um_I.iw[11] ;
 wire \top_I.branch[5].block[14].um_I.iw[12] ;
 wire \top_I.branch[5].block[14].um_I.iw[13] ;
 wire \top_I.branch[5].block[14].um_I.iw[14] ;
 wire \top_I.branch[5].block[14].um_I.iw[15] ;
 wire \top_I.branch[5].block[14].um_I.iw[16] ;
 wire \top_I.branch[5].block[14].um_I.iw[17] ;
 wire \top_I.branch[5].block[14].um_I.iw[1] ;
 wire \top_I.branch[5].block[14].um_I.iw[2] ;
 wire \top_I.branch[5].block[14].um_I.iw[3] ;
 wire \top_I.branch[5].block[14].um_I.iw[4] ;
 wire \top_I.branch[5].block[14].um_I.iw[5] ;
 wire \top_I.branch[5].block[14].um_I.iw[6] ;
 wire \top_I.branch[5].block[14].um_I.iw[7] ;
 wire \top_I.branch[5].block[14].um_I.iw[8] ;
 wire \top_I.branch[5].block[14].um_I.iw[9] ;
 wire \top_I.branch[5].block[14].um_I.k_zero ;
 wire \top_I.branch[5].block[14].um_I.pg_vdd ;
 wire \top_I.branch[5].block[15].um_I.ana[0] ;
 wire \top_I.branch[5].block[15].um_I.ana[1] ;
 wire \top_I.branch[5].block[15].um_I.ana[2] ;
 wire \top_I.branch[5].block[15].um_I.ana[3] ;
 wire \top_I.branch[5].block[15].um_I.ana[4] ;
 wire \top_I.branch[5].block[15].um_I.ana[5] ;
 wire \top_I.branch[5].block[15].um_I.ana[6] ;
 wire \top_I.branch[5].block[15].um_I.ana[7] ;
 wire \top_I.branch[5].block[15].um_I.clk ;
 wire \top_I.branch[5].block[15].um_I.ena ;
 wire \top_I.branch[5].block[15].um_I.iw[10] ;
 wire \top_I.branch[5].block[15].um_I.iw[11] ;
 wire \top_I.branch[5].block[15].um_I.iw[12] ;
 wire \top_I.branch[5].block[15].um_I.iw[13] ;
 wire \top_I.branch[5].block[15].um_I.iw[14] ;
 wire \top_I.branch[5].block[15].um_I.iw[15] ;
 wire \top_I.branch[5].block[15].um_I.iw[16] ;
 wire \top_I.branch[5].block[15].um_I.iw[17] ;
 wire \top_I.branch[5].block[15].um_I.iw[1] ;
 wire \top_I.branch[5].block[15].um_I.iw[2] ;
 wire \top_I.branch[5].block[15].um_I.iw[3] ;
 wire \top_I.branch[5].block[15].um_I.iw[4] ;
 wire \top_I.branch[5].block[15].um_I.iw[5] ;
 wire \top_I.branch[5].block[15].um_I.iw[6] ;
 wire \top_I.branch[5].block[15].um_I.iw[7] ;
 wire \top_I.branch[5].block[15].um_I.iw[8] ;
 wire \top_I.branch[5].block[15].um_I.iw[9] ;
 wire \top_I.branch[5].block[15].um_I.k_zero ;
 wire \top_I.branch[5].block[15].um_I.pg_vdd ;
 wire \top_I.branch[5].block[1].um_I.ana[0] ;
 wire \top_I.branch[5].block[1].um_I.ana[1] ;
 wire \top_I.branch[5].block[1].um_I.ana[2] ;
 wire \top_I.branch[5].block[1].um_I.ana[3] ;
 wire \top_I.branch[5].block[1].um_I.ana[4] ;
 wire \top_I.branch[5].block[1].um_I.ana[5] ;
 wire \top_I.branch[5].block[1].um_I.ana[6] ;
 wire \top_I.branch[5].block[1].um_I.ana[7] ;
 wire \top_I.branch[5].block[1].um_I.clk ;
 wire \top_I.branch[5].block[1].um_I.ena ;
 wire \top_I.branch[5].block[1].um_I.iw[10] ;
 wire \top_I.branch[5].block[1].um_I.iw[11] ;
 wire \top_I.branch[5].block[1].um_I.iw[12] ;
 wire \top_I.branch[5].block[1].um_I.iw[13] ;
 wire \top_I.branch[5].block[1].um_I.iw[14] ;
 wire \top_I.branch[5].block[1].um_I.iw[15] ;
 wire \top_I.branch[5].block[1].um_I.iw[16] ;
 wire \top_I.branch[5].block[1].um_I.iw[17] ;
 wire \top_I.branch[5].block[1].um_I.iw[1] ;
 wire \top_I.branch[5].block[1].um_I.iw[2] ;
 wire \top_I.branch[5].block[1].um_I.iw[3] ;
 wire \top_I.branch[5].block[1].um_I.iw[4] ;
 wire \top_I.branch[5].block[1].um_I.iw[5] ;
 wire \top_I.branch[5].block[1].um_I.iw[6] ;
 wire \top_I.branch[5].block[1].um_I.iw[7] ;
 wire \top_I.branch[5].block[1].um_I.iw[8] ;
 wire \top_I.branch[5].block[1].um_I.iw[9] ;
 wire \top_I.branch[5].block[1].um_I.k_zero ;
 wire \top_I.branch[5].block[1].um_I.pg_vdd ;
 wire \top_I.branch[5].block[2].um_I.ana[0] ;
 wire \top_I.branch[5].block[2].um_I.ana[1] ;
 wire \top_I.branch[5].block[2].um_I.ana[2] ;
 wire \top_I.branch[5].block[2].um_I.ana[3] ;
 wire \top_I.branch[5].block[2].um_I.ana[4] ;
 wire \top_I.branch[5].block[2].um_I.ana[5] ;
 wire \top_I.branch[5].block[2].um_I.ana[6] ;
 wire \top_I.branch[5].block[2].um_I.ana[7] ;
 wire \top_I.branch[5].block[2].um_I.clk ;
 wire \top_I.branch[5].block[2].um_I.ena ;
 wire \top_I.branch[5].block[2].um_I.iw[10] ;
 wire \top_I.branch[5].block[2].um_I.iw[11] ;
 wire \top_I.branch[5].block[2].um_I.iw[12] ;
 wire \top_I.branch[5].block[2].um_I.iw[13] ;
 wire \top_I.branch[5].block[2].um_I.iw[14] ;
 wire \top_I.branch[5].block[2].um_I.iw[15] ;
 wire \top_I.branch[5].block[2].um_I.iw[16] ;
 wire \top_I.branch[5].block[2].um_I.iw[17] ;
 wire \top_I.branch[5].block[2].um_I.iw[1] ;
 wire \top_I.branch[5].block[2].um_I.iw[2] ;
 wire \top_I.branch[5].block[2].um_I.iw[3] ;
 wire \top_I.branch[5].block[2].um_I.iw[4] ;
 wire \top_I.branch[5].block[2].um_I.iw[5] ;
 wire \top_I.branch[5].block[2].um_I.iw[6] ;
 wire \top_I.branch[5].block[2].um_I.iw[7] ;
 wire \top_I.branch[5].block[2].um_I.iw[8] ;
 wire \top_I.branch[5].block[2].um_I.iw[9] ;
 wire \top_I.branch[5].block[2].um_I.k_zero ;
 wire \top_I.branch[5].block[2].um_I.pg_vdd ;
 wire \top_I.branch[5].block[3].um_I.ana[0] ;
 wire \top_I.branch[5].block[3].um_I.ana[1] ;
 wire \top_I.branch[5].block[3].um_I.ana[2] ;
 wire \top_I.branch[5].block[3].um_I.ana[3] ;
 wire \top_I.branch[5].block[3].um_I.ana[4] ;
 wire \top_I.branch[5].block[3].um_I.ana[5] ;
 wire \top_I.branch[5].block[3].um_I.ana[6] ;
 wire \top_I.branch[5].block[3].um_I.ana[7] ;
 wire \top_I.branch[5].block[3].um_I.clk ;
 wire \top_I.branch[5].block[3].um_I.ena ;
 wire \top_I.branch[5].block[3].um_I.iw[10] ;
 wire \top_I.branch[5].block[3].um_I.iw[11] ;
 wire \top_I.branch[5].block[3].um_I.iw[12] ;
 wire \top_I.branch[5].block[3].um_I.iw[13] ;
 wire \top_I.branch[5].block[3].um_I.iw[14] ;
 wire \top_I.branch[5].block[3].um_I.iw[15] ;
 wire \top_I.branch[5].block[3].um_I.iw[16] ;
 wire \top_I.branch[5].block[3].um_I.iw[17] ;
 wire \top_I.branch[5].block[3].um_I.iw[1] ;
 wire \top_I.branch[5].block[3].um_I.iw[2] ;
 wire \top_I.branch[5].block[3].um_I.iw[3] ;
 wire \top_I.branch[5].block[3].um_I.iw[4] ;
 wire \top_I.branch[5].block[3].um_I.iw[5] ;
 wire \top_I.branch[5].block[3].um_I.iw[6] ;
 wire \top_I.branch[5].block[3].um_I.iw[7] ;
 wire \top_I.branch[5].block[3].um_I.iw[8] ;
 wire \top_I.branch[5].block[3].um_I.iw[9] ;
 wire \top_I.branch[5].block[3].um_I.k_zero ;
 wire \top_I.branch[5].block[3].um_I.pg_vdd ;
 wire \top_I.branch[5].block[4].um_I.ana[0] ;
 wire \top_I.branch[5].block[4].um_I.ana[1] ;
 wire \top_I.branch[5].block[4].um_I.ana[2] ;
 wire \top_I.branch[5].block[4].um_I.ana[3] ;
 wire \top_I.branch[5].block[4].um_I.ana[4] ;
 wire \top_I.branch[5].block[4].um_I.ana[5] ;
 wire \top_I.branch[5].block[4].um_I.ana[6] ;
 wire \top_I.branch[5].block[4].um_I.ana[7] ;
 wire \top_I.branch[5].block[4].um_I.clk ;
 wire \top_I.branch[5].block[4].um_I.ena ;
 wire \top_I.branch[5].block[4].um_I.iw[10] ;
 wire \top_I.branch[5].block[4].um_I.iw[11] ;
 wire \top_I.branch[5].block[4].um_I.iw[12] ;
 wire \top_I.branch[5].block[4].um_I.iw[13] ;
 wire \top_I.branch[5].block[4].um_I.iw[14] ;
 wire \top_I.branch[5].block[4].um_I.iw[15] ;
 wire \top_I.branch[5].block[4].um_I.iw[16] ;
 wire \top_I.branch[5].block[4].um_I.iw[17] ;
 wire \top_I.branch[5].block[4].um_I.iw[1] ;
 wire \top_I.branch[5].block[4].um_I.iw[2] ;
 wire \top_I.branch[5].block[4].um_I.iw[3] ;
 wire \top_I.branch[5].block[4].um_I.iw[4] ;
 wire \top_I.branch[5].block[4].um_I.iw[5] ;
 wire \top_I.branch[5].block[4].um_I.iw[6] ;
 wire \top_I.branch[5].block[4].um_I.iw[7] ;
 wire \top_I.branch[5].block[4].um_I.iw[8] ;
 wire \top_I.branch[5].block[4].um_I.iw[9] ;
 wire \top_I.branch[5].block[4].um_I.k_zero ;
 wire \top_I.branch[5].block[4].um_I.pg_vdd ;
 wire \top_I.branch[5].block[5].um_I.ana[0] ;
 wire \top_I.branch[5].block[5].um_I.ana[1] ;
 wire \top_I.branch[5].block[5].um_I.ana[2] ;
 wire \top_I.branch[5].block[5].um_I.ana[3] ;
 wire \top_I.branch[5].block[5].um_I.ana[4] ;
 wire \top_I.branch[5].block[5].um_I.ana[5] ;
 wire \top_I.branch[5].block[5].um_I.ana[6] ;
 wire \top_I.branch[5].block[5].um_I.ana[7] ;
 wire \top_I.branch[5].block[5].um_I.clk ;
 wire \top_I.branch[5].block[5].um_I.ena ;
 wire \top_I.branch[5].block[5].um_I.iw[10] ;
 wire \top_I.branch[5].block[5].um_I.iw[11] ;
 wire \top_I.branch[5].block[5].um_I.iw[12] ;
 wire \top_I.branch[5].block[5].um_I.iw[13] ;
 wire \top_I.branch[5].block[5].um_I.iw[14] ;
 wire \top_I.branch[5].block[5].um_I.iw[15] ;
 wire \top_I.branch[5].block[5].um_I.iw[16] ;
 wire \top_I.branch[5].block[5].um_I.iw[17] ;
 wire \top_I.branch[5].block[5].um_I.iw[1] ;
 wire \top_I.branch[5].block[5].um_I.iw[2] ;
 wire \top_I.branch[5].block[5].um_I.iw[3] ;
 wire \top_I.branch[5].block[5].um_I.iw[4] ;
 wire \top_I.branch[5].block[5].um_I.iw[5] ;
 wire \top_I.branch[5].block[5].um_I.iw[6] ;
 wire \top_I.branch[5].block[5].um_I.iw[7] ;
 wire \top_I.branch[5].block[5].um_I.iw[8] ;
 wire \top_I.branch[5].block[5].um_I.iw[9] ;
 wire \top_I.branch[5].block[5].um_I.k_zero ;
 wire \top_I.branch[5].block[5].um_I.pg_vdd ;
 wire \top_I.branch[5].block[6].um_I.ana[0] ;
 wire \top_I.branch[5].block[6].um_I.ana[1] ;
 wire \top_I.branch[5].block[6].um_I.ana[2] ;
 wire \top_I.branch[5].block[6].um_I.ana[3] ;
 wire \top_I.branch[5].block[6].um_I.ana[4] ;
 wire \top_I.branch[5].block[6].um_I.ana[5] ;
 wire \top_I.branch[5].block[6].um_I.ana[6] ;
 wire \top_I.branch[5].block[6].um_I.ana[7] ;
 wire \top_I.branch[5].block[6].um_I.clk ;
 wire \top_I.branch[5].block[6].um_I.ena ;
 wire \top_I.branch[5].block[6].um_I.iw[10] ;
 wire \top_I.branch[5].block[6].um_I.iw[11] ;
 wire \top_I.branch[5].block[6].um_I.iw[12] ;
 wire \top_I.branch[5].block[6].um_I.iw[13] ;
 wire \top_I.branch[5].block[6].um_I.iw[14] ;
 wire \top_I.branch[5].block[6].um_I.iw[15] ;
 wire \top_I.branch[5].block[6].um_I.iw[16] ;
 wire \top_I.branch[5].block[6].um_I.iw[17] ;
 wire \top_I.branch[5].block[6].um_I.iw[1] ;
 wire \top_I.branch[5].block[6].um_I.iw[2] ;
 wire \top_I.branch[5].block[6].um_I.iw[3] ;
 wire \top_I.branch[5].block[6].um_I.iw[4] ;
 wire \top_I.branch[5].block[6].um_I.iw[5] ;
 wire \top_I.branch[5].block[6].um_I.iw[6] ;
 wire \top_I.branch[5].block[6].um_I.iw[7] ;
 wire \top_I.branch[5].block[6].um_I.iw[8] ;
 wire \top_I.branch[5].block[6].um_I.iw[9] ;
 wire \top_I.branch[5].block[6].um_I.k_zero ;
 wire \top_I.branch[5].block[6].um_I.pg_vdd ;
 wire \top_I.branch[5].block[7].um_I.ana[0] ;
 wire \top_I.branch[5].block[7].um_I.ana[1] ;
 wire \top_I.branch[5].block[7].um_I.ana[2] ;
 wire \top_I.branch[5].block[7].um_I.ana[3] ;
 wire \top_I.branch[5].block[7].um_I.ana[4] ;
 wire \top_I.branch[5].block[7].um_I.ana[5] ;
 wire \top_I.branch[5].block[7].um_I.ana[6] ;
 wire \top_I.branch[5].block[7].um_I.ana[7] ;
 wire \top_I.branch[5].block[7].um_I.clk ;
 wire \top_I.branch[5].block[7].um_I.ena ;
 wire \top_I.branch[5].block[7].um_I.iw[10] ;
 wire \top_I.branch[5].block[7].um_I.iw[11] ;
 wire \top_I.branch[5].block[7].um_I.iw[12] ;
 wire \top_I.branch[5].block[7].um_I.iw[13] ;
 wire \top_I.branch[5].block[7].um_I.iw[14] ;
 wire \top_I.branch[5].block[7].um_I.iw[15] ;
 wire \top_I.branch[5].block[7].um_I.iw[16] ;
 wire \top_I.branch[5].block[7].um_I.iw[17] ;
 wire \top_I.branch[5].block[7].um_I.iw[1] ;
 wire \top_I.branch[5].block[7].um_I.iw[2] ;
 wire \top_I.branch[5].block[7].um_I.iw[3] ;
 wire \top_I.branch[5].block[7].um_I.iw[4] ;
 wire \top_I.branch[5].block[7].um_I.iw[5] ;
 wire \top_I.branch[5].block[7].um_I.iw[6] ;
 wire \top_I.branch[5].block[7].um_I.iw[7] ;
 wire \top_I.branch[5].block[7].um_I.iw[8] ;
 wire \top_I.branch[5].block[7].um_I.iw[9] ;
 wire \top_I.branch[5].block[7].um_I.k_zero ;
 wire \top_I.branch[5].block[7].um_I.pg_vdd ;
 wire \top_I.branch[5].block[8].um_I.ana[0] ;
 wire \top_I.branch[5].block[8].um_I.ana[1] ;
 wire \top_I.branch[5].block[8].um_I.ana[2] ;
 wire \top_I.branch[5].block[8].um_I.ana[3] ;
 wire \top_I.branch[5].block[8].um_I.ana[4] ;
 wire \top_I.branch[5].block[8].um_I.ana[5] ;
 wire \top_I.branch[5].block[8].um_I.ana[6] ;
 wire \top_I.branch[5].block[8].um_I.ana[7] ;
 wire \top_I.branch[5].block[8].um_I.clk ;
 wire \top_I.branch[5].block[8].um_I.ena ;
 wire \top_I.branch[5].block[8].um_I.iw[10] ;
 wire \top_I.branch[5].block[8].um_I.iw[11] ;
 wire \top_I.branch[5].block[8].um_I.iw[12] ;
 wire \top_I.branch[5].block[8].um_I.iw[13] ;
 wire \top_I.branch[5].block[8].um_I.iw[14] ;
 wire \top_I.branch[5].block[8].um_I.iw[15] ;
 wire \top_I.branch[5].block[8].um_I.iw[16] ;
 wire \top_I.branch[5].block[8].um_I.iw[17] ;
 wire \top_I.branch[5].block[8].um_I.iw[1] ;
 wire \top_I.branch[5].block[8].um_I.iw[2] ;
 wire \top_I.branch[5].block[8].um_I.iw[3] ;
 wire \top_I.branch[5].block[8].um_I.iw[4] ;
 wire \top_I.branch[5].block[8].um_I.iw[5] ;
 wire \top_I.branch[5].block[8].um_I.iw[6] ;
 wire \top_I.branch[5].block[8].um_I.iw[7] ;
 wire \top_I.branch[5].block[8].um_I.iw[8] ;
 wire \top_I.branch[5].block[8].um_I.iw[9] ;
 wire \top_I.branch[5].block[8].um_I.k_zero ;
 wire \top_I.branch[5].block[8].um_I.pg_vdd ;
 wire \top_I.branch[5].block[9].um_I.ana[0] ;
 wire \top_I.branch[5].block[9].um_I.ana[1] ;
 wire \top_I.branch[5].block[9].um_I.ana[2] ;
 wire \top_I.branch[5].block[9].um_I.ana[3] ;
 wire \top_I.branch[5].block[9].um_I.ana[4] ;
 wire \top_I.branch[5].block[9].um_I.ana[5] ;
 wire \top_I.branch[5].block[9].um_I.ana[6] ;
 wire \top_I.branch[5].block[9].um_I.ana[7] ;
 wire \top_I.branch[5].block[9].um_I.clk ;
 wire \top_I.branch[5].block[9].um_I.ena ;
 wire \top_I.branch[5].block[9].um_I.iw[10] ;
 wire \top_I.branch[5].block[9].um_I.iw[11] ;
 wire \top_I.branch[5].block[9].um_I.iw[12] ;
 wire \top_I.branch[5].block[9].um_I.iw[13] ;
 wire \top_I.branch[5].block[9].um_I.iw[14] ;
 wire \top_I.branch[5].block[9].um_I.iw[15] ;
 wire \top_I.branch[5].block[9].um_I.iw[16] ;
 wire \top_I.branch[5].block[9].um_I.iw[17] ;
 wire \top_I.branch[5].block[9].um_I.iw[1] ;
 wire \top_I.branch[5].block[9].um_I.iw[2] ;
 wire \top_I.branch[5].block[9].um_I.iw[3] ;
 wire \top_I.branch[5].block[9].um_I.iw[4] ;
 wire \top_I.branch[5].block[9].um_I.iw[5] ;
 wire \top_I.branch[5].block[9].um_I.iw[6] ;
 wire \top_I.branch[5].block[9].um_I.iw[7] ;
 wire \top_I.branch[5].block[9].um_I.iw[8] ;
 wire \top_I.branch[5].block[9].um_I.iw[9] ;
 wire \top_I.branch[5].block[9].um_I.k_zero ;
 wire \top_I.branch[5].block[9].um_I.pg_vdd ;
 wire \top_I.branch[5].l_addr[0] ;
 wire \top_I.branch[5].l_addr[1] ;
 wire \top_I.branch[6].block[0].um_I.ana[0] ;
 wire \top_I.branch[6].block[0].um_I.ana[1] ;
 wire \top_I.branch[6].block[0].um_I.ana[2] ;
 wire \top_I.branch[6].block[0].um_I.ana[3] ;
 wire \top_I.branch[6].block[0].um_I.ana[4] ;
 wire \top_I.branch[6].block[0].um_I.ana[5] ;
 wire \top_I.branch[6].block[0].um_I.ana[6] ;
 wire \top_I.branch[6].block[0].um_I.ana[7] ;
 wire \top_I.branch[6].block[0].um_I.clk ;
 wire \top_I.branch[6].block[0].um_I.ena ;
 wire \top_I.branch[6].block[0].um_I.iw[10] ;
 wire \top_I.branch[6].block[0].um_I.iw[11] ;
 wire \top_I.branch[6].block[0].um_I.iw[12] ;
 wire \top_I.branch[6].block[0].um_I.iw[13] ;
 wire \top_I.branch[6].block[0].um_I.iw[14] ;
 wire \top_I.branch[6].block[0].um_I.iw[15] ;
 wire \top_I.branch[6].block[0].um_I.iw[16] ;
 wire \top_I.branch[6].block[0].um_I.iw[17] ;
 wire \top_I.branch[6].block[0].um_I.iw[1] ;
 wire \top_I.branch[6].block[0].um_I.iw[2] ;
 wire \top_I.branch[6].block[0].um_I.iw[3] ;
 wire \top_I.branch[6].block[0].um_I.iw[4] ;
 wire \top_I.branch[6].block[0].um_I.iw[5] ;
 wire \top_I.branch[6].block[0].um_I.iw[6] ;
 wire \top_I.branch[6].block[0].um_I.iw[7] ;
 wire \top_I.branch[6].block[0].um_I.iw[8] ;
 wire \top_I.branch[6].block[0].um_I.iw[9] ;
 wire \top_I.branch[6].block[0].um_I.k_zero ;
 wire \top_I.branch[6].block[0].um_I.pg_vdd ;
 wire \top_I.branch[6].block[10].um_I.ana[0] ;
 wire \top_I.branch[6].block[10].um_I.ana[1] ;
 wire \top_I.branch[6].block[10].um_I.ana[2] ;
 wire \top_I.branch[6].block[10].um_I.ana[3] ;
 wire \top_I.branch[6].block[10].um_I.ana[4] ;
 wire \top_I.branch[6].block[10].um_I.ana[5] ;
 wire \top_I.branch[6].block[10].um_I.ana[6] ;
 wire \top_I.branch[6].block[10].um_I.ana[7] ;
 wire \top_I.branch[6].block[10].um_I.clk ;
 wire \top_I.branch[6].block[10].um_I.ena ;
 wire \top_I.branch[6].block[10].um_I.iw[10] ;
 wire \top_I.branch[6].block[10].um_I.iw[11] ;
 wire \top_I.branch[6].block[10].um_I.iw[12] ;
 wire \top_I.branch[6].block[10].um_I.iw[13] ;
 wire \top_I.branch[6].block[10].um_I.iw[14] ;
 wire \top_I.branch[6].block[10].um_I.iw[15] ;
 wire \top_I.branch[6].block[10].um_I.iw[16] ;
 wire \top_I.branch[6].block[10].um_I.iw[17] ;
 wire \top_I.branch[6].block[10].um_I.iw[1] ;
 wire \top_I.branch[6].block[10].um_I.iw[2] ;
 wire \top_I.branch[6].block[10].um_I.iw[3] ;
 wire \top_I.branch[6].block[10].um_I.iw[4] ;
 wire \top_I.branch[6].block[10].um_I.iw[5] ;
 wire \top_I.branch[6].block[10].um_I.iw[6] ;
 wire \top_I.branch[6].block[10].um_I.iw[7] ;
 wire \top_I.branch[6].block[10].um_I.iw[8] ;
 wire \top_I.branch[6].block[10].um_I.iw[9] ;
 wire \top_I.branch[6].block[10].um_I.k_zero ;
 wire \top_I.branch[6].block[10].um_I.pg_vdd ;
 wire \top_I.branch[6].block[11].um_I.ana[0] ;
 wire \top_I.branch[6].block[11].um_I.ana[1] ;
 wire \top_I.branch[6].block[11].um_I.ana[2] ;
 wire \top_I.branch[6].block[11].um_I.ana[3] ;
 wire \top_I.branch[6].block[11].um_I.ana[4] ;
 wire \top_I.branch[6].block[11].um_I.ana[5] ;
 wire \top_I.branch[6].block[11].um_I.ana[6] ;
 wire \top_I.branch[6].block[11].um_I.ana[7] ;
 wire \top_I.branch[6].block[11].um_I.clk ;
 wire \top_I.branch[6].block[11].um_I.ena ;
 wire \top_I.branch[6].block[11].um_I.iw[10] ;
 wire \top_I.branch[6].block[11].um_I.iw[11] ;
 wire \top_I.branch[6].block[11].um_I.iw[12] ;
 wire \top_I.branch[6].block[11].um_I.iw[13] ;
 wire \top_I.branch[6].block[11].um_I.iw[14] ;
 wire \top_I.branch[6].block[11].um_I.iw[15] ;
 wire \top_I.branch[6].block[11].um_I.iw[16] ;
 wire \top_I.branch[6].block[11].um_I.iw[17] ;
 wire \top_I.branch[6].block[11].um_I.iw[1] ;
 wire \top_I.branch[6].block[11].um_I.iw[2] ;
 wire \top_I.branch[6].block[11].um_I.iw[3] ;
 wire \top_I.branch[6].block[11].um_I.iw[4] ;
 wire \top_I.branch[6].block[11].um_I.iw[5] ;
 wire \top_I.branch[6].block[11].um_I.iw[6] ;
 wire \top_I.branch[6].block[11].um_I.iw[7] ;
 wire \top_I.branch[6].block[11].um_I.iw[8] ;
 wire \top_I.branch[6].block[11].um_I.iw[9] ;
 wire \top_I.branch[6].block[11].um_I.k_zero ;
 wire \top_I.branch[6].block[11].um_I.pg_vdd ;
 wire \top_I.branch[6].block[12].um_I.ana[0] ;
 wire \top_I.branch[6].block[12].um_I.ana[1] ;
 wire \top_I.branch[6].block[12].um_I.ana[2] ;
 wire \top_I.branch[6].block[12].um_I.ana[3] ;
 wire \top_I.branch[6].block[12].um_I.ana[4] ;
 wire \top_I.branch[6].block[12].um_I.ana[5] ;
 wire \top_I.branch[6].block[12].um_I.ana[6] ;
 wire \top_I.branch[6].block[12].um_I.ana[7] ;
 wire \top_I.branch[6].block[12].um_I.clk ;
 wire \top_I.branch[6].block[12].um_I.ena ;
 wire \top_I.branch[6].block[12].um_I.iw[10] ;
 wire \top_I.branch[6].block[12].um_I.iw[11] ;
 wire \top_I.branch[6].block[12].um_I.iw[12] ;
 wire \top_I.branch[6].block[12].um_I.iw[13] ;
 wire \top_I.branch[6].block[12].um_I.iw[14] ;
 wire \top_I.branch[6].block[12].um_I.iw[15] ;
 wire \top_I.branch[6].block[12].um_I.iw[16] ;
 wire \top_I.branch[6].block[12].um_I.iw[17] ;
 wire \top_I.branch[6].block[12].um_I.iw[1] ;
 wire \top_I.branch[6].block[12].um_I.iw[2] ;
 wire \top_I.branch[6].block[12].um_I.iw[3] ;
 wire \top_I.branch[6].block[12].um_I.iw[4] ;
 wire \top_I.branch[6].block[12].um_I.iw[5] ;
 wire \top_I.branch[6].block[12].um_I.iw[6] ;
 wire \top_I.branch[6].block[12].um_I.iw[7] ;
 wire \top_I.branch[6].block[12].um_I.iw[8] ;
 wire \top_I.branch[6].block[12].um_I.iw[9] ;
 wire \top_I.branch[6].block[12].um_I.k_zero ;
 wire \top_I.branch[6].block[12].um_I.pg_vdd ;
 wire \top_I.branch[6].block[13].um_I.ana[0] ;
 wire \top_I.branch[6].block[13].um_I.ana[1] ;
 wire \top_I.branch[6].block[13].um_I.ana[2] ;
 wire \top_I.branch[6].block[13].um_I.ana[3] ;
 wire \top_I.branch[6].block[13].um_I.ana[4] ;
 wire \top_I.branch[6].block[13].um_I.ana[5] ;
 wire \top_I.branch[6].block[13].um_I.ana[6] ;
 wire \top_I.branch[6].block[13].um_I.ana[7] ;
 wire \top_I.branch[6].block[13].um_I.clk ;
 wire \top_I.branch[6].block[13].um_I.ena ;
 wire \top_I.branch[6].block[13].um_I.iw[10] ;
 wire \top_I.branch[6].block[13].um_I.iw[11] ;
 wire \top_I.branch[6].block[13].um_I.iw[12] ;
 wire \top_I.branch[6].block[13].um_I.iw[13] ;
 wire \top_I.branch[6].block[13].um_I.iw[14] ;
 wire \top_I.branch[6].block[13].um_I.iw[15] ;
 wire \top_I.branch[6].block[13].um_I.iw[16] ;
 wire \top_I.branch[6].block[13].um_I.iw[17] ;
 wire \top_I.branch[6].block[13].um_I.iw[1] ;
 wire \top_I.branch[6].block[13].um_I.iw[2] ;
 wire \top_I.branch[6].block[13].um_I.iw[3] ;
 wire \top_I.branch[6].block[13].um_I.iw[4] ;
 wire \top_I.branch[6].block[13].um_I.iw[5] ;
 wire \top_I.branch[6].block[13].um_I.iw[6] ;
 wire \top_I.branch[6].block[13].um_I.iw[7] ;
 wire \top_I.branch[6].block[13].um_I.iw[8] ;
 wire \top_I.branch[6].block[13].um_I.iw[9] ;
 wire \top_I.branch[6].block[13].um_I.k_zero ;
 wire \top_I.branch[6].block[13].um_I.pg_vdd ;
 wire \top_I.branch[6].block[14].um_I.ana[0] ;
 wire \top_I.branch[6].block[14].um_I.ana[1] ;
 wire \top_I.branch[6].block[14].um_I.ana[2] ;
 wire \top_I.branch[6].block[14].um_I.ana[3] ;
 wire \top_I.branch[6].block[14].um_I.ana[4] ;
 wire \top_I.branch[6].block[14].um_I.ana[5] ;
 wire \top_I.branch[6].block[14].um_I.ana[6] ;
 wire \top_I.branch[6].block[14].um_I.ana[7] ;
 wire \top_I.branch[6].block[14].um_I.clk ;
 wire \top_I.branch[6].block[14].um_I.ena ;
 wire \top_I.branch[6].block[14].um_I.iw[10] ;
 wire \top_I.branch[6].block[14].um_I.iw[11] ;
 wire \top_I.branch[6].block[14].um_I.iw[12] ;
 wire \top_I.branch[6].block[14].um_I.iw[13] ;
 wire \top_I.branch[6].block[14].um_I.iw[14] ;
 wire \top_I.branch[6].block[14].um_I.iw[15] ;
 wire \top_I.branch[6].block[14].um_I.iw[16] ;
 wire \top_I.branch[6].block[14].um_I.iw[17] ;
 wire \top_I.branch[6].block[14].um_I.iw[1] ;
 wire \top_I.branch[6].block[14].um_I.iw[2] ;
 wire \top_I.branch[6].block[14].um_I.iw[3] ;
 wire \top_I.branch[6].block[14].um_I.iw[4] ;
 wire \top_I.branch[6].block[14].um_I.iw[5] ;
 wire \top_I.branch[6].block[14].um_I.iw[6] ;
 wire \top_I.branch[6].block[14].um_I.iw[7] ;
 wire \top_I.branch[6].block[14].um_I.iw[8] ;
 wire \top_I.branch[6].block[14].um_I.iw[9] ;
 wire \top_I.branch[6].block[14].um_I.k_zero ;
 wire \top_I.branch[6].block[14].um_I.pg_vdd ;
 wire \top_I.branch[6].block[15].um_I.ana[0] ;
 wire \top_I.branch[6].block[15].um_I.ana[1] ;
 wire \top_I.branch[6].block[15].um_I.ana[2] ;
 wire \top_I.branch[6].block[15].um_I.ana[3] ;
 wire \top_I.branch[6].block[15].um_I.ana[4] ;
 wire \top_I.branch[6].block[15].um_I.ana[5] ;
 wire \top_I.branch[6].block[15].um_I.ana[6] ;
 wire \top_I.branch[6].block[15].um_I.ana[7] ;
 wire \top_I.branch[6].block[15].um_I.clk ;
 wire \top_I.branch[6].block[15].um_I.ena ;
 wire \top_I.branch[6].block[15].um_I.iw[10] ;
 wire \top_I.branch[6].block[15].um_I.iw[11] ;
 wire \top_I.branch[6].block[15].um_I.iw[12] ;
 wire \top_I.branch[6].block[15].um_I.iw[13] ;
 wire \top_I.branch[6].block[15].um_I.iw[14] ;
 wire \top_I.branch[6].block[15].um_I.iw[15] ;
 wire \top_I.branch[6].block[15].um_I.iw[16] ;
 wire \top_I.branch[6].block[15].um_I.iw[17] ;
 wire \top_I.branch[6].block[15].um_I.iw[1] ;
 wire \top_I.branch[6].block[15].um_I.iw[2] ;
 wire \top_I.branch[6].block[15].um_I.iw[3] ;
 wire \top_I.branch[6].block[15].um_I.iw[4] ;
 wire \top_I.branch[6].block[15].um_I.iw[5] ;
 wire \top_I.branch[6].block[15].um_I.iw[6] ;
 wire \top_I.branch[6].block[15].um_I.iw[7] ;
 wire \top_I.branch[6].block[15].um_I.iw[8] ;
 wire \top_I.branch[6].block[15].um_I.iw[9] ;
 wire \top_I.branch[6].block[15].um_I.k_zero ;
 wire \top_I.branch[6].block[15].um_I.pg_vdd ;
 wire \top_I.branch[6].block[1].um_I.ana[0] ;
 wire \top_I.branch[6].block[1].um_I.ana[1] ;
 wire \top_I.branch[6].block[1].um_I.ana[2] ;
 wire \top_I.branch[6].block[1].um_I.ana[3] ;
 wire \top_I.branch[6].block[1].um_I.ana[4] ;
 wire \top_I.branch[6].block[1].um_I.ana[5] ;
 wire \top_I.branch[6].block[1].um_I.ana[6] ;
 wire \top_I.branch[6].block[1].um_I.ana[7] ;
 wire \top_I.branch[6].block[1].um_I.clk ;
 wire \top_I.branch[6].block[1].um_I.ena ;
 wire \top_I.branch[6].block[1].um_I.iw[10] ;
 wire \top_I.branch[6].block[1].um_I.iw[11] ;
 wire \top_I.branch[6].block[1].um_I.iw[12] ;
 wire \top_I.branch[6].block[1].um_I.iw[13] ;
 wire \top_I.branch[6].block[1].um_I.iw[14] ;
 wire \top_I.branch[6].block[1].um_I.iw[15] ;
 wire \top_I.branch[6].block[1].um_I.iw[16] ;
 wire \top_I.branch[6].block[1].um_I.iw[17] ;
 wire \top_I.branch[6].block[1].um_I.iw[1] ;
 wire \top_I.branch[6].block[1].um_I.iw[2] ;
 wire \top_I.branch[6].block[1].um_I.iw[3] ;
 wire \top_I.branch[6].block[1].um_I.iw[4] ;
 wire \top_I.branch[6].block[1].um_I.iw[5] ;
 wire \top_I.branch[6].block[1].um_I.iw[6] ;
 wire \top_I.branch[6].block[1].um_I.iw[7] ;
 wire \top_I.branch[6].block[1].um_I.iw[8] ;
 wire \top_I.branch[6].block[1].um_I.iw[9] ;
 wire \top_I.branch[6].block[1].um_I.k_zero ;
 wire \top_I.branch[6].block[1].um_I.pg_vdd ;
 wire \top_I.branch[6].block[2].um_I.ana[0] ;
 wire \top_I.branch[6].block[2].um_I.ana[1] ;
 wire \top_I.branch[6].block[2].um_I.ana[2] ;
 wire \top_I.branch[6].block[2].um_I.ana[3] ;
 wire \top_I.branch[6].block[2].um_I.ana[4] ;
 wire \top_I.branch[6].block[2].um_I.ana[5] ;
 wire \top_I.branch[6].block[2].um_I.ana[6] ;
 wire \top_I.branch[6].block[2].um_I.ana[7] ;
 wire \top_I.branch[6].block[2].um_I.clk ;
 wire \top_I.branch[6].block[2].um_I.ena ;
 wire \top_I.branch[6].block[2].um_I.iw[10] ;
 wire \top_I.branch[6].block[2].um_I.iw[11] ;
 wire \top_I.branch[6].block[2].um_I.iw[12] ;
 wire \top_I.branch[6].block[2].um_I.iw[13] ;
 wire \top_I.branch[6].block[2].um_I.iw[14] ;
 wire \top_I.branch[6].block[2].um_I.iw[15] ;
 wire \top_I.branch[6].block[2].um_I.iw[16] ;
 wire \top_I.branch[6].block[2].um_I.iw[17] ;
 wire \top_I.branch[6].block[2].um_I.iw[1] ;
 wire \top_I.branch[6].block[2].um_I.iw[2] ;
 wire \top_I.branch[6].block[2].um_I.iw[3] ;
 wire \top_I.branch[6].block[2].um_I.iw[4] ;
 wire \top_I.branch[6].block[2].um_I.iw[5] ;
 wire \top_I.branch[6].block[2].um_I.iw[6] ;
 wire \top_I.branch[6].block[2].um_I.iw[7] ;
 wire \top_I.branch[6].block[2].um_I.iw[8] ;
 wire \top_I.branch[6].block[2].um_I.iw[9] ;
 wire \top_I.branch[6].block[2].um_I.k_zero ;
 wire \top_I.branch[6].block[2].um_I.pg_vdd ;
 wire \top_I.branch[6].block[3].um_I.ana[0] ;
 wire \top_I.branch[6].block[3].um_I.ana[1] ;
 wire \top_I.branch[6].block[3].um_I.ana[2] ;
 wire \top_I.branch[6].block[3].um_I.ana[3] ;
 wire \top_I.branch[6].block[3].um_I.ana[4] ;
 wire \top_I.branch[6].block[3].um_I.ana[5] ;
 wire \top_I.branch[6].block[3].um_I.ana[6] ;
 wire \top_I.branch[6].block[3].um_I.ana[7] ;
 wire \top_I.branch[6].block[3].um_I.clk ;
 wire \top_I.branch[6].block[3].um_I.ena ;
 wire \top_I.branch[6].block[3].um_I.iw[10] ;
 wire \top_I.branch[6].block[3].um_I.iw[11] ;
 wire \top_I.branch[6].block[3].um_I.iw[12] ;
 wire \top_I.branch[6].block[3].um_I.iw[13] ;
 wire \top_I.branch[6].block[3].um_I.iw[14] ;
 wire \top_I.branch[6].block[3].um_I.iw[15] ;
 wire \top_I.branch[6].block[3].um_I.iw[16] ;
 wire \top_I.branch[6].block[3].um_I.iw[17] ;
 wire \top_I.branch[6].block[3].um_I.iw[1] ;
 wire \top_I.branch[6].block[3].um_I.iw[2] ;
 wire \top_I.branch[6].block[3].um_I.iw[3] ;
 wire \top_I.branch[6].block[3].um_I.iw[4] ;
 wire \top_I.branch[6].block[3].um_I.iw[5] ;
 wire \top_I.branch[6].block[3].um_I.iw[6] ;
 wire \top_I.branch[6].block[3].um_I.iw[7] ;
 wire \top_I.branch[6].block[3].um_I.iw[8] ;
 wire \top_I.branch[6].block[3].um_I.iw[9] ;
 wire \top_I.branch[6].block[3].um_I.k_zero ;
 wire \top_I.branch[6].block[3].um_I.pg_vdd ;
 wire \top_I.branch[6].block[4].um_I.ana[0] ;
 wire \top_I.branch[6].block[4].um_I.ana[1] ;
 wire \top_I.branch[6].block[4].um_I.ana[2] ;
 wire \top_I.branch[6].block[4].um_I.ana[3] ;
 wire \top_I.branch[6].block[4].um_I.ana[4] ;
 wire \top_I.branch[6].block[4].um_I.ana[5] ;
 wire \top_I.branch[6].block[4].um_I.ana[6] ;
 wire \top_I.branch[6].block[4].um_I.ana[7] ;
 wire \top_I.branch[6].block[4].um_I.clk ;
 wire \top_I.branch[6].block[4].um_I.ena ;
 wire \top_I.branch[6].block[4].um_I.iw[10] ;
 wire \top_I.branch[6].block[4].um_I.iw[11] ;
 wire \top_I.branch[6].block[4].um_I.iw[12] ;
 wire \top_I.branch[6].block[4].um_I.iw[13] ;
 wire \top_I.branch[6].block[4].um_I.iw[14] ;
 wire \top_I.branch[6].block[4].um_I.iw[15] ;
 wire \top_I.branch[6].block[4].um_I.iw[16] ;
 wire \top_I.branch[6].block[4].um_I.iw[17] ;
 wire \top_I.branch[6].block[4].um_I.iw[1] ;
 wire \top_I.branch[6].block[4].um_I.iw[2] ;
 wire \top_I.branch[6].block[4].um_I.iw[3] ;
 wire \top_I.branch[6].block[4].um_I.iw[4] ;
 wire \top_I.branch[6].block[4].um_I.iw[5] ;
 wire \top_I.branch[6].block[4].um_I.iw[6] ;
 wire \top_I.branch[6].block[4].um_I.iw[7] ;
 wire \top_I.branch[6].block[4].um_I.iw[8] ;
 wire \top_I.branch[6].block[4].um_I.iw[9] ;
 wire \top_I.branch[6].block[4].um_I.k_zero ;
 wire \top_I.branch[6].block[4].um_I.pg_vdd ;
 wire \top_I.branch[6].block[5].um_I.ana[0] ;
 wire \top_I.branch[6].block[5].um_I.ana[1] ;
 wire \top_I.branch[6].block[5].um_I.ana[2] ;
 wire \top_I.branch[6].block[5].um_I.ana[3] ;
 wire \top_I.branch[6].block[5].um_I.ana[4] ;
 wire \top_I.branch[6].block[5].um_I.ana[5] ;
 wire \top_I.branch[6].block[5].um_I.ana[6] ;
 wire \top_I.branch[6].block[5].um_I.ana[7] ;
 wire \top_I.branch[6].block[5].um_I.clk ;
 wire \top_I.branch[6].block[5].um_I.ena ;
 wire \top_I.branch[6].block[5].um_I.iw[10] ;
 wire \top_I.branch[6].block[5].um_I.iw[11] ;
 wire \top_I.branch[6].block[5].um_I.iw[12] ;
 wire \top_I.branch[6].block[5].um_I.iw[13] ;
 wire \top_I.branch[6].block[5].um_I.iw[14] ;
 wire \top_I.branch[6].block[5].um_I.iw[15] ;
 wire \top_I.branch[6].block[5].um_I.iw[16] ;
 wire \top_I.branch[6].block[5].um_I.iw[17] ;
 wire \top_I.branch[6].block[5].um_I.iw[1] ;
 wire \top_I.branch[6].block[5].um_I.iw[2] ;
 wire \top_I.branch[6].block[5].um_I.iw[3] ;
 wire \top_I.branch[6].block[5].um_I.iw[4] ;
 wire \top_I.branch[6].block[5].um_I.iw[5] ;
 wire \top_I.branch[6].block[5].um_I.iw[6] ;
 wire \top_I.branch[6].block[5].um_I.iw[7] ;
 wire \top_I.branch[6].block[5].um_I.iw[8] ;
 wire \top_I.branch[6].block[5].um_I.iw[9] ;
 wire \top_I.branch[6].block[5].um_I.k_zero ;
 wire \top_I.branch[6].block[5].um_I.pg_vdd ;
 wire \top_I.branch[6].block[6].um_I.ana[0] ;
 wire \top_I.branch[6].block[6].um_I.ana[1] ;
 wire \top_I.branch[6].block[6].um_I.ana[2] ;
 wire \top_I.branch[6].block[6].um_I.ana[3] ;
 wire \top_I.branch[6].block[6].um_I.ana[4] ;
 wire \top_I.branch[6].block[6].um_I.ana[5] ;
 wire \top_I.branch[6].block[6].um_I.ana[6] ;
 wire \top_I.branch[6].block[6].um_I.ana[7] ;
 wire \top_I.branch[6].block[6].um_I.clk ;
 wire \top_I.branch[6].block[6].um_I.ena ;
 wire \top_I.branch[6].block[6].um_I.iw[10] ;
 wire \top_I.branch[6].block[6].um_I.iw[11] ;
 wire \top_I.branch[6].block[6].um_I.iw[12] ;
 wire \top_I.branch[6].block[6].um_I.iw[13] ;
 wire \top_I.branch[6].block[6].um_I.iw[14] ;
 wire \top_I.branch[6].block[6].um_I.iw[15] ;
 wire \top_I.branch[6].block[6].um_I.iw[16] ;
 wire \top_I.branch[6].block[6].um_I.iw[17] ;
 wire \top_I.branch[6].block[6].um_I.iw[1] ;
 wire \top_I.branch[6].block[6].um_I.iw[2] ;
 wire \top_I.branch[6].block[6].um_I.iw[3] ;
 wire \top_I.branch[6].block[6].um_I.iw[4] ;
 wire \top_I.branch[6].block[6].um_I.iw[5] ;
 wire \top_I.branch[6].block[6].um_I.iw[6] ;
 wire \top_I.branch[6].block[6].um_I.iw[7] ;
 wire \top_I.branch[6].block[6].um_I.iw[8] ;
 wire \top_I.branch[6].block[6].um_I.iw[9] ;
 wire \top_I.branch[6].block[6].um_I.k_zero ;
 wire \top_I.branch[6].block[6].um_I.pg_vdd ;
 wire \top_I.branch[6].block[7].um_I.ana[0] ;
 wire \top_I.branch[6].block[7].um_I.ana[1] ;
 wire \top_I.branch[6].block[7].um_I.ana[2] ;
 wire \top_I.branch[6].block[7].um_I.ana[3] ;
 wire \top_I.branch[6].block[7].um_I.ana[4] ;
 wire \top_I.branch[6].block[7].um_I.ana[5] ;
 wire \top_I.branch[6].block[7].um_I.ana[6] ;
 wire \top_I.branch[6].block[7].um_I.ana[7] ;
 wire \top_I.branch[6].block[7].um_I.clk ;
 wire \top_I.branch[6].block[7].um_I.ena ;
 wire \top_I.branch[6].block[7].um_I.iw[10] ;
 wire \top_I.branch[6].block[7].um_I.iw[11] ;
 wire \top_I.branch[6].block[7].um_I.iw[12] ;
 wire \top_I.branch[6].block[7].um_I.iw[13] ;
 wire \top_I.branch[6].block[7].um_I.iw[14] ;
 wire \top_I.branch[6].block[7].um_I.iw[15] ;
 wire \top_I.branch[6].block[7].um_I.iw[16] ;
 wire \top_I.branch[6].block[7].um_I.iw[17] ;
 wire \top_I.branch[6].block[7].um_I.iw[1] ;
 wire \top_I.branch[6].block[7].um_I.iw[2] ;
 wire \top_I.branch[6].block[7].um_I.iw[3] ;
 wire \top_I.branch[6].block[7].um_I.iw[4] ;
 wire \top_I.branch[6].block[7].um_I.iw[5] ;
 wire \top_I.branch[6].block[7].um_I.iw[6] ;
 wire \top_I.branch[6].block[7].um_I.iw[7] ;
 wire \top_I.branch[6].block[7].um_I.iw[8] ;
 wire \top_I.branch[6].block[7].um_I.iw[9] ;
 wire \top_I.branch[6].block[7].um_I.k_zero ;
 wire \top_I.branch[6].block[7].um_I.pg_vdd ;
 wire \top_I.branch[6].block[8].um_I.ana[0] ;
 wire \top_I.branch[6].block[8].um_I.ana[1] ;
 wire \top_I.branch[6].block[8].um_I.ana[2] ;
 wire \top_I.branch[6].block[8].um_I.ana[3] ;
 wire \top_I.branch[6].block[8].um_I.ana[4] ;
 wire \top_I.branch[6].block[8].um_I.ana[5] ;
 wire \top_I.branch[6].block[8].um_I.ana[6] ;
 wire \top_I.branch[6].block[8].um_I.ana[7] ;
 wire \top_I.branch[6].block[8].um_I.clk ;
 wire \top_I.branch[6].block[8].um_I.ena ;
 wire \top_I.branch[6].block[8].um_I.iw[10] ;
 wire \top_I.branch[6].block[8].um_I.iw[11] ;
 wire \top_I.branch[6].block[8].um_I.iw[12] ;
 wire \top_I.branch[6].block[8].um_I.iw[13] ;
 wire \top_I.branch[6].block[8].um_I.iw[14] ;
 wire \top_I.branch[6].block[8].um_I.iw[15] ;
 wire \top_I.branch[6].block[8].um_I.iw[16] ;
 wire \top_I.branch[6].block[8].um_I.iw[17] ;
 wire \top_I.branch[6].block[8].um_I.iw[1] ;
 wire \top_I.branch[6].block[8].um_I.iw[2] ;
 wire \top_I.branch[6].block[8].um_I.iw[3] ;
 wire \top_I.branch[6].block[8].um_I.iw[4] ;
 wire \top_I.branch[6].block[8].um_I.iw[5] ;
 wire \top_I.branch[6].block[8].um_I.iw[6] ;
 wire \top_I.branch[6].block[8].um_I.iw[7] ;
 wire \top_I.branch[6].block[8].um_I.iw[8] ;
 wire \top_I.branch[6].block[8].um_I.iw[9] ;
 wire \top_I.branch[6].block[8].um_I.k_zero ;
 wire \top_I.branch[6].block[8].um_I.pg_vdd ;
 wire \top_I.branch[6].block[9].um_I.ana[0] ;
 wire \top_I.branch[6].block[9].um_I.ana[1] ;
 wire \top_I.branch[6].block[9].um_I.ana[2] ;
 wire \top_I.branch[6].block[9].um_I.ana[3] ;
 wire \top_I.branch[6].block[9].um_I.ana[4] ;
 wire \top_I.branch[6].block[9].um_I.ana[5] ;
 wire \top_I.branch[6].block[9].um_I.ana[6] ;
 wire \top_I.branch[6].block[9].um_I.ana[7] ;
 wire \top_I.branch[6].block[9].um_I.clk ;
 wire \top_I.branch[6].block[9].um_I.ena ;
 wire \top_I.branch[6].block[9].um_I.iw[10] ;
 wire \top_I.branch[6].block[9].um_I.iw[11] ;
 wire \top_I.branch[6].block[9].um_I.iw[12] ;
 wire \top_I.branch[6].block[9].um_I.iw[13] ;
 wire \top_I.branch[6].block[9].um_I.iw[14] ;
 wire \top_I.branch[6].block[9].um_I.iw[15] ;
 wire \top_I.branch[6].block[9].um_I.iw[16] ;
 wire \top_I.branch[6].block[9].um_I.iw[17] ;
 wire \top_I.branch[6].block[9].um_I.iw[1] ;
 wire \top_I.branch[6].block[9].um_I.iw[2] ;
 wire \top_I.branch[6].block[9].um_I.iw[3] ;
 wire \top_I.branch[6].block[9].um_I.iw[4] ;
 wire \top_I.branch[6].block[9].um_I.iw[5] ;
 wire \top_I.branch[6].block[9].um_I.iw[6] ;
 wire \top_I.branch[6].block[9].um_I.iw[7] ;
 wire \top_I.branch[6].block[9].um_I.iw[8] ;
 wire \top_I.branch[6].block[9].um_I.iw[9] ;
 wire \top_I.branch[6].block[9].um_I.k_zero ;
 wire \top_I.branch[6].block[9].um_I.pg_vdd ;
 wire \top_I.branch[6].l_addr[0] ;
 wire \top_I.branch[6].l_addr[2] ;
 wire \top_I.branch[7].block[0].um_I.ana[0] ;
 wire \top_I.branch[7].block[0].um_I.ana[1] ;
 wire \top_I.branch[7].block[0].um_I.ana[2] ;
 wire \top_I.branch[7].block[0].um_I.ana[3] ;
 wire \top_I.branch[7].block[0].um_I.ana[4] ;
 wire \top_I.branch[7].block[0].um_I.ana[5] ;
 wire \top_I.branch[7].block[0].um_I.ana[6] ;
 wire \top_I.branch[7].block[0].um_I.ana[7] ;
 wire \top_I.branch[7].block[0].um_I.clk ;
 wire \top_I.branch[7].block[0].um_I.ena ;
 wire \top_I.branch[7].block[0].um_I.iw[10] ;
 wire \top_I.branch[7].block[0].um_I.iw[11] ;
 wire \top_I.branch[7].block[0].um_I.iw[12] ;
 wire \top_I.branch[7].block[0].um_I.iw[13] ;
 wire \top_I.branch[7].block[0].um_I.iw[14] ;
 wire \top_I.branch[7].block[0].um_I.iw[15] ;
 wire \top_I.branch[7].block[0].um_I.iw[16] ;
 wire \top_I.branch[7].block[0].um_I.iw[17] ;
 wire \top_I.branch[7].block[0].um_I.iw[1] ;
 wire \top_I.branch[7].block[0].um_I.iw[2] ;
 wire \top_I.branch[7].block[0].um_I.iw[3] ;
 wire \top_I.branch[7].block[0].um_I.iw[4] ;
 wire \top_I.branch[7].block[0].um_I.iw[5] ;
 wire \top_I.branch[7].block[0].um_I.iw[6] ;
 wire \top_I.branch[7].block[0].um_I.iw[7] ;
 wire \top_I.branch[7].block[0].um_I.iw[8] ;
 wire \top_I.branch[7].block[0].um_I.iw[9] ;
 wire \top_I.branch[7].block[0].um_I.k_zero ;
 wire \top_I.branch[7].block[0].um_I.pg_vdd ;
 wire \top_I.branch[7].block[10].um_I.ana[0] ;
 wire \top_I.branch[7].block[10].um_I.ana[1] ;
 wire \top_I.branch[7].block[10].um_I.ana[2] ;
 wire \top_I.branch[7].block[10].um_I.ana[3] ;
 wire \top_I.branch[7].block[10].um_I.ana[4] ;
 wire \top_I.branch[7].block[10].um_I.ana[5] ;
 wire \top_I.branch[7].block[10].um_I.ana[6] ;
 wire \top_I.branch[7].block[10].um_I.ana[7] ;
 wire \top_I.branch[7].block[10].um_I.clk ;
 wire \top_I.branch[7].block[10].um_I.ena ;
 wire \top_I.branch[7].block[10].um_I.iw[10] ;
 wire \top_I.branch[7].block[10].um_I.iw[11] ;
 wire \top_I.branch[7].block[10].um_I.iw[12] ;
 wire \top_I.branch[7].block[10].um_I.iw[13] ;
 wire \top_I.branch[7].block[10].um_I.iw[14] ;
 wire \top_I.branch[7].block[10].um_I.iw[15] ;
 wire \top_I.branch[7].block[10].um_I.iw[16] ;
 wire \top_I.branch[7].block[10].um_I.iw[17] ;
 wire \top_I.branch[7].block[10].um_I.iw[1] ;
 wire \top_I.branch[7].block[10].um_I.iw[2] ;
 wire \top_I.branch[7].block[10].um_I.iw[3] ;
 wire \top_I.branch[7].block[10].um_I.iw[4] ;
 wire \top_I.branch[7].block[10].um_I.iw[5] ;
 wire \top_I.branch[7].block[10].um_I.iw[6] ;
 wire \top_I.branch[7].block[10].um_I.iw[7] ;
 wire \top_I.branch[7].block[10].um_I.iw[8] ;
 wire \top_I.branch[7].block[10].um_I.iw[9] ;
 wire \top_I.branch[7].block[10].um_I.k_zero ;
 wire \top_I.branch[7].block[10].um_I.pg_vdd ;
 wire \top_I.branch[7].block[11].um_I.ana[0] ;
 wire \top_I.branch[7].block[11].um_I.ana[1] ;
 wire \top_I.branch[7].block[11].um_I.ana[2] ;
 wire \top_I.branch[7].block[11].um_I.ana[3] ;
 wire \top_I.branch[7].block[11].um_I.ana[4] ;
 wire \top_I.branch[7].block[11].um_I.ana[5] ;
 wire \top_I.branch[7].block[11].um_I.ana[6] ;
 wire \top_I.branch[7].block[11].um_I.ana[7] ;
 wire \top_I.branch[7].block[11].um_I.clk ;
 wire \top_I.branch[7].block[11].um_I.ena ;
 wire \top_I.branch[7].block[11].um_I.iw[10] ;
 wire \top_I.branch[7].block[11].um_I.iw[11] ;
 wire \top_I.branch[7].block[11].um_I.iw[12] ;
 wire \top_I.branch[7].block[11].um_I.iw[13] ;
 wire \top_I.branch[7].block[11].um_I.iw[14] ;
 wire \top_I.branch[7].block[11].um_I.iw[15] ;
 wire \top_I.branch[7].block[11].um_I.iw[16] ;
 wire \top_I.branch[7].block[11].um_I.iw[17] ;
 wire \top_I.branch[7].block[11].um_I.iw[1] ;
 wire \top_I.branch[7].block[11].um_I.iw[2] ;
 wire \top_I.branch[7].block[11].um_I.iw[3] ;
 wire \top_I.branch[7].block[11].um_I.iw[4] ;
 wire \top_I.branch[7].block[11].um_I.iw[5] ;
 wire \top_I.branch[7].block[11].um_I.iw[6] ;
 wire \top_I.branch[7].block[11].um_I.iw[7] ;
 wire \top_I.branch[7].block[11].um_I.iw[8] ;
 wire \top_I.branch[7].block[11].um_I.iw[9] ;
 wire \top_I.branch[7].block[11].um_I.k_zero ;
 wire \top_I.branch[7].block[11].um_I.pg_vdd ;
 wire \top_I.branch[7].block[12].um_I.ana[0] ;
 wire \top_I.branch[7].block[12].um_I.ana[1] ;
 wire \top_I.branch[7].block[12].um_I.ana[2] ;
 wire \top_I.branch[7].block[12].um_I.ana[3] ;
 wire \top_I.branch[7].block[12].um_I.ana[4] ;
 wire \top_I.branch[7].block[12].um_I.ana[5] ;
 wire \top_I.branch[7].block[12].um_I.ana[6] ;
 wire \top_I.branch[7].block[12].um_I.ana[7] ;
 wire \top_I.branch[7].block[12].um_I.clk ;
 wire \top_I.branch[7].block[12].um_I.ena ;
 wire \top_I.branch[7].block[12].um_I.iw[10] ;
 wire \top_I.branch[7].block[12].um_I.iw[11] ;
 wire \top_I.branch[7].block[12].um_I.iw[12] ;
 wire \top_I.branch[7].block[12].um_I.iw[13] ;
 wire \top_I.branch[7].block[12].um_I.iw[14] ;
 wire \top_I.branch[7].block[12].um_I.iw[15] ;
 wire \top_I.branch[7].block[12].um_I.iw[16] ;
 wire \top_I.branch[7].block[12].um_I.iw[17] ;
 wire \top_I.branch[7].block[12].um_I.iw[1] ;
 wire \top_I.branch[7].block[12].um_I.iw[2] ;
 wire \top_I.branch[7].block[12].um_I.iw[3] ;
 wire \top_I.branch[7].block[12].um_I.iw[4] ;
 wire \top_I.branch[7].block[12].um_I.iw[5] ;
 wire \top_I.branch[7].block[12].um_I.iw[6] ;
 wire \top_I.branch[7].block[12].um_I.iw[7] ;
 wire \top_I.branch[7].block[12].um_I.iw[8] ;
 wire \top_I.branch[7].block[12].um_I.iw[9] ;
 wire \top_I.branch[7].block[12].um_I.k_zero ;
 wire \top_I.branch[7].block[12].um_I.pg_vdd ;
 wire \top_I.branch[7].block[13].um_I.ana[0] ;
 wire \top_I.branch[7].block[13].um_I.ana[1] ;
 wire \top_I.branch[7].block[13].um_I.ana[2] ;
 wire \top_I.branch[7].block[13].um_I.ana[3] ;
 wire \top_I.branch[7].block[13].um_I.ana[4] ;
 wire \top_I.branch[7].block[13].um_I.ana[5] ;
 wire \top_I.branch[7].block[13].um_I.ana[6] ;
 wire \top_I.branch[7].block[13].um_I.ana[7] ;
 wire \top_I.branch[7].block[13].um_I.clk ;
 wire \top_I.branch[7].block[13].um_I.ena ;
 wire \top_I.branch[7].block[13].um_I.iw[10] ;
 wire \top_I.branch[7].block[13].um_I.iw[11] ;
 wire \top_I.branch[7].block[13].um_I.iw[12] ;
 wire \top_I.branch[7].block[13].um_I.iw[13] ;
 wire \top_I.branch[7].block[13].um_I.iw[14] ;
 wire \top_I.branch[7].block[13].um_I.iw[15] ;
 wire \top_I.branch[7].block[13].um_I.iw[16] ;
 wire \top_I.branch[7].block[13].um_I.iw[17] ;
 wire \top_I.branch[7].block[13].um_I.iw[1] ;
 wire \top_I.branch[7].block[13].um_I.iw[2] ;
 wire \top_I.branch[7].block[13].um_I.iw[3] ;
 wire \top_I.branch[7].block[13].um_I.iw[4] ;
 wire \top_I.branch[7].block[13].um_I.iw[5] ;
 wire \top_I.branch[7].block[13].um_I.iw[6] ;
 wire \top_I.branch[7].block[13].um_I.iw[7] ;
 wire \top_I.branch[7].block[13].um_I.iw[8] ;
 wire \top_I.branch[7].block[13].um_I.iw[9] ;
 wire \top_I.branch[7].block[13].um_I.k_zero ;
 wire \top_I.branch[7].block[13].um_I.pg_vdd ;
 wire \top_I.branch[7].block[14].um_I.ana[0] ;
 wire \top_I.branch[7].block[14].um_I.ana[1] ;
 wire \top_I.branch[7].block[14].um_I.ana[2] ;
 wire \top_I.branch[7].block[14].um_I.ana[3] ;
 wire \top_I.branch[7].block[14].um_I.ana[4] ;
 wire \top_I.branch[7].block[14].um_I.ana[5] ;
 wire \top_I.branch[7].block[14].um_I.ana[6] ;
 wire \top_I.branch[7].block[14].um_I.ana[7] ;
 wire \top_I.branch[7].block[14].um_I.clk ;
 wire \top_I.branch[7].block[14].um_I.ena ;
 wire \top_I.branch[7].block[14].um_I.iw[10] ;
 wire \top_I.branch[7].block[14].um_I.iw[11] ;
 wire \top_I.branch[7].block[14].um_I.iw[12] ;
 wire \top_I.branch[7].block[14].um_I.iw[13] ;
 wire \top_I.branch[7].block[14].um_I.iw[14] ;
 wire \top_I.branch[7].block[14].um_I.iw[15] ;
 wire \top_I.branch[7].block[14].um_I.iw[16] ;
 wire \top_I.branch[7].block[14].um_I.iw[17] ;
 wire \top_I.branch[7].block[14].um_I.iw[1] ;
 wire \top_I.branch[7].block[14].um_I.iw[2] ;
 wire \top_I.branch[7].block[14].um_I.iw[3] ;
 wire \top_I.branch[7].block[14].um_I.iw[4] ;
 wire \top_I.branch[7].block[14].um_I.iw[5] ;
 wire \top_I.branch[7].block[14].um_I.iw[6] ;
 wire \top_I.branch[7].block[14].um_I.iw[7] ;
 wire \top_I.branch[7].block[14].um_I.iw[8] ;
 wire \top_I.branch[7].block[14].um_I.iw[9] ;
 wire \top_I.branch[7].block[14].um_I.k_zero ;
 wire \top_I.branch[7].block[14].um_I.pg_vdd ;
 wire \top_I.branch[7].block[15].um_I.ana[0] ;
 wire \top_I.branch[7].block[15].um_I.ana[1] ;
 wire \top_I.branch[7].block[15].um_I.ana[2] ;
 wire \top_I.branch[7].block[15].um_I.ana[3] ;
 wire \top_I.branch[7].block[15].um_I.ana[4] ;
 wire \top_I.branch[7].block[15].um_I.ana[5] ;
 wire \top_I.branch[7].block[15].um_I.ana[6] ;
 wire \top_I.branch[7].block[15].um_I.ana[7] ;
 wire \top_I.branch[7].block[15].um_I.clk ;
 wire \top_I.branch[7].block[15].um_I.ena ;
 wire \top_I.branch[7].block[15].um_I.iw[10] ;
 wire \top_I.branch[7].block[15].um_I.iw[11] ;
 wire \top_I.branch[7].block[15].um_I.iw[12] ;
 wire \top_I.branch[7].block[15].um_I.iw[13] ;
 wire \top_I.branch[7].block[15].um_I.iw[14] ;
 wire \top_I.branch[7].block[15].um_I.iw[15] ;
 wire \top_I.branch[7].block[15].um_I.iw[16] ;
 wire \top_I.branch[7].block[15].um_I.iw[17] ;
 wire \top_I.branch[7].block[15].um_I.iw[1] ;
 wire \top_I.branch[7].block[15].um_I.iw[2] ;
 wire \top_I.branch[7].block[15].um_I.iw[3] ;
 wire \top_I.branch[7].block[15].um_I.iw[4] ;
 wire \top_I.branch[7].block[15].um_I.iw[5] ;
 wire \top_I.branch[7].block[15].um_I.iw[6] ;
 wire \top_I.branch[7].block[15].um_I.iw[7] ;
 wire \top_I.branch[7].block[15].um_I.iw[8] ;
 wire \top_I.branch[7].block[15].um_I.iw[9] ;
 wire \top_I.branch[7].block[15].um_I.k_zero ;
 wire \top_I.branch[7].block[15].um_I.pg_vdd ;
 wire \top_I.branch[7].block[1].um_I.ana[0] ;
 wire \top_I.branch[7].block[1].um_I.ana[1] ;
 wire \top_I.branch[7].block[1].um_I.ana[2] ;
 wire \top_I.branch[7].block[1].um_I.ana[3] ;
 wire \top_I.branch[7].block[1].um_I.ana[4] ;
 wire \top_I.branch[7].block[1].um_I.ana[5] ;
 wire \top_I.branch[7].block[1].um_I.ana[6] ;
 wire \top_I.branch[7].block[1].um_I.ana[7] ;
 wire \top_I.branch[7].block[1].um_I.clk ;
 wire \top_I.branch[7].block[1].um_I.ena ;
 wire \top_I.branch[7].block[1].um_I.iw[10] ;
 wire \top_I.branch[7].block[1].um_I.iw[11] ;
 wire \top_I.branch[7].block[1].um_I.iw[12] ;
 wire \top_I.branch[7].block[1].um_I.iw[13] ;
 wire \top_I.branch[7].block[1].um_I.iw[14] ;
 wire \top_I.branch[7].block[1].um_I.iw[15] ;
 wire \top_I.branch[7].block[1].um_I.iw[16] ;
 wire \top_I.branch[7].block[1].um_I.iw[17] ;
 wire \top_I.branch[7].block[1].um_I.iw[1] ;
 wire \top_I.branch[7].block[1].um_I.iw[2] ;
 wire \top_I.branch[7].block[1].um_I.iw[3] ;
 wire \top_I.branch[7].block[1].um_I.iw[4] ;
 wire \top_I.branch[7].block[1].um_I.iw[5] ;
 wire \top_I.branch[7].block[1].um_I.iw[6] ;
 wire \top_I.branch[7].block[1].um_I.iw[7] ;
 wire \top_I.branch[7].block[1].um_I.iw[8] ;
 wire \top_I.branch[7].block[1].um_I.iw[9] ;
 wire \top_I.branch[7].block[1].um_I.k_zero ;
 wire \top_I.branch[7].block[1].um_I.pg_vdd ;
 wire \top_I.branch[7].block[2].um_I.ana[0] ;
 wire \top_I.branch[7].block[2].um_I.ana[1] ;
 wire \top_I.branch[7].block[2].um_I.ana[2] ;
 wire \top_I.branch[7].block[2].um_I.ana[3] ;
 wire \top_I.branch[7].block[2].um_I.ana[4] ;
 wire \top_I.branch[7].block[2].um_I.ana[5] ;
 wire \top_I.branch[7].block[2].um_I.ana[6] ;
 wire \top_I.branch[7].block[2].um_I.ana[7] ;
 wire \top_I.branch[7].block[2].um_I.clk ;
 wire \top_I.branch[7].block[2].um_I.ena ;
 wire \top_I.branch[7].block[2].um_I.iw[10] ;
 wire \top_I.branch[7].block[2].um_I.iw[11] ;
 wire \top_I.branch[7].block[2].um_I.iw[12] ;
 wire \top_I.branch[7].block[2].um_I.iw[13] ;
 wire \top_I.branch[7].block[2].um_I.iw[14] ;
 wire \top_I.branch[7].block[2].um_I.iw[15] ;
 wire \top_I.branch[7].block[2].um_I.iw[16] ;
 wire \top_I.branch[7].block[2].um_I.iw[17] ;
 wire \top_I.branch[7].block[2].um_I.iw[1] ;
 wire \top_I.branch[7].block[2].um_I.iw[2] ;
 wire \top_I.branch[7].block[2].um_I.iw[3] ;
 wire \top_I.branch[7].block[2].um_I.iw[4] ;
 wire \top_I.branch[7].block[2].um_I.iw[5] ;
 wire \top_I.branch[7].block[2].um_I.iw[6] ;
 wire \top_I.branch[7].block[2].um_I.iw[7] ;
 wire \top_I.branch[7].block[2].um_I.iw[8] ;
 wire \top_I.branch[7].block[2].um_I.iw[9] ;
 wire \top_I.branch[7].block[2].um_I.k_zero ;
 wire \top_I.branch[7].block[2].um_I.pg_vdd ;
 wire \top_I.branch[7].block[3].um_I.ana[0] ;
 wire \top_I.branch[7].block[3].um_I.ana[1] ;
 wire \top_I.branch[7].block[3].um_I.ana[2] ;
 wire \top_I.branch[7].block[3].um_I.ana[3] ;
 wire \top_I.branch[7].block[3].um_I.ana[4] ;
 wire \top_I.branch[7].block[3].um_I.ana[5] ;
 wire \top_I.branch[7].block[3].um_I.ana[6] ;
 wire \top_I.branch[7].block[3].um_I.ana[7] ;
 wire \top_I.branch[7].block[3].um_I.clk ;
 wire \top_I.branch[7].block[3].um_I.ena ;
 wire \top_I.branch[7].block[3].um_I.iw[10] ;
 wire \top_I.branch[7].block[3].um_I.iw[11] ;
 wire \top_I.branch[7].block[3].um_I.iw[12] ;
 wire \top_I.branch[7].block[3].um_I.iw[13] ;
 wire \top_I.branch[7].block[3].um_I.iw[14] ;
 wire \top_I.branch[7].block[3].um_I.iw[15] ;
 wire \top_I.branch[7].block[3].um_I.iw[16] ;
 wire \top_I.branch[7].block[3].um_I.iw[17] ;
 wire \top_I.branch[7].block[3].um_I.iw[1] ;
 wire \top_I.branch[7].block[3].um_I.iw[2] ;
 wire \top_I.branch[7].block[3].um_I.iw[3] ;
 wire \top_I.branch[7].block[3].um_I.iw[4] ;
 wire \top_I.branch[7].block[3].um_I.iw[5] ;
 wire \top_I.branch[7].block[3].um_I.iw[6] ;
 wire \top_I.branch[7].block[3].um_I.iw[7] ;
 wire \top_I.branch[7].block[3].um_I.iw[8] ;
 wire \top_I.branch[7].block[3].um_I.iw[9] ;
 wire \top_I.branch[7].block[3].um_I.k_zero ;
 wire \top_I.branch[7].block[3].um_I.pg_vdd ;
 wire \top_I.branch[7].block[4].um_I.ana[0] ;
 wire \top_I.branch[7].block[4].um_I.ana[1] ;
 wire \top_I.branch[7].block[4].um_I.ana[2] ;
 wire \top_I.branch[7].block[4].um_I.ana[3] ;
 wire \top_I.branch[7].block[4].um_I.ana[4] ;
 wire \top_I.branch[7].block[4].um_I.ana[5] ;
 wire \top_I.branch[7].block[4].um_I.ana[6] ;
 wire \top_I.branch[7].block[4].um_I.ana[7] ;
 wire \top_I.branch[7].block[4].um_I.clk ;
 wire \top_I.branch[7].block[4].um_I.ena ;
 wire \top_I.branch[7].block[4].um_I.iw[10] ;
 wire \top_I.branch[7].block[4].um_I.iw[11] ;
 wire \top_I.branch[7].block[4].um_I.iw[12] ;
 wire \top_I.branch[7].block[4].um_I.iw[13] ;
 wire \top_I.branch[7].block[4].um_I.iw[14] ;
 wire \top_I.branch[7].block[4].um_I.iw[15] ;
 wire \top_I.branch[7].block[4].um_I.iw[16] ;
 wire \top_I.branch[7].block[4].um_I.iw[17] ;
 wire \top_I.branch[7].block[4].um_I.iw[1] ;
 wire \top_I.branch[7].block[4].um_I.iw[2] ;
 wire \top_I.branch[7].block[4].um_I.iw[3] ;
 wire \top_I.branch[7].block[4].um_I.iw[4] ;
 wire \top_I.branch[7].block[4].um_I.iw[5] ;
 wire \top_I.branch[7].block[4].um_I.iw[6] ;
 wire \top_I.branch[7].block[4].um_I.iw[7] ;
 wire \top_I.branch[7].block[4].um_I.iw[8] ;
 wire \top_I.branch[7].block[4].um_I.iw[9] ;
 wire \top_I.branch[7].block[4].um_I.k_zero ;
 wire \top_I.branch[7].block[4].um_I.pg_vdd ;
 wire \top_I.branch[7].block[5].um_I.ana[0] ;
 wire \top_I.branch[7].block[5].um_I.ana[1] ;
 wire \top_I.branch[7].block[5].um_I.ana[2] ;
 wire \top_I.branch[7].block[5].um_I.ana[3] ;
 wire \top_I.branch[7].block[5].um_I.ana[4] ;
 wire \top_I.branch[7].block[5].um_I.ana[5] ;
 wire \top_I.branch[7].block[5].um_I.ana[6] ;
 wire \top_I.branch[7].block[5].um_I.ana[7] ;
 wire \top_I.branch[7].block[5].um_I.clk ;
 wire \top_I.branch[7].block[5].um_I.ena ;
 wire \top_I.branch[7].block[5].um_I.iw[10] ;
 wire \top_I.branch[7].block[5].um_I.iw[11] ;
 wire \top_I.branch[7].block[5].um_I.iw[12] ;
 wire \top_I.branch[7].block[5].um_I.iw[13] ;
 wire \top_I.branch[7].block[5].um_I.iw[14] ;
 wire \top_I.branch[7].block[5].um_I.iw[15] ;
 wire \top_I.branch[7].block[5].um_I.iw[16] ;
 wire \top_I.branch[7].block[5].um_I.iw[17] ;
 wire \top_I.branch[7].block[5].um_I.iw[1] ;
 wire \top_I.branch[7].block[5].um_I.iw[2] ;
 wire \top_I.branch[7].block[5].um_I.iw[3] ;
 wire \top_I.branch[7].block[5].um_I.iw[4] ;
 wire \top_I.branch[7].block[5].um_I.iw[5] ;
 wire \top_I.branch[7].block[5].um_I.iw[6] ;
 wire \top_I.branch[7].block[5].um_I.iw[7] ;
 wire \top_I.branch[7].block[5].um_I.iw[8] ;
 wire \top_I.branch[7].block[5].um_I.iw[9] ;
 wire \top_I.branch[7].block[5].um_I.k_zero ;
 wire \top_I.branch[7].block[5].um_I.pg_vdd ;
 wire \top_I.branch[7].block[6].um_I.ana[0] ;
 wire \top_I.branch[7].block[6].um_I.ana[1] ;
 wire \top_I.branch[7].block[6].um_I.ana[2] ;
 wire \top_I.branch[7].block[6].um_I.ana[3] ;
 wire \top_I.branch[7].block[6].um_I.ana[4] ;
 wire \top_I.branch[7].block[6].um_I.ana[5] ;
 wire \top_I.branch[7].block[6].um_I.ana[6] ;
 wire \top_I.branch[7].block[6].um_I.ana[7] ;
 wire \top_I.branch[7].block[6].um_I.clk ;
 wire \top_I.branch[7].block[6].um_I.ena ;
 wire \top_I.branch[7].block[6].um_I.iw[10] ;
 wire \top_I.branch[7].block[6].um_I.iw[11] ;
 wire \top_I.branch[7].block[6].um_I.iw[12] ;
 wire \top_I.branch[7].block[6].um_I.iw[13] ;
 wire \top_I.branch[7].block[6].um_I.iw[14] ;
 wire \top_I.branch[7].block[6].um_I.iw[15] ;
 wire \top_I.branch[7].block[6].um_I.iw[16] ;
 wire \top_I.branch[7].block[6].um_I.iw[17] ;
 wire \top_I.branch[7].block[6].um_I.iw[1] ;
 wire \top_I.branch[7].block[6].um_I.iw[2] ;
 wire \top_I.branch[7].block[6].um_I.iw[3] ;
 wire \top_I.branch[7].block[6].um_I.iw[4] ;
 wire \top_I.branch[7].block[6].um_I.iw[5] ;
 wire \top_I.branch[7].block[6].um_I.iw[6] ;
 wire \top_I.branch[7].block[6].um_I.iw[7] ;
 wire \top_I.branch[7].block[6].um_I.iw[8] ;
 wire \top_I.branch[7].block[6].um_I.iw[9] ;
 wire \top_I.branch[7].block[6].um_I.k_zero ;
 wire \top_I.branch[7].block[6].um_I.pg_vdd ;
 wire \top_I.branch[7].block[7].um_I.ana[0] ;
 wire \top_I.branch[7].block[7].um_I.ana[1] ;
 wire \top_I.branch[7].block[7].um_I.ana[2] ;
 wire \top_I.branch[7].block[7].um_I.ana[3] ;
 wire \top_I.branch[7].block[7].um_I.ana[4] ;
 wire \top_I.branch[7].block[7].um_I.ana[5] ;
 wire \top_I.branch[7].block[7].um_I.ana[6] ;
 wire \top_I.branch[7].block[7].um_I.ana[7] ;
 wire \top_I.branch[7].block[7].um_I.clk ;
 wire \top_I.branch[7].block[7].um_I.ena ;
 wire \top_I.branch[7].block[7].um_I.iw[10] ;
 wire \top_I.branch[7].block[7].um_I.iw[11] ;
 wire \top_I.branch[7].block[7].um_I.iw[12] ;
 wire \top_I.branch[7].block[7].um_I.iw[13] ;
 wire \top_I.branch[7].block[7].um_I.iw[14] ;
 wire \top_I.branch[7].block[7].um_I.iw[15] ;
 wire \top_I.branch[7].block[7].um_I.iw[16] ;
 wire \top_I.branch[7].block[7].um_I.iw[17] ;
 wire \top_I.branch[7].block[7].um_I.iw[1] ;
 wire \top_I.branch[7].block[7].um_I.iw[2] ;
 wire \top_I.branch[7].block[7].um_I.iw[3] ;
 wire \top_I.branch[7].block[7].um_I.iw[4] ;
 wire \top_I.branch[7].block[7].um_I.iw[5] ;
 wire \top_I.branch[7].block[7].um_I.iw[6] ;
 wire \top_I.branch[7].block[7].um_I.iw[7] ;
 wire \top_I.branch[7].block[7].um_I.iw[8] ;
 wire \top_I.branch[7].block[7].um_I.iw[9] ;
 wire \top_I.branch[7].block[7].um_I.k_zero ;
 wire \top_I.branch[7].block[7].um_I.pg_vdd ;
 wire \top_I.branch[7].block[8].um_I.ana[0] ;
 wire \top_I.branch[7].block[8].um_I.ana[1] ;
 wire \top_I.branch[7].block[8].um_I.ana[2] ;
 wire \top_I.branch[7].block[8].um_I.ana[3] ;
 wire \top_I.branch[7].block[8].um_I.ana[4] ;
 wire \top_I.branch[7].block[8].um_I.ana[5] ;
 wire \top_I.branch[7].block[8].um_I.ana[6] ;
 wire \top_I.branch[7].block[8].um_I.ana[7] ;
 wire \top_I.branch[7].block[8].um_I.clk ;
 wire \top_I.branch[7].block[8].um_I.ena ;
 wire \top_I.branch[7].block[8].um_I.iw[10] ;
 wire \top_I.branch[7].block[8].um_I.iw[11] ;
 wire \top_I.branch[7].block[8].um_I.iw[12] ;
 wire \top_I.branch[7].block[8].um_I.iw[13] ;
 wire \top_I.branch[7].block[8].um_I.iw[14] ;
 wire \top_I.branch[7].block[8].um_I.iw[15] ;
 wire \top_I.branch[7].block[8].um_I.iw[16] ;
 wire \top_I.branch[7].block[8].um_I.iw[17] ;
 wire \top_I.branch[7].block[8].um_I.iw[1] ;
 wire \top_I.branch[7].block[8].um_I.iw[2] ;
 wire \top_I.branch[7].block[8].um_I.iw[3] ;
 wire \top_I.branch[7].block[8].um_I.iw[4] ;
 wire \top_I.branch[7].block[8].um_I.iw[5] ;
 wire \top_I.branch[7].block[8].um_I.iw[6] ;
 wire \top_I.branch[7].block[8].um_I.iw[7] ;
 wire \top_I.branch[7].block[8].um_I.iw[8] ;
 wire \top_I.branch[7].block[8].um_I.iw[9] ;
 wire \top_I.branch[7].block[8].um_I.k_zero ;
 wire \top_I.branch[7].block[8].um_I.pg_vdd ;
 wire \top_I.branch[7].block[9].um_I.ana[0] ;
 wire \top_I.branch[7].block[9].um_I.ana[1] ;
 wire \top_I.branch[7].block[9].um_I.ana[2] ;
 wire \top_I.branch[7].block[9].um_I.ana[3] ;
 wire \top_I.branch[7].block[9].um_I.ana[4] ;
 wire \top_I.branch[7].block[9].um_I.ana[5] ;
 wire \top_I.branch[7].block[9].um_I.ana[6] ;
 wire \top_I.branch[7].block[9].um_I.ana[7] ;
 wire \top_I.branch[7].block[9].um_I.clk ;
 wire \top_I.branch[7].block[9].um_I.ena ;
 wire \top_I.branch[7].block[9].um_I.iw[10] ;
 wire \top_I.branch[7].block[9].um_I.iw[11] ;
 wire \top_I.branch[7].block[9].um_I.iw[12] ;
 wire \top_I.branch[7].block[9].um_I.iw[13] ;
 wire \top_I.branch[7].block[9].um_I.iw[14] ;
 wire \top_I.branch[7].block[9].um_I.iw[15] ;
 wire \top_I.branch[7].block[9].um_I.iw[16] ;
 wire \top_I.branch[7].block[9].um_I.iw[17] ;
 wire \top_I.branch[7].block[9].um_I.iw[1] ;
 wire \top_I.branch[7].block[9].um_I.iw[2] ;
 wire \top_I.branch[7].block[9].um_I.iw[3] ;
 wire \top_I.branch[7].block[9].um_I.iw[4] ;
 wire \top_I.branch[7].block[9].um_I.iw[5] ;
 wire \top_I.branch[7].block[9].um_I.iw[6] ;
 wire \top_I.branch[7].block[9].um_I.iw[7] ;
 wire \top_I.branch[7].block[9].um_I.iw[8] ;
 wire \top_I.branch[7].block[9].um_I.iw[9] ;
 wire \top_I.branch[7].block[9].um_I.k_zero ;
 wire \top_I.branch[7].block[9].um_I.pg_vdd ;
 wire \top_I.branch[7].l_addr[0] ;
 wire \top_I.branch[7].l_addr[2] ;
 wire \top_I.branch[8].block[0].um_I.ana[0] ;
 wire \top_I.branch[8].block[0].um_I.ana[1] ;
 wire \top_I.branch[8].block[0].um_I.ana[2] ;
 wire \top_I.branch[8].block[0].um_I.ana[3] ;
 wire \top_I.branch[8].block[0].um_I.ana[4] ;
 wire \top_I.branch[8].block[0].um_I.ana[5] ;
 wire \top_I.branch[8].block[0].um_I.ana[6] ;
 wire \top_I.branch[8].block[0].um_I.ana[7] ;
 wire \top_I.branch[8].block[0].um_I.clk ;
 wire \top_I.branch[8].block[0].um_I.ena ;
 wire \top_I.branch[8].block[0].um_I.iw[10] ;
 wire \top_I.branch[8].block[0].um_I.iw[11] ;
 wire \top_I.branch[8].block[0].um_I.iw[12] ;
 wire \top_I.branch[8].block[0].um_I.iw[13] ;
 wire \top_I.branch[8].block[0].um_I.iw[14] ;
 wire \top_I.branch[8].block[0].um_I.iw[15] ;
 wire \top_I.branch[8].block[0].um_I.iw[16] ;
 wire \top_I.branch[8].block[0].um_I.iw[17] ;
 wire \top_I.branch[8].block[0].um_I.iw[1] ;
 wire \top_I.branch[8].block[0].um_I.iw[2] ;
 wire \top_I.branch[8].block[0].um_I.iw[3] ;
 wire \top_I.branch[8].block[0].um_I.iw[4] ;
 wire \top_I.branch[8].block[0].um_I.iw[5] ;
 wire \top_I.branch[8].block[0].um_I.iw[6] ;
 wire \top_I.branch[8].block[0].um_I.iw[7] ;
 wire \top_I.branch[8].block[0].um_I.iw[8] ;
 wire \top_I.branch[8].block[0].um_I.iw[9] ;
 wire \top_I.branch[8].block[0].um_I.k_zero ;
 wire \top_I.branch[8].block[0].um_I.pg_vdd ;
 wire \top_I.branch[8].block[10].um_I.ana[0] ;
 wire \top_I.branch[8].block[10].um_I.ana[1] ;
 wire \top_I.branch[8].block[10].um_I.ana[2] ;
 wire \top_I.branch[8].block[10].um_I.ana[3] ;
 wire \top_I.branch[8].block[10].um_I.ana[4] ;
 wire \top_I.branch[8].block[10].um_I.ana[5] ;
 wire \top_I.branch[8].block[10].um_I.ana[6] ;
 wire \top_I.branch[8].block[10].um_I.ana[7] ;
 wire \top_I.branch[8].block[10].um_I.clk ;
 wire \top_I.branch[8].block[10].um_I.ena ;
 wire \top_I.branch[8].block[10].um_I.iw[10] ;
 wire \top_I.branch[8].block[10].um_I.iw[11] ;
 wire \top_I.branch[8].block[10].um_I.iw[12] ;
 wire \top_I.branch[8].block[10].um_I.iw[13] ;
 wire \top_I.branch[8].block[10].um_I.iw[14] ;
 wire \top_I.branch[8].block[10].um_I.iw[15] ;
 wire \top_I.branch[8].block[10].um_I.iw[16] ;
 wire \top_I.branch[8].block[10].um_I.iw[17] ;
 wire \top_I.branch[8].block[10].um_I.iw[1] ;
 wire \top_I.branch[8].block[10].um_I.iw[2] ;
 wire \top_I.branch[8].block[10].um_I.iw[3] ;
 wire \top_I.branch[8].block[10].um_I.iw[4] ;
 wire \top_I.branch[8].block[10].um_I.iw[5] ;
 wire \top_I.branch[8].block[10].um_I.iw[6] ;
 wire \top_I.branch[8].block[10].um_I.iw[7] ;
 wire \top_I.branch[8].block[10].um_I.iw[8] ;
 wire \top_I.branch[8].block[10].um_I.iw[9] ;
 wire \top_I.branch[8].block[10].um_I.k_zero ;
 wire \top_I.branch[8].block[10].um_I.pg_vdd ;
 wire \top_I.branch[8].block[11].um_I.ana[0] ;
 wire \top_I.branch[8].block[11].um_I.ana[1] ;
 wire \top_I.branch[8].block[11].um_I.ana[2] ;
 wire \top_I.branch[8].block[11].um_I.ana[3] ;
 wire \top_I.branch[8].block[11].um_I.ana[4] ;
 wire \top_I.branch[8].block[11].um_I.ana[5] ;
 wire \top_I.branch[8].block[11].um_I.ana[6] ;
 wire \top_I.branch[8].block[11].um_I.ana[7] ;
 wire \top_I.branch[8].block[11].um_I.clk ;
 wire \top_I.branch[8].block[11].um_I.ena ;
 wire \top_I.branch[8].block[11].um_I.iw[10] ;
 wire \top_I.branch[8].block[11].um_I.iw[11] ;
 wire \top_I.branch[8].block[11].um_I.iw[12] ;
 wire \top_I.branch[8].block[11].um_I.iw[13] ;
 wire \top_I.branch[8].block[11].um_I.iw[14] ;
 wire \top_I.branch[8].block[11].um_I.iw[15] ;
 wire \top_I.branch[8].block[11].um_I.iw[16] ;
 wire \top_I.branch[8].block[11].um_I.iw[17] ;
 wire \top_I.branch[8].block[11].um_I.iw[1] ;
 wire \top_I.branch[8].block[11].um_I.iw[2] ;
 wire \top_I.branch[8].block[11].um_I.iw[3] ;
 wire \top_I.branch[8].block[11].um_I.iw[4] ;
 wire \top_I.branch[8].block[11].um_I.iw[5] ;
 wire \top_I.branch[8].block[11].um_I.iw[6] ;
 wire \top_I.branch[8].block[11].um_I.iw[7] ;
 wire \top_I.branch[8].block[11].um_I.iw[8] ;
 wire \top_I.branch[8].block[11].um_I.iw[9] ;
 wire \top_I.branch[8].block[11].um_I.k_zero ;
 wire \top_I.branch[8].block[11].um_I.pg_vdd ;
 wire \top_I.branch[8].block[12].um_I.ana[0] ;
 wire \top_I.branch[8].block[12].um_I.ana[1] ;
 wire \top_I.branch[8].block[12].um_I.ana[2] ;
 wire \top_I.branch[8].block[12].um_I.ana[3] ;
 wire \top_I.branch[8].block[12].um_I.ana[4] ;
 wire \top_I.branch[8].block[12].um_I.ana[5] ;
 wire \top_I.branch[8].block[12].um_I.ana[6] ;
 wire \top_I.branch[8].block[12].um_I.ana[7] ;
 wire \top_I.branch[8].block[12].um_I.clk ;
 wire \top_I.branch[8].block[12].um_I.ena ;
 wire \top_I.branch[8].block[12].um_I.iw[10] ;
 wire \top_I.branch[8].block[12].um_I.iw[11] ;
 wire \top_I.branch[8].block[12].um_I.iw[12] ;
 wire \top_I.branch[8].block[12].um_I.iw[13] ;
 wire \top_I.branch[8].block[12].um_I.iw[14] ;
 wire \top_I.branch[8].block[12].um_I.iw[15] ;
 wire \top_I.branch[8].block[12].um_I.iw[16] ;
 wire \top_I.branch[8].block[12].um_I.iw[17] ;
 wire \top_I.branch[8].block[12].um_I.iw[1] ;
 wire \top_I.branch[8].block[12].um_I.iw[2] ;
 wire \top_I.branch[8].block[12].um_I.iw[3] ;
 wire \top_I.branch[8].block[12].um_I.iw[4] ;
 wire \top_I.branch[8].block[12].um_I.iw[5] ;
 wire \top_I.branch[8].block[12].um_I.iw[6] ;
 wire \top_I.branch[8].block[12].um_I.iw[7] ;
 wire \top_I.branch[8].block[12].um_I.iw[8] ;
 wire \top_I.branch[8].block[12].um_I.iw[9] ;
 wire \top_I.branch[8].block[12].um_I.k_zero ;
 wire \top_I.branch[8].block[12].um_I.pg_vdd ;
 wire \top_I.branch[8].block[13].um_I.ana[0] ;
 wire \top_I.branch[8].block[13].um_I.ana[1] ;
 wire \top_I.branch[8].block[13].um_I.ana[2] ;
 wire \top_I.branch[8].block[13].um_I.ana[3] ;
 wire \top_I.branch[8].block[13].um_I.ana[4] ;
 wire \top_I.branch[8].block[13].um_I.ana[5] ;
 wire \top_I.branch[8].block[13].um_I.ana[6] ;
 wire \top_I.branch[8].block[13].um_I.ana[7] ;
 wire \top_I.branch[8].block[13].um_I.clk ;
 wire \top_I.branch[8].block[13].um_I.ena ;
 wire \top_I.branch[8].block[13].um_I.iw[10] ;
 wire \top_I.branch[8].block[13].um_I.iw[11] ;
 wire \top_I.branch[8].block[13].um_I.iw[12] ;
 wire \top_I.branch[8].block[13].um_I.iw[13] ;
 wire \top_I.branch[8].block[13].um_I.iw[14] ;
 wire \top_I.branch[8].block[13].um_I.iw[15] ;
 wire \top_I.branch[8].block[13].um_I.iw[16] ;
 wire \top_I.branch[8].block[13].um_I.iw[17] ;
 wire \top_I.branch[8].block[13].um_I.iw[1] ;
 wire \top_I.branch[8].block[13].um_I.iw[2] ;
 wire \top_I.branch[8].block[13].um_I.iw[3] ;
 wire \top_I.branch[8].block[13].um_I.iw[4] ;
 wire \top_I.branch[8].block[13].um_I.iw[5] ;
 wire \top_I.branch[8].block[13].um_I.iw[6] ;
 wire \top_I.branch[8].block[13].um_I.iw[7] ;
 wire \top_I.branch[8].block[13].um_I.iw[8] ;
 wire \top_I.branch[8].block[13].um_I.iw[9] ;
 wire \top_I.branch[8].block[13].um_I.k_zero ;
 wire \top_I.branch[8].block[13].um_I.pg_vdd ;
 wire \top_I.branch[8].block[14].um_I.ana[0] ;
 wire \top_I.branch[8].block[14].um_I.ana[1] ;
 wire \top_I.branch[8].block[14].um_I.ana[2] ;
 wire \top_I.branch[8].block[14].um_I.ana[3] ;
 wire \top_I.branch[8].block[14].um_I.ana[4] ;
 wire \top_I.branch[8].block[14].um_I.ana[5] ;
 wire \top_I.branch[8].block[14].um_I.ana[6] ;
 wire \top_I.branch[8].block[14].um_I.ana[7] ;
 wire \top_I.branch[8].block[14].um_I.clk ;
 wire \top_I.branch[8].block[14].um_I.ena ;
 wire \top_I.branch[8].block[14].um_I.iw[10] ;
 wire \top_I.branch[8].block[14].um_I.iw[11] ;
 wire \top_I.branch[8].block[14].um_I.iw[12] ;
 wire \top_I.branch[8].block[14].um_I.iw[13] ;
 wire \top_I.branch[8].block[14].um_I.iw[14] ;
 wire \top_I.branch[8].block[14].um_I.iw[15] ;
 wire \top_I.branch[8].block[14].um_I.iw[16] ;
 wire \top_I.branch[8].block[14].um_I.iw[17] ;
 wire \top_I.branch[8].block[14].um_I.iw[1] ;
 wire \top_I.branch[8].block[14].um_I.iw[2] ;
 wire \top_I.branch[8].block[14].um_I.iw[3] ;
 wire \top_I.branch[8].block[14].um_I.iw[4] ;
 wire \top_I.branch[8].block[14].um_I.iw[5] ;
 wire \top_I.branch[8].block[14].um_I.iw[6] ;
 wire \top_I.branch[8].block[14].um_I.iw[7] ;
 wire \top_I.branch[8].block[14].um_I.iw[8] ;
 wire \top_I.branch[8].block[14].um_I.iw[9] ;
 wire \top_I.branch[8].block[14].um_I.k_zero ;
 wire \top_I.branch[8].block[14].um_I.pg_vdd ;
 wire \top_I.branch[8].block[15].um_I.ana[0] ;
 wire \top_I.branch[8].block[15].um_I.ana[1] ;
 wire \top_I.branch[8].block[15].um_I.ana[2] ;
 wire \top_I.branch[8].block[15].um_I.ana[3] ;
 wire \top_I.branch[8].block[15].um_I.ana[4] ;
 wire \top_I.branch[8].block[15].um_I.ana[5] ;
 wire \top_I.branch[8].block[15].um_I.ana[6] ;
 wire \top_I.branch[8].block[15].um_I.ana[7] ;
 wire \top_I.branch[8].block[15].um_I.clk ;
 wire \top_I.branch[8].block[15].um_I.ena ;
 wire \top_I.branch[8].block[15].um_I.iw[10] ;
 wire \top_I.branch[8].block[15].um_I.iw[11] ;
 wire \top_I.branch[8].block[15].um_I.iw[12] ;
 wire \top_I.branch[8].block[15].um_I.iw[13] ;
 wire \top_I.branch[8].block[15].um_I.iw[14] ;
 wire \top_I.branch[8].block[15].um_I.iw[15] ;
 wire \top_I.branch[8].block[15].um_I.iw[16] ;
 wire \top_I.branch[8].block[15].um_I.iw[17] ;
 wire \top_I.branch[8].block[15].um_I.iw[1] ;
 wire \top_I.branch[8].block[15].um_I.iw[2] ;
 wire \top_I.branch[8].block[15].um_I.iw[3] ;
 wire \top_I.branch[8].block[15].um_I.iw[4] ;
 wire \top_I.branch[8].block[15].um_I.iw[5] ;
 wire \top_I.branch[8].block[15].um_I.iw[6] ;
 wire \top_I.branch[8].block[15].um_I.iw[7] ;
 wire \top_I.branch[8].block[15].um_I.iw[8] ;
 wire \top_I.branch[8].block[15].um_I.iw[9] ;
 wire \top_I.branch[8].block[15].um_I.k_zero ;
 wire \top_I.branch[8].block[15].um_I.pg_vdd ;
 wire \top_I.branch[8].block[1].um_I.ana[0] ;
 wire \top_I.branch[8].block[1].um_I.ana[1] ;
 wire \top_I.branch[8].block[1].um_I.ana[2] ;
 wire \top_I.branch[8].block[1].um_I.ana[3] ;
 wire \top_I.branch[8].block[1].um_I.ana[4] ;
 wire \top_I.branch[8].block[1].um_I.ana[5] ;
 wire \top_I.branch[8].block[1].um_I.ana[6] ;
 wire \top_I.branch[8].block[1].um_I.ana[7] ;
 wire \top_I.branch[8].block[1].um_I.clk ;
 wire \top_I.branch[8].block[1].um_I.ena ;
 wire \top_I.branch[8].block[1].um_I.iw[10] ;
 wire \top_I.branch[8].block[1].um_I.iw[11] ;
 wire \top_I.branch[8].block[1].um_I.iw[12] ;
 wire \top_I.branch[8].block[1].um_I.iw[13] ;
 wire \top_I.branch[8].block[1].um_I.iw[14] ;
 wire \top_I.branch[8].block[1].um_I.iw[15] ;
 wire \top_I.branch[8].block[1].um_I.iw[16] ;
 wire \top_I.branch[8].block[1].um_I.iw[17] ;
 wire \top_I.branch[8].block[1].um_I.iw[1] ;
 wire \top_I.branch[8].block[1].um_I.iw[2] ;
 wire \top_I.branch[8].block[1].um_I.iw[3] ;
 wire \top_I.branch[8].block[1].um_I.iw[4] ;
 wire \top_I.branch[8].block[1].um_I.iw[5] ;
 wire \top_I.branch[8].block[1].um_I.iw[6] ;
 wire \top_I.branch[8].block[1].um_I.iw[7] ;
 wire \top_I.branch[8].block[1].um_I.iw[8] ;
 wire \top_I.branch[8].block[1].um_I.iw[9] ;
 wire \top_I.branch[8].block[1].um_I.k_zero ;
 wire \top_I.branch[8].block[1].um_I.pg_vdd ;
 wire \top_I.branch[8].block[2].um_I.ana[0] ;
 wire \top_I.branch[8].block[2].um_I.ana[1] ;
 wire \top_I.branch[8].block[2].um_I.ana[2] ;
 wire \top_I.branch[8].block[2].um_I.ana[3] ;
 wire \top_I.branch[8].block[2].um_I.ana[4] ;
 wire \top_I.branch[8].block[2].um_I.ana[5] ;
 wire \top_I.branch[8].block[2].um_I.ana[6] ;
 wire \top_I.branch[8].block[2].um_I.ana[7] ;
 wire \top_I.branch[8].block[2].um_I.clk ;
 wire \top_I.branch[8].block[2].um_I.ena ;
 wire \top_I.branch[8].block[2].um_I.iw[10] ;
 wire \top_I.branch[8].block[2].um_I.iw[11] ;
 wire \top_I.branch[8].block[2].um_I.iw[12] ;
 wire \top_I.branch[8].block[2].um_I.iw[13] ;
 wire \top_I.branch[8].block[2].um_I.iw[14] ;
 wire \top_I.branch[8].block[2].um_I.iw[15] ;
 wire \top_I.branch[8].block[2].um_I.iw[16] ;
 wire \top_I.branch[8].block[2].um_I.iw[17] ;
 wire \top_I.branch[8].block[2].um_I.iw[1] ;
 wire \top_I.branch[8].block[2].um_I.iw[2] ;
 wire \top_I.branch[8].block[2].um_I.iw[3] ;
 wire \top_I.branch[8].block[2].um_I.iw[4] ;
 wire \top_I.branch[8].block[2].um_I.iw[5] ;
 wire \top_I.branch[8].block[2].um_I.iw[6] ;
 wire \top_I.branch[8].block[2].um_I.iw[7] ;
 wire \top_I.branch[8].block[2].um_I.iw[8] ;
 wire \top_I.branch[8].block[2].um_I.iw[9] ;
 wire \top_I.branch[8].block[2].um_I.k_zero ;
 wire \top_I.branch[8].block[2].um_I.pg_vdd ;
 wire \top_I.branch[8].block[3].um_I.ana[0] ;
 wire \top_I.branch[8].block[3].um_I.ana[1] ;
 wire \top_I.branch[8].block[3].um_I.ana[2] ;
 wire \top_I.branch[8].block[3].um_I.ana[3] ;
 wire \top_I.branch[8].block[3].um_I.ana[4] ;
 wire \top_I.branch[8].block[3].um_I.ana[5] ;
 wire \top_I.branch[8].block[3].um_I.ana[6] ;
 wire \top_I.branch[8].block[3].um_I.ana[7] ;
 wire \top_I.branch[8].block[3].um_I.clk ;
 wire \top_I.branch[8].block[3].um_I.ena ;
 wire \top_I.branch[8].block[3].um_I.iw[10] ;
 wire \top_I.branch[8].block[3].um_I.iw[11] ;
 wire \top_I.branch[8].block[3].um_I.iw[12] ;
 wire \top_I.branch[8].block[3].um_I.iw[13] ;
 wire \top_I.branch[8].block[3].um_I.iw[14] ;
 wire \top_I.branch[8].block[3].um_I.iw[15] ;
 wire \top_I.branch[8].block[3].um_I.iw[16] ;
 wire \top_I.branch[8].block[3].um_I.iw[17] ;
 wire \top_I.branch[8].block[3].um_I.iw[1] ;
 wire \top_I.branch[8].block[3].um_I.iw[2] ;
 wire \top_I.branch[8].block[3].um_I.iw[3] ;
 wire \top_I.branch[8].block[3].um_I.iw[4] ;
 wire \top_I.branch[8].block[3].um_I.iw[5] ;
 wire \top_I.branch[8].block[3].um_I.iw[6] ;
 wire \top_I.branch[8].block[3].um_I.iw[7] ;
 wire \top_I.branch[8].block[3].um_I.iw[8] ;
 wire \top_I.branch[8].block[3].um_I.iw[9] ;
 wire \top_I.branch[8].block[3].um_I.k_zero ;
 wire \top_I.branch[8].block[3].um_I.pg_vdd ;
 wire \top_I.branch[8].block[4].um_I.ana[0] ;
 wire \top_I.branch[8].block[4].um_I.ana[1] ;
 wire \top_I.branch[8].block[4].um_I.ana[2] ;
 wire \top_I.branch[8].block[4].um_I.ana[3] ;
 wire \top_I.branch[8].block[4].um_I.ana[4] ;
 wire \top_I.branch[8].block[4].um_I.ana[5] ;
 wire \top_I.branch[8].block[4].um_I.ana[6] ;
 wire \top_I.branch[8].block[4].um_I.ana[7] ;
 wire \top_I.branch[8].block[4].um_I.clk ;
 wire \top_I.branch[8].block[4].um_I.ena ;
 wire \top_I.branch[8].block[4].um_I.iw[10] ;
 wire \top_I.branch[8].block[4].um_I.iw[11] ;
 wire \top_I.branch[8].block[4].um_I.iw[12] ;
 wire \top_I.branch[8].block[4].um_I.iw[13] ;
 wire \top_I.branch[8].block[4].um_I.iw[14] ;
 wire \top_I.branch[8].block[4].um_I.iw[15] ;
 wire \top_I.branch[8].block[4].um_I.iw[16] ;
 wire \top_I.branch[8].block[4].um_I.iw[17] ;
 wire \top_I.branch[8].block[4].um_I.iw[1] ;
 wire \top_I.branch[8].block[4].um_I.iw[2] ;
 wire \top_I.branch[8].block[4].um_I.iw[3] ;
 wire \top_I.branch[8].block[4].um_I.iw[4] ;
 wire \top_I.branch[8].block[4].um_I.iw[5] ;
 wire \top_I.branch[8].block[4].um_I.iw[6] ;
 wire \top_I.branch[8].block[4].um_I.iw[7] ;
 wire \top_I.branch[8].block[4].um_I.iw[8] ;
 wire \top_I.branch[8].block[4].um_I.iw[9] ;
 wire \top_I.branch[8].block[4].um_I.k_zero ;
 wire \top_I.branch[8].block[4].um_I.pg_vdd ;
 wire \top_I.branch[8].block[5].um_I.ana[0] ;
 wire \top_I.branch[8].block[5].um_I.ana[1] ;
 wire \top_I.branch[8].block[5].um_I.ana[2] ;
 wire \top_I.branch[8].block[5].um_I.ana[3] ;
 wire \top_I.branch[8].block[5].um_I.ana[4] ;
 wire \top_I.branch[8].block[5].um_I.ana[5] ;
 wire \top_I.branch[8].block[5].um_I.ana[6] ;
 wire \top_I.branch[8].block[5].um_I.ana[7] ;
 wire \top_I.branch[8].block[5].um_I.clk ;
 wire \top_I.branch[8].block[5].um_I.ena ;
 wire \top_I.branch[8].block[5].um_I.iw[10] ;
 wire \top_I.branch[8].block[5].um_I.iw[11] ;
 wire \top_I.branch[8].block[5].um_I.iw[12] ;
 wire \top_I.branch[8].block[5].um_I.iw[13] ;
 wire \top_I.branch[8].block[5].um_I.iw[14] ;
 wire \top_I.branch[8].block[5].um_I.iw[15] ;
 wire \top_I.branch[8].block[5].um_I.iw[16] ;
 wire \top_I.branch[8].block[5].um_I.iw[17] ;
 wire \top_I.branch[8].block[5].um_I.iw[1] ;
 wire \top_I.branch[8].block[5].um_I.iw[2] ;
 wire \top_I.branch[8].block[5].um_I.iw[3] ;
 wire \top_I.branch[8].block[5].um_I.iw[4] ;
 wire \top_I.branch[8].block[5].um_I.iw[5] ;
 wire \top_I.branch[8].block[5].um_I.iw[6] ;
 wire \top_I.branch[8].block[5].um_I.iw[7] ;
 wire \top_I.branch[8].block[5].um_I.iw[8] ;
 wire \top_I.branch[8].block[5].um_I.iw[9] ;
 wire \top_I.branch[8].block[5].um_I.k_zero ;
 wire \top_I.branch[8].block[5].um_I.pg_vdd ;
 wire \top_I.branch[8].block[6].um_I.ana[0] ;
 wire \top_I.branch[8].block[6].um_I.ana[1] ;
 wire \top_I.branch[8].block[6].um_I.ana[2] ;
 wire \top_I.branch[8].block[6].um_I.ana[3] ;
 wire \top_I.branch[8].block[6].um_I.ana[4] ;
 wire \top_I.branch[8].block[6].um_I.ana[5] ;
 wire \top_I.branch[8].block[6].um_I.ana[6] ;
 wire \top_I.branch[8].block[6].um_I.ana[7] ;
 wire \top_I.branch[8].block[6].um_I.clk ;
 wire \top_I.branch[8].block[6].um_I.ena ;
 wire \top_I.branch[8].block[6].um_I.iw[10] ;
 wire \top_I.branch[8].block[6].um_I.iw[11] ;
 wire \top_I.branch[8].block[6].um_I.iw[12] ;
 wire \top_I.branch[8].block[6].um_I.iw[13] ;
 wire \top_I.branch[8].block[6].um_I.iw[14] ;
 wire \top_I.branch[8].block[6].um_I.iw[15] ;
 wire \top_I.branch[8].block[6].um_I.iw[16] ;
 wire \top_I.branch[8].block[6].um_I.iw[17] ;
 wire \top_I.branch[8].block[6].um_I.iw[1] ;
 wire \top_I.branch[8].block[6].um_I.iw[2] ;
 wire \top_I.branch[8].block[6].um_I.iw[3] ;
 wire \top_I.branch[8].block[6].um_I.iw[4] ;
 wire \top_I.branch[8].block[6].um_I.iw[5] ;
 wire \top_I.branch[8].block[6].um_I.iw[6] ;
 wire \top_I.branch[8].block[6].um_I.iw[7] ;
 wire \top_I.branch[8].block[6].um_I.iw[8] ;
 wire \top_I.branch[8].block[6].um_I.iw[9] ;
 wire \top_I.branch[8].block[6].um_I.k_zero ;
 wire \top_I.branch[8].block[6].um_I.pg_vdd ;
 wire \top_I.branch[8].block[7].um_I.ana[0] ;
 wire \top_I.branch[8].block[7].um_I.ana[1] ;
 wire \top_I.branch[8].block[7].um_I.ana[2] ;
 wire \top_I.branch[8].block[7].um_I.ana[3] ;
 wire \top_I.branch[8].block[7].um_I.ana[4] ;
 wire \top_I.branch[8].block[7].um_I.ana[5] ;
 wire \top_I.branch[8].block[7].um_I.ana[6] ;
 wire \top_I.branch[8].block[7].um_I.ana[7] ;
 wire \top_I.branch[8].block[7].um_I.clk ;
 wire \top_I.branch[8].block[7].um_I.ena ;
 wire \top_I.branch[8].block[7].um_I.iw[10] ;
 wire \top_I.branch[8].block[7].um_I.iw[11] ;
 wire \top_I.branch[8].block[7].um_I.iw[12] ;
 wire \top_I.branch[8].block[7].um_I.iw[13] ;
 wire \top_I.branch[8].block[7].um_I.iw[14] ;
 wire \top_I.branch[8].block[7].um_I.iw[15] ;
 wire \top_I.branch[8].block[7].um_I.iw[16] ;
 wire \top_I.branch[8].block[7].um_I.iw[17] ;
 wire \top_I.branch[8].block[7].um_I.iw[1] ;
 wire \top_I.branch[8].block[7].um_I.iw[2] ;
 wire \top_I.branch[8].block[7].um_I.iw[3] ;
 wire \top_I.branch[8].block[7].um_I.iw[4] ;
 wire \top_I.branch[8].block[7].um_I.iw[5] ;
 wire \top_I.branch[8].block[7].um_I.iw[6] ;
 wire \top_I.branch[8].block[7].um_I.iw[7] ;
 wire \top_I.branch[8].block[7].um_I.iw[8] ;
 wire \top_I.branch[8].block[7].um_I.iw[9] ;
 wire \top_I.branch[8].block[7].um_I.k_zero ;
 wire \top_I.branch[8].block[7].um_I.pg_vdd ;
 wire \top_I.branch[8].block[8].um_I.ana[0] ;
 wire \top_I.branch[8].block[8].um_I.ana[1] ;
 wire \top_I.branch[8].block[8].um_I.ana[2] ;
 wire \top_I.branch[8].block[8].um_I.ana[3] ;
 wire \top_I.branch[8].block[8].um_I.ana[4] ;
 wire \top_I.branch[8].block[8].um_I.ana[5] ;
 wire \top_I.branch[8].block[8].um_I.ana[6] ;
 wire \top_I.branch[8].block[8].um_I.ana[7] ;
 wire \top_I.branch[8].block[8].um_I.clk ;
 wire \top_I.branch[8].block[8].um_I.ena ;
 wire \top_I.branch[8].block[8].um_I.iw[10] ;
 wire \top_I.branch[8].block[8].um_I.iw[11] ;
 wire \top_I.branch[8].block[8].um_I.iw[12] ;
 wire \top_I.branch[8].block[8].um_I.iw[13] ;
 wire \top_I.branch[8].block[8].um_I.iw[14] ;
 wire \top_I.branch[8].block[8].um_I.iw[15] ;
 wire \top_I.branch[8].block[8].um_I.iw[16] ;
 wire \top_I.branch[8].block[8].um_I.iw[17] ;
 wire \top_I.branch[8].block[8].um_I.iw[1] ;
 wire \top_I.branch[8].block[8].um_I.iw[2] ;
 wire \top_I.branch[8].block[8].um_I.iw[3] ;
 wire \top_I.branch[8].block[8].um_I.iw[4] ;
 wire \top_I.branch[8].block[8].um_I.iw[5] ;
 wire \top_I.branch[8].block[8].um_I.iw[6] ;
 wire \top_I.branch[8].block[8].um_I.iw[7] ;
 wire \top_I.branch[8].block[8].um_I.iw[8] ;
 wire \top_I.branch[8].block[8].um_I.iw[9] ;
 wire \top_I.branch[8].block[8].um_I.k_zero ;
 wire \top_I.branch[8].block[8].um_I.pg_vdd ;
 wire \top_I.branch[8].block[9].um_I.ana[0] ;
 wire \top_I.branch[8].block[9].um_I.ana[1] ;
 wire \top_I.branch[8].block[9].um_I.ana[2] ;
 wire \top_I.branch[8].block[9].um_I.ana[3] ;
 wire \top_I.branch[8].block[9].um_I.ana[4] ;
 wire \top_I.branch[8].block[9].um_I.ana[5] ;
 wire \top_I.branch[8].block[9].um_I.ana[6] ;
 wire \top_I.branch[8].block[9].um_I.ana[7] ;
 wire \top_I.branch[8].block[9].um_I.clk ;
 wire \top_I.branch[8].block[9].um_I.ena ;
 wire \top_I.branch[8].block[9].um_I.iw[10] ;
 wire \top_I.branch[8].block[9].um_I.iw[11] ;
 wire \top_I.branch[8].block[9].um_I.iw[12] ;
 wire \top_I.branch[8].block[9].um_I.iw[13] ;
 wire \top_I.branch[8].block[9].um_I.iw[14] ;
 wire \top_I.branch[8].block[9].um_I.iw[15] ;
 wire \top_I.branch[8].block[9].um_I.iw[16] ;
 wire \top_I.branch[8].block[9].um_I.iw[17] ;
 wire \top_I.branch[8].block[9].um_I.iw[1] ;
 wire \top_I.branch[8].block[9].um_I.iw[2] ;
 wire \top_I.branch[8].block[9].um_I.iw[3] ;
 wire \top_I.branch[8].block[9].um_I.iw[4] ;
 wire \top_I.branch[8].block[9].um_I.iw[5] ;
 wire \top_I.branch[8].block[9].um_I.iw[6] ;
 wire \top_I.branch[8].block[9].um_I.iw[7] ;
 wire \top_I.branch[8].block[9].um_I.iw[8] ;
 wire \top_I.branch[8].block[9].um_I.iw[9] ;
 wire \top_I.branch[8].block[9].um_I.k_zero ;
 wire \top_I.branch[8].block[9].um_I.pg_vdd ;
 wire \top_I.branch[8].l_addr[0] ;
 wire \top_I.branch[8].l_addr[2] ;
 wire \top_I.branch[9].block[0].um_I.ana[0] ;
 wire \top_I.branch[9].block[0].um_I.ana[1] ;
 wire \top_I.branch[9].block[0].um_I.ana[2] ;
 wire \top_I.branch[9].block[0].um_I.ana[3] ;
 wire \top_I.branch[9].block[0].um_I.ana[4] ;
 wire \top_I.branch[9].block[0].um_I.ana[5] ;
 wire \top_I.branch[9].block[0].um_I.ana[6] ;
 wire \top_I.branch[9].block[0].um_I.ana[7] ;
 wire \top_I.branch[9].block[0].um_I.clk ;
 wire \top_I.branch[9].block[0].um_I.ena ;
 wire \top_I.branch[9].block[0].um_I.iw[10] ;
 wire \top_I.branch[9].block[0].um_I.iw[11] ;
 wire \top_I.branch[9].block[0].um_I.iw[12] ;
 wire \top_I.branch[9].block[0].um_I.iw[13] ;
 wire \top_I.branch[9].block[0].um_I.iw[14] ;
 wire \top_I.branch[9].block[0].um_I.iw[15] ;
 wire \top_I.branch[9].block[0].um_I.iw[16] ;
 wire \top_I.branch[9].block[0].um_I.iw[17] ;
 wire \top_I.branch[9].block[0].um_I.iw[1] ;
 wire \top_I.branch[9].block[0].um_I.iw[2] ;
 wire \top_I.branch[9].block[0].um_I.iw[3] ;
 wire \top_I.branch[9].block[0].um_I.iw[4] ;
 wire \top_I.branch[9].block[0].um_I.iw[5] ;
 wire \top_I.branch[9].block[0].um_I.iw[6] ;
 wire \top_I.branch[9].block[0].um_I.iw[7] ;
 wire \top_I.branch[9].block[0].um_I.iw[8] ;
 wire \top_I.branch[9].block[0].um_I.iw[9] ;
 wire \top_I.branch[9].block[0].um_I.k_zero ;
 wire \top_I.branch[9].block[0].um_I.pg_vdd ;
 wire \top_I.branch[9].block[10].um_I.ana[0] ;
 wire \top_I.branch[9].block[10].um_I.ana[1] ;
 wire \top_I.branch[9].block[10].um_I.ana[2] ;
 wire \top_I.branch[9].block[10].um_I.ana[3] ;
 wire \top_I.branch[9].block[10].um_I.ana[4] ;
 wire \top_I.branch[9].block[10].um_I.ana[5] ;
 wire \top_I.branch[9].block[10].um_I.ana[6] ;
 wire \top_I.branch[9].block[10].um_I.ana[7] ;
 wire \top_I.branch[9].block[10].um_I.clk ;
 wire \top_I.branch[9].block[10].um_I.ena ;
 wire \top_I.branch[9].block[10].um_I.iw[10] ;
 wire \top_I.branch[9].block[10].um_I.iw[11] ;
 wire \top_I.branch[9].block[10].um_I.iw[12] ;
 wire \top_I.branch[9].block[10].um_I.iw[13] ;
 wire \top_I.branch[9].block[10].um_I.iw[14] ;
 wire \top_I.branch[9].block[10].um_I.iw[15] ;
 wire \top_I.branch[9].block[10].um_I.iw[16] ;
 wire \top_I.branch[9].block[10].um_I.iw[17] ;
 wire \top_I.branch[9].block[10].um_I.iw[1] ;
 wire \top_I.branch[9].block[10].um_I.iw[2] ;
 wire \top_I.branch[9].block[10].um_I.iw[3] ;
 wire \top_I.branch[9].block[10].um_I.iw[4] ;
 wire \top_I.branch[9].block[10].um_I.iw[5] ;
 wire \top_I.branch[9].block[10].um_I.iw[6] ;
 wire \top_I.branch[9].block[10].um_I.iw[7] ;
 wire \top_I.branch[9].block[10].um_I.iw[8] ;
 wire \top_I.branch[9].block[10].um_I.iw[9] ;
 wire \top_I.branch[9].block[10].um_I.k_zero ;
 wire \top_I.branch[9].block[10].um_I.pg_vdd ;
 wire \top_I.branch[9].block[11].um_I.ana[0] ;
 wire \top_I.branch[9].block[11].um_I.ana[1] ;
 wire \top_I.branch[9].block[11].um_I.ana[2] ;
 wire \top_I.branch[9].block[11].um_I.ana[3] ;
 wire \top_I.branch[9].block[11].um_I.ana[4] ;
 wire \top_I.branch[9].block[11].um_I.ana[5] ;
 wire \top_I.branch[9].block[11].um_I.ana[6] ;
 wire \top_I.branch[9].block[11].um_I.ana[7] ;
 wire \top_I.branch[9].block[11].um_I.clk ;
 wire \top_I.branch[9].block[11].um_I.ena ;
 wire \top_I.branch[9].block[11].um_I.iw[10] ;
 wire \top_I.branch[9].block[11].um_I.iw[11] ;
 wire \top_I.branch[9].block[11].um_I.iw[12] ;
 wire \top_I.branch[9].block[11].um_I.iw[13] ;
 wire \top_I.branch[9].block[11].um_I.iw[14] ;
 wire \top_I.branch[9].block[11].um_I.iw[15] ;
 wire \top_I.branch[9].block[11].um_I.iw[16] ;
 wire \top_I.branch[9].block[11].um_I.iw[17] ;
 wire \top_I.branch[9].block[11].um_I.iw[1] ;
 wire \top_I.branch[9].block[11].um_I.iw[2] ;
 wire \top_I.branch[9].block[11].um_I.iw[3] ;
 wire \top_I.branch[9].block[11].um_I.iw[4] ;
 wire \top_I.branch[9].block[11].um_I.iw[5] ;
 wire \top_I.branch[9].block[11].um_I.iw[6] ;
 wire \top_I.branch[9].block[11].um_I.iw[7] ;
 wire \top_I.branch[9].block[11].um_I.iw[8] ;
 wire \top_I.branch[9].block[11].um_I.iw[9] ;
 wire \top_I.branch[9].block[11].um_I.k_zero ;
 wire \top_I.branch[9].block[11].um_I.pg_vdd ;
 wire \top_I.branch[9].block[12].um_I.ana[0] ;
 wire \top_I.branch[9].block[12].um_I.ana[1] ;
 wire \top_I.branch[9].block[12].um_I.ana[2] ;
 wire \top_I.branch[9].block[12].um_I.ana[3] ;
 wire \top_I.branch[9].block[12].um_I.ana[4] ;
 wire \top_I.branch[9].block[12].um_I.ana[5] ;
 wire \top_I.branch[9].block[12].um_I.ana[6] ;
 wire \top_I.branch[9].block[12].um_I.ana[7] ;
 wire \top_I.branch[9].block[12].um_I.clk ;
 wire \top_I.branch[9].block[12].um_I.ena ;
 wire \top_I.branch[9].block[12].um_I.iw[10] ;
 wire \top_I.branch[9].block[12].um_I.iw[11] ;
 wire \top_I.branch[9].block[12].um_I.iw[12] ;
 wire \top_I.branch[9].block[12].um_I.iw[13] ;
 wire \top_I.branch[9].block[12].um_I.iw[14] ;
 wire \top_I.branch[9].block[12].um_I.iw[15] ;
 wire \top_I.branch[9].block[12].um_I.iw[16] ;
 wire \top_I.branch[9].block[12].um_I.iw[17] ;
 wire \top_I.branch[9].block[12].um_I.iw[1] ;
 wire \top_I.branch[9].block[12].um_I.iw[2] ;
 wire \top_I.branch[9].block[12].um_I.iw[3] ;
 wire \top_I.branch[9].block[12].um_I.iw[4] ;
 wire \top_I.branch[9].block[12].um_I.iw[5] ;
 wire \top_I.branch[9].block[12].um_I.iw[6] ;
 wire \top_I.branch[9].block[12].um_I.iw[7] ;
 wire \top_I.branch[9].block[12].um_I.iw[8] ;
 wire \top_I.branch[9].block[12].um_I.iw[9] ;
 wire \top_I.branch[9].block[12].um_I.k_zero ;
 wire \top_I.branch[9].block[12].um_I.pg_vdd ;
 wire \top_I.branch[9].block[13].um_I.ana[0] ;
 wire \top_I.branch[9].block[13].um_I.ana[1] ;
 wire \top_I.branch[9].block[13].um_I.ana[2] ;
 wire \top_I.branch[9].block[13].um_I.ana[3] ;
 wire \top_I.branch[9].block[13].um_I.ana[4] ;
 wire \top_I.branch[9].block[13].um_I.ana[5] ;
 wire \top_I.branch[9].block[13].um_I.ana[6] ;
 wire \top_I.branch[9].block[13].um_I.ana[7] ;
 wire \top_I.branch[9].block[13].um_I.clk ;
 wire \top_I.branch[9].block[13].um_I.ena ;
 wire \top_I.branch[9].block[13].um_I.iw[10] ;
 wire \top_I.branch[9].block[13].um_I.iw[11] ;
 wire \top_I.branch[9].block[13].um_I.iw[12] ;
 wire \top_I.branch[9].block[13].um_I.iw[13] ;
 wire \top_I.branch[9].block[13].um_I.iw[14] ;
 wire \top_I.branch[9].block[13].um_I.iw[15] ;
 wire \top_I.branch[9].block[13].um_I.iw[16] ;
 wire \top_I.branch[9].block[13].um_I.iw[17] ;
 wire \top_I.branch[9].block[13].um_I.iw[1] ;
 wire \top_I.branch[9].block[13].um_I.iw[2] ;
 wire \top_I.branch[9].block[13].um_I.iw[3] ;
 wire \top_I.branch[9].block[13].um_I.iw[4] ;
 wire \top_I.branch[9].block[13].um_I.iw[5] ;
 wire \top_I.branch[9].block[13].um_I.iw[6] ;
 wire \top_I.branch[9].block[13].um_I.iw[7] ;
 wire \top_I.branch[9].block[13].um_I.iw[8] ;
 wire \top_I.branch[9].block[13].um_I.iw[9] ;
 wire \top_I.branch[9].block[13].um_I.k_zero ;
 wire \top_I.branch[9].block[13].um_I.pg_vdd ;
 wire \top_I.branch[9].block[14].um_I.ana[0] ;
 wire \top_I.branch[9].block[14].um_I.ana[1] ;
 wire \top_I.branch[9].block[14].um_I.ana[2] ;
 wire \top_I.branch[9].block[14].um_I.ana[3] ;
 wire \top_I.branch[9].block[14].um_I.ana[4] ;
 wire \top_I.branch[9].block[14].um_I.ana[5] ;
 wire \top_I.branch[9].block[14].um_I.ana[6] ;
 wire \top_I.branch[9].block[14].um_I.ana[7] ;
 wire \top_I.branch[9].block[14].um_I.clk ;
 wire \top_I.branch[9].block[14].um_I.ena ;
 wire \top_I.branch[9].block[14].um_I.iw[10] ;
 wire \top_I.branch[9].block[14].um_I.iw[11] ;
 wire \top_I.branch[9].block[14].um_I.iw[12] ;
 wire \top_I.branch[9].block[14].um_I.iw[13] ;
 wire \top_I.branch[9].block[14].um_I.iw[14] ;
 wire \top_I.branch[9].block[14].um_I.iw[15] ;
 wire \top_I.branch[9].block[14].um_I.iw[16] ;
 wire \top_I.branch[9].block[14].um_I.iw[17] ;
 wire \top_I.branch[9].block[14].um_I.iw[1] ;
 wire \top_I.branch[9].block[14].um_I.iw[2] ;
 wire \top_I.branch[9].block[14].um_I.iw[3] ;
 wire \top_I.branch[9].block[14].um_I.iw[4] ;
 wire \top_I.branch[9].block[14].um_I.iw[5] ;
 wire \top_I.branch[9].block[14].um_I.iw[6] ;
 wire \top_I.branch[9].block[14].um_I.iw[7] ;
 wire \top_I.branch[9].block[14].um_I.iw[8] ;
 wire \top_I.branch[9].block[14].um_I.iw[9] ;
 wire \top_I.branch[9].block[14].um_I.k_zero ;
 wire \top_I.branch[9].block[14].um_I.pg_vdd ;
 wire \top_I.branch[9].block[15].um_I.ana[0] ;
 wire \top_I.branch[9].block[15].um_I.ana[1] ;
 wire \top_I.branch[9].block[15].um_I.ana[2] ;
 wire \top_I.branch[9].block[15].um_I.ana[3] ;
 wire \top_I.branch[9].block[15].um_I.ana[4] ;
 wire \top_I.branch[9].block[15].um_I.ana[5] ;
 wire \top_I.branch[9].block[15].um_I.ana[6] ;
 wire \top_I.branch[9].block[15].um_I.ana[7] ;
 wire \top_I.branch[9].block[15].um_I.clk ;
 wire \top_I.branch[9].block[15].um_I.ena ;
 wire \top_I.branch[9].block[15].um_I.iw[10] ;
 wire \top_I.branch[9].block[15].um_I.iw[11] ;
 wire \top_I.branch[9].block[15].um_I.iw[12] ;
 wire \top_I.branch[9].block[15].um_I.iw[13] ;
 wire \top_I.branch[9].block[15].um_I.iw[14] ;
 wire \top_I.branch[9].block[15].um_I.iw[15] ;
 wire \top_I.branch[9].block[15].um_I.iw[16] ;
 wire \top_I.branch[9].block[15].um_I.iw[17] ;
 wire \top_I.branch[9].block[15].um_I.iw[1] ;
 wire \top_I.branch[9].block[15].um_I.iw[2] ;
 wire \top_I.branch[9].block[15].um_I.iw[3] ;
 wire \top_I.branch[9].block[15].um_I.iw[4] ;
 wire \top_I.branch[9].block[15].um_I.iw[5] ;
 wire \top_I.branch[9].block[15].um_I.iw[6] ;
 wire \top_I.branch[9].block[15].um_I.iw[7] ;
 wire \top_I.branch[9].block[15].um_I.iw[8] ;
 wire \top_I.branch[9].block[15].um_I.iw[9] ;
 wire \top_I.branch[9].block[15].um_I.k_zero ;
 wire \top_I.branch[9].block[15].um_I.pg_vdd ;
 wire \top_I.branch[9].block[1].um_I.ana[0] ;
 wire \top_I.branch[9].block[1].um_I.ana[1] ;
 wire \top_I.branch[9].block[1].um_I.ana[2] ;
 wire \top_I.branch[9].block[1].um_I.ana[3] ;
 wire \top_I.branch[9].block[1].um_I.ana[4] ;
 wire \top_I.branch[9].block[1].um_I.ana[5] ;
 wire \top_I.branch[9].block[1].um_I.ana[6] ;
 wire \top_I.branch[9].block[1].um_I.ana[7] ;
 wire \top_I.branch[9].block[1].um_I.clk ;
 wire \top_I.branch[9].block[1].um_I.ena ;
 wire \top_I.branch[9].block[1].um_I.iw[10] ;
 wire \top_I.branch[9].block[1].um_I.iw[11] ;
 wire \top_I.branch[9].block[1].um_I.iw[12] ;
 wire \top_I.branch[9].block[1].um_I.iw[13] ;
 wire \top_I.branch[9].block[1].um_I.iw[14] ;
 wire \top_I.branch[9].block[1].um_I.iw[15] ;
 wire \top_I.branch[9].block[1].um_I.iw[16] ;
 wire \top_I.branch[9].block[1].um_I.iw[17] ;
 wire \top_I.branch[9].block[1].um_I.iw[1] ;
 wire \top_I.branch[9].block[1].um_I.iw[2] ;
 wire \top_I.branch[9].block[1].um_I.iw[3] ;
 wire \top_I.branch[9].block[1].um_I.iw[4] ;
 wire \top_I.branch[9].block[1].um_I.iw[5] ;
 wire \top_I.branch[9].block[1].um_I.iw[6] ;
 wire \top_I.branch[9].block[1].um_I.iw[7] ;
 wire \top_I.branch[9].block[1].um_I.iw[8] ;
 wire \top_I.branch[9].block[1].um_I.iw[9] ;
 wire \top_I.branch[9].block[1].um_I.k_zero ;
 wire \top_I.branch[9].block[1].um_I.pg_vdd ;
 wire \top_I.branch[9].block[2].um_I.ana[0] ;
 wire \top_I.branch[9].block[2].um_I.ana[1] ;
 wire \top_I.branch[9].block[2].um_I.ana[2] ;
 wire \top_I.branch[9].block[2].um_I.ana[3] ;
 wire \top_I.branch[9].block[2].um_I.ana[4] ;
 wire \top_I.branch[9].block[2].um_I.ana[5] ;
 wire \top_I.branch[9].block[2].um_I.ana[6] ;
 wire \top_I.branch[9].block[2].um_I.ana[7] ;
 wire \top_I.branch[9].block[2].um_I.clk ;
 wire \top_I.branch[9].block[2].um_I.ena ;
 wire \top_I.branch[9].block[2].um_I.iw[10] ;
 wire \top_I.branch[9].block[2].um_I.iw[11] ;
 wire \top_I.branch[9].block[2].um_I.iw[12] ;
 wire \top_I.branch[9].block[2].um_I.iw[13] ;
 wire \top_I.branch[9].block[2].um_I.iw[14] ;
 wire \top_I.branch[9].block[2].um_I.iw[15] ;
 wire \top_I.branch[9].block[2].um_I.iw[16] ;
 wire \top_I.branch[9].block[2].um_I.iw[17] ;
 wire \top_I.branch[9].block[2].um_I.iw[1] ;
 wire \top_I.branch[9].block[2].um_I.iw[2] ;
 wire \top_I.branch[9].block[2].um_I.iw[3] ;
 wire \top_I.branch[9].block[2].um_I.iw[4] ;
 wire \top_I.branch[9].block[2].um_I.iw[5] ;
 wire \top_I.branch[9].block[2].um_I.iw[6] ;
 wire \top_I.branch[9].block[2].um_I.iw[7] ;
 wire \top_I.branch[9].block[2].um_I.iw[8] ;
 wire \top_I.branch[9].block[2].um_I.iw[9] ;
 wire \top_I.branch[9].block[2].um_I.k_zero ;
 wire \top_I.branch[9].block[2].um_I.pg_vdd ;
 wire \top_I.branch[9].block[3].um_I.ana[0] ;
 wire \top_I.branch[9].block[3].um_I.ana[1] ;
 wire \top_I.branch[9].block[3].um_I.ana[2] ;
 wire \top_I.branch[9].block[3].um_I.ana[3] ;
 wire \top_I.branch[9].block[3].um_I.ana[4] ;
 wire \top_I.branch[9].block[3].um_I.ana[5] ;
 wire \top_I.branch[9].block[3].um_I.ana[6] ;
 wire \top_I.branch[9].block[3].um_I.ana[7] ;
 wire \top_I.branch[9].block[3].um_I.clk ;
 wire \top_I.branch[9].block[3].um_I.ena ;
 wire \top_I.branch[9].block[3].um_I.iw[10] ;
 wire \top_I.branch[9].block[3].um_I.iw[11] ;
 wire \top_I.branch[9].block[3].um_I.iw[12] ;
 wire \top_I.branch[9].block[3].um_I.iw[13] ;
 wire \top_I.branch[9].block[3].um_I.iw[14] ;
 wire \top_I.branch[9].block[3].um_I.iw[15] ;
 wire \top_I.branch[9].block[3].um_I.iw[16] ;
 wire \top_I.branch[9].block[3].um_I.iw[17] ;
 wire \top_I.branch[9].block[3].um_I.iw[1] ;
 wire \top_I.branch[9].block[3].um_I.iw[2] ;
 wire \top_I.branch[9].block[3].um_I.iw[3] ;
 wire \top_I.branch[9].block[3].um_I.iw[4] ;
 wire \top_I.branch[9].block[3].um_I.iw[5] ;
 wire \top_I.branch[9].block[3].um_I.iw[6] ;
 wire \top_I.branch[9].block[3].um_I.iw[7] ;
 wire \top_I.branch[9].block[3].um_I.iw[8] ;
 wire \top_I.branch[9].block[3].um_I.iw[9] ;
 wire \top_I.branch[9].block[3].um_I.k_zero ;
 wire \top_I.branch[9].block[3].um_I.pg_vdd ;
 wire \top_I.branch[9].block[4].um_I.ana[0] ;
 wire \top_I.branch[9].block[4].um_I.ana[1] ;
 wire \top_I.branch[9].block[4].um_I.ana[2] ;
 wire \top_I.branch[9].block[4].um_I.ana[3] ;
 wire \top_I.branch[9].block[4].um_I.ana[4] ;
 wire \top_I.branch[9].block[4].um_I.ana[5] ;
 wire \top_I.branch[9].block[4].um_I.ana[6] ;
 wire \top_I.branch[9].block[4].um_I.ana[7] ;
 wire \top_I.branch[9].block[4].um_I.clk ;
 wire \top_I.branch[9].block[4].um_I.ena ;
 wire \top_I.branch[9].block[4].um_I.iw[10] ;
 wire \top_I.branch[9].block[4].um_I.iw[11] ;
 wire \top_I.branch[9].block[4].um_I.iw[12] ;
 wire \top_I.branch[9].block[4].um_I.iw[13] ;
 wire \top_I.branch[9].block[4].um_I.iw[14] ;
 wire \top_I.branch[9].block[4].um_I.iw[15] ;
 wire \top_I.branch[9].block[4].um_I.iw[16] ;
 wire \top_I.branch[9].block[4].um_I.iw[17] ;
 wire \top_I.branch[9].block[4].um_I.iw[1] ;
 wire \top_I.branch[9].block[4].um_I.iw[2] ;
 wire \top_I.branch[9].block[4].um_I.iw[3] ;
 wire \top_I.branch[9].block[4].um_I.iw[4] ;
 wire \top_I.branch[9].block[4].um_I.iw[5] ;
 wire \top_I.branch[9].block[4].um_I.iw[6] ;
 wire \top_I.branch[9].block[4].um_I.iw[7] ;
 wire \top_I.branch[9].block[4].um_I.iw[8] ;
 wire \top_I.branch[9].block[4].um_I.iw[9] ;
 wire \top_I.branch[9].block[4].um_I.k_zero ;
 wire \top_I.branch[9].block[4].um_I.pg_vdd ;
 wire \top_I.branch[9].block[5].um_I.ana[0] ;
 wire \top_I.branch[9].block[5].um_I.ana[1] ;
 wire \top_I.branch[9].block[5].um_I.ana[2] ;
 wire \top_I.branch[9].block[5].um_I.ana[3] ;
 wire \top_I.branch[9].block[5].um_I.ana[4] ;
 wire \top_I.branch[9].block[5].um_I.ana[5] ;
 wire \top_I.branch[9].block[5].um_I.ana[6] ;
 wire \top_I.branch[9].block[5].um_I.ana[7] ;
 wire \top_I.branch[9].block[5].um_I.clk ;
 wire \top_I.branch[9].block[5].um_I.ena ;
 wire \top_I.branch[9].block[5].um_I.iw[10] ;
 wire \top_I.branch[9].block[5].um_I.iw[11] ;
 wire \top_I.branch[9].block[5].um_I.iw[12] ;
 wire \top_I.branch[9].block[5].um_I.iw[13] ;
 wire \top_I.branch[9].block[5].um_I.iw[14] ;
 wire \top_I.branch[9].block[5].um_I.iw[15] ;
 wire \top_I.branch[9].block[5].um_I.iw[16] ;
 wire \top_I.branch[9].block[5].um_I.iw[17] ;
 wire \top_I.branch[9].block[5].um_I.iw[1] ;
 wire \top_I.branch[9].block[5].um_I.iw[2] ;
 wire \top_I.branch[9].block[5].um_I.iw[3] ;
 wire \top_I.branch[9].block[5].um_I.iw[4] ;
 wire \top_I.branch[9].block[5].um_I.iw[5] ;
 wire \top_I.branch[9].block[5].um_I.iw[6] ;
 wire \top_I.branch[9].block[5].um_I.iw[7] ;
 wire \top_I.branch[9].block[5].um_I.iw[8] ;
 wire \top_I.branch[9].block[5].um_I.iw[9] ;
 wire \top_I.branch[9].block[5].um_I.k_zero ;
 wire \top_I.branch[9].block[5].um_I.pg_vdd ;
 wire \top_I.branch[9].block[6].um_I.ana[0] ;
 wire \top_I.branch[9].block[6].um_I.ana[1] ;
 wire \top_I.branch[9].block[6].um_I.ana[2] ;
 wire \top_I.branch[9].block[6].um_I.ana[3] ;
 wire \top_I.branch[9].block[6].um_I.ana[4] ;
 wire \top_I.branch[9].block[6].um_I.ana[5] ;
 wire \top_I.branch[9].block[6].um_I.ana[6] ;
 wire \top_I.branch[9].block[6].um_I.ana[7] ;
 wire \top_I.branch[9].block[6].um_I.clk ;
 wire \top_I.branch[9].block[6].um_I.ena ;
 wire \top_I.branch[9].block[6].um_I.iw[10] ;
 wire \top_I.branch[9].block[6].um_I.iw[11] ;
 wire \top_I.branch[9].block[6].um_I.iw[12] ;
 wire \top_I.branch[9].block[6].um_I.iw[13] ;
 wire \top_I.branch[9].block[6].um_I.iw[14] ;
 wire \top_I.branch[9].block[6].um_I.iw[15] ;
 wire \top_I.branch[9].block[6].um_I.iw[16] ;
 wire \top_I.branch[9].block[6].um_I.iw[17] ;
 wire \top_I.branch[9].block[6].um_I.iw[1] ;
 wire \top_I.branch[9].block[6].um_I.iw[2] ;
 wire \top_I.branch[9].block[6].um_I.iw[3] ;
 wire \top_I.branch[9].block[6].um_I.iw[4] ;
 wire \top_I.branch[9].block[6].um_I.iw[5] ;
 wire \top_I.branch[9].block[6].um_I.iw[6] ;
 wire \top_I.branch[9].block[6].um_I.iw[7] ;
 wire \top_I.branch[9].block[6].um_I.iw[8] ;
 wire \top_I.branch[9].block[6].um_I.iw[9] ;
 wire \top_I.branch[9].block[6].um_I.k_zero ;
 wire \top_I.branch[9].block[6].um_I.pg_vdd ;
 wire \top_I.branch[9].block[7].um_I.ana[0] ;
 wire \top_I.branch[9].block[7].um_I.ana[1] ;
 wire \top_I.branch[9].block[7].um_I.ana[2] ;
 wire \top_I.branch[9].block[7].um_I.ana[3] ;
 wire \top_I.branch[9].block[7].um_I.ana[4] ;
 wire \top_I.branch[9].block[7].um_I.ana[5] ;
 wire \top_I.branch[9].block[7].um_I.ana[6] ;
 wire \top_I.branch[9].block[7].um_I.ana[7] ;
 wire \top_I.branch[9].block[7].um_I.clk ;
 wire \top_I.branch[9].block[7].um_I.ena ;
 wire \top_I.branch[9].block[7].um_I.iw[10] ;
 wire \top_I.branch[9].block[7].um_I.iw[11] ;
 wire \top_I.branch[9].block[7].um_I.iw[12] ;
 wire \top_I.branch[9].block[7].um_I.iw[13] ;
 wire \top_I.branch[9].block[7].um_I.iw[14] ;
 wire \top_I.branch[9].block[7].um_I.iw[15] ;
 wire \top_I.branch[9].block[7].um_I.iw[16] ;
 wire \top_I.branch[9].block[7].um_I.iw[17] ;
 wire \top_I.branch[9].block[7].um_I.iw[1] ;
 wire \top_I.branch[9].block[7].um_I.iw[2] ;
 wire \top_I.branch[9].block[7].um_I.iw[3] ;
 wire \top_I.branch[9].block[7].um_I.iw[4] ;
 wire \top_I.branch[9].block[7].um_I.iw[5] ;
 wire \top_I.branch[9].block[7].um_I.iw[6] ;
 wire \top_I.branch[9].block[7].um_I.iw[7] ;
 wire \top_I.branch[9].block[7].um_I.iw[8] ;
 wire \top_I.branch[9].block[7].um_I.iw[9] ;
 wire \top_I.branch[9].block[7].um_I.k_zero ;
 wire \top_I.branch[9].block[7].um_I.pg_vdd ;
 wire \top_I.branch[9].block[8].um_I.ana[0] ;
 wire \top_I.branch[9].block[8].um_I.ana[1] ;
 wire \top_I.branch[9].block[8].um_I.ana[2] ;
 wire \top_I.branch[9].block[8].um_I.ana[3] ;
 wire \top_I.branch[9].block[8].um_I.ana[4] ;
 wire \top_I.branch[9].block[8].um_I.ana[5] ;
 wire \top_I.branch[9].block[8].um_I.ana[6] ;
 wire \top_I.branch[9].block[8].um_I.ana[7] ;
 wire \top_I.branch[9].block[8].um_I.clk ;
 wire \top_I.branch[9].block[8].um_I.ena ;
 wire \top_I.branch[9].block[8].um_I.iw[10] ;
 wire \top_I.branch[9].block[8].um_I.iw[11] ;
 wire \top_I.branch[9].block[8].um_I.iw[12] ;
 wire \top_I.branch[9].block[8].um_I.iw[13] ;
 wire \top_I.branch[9].block[8].um_I.iw[14] ;
 wire \top_I.branch[9].block[8].um_I.iw[15] ;
 wire \top_I.branch[9].block[8].um_I.iw[16] ;
 wire \top_I.branch[9].block[8].um_I.iw[17] ;
 wire \top_I.branch[9].block[8].um_I.iw[1] ;
 wire \top_I.branch[9].block[8].um_I.iw[2] ;
 wire \top_I.branch[9].block[8].um_I.iw[3] ;
 wire \top_I.branch[9].block[8].um_I.iw[4] ;
 wire \top_I.branch[9].block[8].um_I.iw[5] ;
 wire \top_I.branch[9].block[8].um_I.iw[6] ;
 wire \top_I.branch[9].block[8].um_I.iw[7] ;
 wire \top_I.branch[9].block[8].um_I.iw[8] ;
 wire \top_I.branch[9].block[8].um_I.iw[9] ;
 wire \top_I.branch[9].block[8].um_I.k_zero ;
 wire \top_I.branch[9].block[8].um_I.pg_vdd ;
 wire \top_I.branch[9].block[9].um_I.ana[0] ;
 wire \top_I.branch[9].block[9].um_I.ana[1] ;
 wire \top_I.branch[9].block[9].um_I.ana[2] ;
 wire \top_I.branch[9].block[9].um_I.ana[3] ;
 wire \top_I.branch[9].block[9].um_I.ana[4] ;
 wire \top_I.branch[9].block[9].um_I.ana[5] ;
 wire \top_I.branch[9].block[9].um_I.ana[6] ;
 wire \top_I.branch[9].block[9].um_I.ana[7] ;
 wire \top_I.branch[9].block[9].um_I.clk ;
 wire \top_I.branch[9].block[9].um_I.ena ;
 wire \top_I.branch[9].block[9].um_I.iw[10] ;
 wire \top_I.branch[9].block[9].um_I.iw[11] ;
 wire \top_I.branch[9].block[9].um_I.iw[12] ;
 wire \top_I.branch[9].block[9].um_I.iw[13] ;
 wire \top_I.branch[9].block[9].um_I.iw[14] ;
 wire \top_I.branch[9].block[9].um_I.iw[15] ;
 wire \top_I.branch[9].block[9].um_I.iw[16] ;
 wire \top_I.branch[9].block[9].um_I.iw[17] ;
 wire \top_I.branch[9].block[9].um_I.iw[1] ;
 wire \top_I.branch[9].block[9].um_I.iw[2] ;
 wire \top_I.branch[9].block[9].um_I.iw[3] ;
 wire \top_I.branch[9].block[9].um_I.iw[4] ;
 wire \top_I.branch[9].block[9].um_I.iw[5] ;
 wire \top_I.branch[9].block[9].um_I.iw[6] ;
 wire \top_I.branch[9].block[9].um_I.iw[7] ;
 wire \top_I.branch[9].block[9].um_I.iw[8] ;
 wire \top_I.branch[9].block[9].um_I.iw[9] ;
 wire \top_I.branch[9].block[9].um_I.k_zero ;
 wire \top_I.branch[9].block[9].um_I.pg_vdd ;
 wire \top_I.branch[9].l_addr[0] ;
 wire \top_I.branch[9].l_addr[2] ;

 tt_pg_vdd_1 \top_I.branch[0].block[0].um_I.block_0_0.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[0].block[0].um_I.block_0_0.vpwr ),
    .ctrl(\top_I.branch[0].block[0].um_I.pg_vdd ));
 tt_um_chip_rom \top_I.branch[0].block[0].um_I.block_0_0.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[0].block[0].um_I.block_0_0.vpwr ),
    .clk(\top_I.branch[0].block[0].um_I.clk ),
    .ena(\top_I.branch[0].block[0].um_I.ena ),
    .rst_n(\top_I.branch[0].block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].block[0].um_I.iw[9] ,
    \top_I.branch[0].block[0].um_I.iw[8] ,
    \top_I.branch[0].block[0].um_I.iw[7] ,
    \top_I.branch[0].block[0].um_I.iw[6] ,
    \top_I.branch[0].block[0].um_I.iw[5] ,
    \top_I.branch[0].block[0].um_I.iw[4] ,
    \top_I.branch[0].block[0].um_I.iw[3] ,
    \top_I.branch[0].block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].block[0].um_I.iw[17] ,
    \top_I.branch[0].block[0].um_I.iw[16] ,
    \top_I.branch[0].block[0].um_I.iw[15] ,
    \top_I.branch[0].block[0].um_I.iw[14] ,
    \top_I.branch[0].block[0].um_I.iw[13] ,
    \top_I.branch[0].block[0].um_I.iw[12] ,
    \top_I.branch[0].block[0].um_I.iw[11] ,
    \top_I.branch[0].block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].block[0].um_I.ow[23] ,
    \top_I.branch[0].block[0].um_I.ow[22] ,
    \top_I.branch[0].block[0].um_I.ow[21] ,
    \top_I.branch[0].block[0].um_I.ow[20] ,
    \top_I.branch[0].block[0].um_I.ow[19] ,
    \top_I.branch[0].block[0].um_I.ow[18] ,
    \top_I.branch[0].block[0].um_I.ow[17] ,
    \top_I.branch[0].block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].block[0].um_I.ow[15] ,
    \top_I.branch[0].block[0].um_I.ow[14] ,
    \top_I.branch[0].block[0].um_I.ow[13] ,
    \top_I.branch[0].block[0].um_I.ow[12] ,
    \top_I.branch[0].block[0].um_I.ow[11] ,
    \top_I.branch[0].block[0].um_I.ow[10] ,
    \top_I.branch[0].block[0].um_I.ow[9] ,
    \top_I.branch[0].block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].block[0].um_I.ow[7] ,
    \top_I.branch[0].block[0].um_I.ow[6] ,
    \top_I.branch[0].block[0].um_I.ow[5] ,
    \top_I.branch[0].block[0].um_I.ow[4] ,
    \top_I.branch[0].block[0].um_I.ow[3] ,
    \top_I.branch[0].block[0].um_I.ow[2] ,
    \top_I.branch[0].block[0].um_I.ow[1] ,
    \top_I.branch[0].block[0].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[0].block[1].um_I.block_0_1.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[0].block[1].um_I.block_0_1.vpwr ),
    .ctrl(\top_I.branch[0].block[1].um_I.pg_vdd ));
 tt_um_factory_test \top_I.branch[0].block[1].um_I.block_0_1.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[0].block[1].um_I.block_0_1.vpwr ),
    .clk(\top_I.branch[0].block[1].um_I.clk ),
    .ena(\top_I.branch[0].block[1].um_I.ena ),
    .rst_n(\top_I.branch[0].block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[0].block[1].um_I.iw[9] ,
    \top_I.branch[0].block[1].um_I.iw[8] ,
    \top_I.branch[0].block[1].um_I.iw[7] ,
    \top_I.branch[0].block[1].um_I.iw[6] ,
    \top_I.branch[0].block[1].um_I.iw[5] ,
    \top_I.branch[0].block[1].um_I.iw[4] ,
    \top_I.branch[0].block[1].um_I.iw[3] ,
    \top_I.branch[0].block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[0].block[1].um_I.iw[17] ,
    \top_I.branch[0].block[1].um_I.iw[16] ,
    \top_I.branch[0].block[1].um_I.iw[15] ,
    \top_I.branch[0].block[1].um_I.iw[14] ,
    \top_I.branch[0].block[1].um_I.iw[13] ,
    \top_I.branch[0].block[1].um_I.iw[12] ,
    \top_I.branch[0].block[1].um_I.iw[11] ,
    \top_I.branch[0].block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[0].block[1].um_I.ow[23] ,
    \top_I.branch[0].block[1].um_I.ow[22] ,
    \top_I.branch[0].block[1].um_I.ow[21] ,
    \top_I.branch[0].block[1].um_I.ow[20] ,
    \top_I.branch[0].block[1].um_I.ow[19] ,
    \top_I.branch[0].block[1].um_I.ow[18] ,
    \top_I.branch[0].block[1].um_I.ow[17] ,
    \top_I.branch[0].block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[0].block[1].um_I.ow[15] ,
    \top_I.branch[0].block[1].um_I.ow[14] ,
    \top_I.branch[0].block[1].um_I.ow[13] ,
    \top_I.branch[0].block[1].um_I.ow[12] ,
    \top_I.branch[0].block[1].um_I.ow[11] ,
    \top_I.branch[0].block[1].um_I.ow[10] ,
    \top_I.branch[0].block[1].um_I.ow[9] ,
    \top_I.branch[0].block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[0].block[1].um_I.ow[7] ,
    \top_I.branch[0].block[1].um_I.ow[6] ,
    \top_I.branch[0].block[1].um_I.ow[5] ,
    \top_I.branch[0].block[1].um_I.ow[4] ,
    \top_I.branch[0].block[1].um_I.ow[3] ,
    \top_I.branch[0].block[1].um_I.ow[2] ,
    \top_I.branch[0].block[1].um_I.ow[1] ,
    \top_I.branch[0].block[1].um_I.ow[0] }));
 tt_mux \top_I.branch[0].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[0].l_k_one ),
    .k_zero(\top_I.branch[0].l_addr[0] ),
    .addr({\top_I.branch[0].l_addr[0] ,
    \top_I.branch[0].l_addr[0] ,
    \top_I.branch[0].l_addr[0] ,
    \top_I.branch[0].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[0].block[15].um_I.ena ,
    \top_I.branch[0].block[14].um_I.ena ,
    \top_I.branch[0].block[13].um_I.ena ,
    \top_I.branch[0].block[12].um_I.ena ,
    \top_I.branch[0].block[11].um_I.ena ,
    \top_I.branch[0].block[10].um_I.ena ,
    \top_I.branch[0].block[9].um_I.ena ,
    \top_I.branch[0].block[8].um_I.ena ,
    \top_I.branch[0].block[7].um_I.ena ,
    \top_I.branch[0].block[6].um_I.ena ,
    \top_I.branch[0].block[5].um_I.ena ,
    \top_I.branch[0].block[4].um_I.ena ,
    \top_I.branch[0].block[3].um_I.ena ,
    \top_I.branch[0].block[2].um_I.ena ,
    \top_I.branch[0].block[1].um_I.ena ,
    \top_I.branch[0].block[0].um_I.ena }),
    .um_iw({\top_I.branch[0].block[15].um_I.iw[17] ,
    \top_I.branch[0].block[15].um_I.iw[16] ,
    \top_I.branch[0].block[15].um_I.iw[15] ,
    \top_I.branch[0].block[15].um_I.iw[14] ,
    \top_I.branch[0].block[15].um_I.iw[13] ,
    \top_I.branch[0].block[15].um_I.iw[12] ,
    \top_I.branch[0].block[15].um_I.iw[11] ,
    \top_I.branch[0].block[15].um_I.iw[10] ,
    \top_I.branch[0].block[15].um_I.iw[9] ,
    \top_I.branch[0].block[15].um_I.iw[8] ,
    \top_I.branch[0].block[15].um_I.iw[7] ,
    \top_I.branch[0].block[15].um_I.iw[6] ,
    \top_I.branch[0].block[15].um_I.iw[5] ,
    \top_I.branch[0].block[15].um_I.iw[4] ,
    \top_I.branch[0].block[15].um_I.iw[3] ,
    \top_I.branch[0].block[15].um_I.iw[2] ,
    \top_I.branch[0].block[15].um_I.iw[1] ,
    \top_I.branch[0].block[15].um_I.clk ,
    \top_I.branch[0].block[14].um_I.iw[17] ,
    \top_I.branch[0].block[14].um_I.iw[16] ,
    \top_I.branch[0].block[14].um_I.iw[15] ,
    \top_I.branch[0].block[14].um_I.iw[14] ,
    \top_I.branch[0].block[14].um_I.iw[13] ,
    \top_I.branch[0].block[14].um_I.iw[12] ,
    \top_I.branch[0].block[14].um_I.iw[11] ,
    \top_I.branch[0].block[14].um_I.iw[10] ,
    \top_I.branch[0].block[14].um_I.iw[9] ,
    \top_I.branch[0].block[14].um_I.iw[8] ,
    \top_I.branch[0].block[14].um_I.iw[7] ,
    \top_I.branch[0].block[14].um_I.iw[6] ,
    \top_I.branch[0].block[14].um_I.iw[5] ,
    \top_I.branch[0].block[14].um_I.iw[4] ,
    \top_I.branch[0].block[14].um_I.iw[3] ,
    \top_I.branch[0].block[14].um_I.iw[2] ,
    \top_I.branch[0].block[14].um_I.iw[1] ,
    \top_I.branch[0].block[14].um_I.clk ,
    \top_I.branch[0].block[13].um_I.iw[17] ,
    \top_I.branch[0].block[13].um_I.iw[16] ,
    \top_I.branch[0].block[13].um_I.iw[15] ,
    \top_I.branch[0].block[13].um_I.iw[14] ,
    \top_I.branch[0].block[13].um_I.iw[13] ,
    \top_I.branch[0].block[13].um_I.iw[12] ,
    \top_I.branch[0].block[13].um_I.iw[11] ,
    \top_I.branch[0].block[13].um_I.iw[10] ,
    \top_I.branch[0].block[13].um_I.iw[9] ,
    \top_I.branch[0].block[13].um_I.iw[8] ,
    \top_I.branch[0].block[13].um_I.iw[7] ,
    \top_I.branch[0].block[13].um_I.iw[6] ,
    \top_I.branch[0].block[13].um_I.iw[5] ,
    \top_I.branch[0].block[13].um_I.iw[4] ,
    \top_I.branch[0].block[13].um_I.iw[3] ,
    \top_I.branch[0].block[13].um_I.iw[2] ,
    \top_I.branch[0].block[13].um_I.iw[1] ,
    \top_I.branch[0].block[13].um_I.clk ,
    \top_I.branch[0].block[12].um_I.iw[17] ,
    \top_I.branch[0].block[12].um_I.iw[16] ,
    \top_I.branch[0].block[12].um_I.iw[15] ,
    \top_I.branch[0].block[12].um_I.iw[14] ,
    \top_I.branch[0].block[12].um_I.iw[13] ,
    \top_I.branch[0].block[12].um_I.iw[12] ,
    \top_I.branch[0].block[12].um_I.iw[11] ,
    \top_I.branch[0].block[12].um_I.iw[10] ,
    \top_I.branch[0].block[12].um_I.iw[9] ,
    \top_I.branch[0].block[12].um_I.iw[8] ,
    \top_I.branch[0].block[12].um_I.iw[7] ,
    \top_I.branch[0].block[12].um_I.iw[6] ,
    \top_I.branch[0].block[12].um_I.iw[5] ,
    \top_I.branch[0].block[12].um_I.iw[4] ,
    \top_I.branch[0].block[12].um_I.iw[3] ,
    \top_I.branch[0].block[12].um_I.iw[2] ,
    \top_I.branch[0].block[12].um_I.iw[1] ,
    \top_I.branch[0].block[12].um_I.clk ,
    \top_I.branch[0].block[11].um_I.iw[17] ,
    \top_I.branch[0].block[11].um_I.iw[16] ,
    \top_I.branch[0].block[11].um_I.iw[15] ,
    \top_I.branch[0].block[11].um_I.iw[14] ,
    \top_I.branch[0].block[11].um_I.iw[13] ,
    \top_I.branch[0].block[11].um_I.iw[12] ,
    \top_I.branch[0].block[11].um_I.iw[11] ,
    \top_I.branch[0].block[11].um_I.iw[10] ,
    \top_I.branch[0].block[11].um_I.iw[9] ,
    \top_I.branch[0].block[11].um_I.iw[8] ,
    \top_I.branch[0].block[11].um_I.iw[7] ,
    \top_I.branch[0].block[11].um_I.iw[6] ,
    \top_I.branch[0].block[11].um_I.iw[5] ,
    \top_I.branch[0].block[11].um_I.iw[4] ,
    \top_I.branch[0].block[11].um_I.iw[3] ,
    \top_I.branch[0].block[11].um_I.iw[2] ,
    \top_I.branch[0].block[11].um_I.iw[1] ,
    \top_I.branch[0].block[11].um_I.clk ,
    \top_I.branch[0].block[10].um_I.iw[17] ,
    \top_I.branch[0].block[10].um_I.iw[16] ,
    \top_I.branch[0].block[10].um_I.iw[15] ,
    \top_I.branch[0].block[10].um_I.iw[14] ,
    \top_I.branch[0].block[10].um_I.iw[13] ,
    \top_I.branch[0].block[10].um_I.iw[12] ,
    \top_I.branch[0].block[10].um_I.iw[11] ,
    \top_I.branch[0].block[10].um_I.iw[10] ,
    \top_I.branch[0].block[10].um_I.iw[9] ,
    \top_I.branch[0].block[10].um_I.iw[8] ,
    \top_I.branch[0].block[10].um_I.iw[7] ,
    \top_I.branch[0].block[10].um_I.iw[6] ,
    \top_I.branch[0].block[10].um_I.iw[5] ,
    \top_I.branch[0].block[10].um_I.iw[4] ,
    \top_I.branch[0].block[10].um_I.iw[3] ,
    \top_I.branch[0].block[10].um_I.iw[2] ,
    \top_I.branch[0].block[10].um_I.iw[1] ,
    \top_I.branch[0].block[10].um_I.clk ,
    \top_I.branch[0].block[9].um_I.iw[17] ,
    \top_I.branch[0].block[9].um_I.iw[16] ,
    \top_I.branch[0].block[9].um_I.iw[15] ,
    \top_I.branch[0].block[9].um_I.iw[14] ,
    \top_I.branch[0].block[9].um_I.iw[13] ,
    \top_I.branch[0].block[9].um_I.iw[12] ,
    \top_I.branch[0].block[9].um_I.iw[11] ,
    \top_I.branch[0].block[9].um_I.iw[10] ,
    \top_I.branch[0].block[9].um_I.iw[9] ,
    \top_I.branch[0].block[9].um_I.iw[8] ,
    \top_I.branch[0].block[9].um_I.iw[7] ,
    \top_I.branch[0].block[9].um_I.iw[6] ,
    \top_I.branch[0].block[9].um_I.iw[5] ,
    \top_I.branch[0].block[9].um_I.iw[4] ,
    \top_I.branch[0].block[9].um_I.iw[3] ,
    \top_I.branch[0].block[9].um_I.iw[2] ,
    \top_I.branch[0].block[9].um_I.iw[1] ,
    \top_I.branch[0].block[9].um_I.clk ,
    \top_I.branch[0].block[8].um_I.iw[17] ,
    \top_I.branch[0].block[8].um_I.iw[16] ,
    \top_I.branch[0].block[8].um_I.iw[15] ,
    \top_I.branch[0].block[8].um_I.iw[14] ,
    \top_I.branch[0].block[8].um_I.iw[13] ,
    \top_I.branch[0].block[8].um_I.iw[12] ,
    \top_I.branch[0].block[8].um_I.iw[11] ,
    \top_I.branch[0].block[8].um_I.iw[10] ,
    \top_I.branch[0].block[8].um_I.iw[9] ,
    \top_I.branch[0].block[8].um_I.iw[8] ,
    \top_I.branch[0].block[8].um_I.iw[7] ,
    \top_I.branch[0].block[8].um_I.iw[6] ,
    \top_I.branch[0].block[8].um_I.iw[5] ,
    \top_I.branch[0].block[8].um_I.iw[4] ,
    \top_I.branch[0].block[8].um_I.iw[3] ,
    \top_I.branch[0].block[8].um_I.iw[2] ,
    \top_I.branch[0].block[8].um_I.iw[1] ,
    \top_I.branch[0].block[8].um_I.clk ,
    \top_I.branch[0].block[7].um_I.iw[17] ,
    \top_I.branch[0].block[7].um_I.iw[16] ,
    \top_I.branch[0].block[7].um_I.iw[15] ,
    \top_I.branch[0].block[7].um_I.iw[14] ,
    \top_I.branch[0].block[7].um_I.iw[13] ,
    \top_I.branch[0].block[7].um_I.iw[12] ,
    \top_I.branch[0].block[7].um_I.iw[11] ,
    \top_I.branch[0].block[7].um_I.iw[10] ,
    \top_I.branch[0].block[7].um_I.iw[9] ,
    \top_I.branch[0].block[7].um_I.iw[8] ,
    \top_I.branch[0].block[7].um_I.iw[7] ,
    \top_I.branch[0].block[7].um_I.iw[6] ,
    \top_I.branch[0].block[7].um_I.iw[5] ,
    \top_I.branch[0].block[7].um_I.iw[4] ,
    \top_I.branch[0].block[7].um_I.iw[3] ,
    \top_I.branch[0].block[7].um_I.iw[2] ,
    \top_I.branch[0].block[7].um_I.iw[1] ,
    \top_I.branch[0].block[7].um_I.clk ,
    \top_I.branch[0].block[6].um_I.iw[17] ,
    \top_I.branch[0].block[6].um_I.iw[16] ,
    \top_I.branch[0].block[6].um_I.iw[15] ,
    \top_I.branch[0].block[6].um_I.iw[14] ,
    \top_I.branch[0].block[6].um_I.iw[13] ,
    \top_I.branch[0].block[6].um_I.iw[12] ,
    \top_I.branch[0].block[6].um_I.iw[11] ,
    \top_I.branch[0].block[6].um_I.iw[10] ,
    \top_I.branch[0].block[6].um_I.iw[9] ,
    \top_I.branch[0].block[6].um_I.iw[8] ,
    \top_I.branch[0].block[6].um_I.iw[7] ,
    \top_I.branch[0].block[6].um_I.iw[6] ,
    \top_I.branch[0].block[6].um_I.iw[5] ,
    \top_I.branch[0].block[6].um_I.iw[4] ,
    \top_I.branch[0].block[6].um_I.iw[3] ,
    \top_I.branch[0].block[6].um_I.iw[2] ,
    \top_I.branch[0].block[6].um_I.iw[1] ,
    \top_I.branch[0].block[6].um_I.clk ,
    \top_I.branch[0].block[5].um_I.iw[17] ,
    \top_I.branch[0].block[5].um_I.iw[16] ,
    \top_I.branch[0].block[5].um_I.iw[15] ,
    \top_I.branch[0].block[5].um_I.iw[14] ,
    \top_I.branch[0].block[5].um_I.iw[13] ,
    \top_I.branch[0].block[5].um_I.iw[12] ,
    \top_I.branch[0].block[5].um_I.iw[11] ,
    \top_I.branch[0].block[5].um_I.iw[10] ,
    \top_I.branch[0].block[5].um_I.iw[9] ,
    \top_I.branch[0].block[5].um_I.iw[8] ,
    \top_I.branch[0].block[5].um_I.iw[7] ,
    \top_I.branch[0].block[5].um_I.iw[6] ,
    \top_I.branch[0].block[5].um_I.iw[5] ,
    \top_I.branch[0].block[5].um_I.iw[4] ,
    \top_I.branch[0].block[5].um_I.iw[3] ,
    \top_I.branch[0].block[5].um_I.iw[2] ,
    \top_I.branch[0].block[5].um_I.iw[1] ,
    \top_I.branch[0].block[5].um_I.clk ,
    \top_I.branch[0].block[4].um_I.iw[17] ,
    \top_I.branch[0].block[4].um_I.iw[16] ,
    \top_I.branch[0].block[4].um_I.iw[15] ,
    \top_I.branch[0].block[4].um_I.iw[14] ,
    \top_I.branch[0].block[4].um_I.iw[13] ,
    \top_I.branch[0].block[4].um_I.iw[12] ,
    \top_I.branch[0].block[4].um_I.iw[11] ,
    \top_I.branch[0].block[4].um_I.iw[10] ,
    \top_I.branch[0].block[4].um_I.iw[9] ,
    \top_I.branch[0].block[4].um_I.iw[8] ,
    \top_I.branch[0].block[4].um_I.iw[7] ,
    \top_I.branch[0].block[4].um_I.iw[6] ,
    \top_I.branch[0].block[4].um_I.iw[5] ,
    \top_I.branch[0].block[4].um_I.iw[4] ,
    \top_I.branch[0].block[4].um_I.iw[3] ,
    \top_I.branch[0].block[4].um_I.iw[2] ,
    \top_I.branch[0].block[4].um_I.iw[1] ,
    \top_I.branch[0].block[4].um_I.clk ,
    \top_I.branch[0].block[3].um_I.iw[17] ,
    \top_I.branch[0].block[3].um_I.iw[16] ,
    \top_I.branch[0].block[3].um_I.iw[15] ,
    \top_I.branch[0].block[3].um_I.iw[14] ,
    \top_I.branch[0].block[3].um_I.iw[13] ,
    \top_I.branch[0].block[3].um_I.iw[12] ,
    \top_I.branch[0].block[3].um_I.iw[11] ,
    \top_I.branch[0].block[3].um_I.iw[10] ,
    \top_I.branch[0].block[3].um_I.iw[9] ,
    \top_I.branch[0].block[3].um_I.iw[8] ,
    \top_I.branch[0].block[3].um_I.iw[7] ,
    \top_I.branch[0].block[3].um_I.iw[6] ,
    \top_I.branch[0].block[3].um_I.iw[5] ,
    \top_I.branch[0].block[3].um_I.iw[4] ,
    \top_I.branch[0].block[3].um_I.iw[3] ,
    \top_I.branch[0].block[3].um_I.iw[2] ,
    \top_I.branch[0].block[3].um_I.iw[1] ,
    \top_I.branch[0].block[3].um_I.clk ,
    \top_I.branch[0].block[2].um_I.iw[17] ,
    \top_I.branch[0].block[2].um_I.iw[16] ,
    \top_I.branch[0].block[2].um_I.iw[15] ,
    \top_I.branch[0].block[2].um_I.iw[14] ,
    \top_I.branch[0].block[2].um_I.iw[13] ,
    \top_I.branch[0].block[2].um_I.iw[12] ,
    \top_I.branch[0].block[2].um_I.iw[11] ,
    \top_I.branch[0].block[2].um_I.iw[10] ,
    \top_I.branch[0].block[2].um_I.iw[9] ,
    \top_I.branch[0].block[2].um_I.iw[8] ,
    \top_I.branch[0].block[2].um_I.iw[7] ,
    \top_I.branch[0].block[2].um_I.iw[6] ,
    \top_I.branch[0].block[2].um_I.iw[5] ,
    \top_I.branch[0].block[2].um_I.iw[4] ,
    \top_I.branch[0].block[2].um_I.iw[3] ,
    \top_I.branch[0].block[2].um_I.iw[2] ,
    \top_I.branch[0].block[2].um_I.iw[1] ,
    \top_I.branch[0].block[2].um_I.clk ,
    \top_I.branch[0].block[1].um_I.iw[17] ,
    \top_I.branch[0].block[1].um_I.iw[16] ,
    \top_I.branch[0].block[1].um_I.iw[15] ,
    \top_I.branch[0].block[1].um_I.iw[14] ,
    \top_I.branch[0].block[1].um_I.iw[13] ,
    \top_I.branch[0].block[1].um_I.iw[12] ,
    \top_I.branch[0].block[1].um_I.iw[11] ,
    \top_I.branch[0].block[1].um_I.iw[10] ,
    \top_I.branch[0].block[1].um_I.iw[9] ,
    \top_I.branch[0].block[1].um_I.iw[8] ,
    \top_I.branch[0].block[1].um_I.iw[7] ,
    \top_I.branch[0].block[1].um_I.iw[6] ,
    \top_I.branch[0].block[1].um_I.iw[5] ,
    \top_I.branch[0].block[1].um_I.iw[4] ,
    \top_I.branch[0].block[1].um_I.iw[3] ,
    \top_I.branch[0].block[1].um_I.iw[2] ,
    \top_I.branch[0].block[1].um_I.iw[1] ,
    \top_I.branch[0].block[1].um_I.clk ,
    \top_I.branch[0].block[0].um_I.iw[17] ,
    \top_I.branch[0].block[0].um_I.iw[16] ,
    \top_I.branch[0].block[0].um_I.iw[15] ,
    \top_I.branch[0].block[0].um_I.iw[14] ,
    \top_I.branch[0].block[0].um_I.iw[13] ,
    \top_I.branch[0].block[0].um_I.iw[12] ,
    \top_I.branch[0].block[0].um_I.iw[11] ,
    \top_I.branch[0].block[0].um_I.iw[10] ,
    \top_I.branch[0].block[0].um_I.iw[9] ,
    \top_I.branch[0].block[0].um_I.iw[8] ,
    \top_I.branch[0].block[0].um_I.iw[7] ,
    \top_I.branch[0].block[0].um_I.iw[6] ,
    \top_I.branch[0].block[0].um_I.iw[5] ,
    \top_I.branch[0].block[0].um_I.iw[4] ,
    \top_I.branch[0].block[0].um_I.iw[3] ,
    \top_I.branch[0].block[0].um_I.iw[2] ,
    \top_I.branch[0].block[0].um_I.iw[1] ,
    \top_I.branch[0].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[1].um_I.k_zero ,
    \top_I.branch[0].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[15].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[14].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[13].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[12].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[11].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[10].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[9].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[8].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[7].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[6].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[5].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[4].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[3].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[2].um_I.k_zero ,
    \top_I.branch[0].block[1].um_I.ow[23] ,
    \top_I.branch[0].block[1].um_I.ow[22] ,
    \top_I.branch[0].block[1].um_I.ow[21] ,
    \top_I.branch[0].block[1].um_I.ow[20] ,
    \top_I.branch[0].block[1].um_I.ow[19] ,
    \top_I.branch[0].block[1].um_I.ow[18] ,
    \top_I.branch[0].block[1].um_I.ow[17] ,
    \top_I.branch[0].block[1].um_I.ow[16] ,
    \top_I.branch[0].block[1].um_I.ow[15] ,
    \top_I.branch[0].block[1].um_I.ow[14] ,
    \top_I.branch[0].block[1].um_I.ow[13] ,
    \top_I.branch[0].block[1].um_I.ow[12] ,
    \top_I.branch[0].block[1].um_I.ow[11] ,
    \top_I.branch[0].block[1].um_I.ow[10] ,
    \top_I.branch[0].block[1].um_I.ow[9] ,
    \top_I.branch[0].block[1].um_I.ow[8] ,
    \top_I.branch[0].block[1].um_I.ow[7] ,
    \top_I.branch[0].block[1].um_I.ow[6] ,
    \top_I.branch[0].block[1].um_I.ow[5] ,
    \top_I.branch[0].block[1].um_I.ow[4] ,
    \top_I.branch[0].block[1].um_I.ow[3] ,
    \top_I.branch[0].block[1].um_I.ow[2] ,
    \top_I.branch[0].block[1].um_I.ow[1] ,
    \top_I.branch[0].block[1].um_I.ow[0] ,
    \top_I.branch[0].block[0].um_I.ow[23] ,
    \top_I.branch[0].block[0].um_I.ow[22] ,
    \top_I.branch[0].block[0].um_I.ow[21] ,
    \top_I.branch[0].block[0].um_I.ow[20] ,
    \top_I.branch[0].block[0].um_I.ow[19] ,
    \top_I.branch[0].block[0].um_I.ow[18] ,
    \top_I.branch[0].block[0].um_I.ow[17] ,
    \top_I.branch[0].block[0].um_I.ow[16] ,
    \top_I.branch[0].block[0].um_I.ow[15] ,
    \top_I.branch[0].block[0].um_I.ow[14] ,
    \top_I.branch[0].block[0].um_I.ow[13] ,
    \top_I.branch[0].block[0].um_I.ow[12] ,
    \top_I.branch[0].block[0].um_I.ow[11] ,
    \top_I.branch[0].block[0].um_I.ow[10] ,
    \top_I.branch[0].block[0].um_I.ow[9] ,
    \top_I.branch[0].block[0].um_I.ow[8] ,
    \top_I.branch[0].block[0].um_I.ow[7] ,
    \top_I.branch[0].block[0].um_I.ow[6] ,
    \top_I.branch[0].block[0].um_I.ow[5] ,
    \top_I.branch[0].block[0].um_I.ow[4] ,
    \top_I.branch[0].block[0].um_I.ow[3] ,
    \top_I.branch[0].block[0].um_I.ow[2] ,
    \top_I.branch[0].block[0].um_I.ow[1] ,
    \top_I.branch[0].block[0].um_I.ow[0] }),
    .um_pg_vdd({\top_I.branch[0].block[15].um_I.pg_vdd ,
    \top_I.branch[0].block[14].um_I.pg_vdd ,
    \top_I.branch[0].block[13].um_I.pg_vdd ,
    \top_I.branch[0].block[12].um_I.pg_vdd ,
    \top_I.branch[0].block[11].um_I.pg_vdd ,
    \top_I.branch[0].block[10].um_I.pg_vdd ,
    \top_I.branch[0].block[9].um_I.pg_vdd ,
    \top_I.branch[0].block[8].um_I.pg_vdd ,
    \top_I.branch[0].block[7].um_I.pg_vdd ,
    \top_I.branch[0].block[6].um_I.pg_vdd ,
    \top_I.branch[0].block[5].um_I.pg_vdd ,
    \top_I.branch[0].block[4].um_I.pg_vdd ,
    \top_I.branch[0].block[3].um_I.pg_vdd ,
    \top_I.branch[0].block[2].um_I.pg_vdd ,
    \top_I.branch[0].block[1].um_I.pg_vdd ,
    \top_I.branch[0].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[10].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[10].l_addr[0] ),
    .k_zero(\top_I.branch[10].l_addr[1] ),
    .addr({\top_I.branch[10].l_addr[1] ,
    \top_I.branch[10].l_addr[0] ,
    \top_I.branch[10].l_addr[1] ,
    \top_I.branch[10].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[10].block[15].um_I.ena ,
    \top_I.branch[10].block[14].um_I.ena ,
    \top_I.branch[10].block[13].um_I.ena ,
    \top_I.branch[10].block[12].um_I.ena ,
    \top_I.branch[10].block[11].um_I.ena ,
    \top_I.branch[10].block[10].um_I.ena ,
    \top_I.branch[10].block[9].um_I.ena ,
    \top_I.branch[10].block[8].um_I.ena ,
    \top_I.branch[10].block[7].um_I.ena ,
    \top_I.branch[10].block[6].um_I.ena ,
    \top_I.branch[10].block[5].um_I.ena ,
    \top_I.branch[10].block[4].um_I.ena ,
    \top_I.branch[10].block[3].um_I.ena ,
    \top_I.branch[10].block[2].um_I.ena ,
    \top_I.branch[10].block[1].um_I.ena ,
    \top_I.branch[10].block[0].um_I.ena }),
    .um_iw({\top_I.branch[10].block[15].um_I.iw[17] ,
    \top_I.branch[10].block[15].um_I.iw[16] ,
    \top_I.branch[10].block[15].um_I.iw[15] ,
    \top_I.branch[10].block[15].um_I.iw[14] ,
    \top_I.branch[10].block[15].um_I.iw[13] ,
    \top_I.branch[10].block[15].um_I.iw[12] ,
    \top_I.branch[10].block[15].um_I.iw[11] ,
    \top_I.branch[10].block[15].um_I.iw[10] ,
    \top_I.branch[10].block[15].um_I.iw[9] ,
    \top_I.branch[10].block[15].um_I.iw[8] ,
    \top_I.branch[10].block[15].um_I.iw[7] ,
    \top_I.branch[10].block[15].um_I.iw[6] ,
    \top_I.branch[10].block[15].um_I.iw[5] ,
    \top_I.branch[10].block[15].um_I.iw[4] ,
    \top_I.branch[10].block[15].um_I.iw[3] ,
    \top_I.branch[10].block[15].um_I.iw[2] ,
    \top_I.branch[10].block[15].um_I.iw[1] ,
    \top_I.branch[10].block[15].um_I.clk ,
    \top_I.branch[10].block[14].um_I.iw[17] ,
    \top_I.branch[10].block[14].um_I.iw[16] ,
    \top_I.branch[10].block[14].um_I.iw[15] ,
    \top_I.branch[10].block[14].um_I.iw[14] ,
    \top_I.branch[10].block[14].um_I.iw[13] ,
    \top_I.branch[10].block[14].um_I.iw[12] ,
    \top_I.branch[10].block[14].um_I.iw[11] ,
    \top_I.branch[10].block[14].um_I.iw[10] ,
    \top_I.branch[10].block[14].um_I.iw[9] ,
    \top_I.branch[10].block[14].um_I.iw[8] ,
    \top_I.branch[10].block[14].um_I.iw[7] ,
    \top_I.branch[10].block[14].um_I.iw[6] ,
    \top_I.branch[10].block[14].um_I.iw[5] ,
    \top_I.branch[10].block[14].um_I.iw[4] ,
    \top_I.branch[10].block[14].um_I.iw[3] ,
    \top_I.branch[10].block[14].um_I.iw[2] ,
    \top_I.branch[10].block[14].um_I.iw[1] ,
    \top_I.branch[10].block[14].um_I.clk ,
    \top_I.branch[10].block[13].um_I.iw[17] ,
    \top_I.branch[10].block[13].um_I.iw[16] ,
    \top_I.branch[10].block[13].um_I.iw[15] ,
    \top_I.branch[10].block[13].um_I.iw[14] ,
    \top_I.branch[10].block[13].um_I.iw[13] ,
    \top_I.branch[10].block[13].um_I.iw[12] ,
    \top_I.branch[10].block[13].um_I.iw[11] ,
    \top_I.branch[10].block[13].um_I.iw[10] ,
    \top_I.branch[10].block[13].um_I.iw[9] ,
    \top_I.branch[10].block[13].um_I.iw[8] ,
    \top_I.branch[10].block[13].um_I.iw[7] ,
    \top_I.branch[10].block[13].um_I.iw[6] ,
    \top_I.branch[10].block[13].um_I.iw[5] ,
    \top_I.branch[10].block[13].um_I.iw[4] ,
    \top_I.branch[10].block[13].um_I.iw[3] ,
    \top_I.branch[10].block[13].um_I.iw[2] ,
    \top_I.branch[10].block[13].um_I.iw[1] ,
    \top_I.branch[10].block[13].um_I.clk ,
    \top_I.branch[10].block[12].um_I.iw[17] ,
    \top_I.branch[10].block[12].um_I.iw[16] ,
    \top_I.branch[10].block[12].um_I.iw[15] ,
    \top_I.branch[10].block[12].um_I.iw[14] ,
    \top_I.branch[10].block[12].um_I.iw[13] ,
    \top_I.branch[10].block[12].um_I.iw[12] ,
    \top_I.branch[10].block[12].um_I.iw[11] ,
    \top_I.branch[10].block[12].um_I.iw[10] ,
    \top_I.branch[10].block[12].um_I.iw[9] ,
    \top_I.branch[10].block[12].um_I.iw[8] ,
    \top_I.branch[10].block[12].um_I.iw[7] ,
    \top_I.branch[10].block[12].um_I.iw[6] ,
    \top_I.branch[10].block[12].um_I.iw[5] ,
    \top_I.branch[10].block[12].um_I.iw[4] ,
    \top_I.branch[10].block[12].um_I.iw[3] ,
    \top_I.branch[10].block[12].um_I.iw[2] ,
    \top_I.branch[10].block[12].um_I.iw[1] ,
    \top_I.branch[10].block[12].um_I.clk ,
    \top_I.branch[10].block[11].um_I.iw[17] ,
    \top_I.branch[10].block[11].um_I.iw[16] ,
    \top_I.branch[10].block[11].um_I.iw[15] ,
    \top_I.branch[10].block[11].um_I.iw[14] ,
    \top_I.branch[10].block[11].um_I.iw[13] ,
    \top_I.branch[10].block[11].um_I.iw[12] ,
    \top_I.branch[10].block[11].um_I.iw[11] ,
    \top_I.branch[10].block[11].um_I.iw[10] ,
    \top_I.branch[10].block[11].um_I.iw[9] ,
    \top_I.branch[10].block[11].um_I.iw[8] ,
    \top_I.branch[10].block[11].um_I.iw[7] ,
    \top_I.branch[10].block[11].um_I.iw[6] ,
    \top_I.branch[10].block[11].um_I.iw[5] ,
    \top_I.branch[10].block[11].um_I.iw[4] ,
    \top_I.branch[10].block[11].um_I.iw[3] ,
    \top_I.branch[10].block[11].um_I.iw[2] ,
    \top_I.branch[10].block[11].um_I.iw[1] ,
    \top_I.branch[10].block[11].um_I.clk ,
    \top_I.branch[10].block[10].um_I.iw[17] ,
    \top_I.branch[10].block[10].um_I.iw[16] ,
    \top_I.branch[10].block[10].um_I.iw[15] ,
    \top_I.branch[10].block[10].um_I.iw[14] ,
    \top_I.branch[10].block[10].um_I.iw[13] ,
    \top_I.branch[10].block[10].um_I.iw[12] ,
    \top_I.branch[10].block[10].um_I.iw[11] ,
    \top_I.branch[10].block[10].um_I.iw[10] ,
    \top_I.branch[10].block[10].um_I.iw[9] ,
    \top_I.branch[10].block[10].um_I.iw[8] ,
    \top_I.branch[10].block[10].um_I.iw[7] ,
    \top_I.branch[10].block[10].um_I.iw[6] ,
    \top_I.branch[10].block[10].um_I.iw[5] ,
    \top_I.branch[10].block[10].um_I.iw[4] ,
    \top_I.branch[10].block[10].um_I.iw[3] ,
    \top_I.branch[10].block[10].um_I.iw[2] ,
    \top_I.branch[10].block[10].um_I.iw[1] ,
    \top_I.branch[10].block[10].um_I.clk ,
    \top_I.branch[10].block[9].um_I.iw[17] ,
    \top_I.branch[10].block[9].um_I.iw[16] ,
    \top_I.branch[10].block[9].um_I.iw[15] ,
    \top_I.branch[10].block[9].um_I.iw[14] ,
    \top_I.branch[10].block[9].um_I.iw[13] ,
    \top_I.branch[10].block[9].um_I.iw[12] ,
    \top_I.branch[10].block[9].um_I.iw[11] ,
    \top_I.branch[10].block[9].um_I.iw[10] ,
    \top_I.branch[10].block[9].um_I.iw[9] ,
    \top_I.branch[10].block[9].um_I.iw[8] ,
    \top_I.branch[10].block[9].um_I.iw[7] ,
    \top_I.branch[10].block[9].um_I.iw[6] ,
    \top_I.branch[10].block[9].um_I.iw[5] ,
    \top_I.branch[10].block[9].um_I.iw[4] ,
    \top_I.branch[10].block[9].um_I.iw[3] ,
    \top_I.branch[10].block[9].um_I.iw[2] ,
    \top_I.branch[10].block[9].um_I.iw[1] ,
    \top_I.branch[10].block[9].um_I.clk ,
    \top_I.branch[10].block[8].um_I.iw[17] ,
    \top_I.branch[10].block[8].um_I.iw[16] ,
    \top_I.branch[10].block[8].um_I.iw[15] ,
    \top_I.branch[10].block[8].um_I.iw[14] ,
    \top_I.branch[10].block[8].um_I.iw[13] ,
    \top_I.branch[10].block[8].um_I.iw[12] ,
    \top_I.branch[10].block[8].um_I.iw[11] ,
    \top_I.branch[10].block[8].um_I.iw[10] ,
    \top_I.branch[10].block[8].um_I.iw[9] ,
    \top_I.branch[10].block[8].um_I.iw[8] ,
    \top_I.branch[10].block[8].um_I.iw[7] ,
    \top_I.branch[10].block[8].um_I.iw[6] ,
    \top_I.branch[10].block[8].um_I.iw[5] ,
    \top_I.branch[10].block[8].um_I.iw[4] ,
    \top_I.branch[10].block[8].um_I.iw[3] ,
    \top_I.branch[10].block[8].um_I.iw[2] ,
    \top_I.branch[10].block[8].um_I.iw[1] ,
    \top_I.branch[10].block[8].um_I.clk ,
    \top_I.branch[10].block[7].um_I.iw[17] ,
    \top_I.branch[10].block[7].um_I.iw[16] ,
    \top_I.branch[10].block[7].um_I.iw[15] ,
    \top_I.branch[10].block[7].um_I.iw[14] ,
    \top_I.branch[10].block[7].um_I.iw[13] ,
    \top_I.branch[10].block[7].um_I.iw[12] ,
    \top_I.branch[10].block[7].um_I.iw[11] ,
    \top_I.branch[10].block[7].um_I.iw[10] ,
    \top_I.branch[10].block[7].um_I.iw[9] ,
    \top_I.branch[10].block[7].um_I.iw[8] ,
    \top_I.branch[10].block[7].um_I.iw[7] ,
    \top_I.branch[10].block[7].um_I.iw[6] ,
    \top_I.branch[10].block[7].um_I.iw[5] ,
    \top_I.branch[10].block[7].um_I.iw[4] ,
    \top_I.branch[10].block[7].um_I.iw[3] ,
    \top_I.branch[10].block[7].um_I.iw[2] ,
    \top_I.branch[10].block[7].um_I.iw[1] ,
    \top_I.branch[10].block[7].um_I.clk ,
    \top_I.branch[10].block[6].um_I.iw[17] ,
    \top_I.branch[10].block[6].um_I.iw[16] ,
    \top_I.branch[10].block[6].um_I.iw[15] ,
    \top_I.branch[10].block[6].um_I.iw[14] ,
    \top_I.branch[10].block[6].um_I.iw[13] ,
    \top_I.branch[10].block[6].um_I.iw[12] ,
    \top_I.branch[10].block[6].um_I.iw[11] ,
    \top_I.branch[10].block[6].um_I.iw[10] ,
    \top_I.branch[10].block[6].um_I.iw[9] ,
    \top_I.branch[10].block[6].um_I.iw[8] ,
    \top_I.branch[10].block[6].um_I.iw[7] ,
    \top_I.branch[10].block[6].um_I.iw[6] ,
    \top_I.branch[10].block[6].um_I.iw[5] ,
    \top_I.branch[10].block[6].um_I.iw[4] ,
    \top_I.branch[10].block[6].um_I.iw[3] ,
    \top_I.branch[10].block[6].um_I.iw[2] ,
    \top_I.branch[10].block[6].um_I.iw[1] ,
    \top_I.branch[10].block[6].um_I.clk ,
    \top_I.branch[10].block[5].um_I.iw[17] ,
    \top_I.branch[10].block[5].um_I.iw[16] ,
    \top_I.branch[10].block[5].um_I.iw[15] ,
    \top_I.branch[10].block[5].um_I.iw[14] ,
    \top_I.branch[10].block[5].um_I.iw[13] ,
    \top_I.branch[10].block[5].um_I.iw[12] ,
    \top_I.branch[10].block[5].um_I.iw[11] ,
    \top_I.branch[10].block[5].um_I.iw[10] ,
    \top_I.branch[10].block[5].um_I.iw[9] ,
    \top_I.branch[10].block[5].um_I.iw[8] ,
    \top_I.branch[10].block[5].um_I.iw[7] ,
    \top_I.branch[10].block[5].um_I.iw[6] ,
    \top_I.branch[10].block[5].um_I.iw[5] ,
    \top_I.branch[10].block[5].um_I.iw[4] ,
    \top_I.branch[10].block[5].um_I.iw[3] ,
    \top_I.branch[10].block[5].um_I.iw[2] ,
    \top_I.branch[10].block[5].um_I.iw[1] ,
    \top_I.branch[10].block[5].um_I.clk ,
    \top_I.branch[10].block[4].um_I.iw[17] ,
    \top_I.branch[10].block[4].um_I.iw[16] ,
    \top_I.branch[10].block[4].um_I.iw[15] ,
    \top_I.branch[10].block[4].um_I.iw[14] ,
    \top_I.branch[10].block[4].um_I.iw[13] ,
    \top_I.branch[10].block[4].um_I.iw[12] ,
    \top_I.branch[10].block[4].um_I.iw[11] ,
    \top_I.branch[10].block[4].um_I.iw[10] ,
    \top_I.branch[10].block[4].um_I.iw[9] ,
    \top_I.branch[10].block[4].um_I.iw[8] ,
    \top_I.branch[10].block[4].um_I.iw[7] ,
    \top_I.branch[10].block[4].um_I.iw[6] ,
    \top_I.branch[10].block[4].um_I.iw[5] ,
    \top_I.branch[10].block[4].um_I.iw[4] ,
    \top_I.branch[10].block[4].um_I.iw[3] ,
    \top_I.branch[10].block[4].um_I.iw[2] ,
    \top_I.branch[10].block[4].um_I.iw[1] ,
    \top_I.branch[10].block[4].um_I.clk ,
    \top_I.branch[10].block[3].um_I.iw[17] ,
    \top_I.branch[10].block[3].um_I.iw[16] ,
    \top_I.branch[10].block[3].um_I.iw[15] ,
    \top_I.branch[10].block[3].um_I.iw[14] ,
    \top_I.branch[10].block[3].um_I.iw[13] ,
    \top_I.branch[10].block[3].um_I.iw[12] ,
    \top_I.branch[10].block[3].um_I.iw[11] ,
    \top_I.branch[10].block[3].um_I.iw[10] ,
    \top_I.branch[10].block[3].um_I.iw[9] ,
    \top_I.branch[10].block[3].um_I.iw[8] ,
    \top_I.branch[10].block[3].um_I.iw[7] ,
    \top_I.branch[10].block[3].um_I.iw[6] ,
    \top_I.branch[10].block[3].um_I.iw[5] ,
    \top_I.branch[10].block[3].um_I.iw[4] ,
    \top_I.branch[10].block[3].um_I.iw[3] ,
    \top_I.branch[10].block[3].um_I.iw[2] ,
    \top_I.branch[10].block[3].um_I.iw[1] ,
    \top_I.branch[10].block[3].um_I.clk ,
    \top_I.branch[10].block[2].um_I.iw[17] ,
    \top_I.branch[10].block[2].um_I.iw[16] ,
    \top_I.branch[10].block[2].um_I.iw[15] ,
    \top_I.branch[10].block[2].um_I.iw[14] ,
    \top_I.branch[10].block[2].um_I.iw[13] ,
    \top_I.branch[10].block[2].um_I.iw[12] ,
    \top_I.branch[10].block[2].um_I.iw[11] ,
    \top_I.branch[10].block[2].um_I.iw[10] ,
    \top_I.branch[10].block[2].um_I.iw[9] ,
    \top_I.branch[10].block[2].um_I.iw[8] ,
    \top_I.branch[10].block[2].um_I.iw[7] ,
    \top_I.branch[10].block[2].um_I.iw[6] ,
    \top_I.branch[10].block[2].um_I.iw[5] ,
    \top_I.branch[10].block[2].um_I.iw[4] ,
    \top_I.branch[10].block[2].um_I.iw[3] ,
    \top_I.branch[10].block[2].um_I.iw[2] ,
    \top_I.branch[10].block[2].um_I.iw[1] ,
    \top_I.branch[10].block[2].um_I.clk ,
    \top_I.branch[10].block[1].um_I.iw[17] ,
    \top_I.branch[10].block[1].um_I.iw[16] ,
    \top_I.branch[10].block[1].um_I.iw[15] ,
    \top_I.branch[10].block[1].um_I.iw[14] ,
    \top_I.branch[10].block[1].um_I.iw[13] ,
    \top_I.branch[10].block[1].um_I.iw[12] ,
    \top_I.branch[10].block[1].um_I.iw[11] ,
    \top_I.branch[10].block[1].um_I.iw[10] ,
    \top_I.branch[10].block[1].um_I.iw[9] ,
    \top_I.branch[10].block[1].um_I.iw[8] ,
    \top_I.branch[10].block[1].um_I.iw[7] ,
    \top_I.branch[10].block[1].um_I.iw[6] ,
    \top_I.branch[10].block[1].um_I.iw[5] ,
    \top_I.branch[10].block[1].um_I.iw[4] ,
    \top_I.branch[10].block[1].um_I.iw[3] ,
    \top_I.branch[10].block[1].um_I.iw[2] ,
    \top_I.branch[10].block[1].um_I.iw[1] ,
    \top_I.branch[10].block[1].um_I.clk ,
    \top_I.branch[10].block[0].um_I.iw[17] ,
    \top_I.branch[10].block[0].um_I.iw[16] ,
    \top_I.branch[10].block[0].um_I.iw[15] ,
    \top_I.branch[10].block[0].um_I.iw[14] ,
    \top_I.branch[10].block[0].um_I.iw[13] ,
    \top_I.branch[10].block[0].um_I.iw[12] ,
    \top_I.branch[10].block[0].um_I.iw[11] ,
    \top_I.branch[10].block[0].um_I.iw[10] ,
    \top_I.branch[10].block[0].um_I.iw[9] ,
    \top_I.branch[10].block[0].um_I.iw[8] ,
    \top_I.branch[10].block[0].um_I.iw[7] ,
    \top_I.branch[10].block[0].um_I.iw[6] ,
    \top_I.branch[10].block[0].um_I.iw[5] ,
    \top_I.branch[10].block[0].um_I.iw[4] ,
    \top_I.branch[10].block[0].um_I.iw[3] ,
    \top_I.branch[10].block[0].um_I.iw[2] ,
    \top_I.branch[10].block[0].um_I.iw[1] ,
    \top_I.branch[10].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[15].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[14].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[13].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[12].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[11].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[10].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[9].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[8].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[7].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[6].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[5].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[4].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[3].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[2].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[1].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero ,
    \top_I.branch[10].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[10].block[15].um_I.pg_vdd ,
    \top_I.branch[10].block[14].um_I.pg_vdd ,
    \top_I.branch[10].block[13].um_I.pg_vdd ,
    \top_I.branch[10].block[12].um_I.pg_vdd ,
    \top_I.branch[10].block[11].um_I.pg_vdd ,
    \top_I.branch[10].block[10].um_I.pg_vdd ,
    \top_I.branch[10].block[9].um_I.pg_vdd ,
    \top_I.branch[10].block[8].um_I.pg_vdd ,
    \top_I.branch[10].block[7].um_I.pg_vdd ,
    \top_I.branch[10].block[6].um_I.pg_vdd ,
    \top_I.branch[10].block[5].um_I.pg_vdd ,
    \top_I.branch[10].block[4].um_I.pg_vdd ,
    \top_I.branch[10].block[3].um_I.pg_vdd ,
    \top_I.branch[10].block[2].um_I.pg_vdd ,
    \top_I.branch[10].block[1].um_I.pg_vdd ,
    \top_I.branch[10].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[11].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[11].l_addr[0] ),
    .k_zero(\top_I.branch[11].l_addr[1] ),
    .addr({\top_I.branch[11].l_addr[1] ,
    \top_I.branch[11].l_addr[0] ,
    \top_I.branch[11].l_addr[1] ,
    \top_I.branch[11].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[11].block[15].um_I.ena ,
    \top_I.branch[11].block[14].um_I.ena ,
    \top_I.branch[11].block[13].um_I.ena ,
    \top_I.branch[11].block[12].um_I.ena ,
    \top_I.branch[11].block[11].um_I.ena ,
    \top_I.branch[11].block[10].um_I.ena ,
    \top_I.branch[11].block[9].um_I.ena ,
    \top_I.branch[11].block[8].um_I.ena ,
    \top_I.branch[11].block[7].um_I.ena ,
    \top_I.branch[11].block[6].um_I.ena ,
    \top_I.branch[11].block[5].um_I.ena ,
    \top_I.branch[11].block[4].um_I.ena ,
    \top_I.branch[11].block[3].um_I.ena ,
    \top_I.branch[11].block[2].um_I.ena ,
    \top_I.branch[11].block[1].um_I.ena ,
    \top_I.branch[11].block[0].um_I.ena }),
    .um_iw({\top_I.branch[11].block[15].um_I.iw[17] ,
    \top_I.branch[11].block[15].um_I.iw[16] ,
    \top_I.branch[11].block[15].um_I.iw[15] ,
    \top_I.branch[11].block[15].um_I.iw[14] ,
    \top_I.branch[11].block[15].um_I.iw[13] ,
    \top_I.branch[11].block[15].um_I.iw[12] ,
    \top_I.branch[11].block[15].um_I.iw[11] ,
    \top_I.branch[11].block[15].um_I.iw[10] ,
    \top_I.branch[11].block[15].um_I.iw[9] ,
    \top_I.branch[11].block[15].um_I.iw[8] ,
    \top_I.branch[11].block[15].um_I.iw[7] ,
    \top_I.branch[11].block[15].um_I.iw[6] ,
    \top_I.branch[11].block[15].um_I.iw[5] ,
    \top_I.branch[11].block[15].um_I.iw[4] ,
    \top_I.branch[11].block[15].um_I.iw[3] ,
    \top_I.branch[11].block[15].um_I.iw[2] ,
    \top_I.branch[11].block[15].um_I.iw[1] ,
    \top_I.branch[11].block[15].um_I.clk ,
    \top_I.branch[11].block[14].um_I.iw[17] ,
    \top_I.branch[11].block[14].um_I.iw[16] ,
    \top_I.branch[11].block[14].um_I.iw[15] ,
    \top_I.branch[11].block[14].um_I.iw[14] ,
    \top_I.branch[11].block[14].um_I.iw[13] ,
    \top_I.branch[11].block[14].um_I.iw[12] ,
    \top_I.branch[11].block[14].um_I.iw[11] ,
    \top_I.branch[11].block[14].um_I.iw[10] ,
    \top_I.branch[11].block[14].um_I.iw[9] ,
    \top_I.branch[11].block[14].um_I.iw[8] ,
    \top_I.branch[11].block[14].um_I.iw[7] ,
    \top_I.branch[11].block[14].um_I.iw[6] ,
    \top_I.branch[11].block[14].um_I.iw[5] ,
    \top_I.branch[11].block[14].um_I.iw[4] ,
    \top_I.branch[11].block[14].um_I.iw[3] ,
    \top_I.branch[11].block[14].um_I.iw[2] ,
    \top_I.branch[11].block[14].um_I.iw[1] ,
    \top_I.branch[11].block[14].um_I.clk ,
    \top_I.branch[11].block[13].um_I.iw[17] ,
    \top_I.branch[11].block[13].um_I.iw[16] ,
    \top_I.branch[11].block[13].um_I.iw[15] ,
    \top_I.branch[11].block[13].um_I.iw[14] ,
    \top_I.branch[11].block[13].um_I.iw[13] ,
    \top_I.branch[11].block[13].um_I.iw[12] ,
    \top_I.branch[11].block[13].um_I.iw[11] ,
    \top_I.branch[11].block[13].um_I.iw[10] ,
    \top_I.branch[11].block[13].um_I.iw[9] ,
    \top_I.branch[11].block[13].um_I.iw[8] ,
    \top_I.branch[11].block[13].um_I.iw[7] ,
    \top_I.branch[11].block[13].um_I.iw[6] ,
    \top_I.branch[11].block[13].um_I.iw[5] ,
    \top_I.branch[11].block[13].um_I.iw[4] ,
    \top_I.branch[11].block[13].um_I.iw[3] ,
    \top_I.branch[11].block[13].um_I.iw[2] ,
    \top_I.branch[11].block[13].um_I.iw[1] ,
    \top_I.branch[11].block[13].um_I.clk ,
    \top_I.branch[11].block[12].um_I.iw[17] ,
    \top_I.branch[11].block[12].um_I.iw[16] ,
    \top_I.branch[11].block[12].um_I.iw[15] ,
    \top_I.branch[11].block[12].um_I.iw[14] ,
    \top_I.branch[11].block[12].um_I.iw[13] ,
    \top_I.branch[11].block[12].um_I.iw[12] ,
    \top_I.branch[11].block[12].um_I.iw[11] ,
    \top_I.branch[11].block[12].um_I.iw[10] ,
    \top_I.branch[11].block[12].um_I.iw[9] ,
    \top_I.branch[11].block[12].um_I.iw[8] ,
    \top_I.branch[11].block[12].um_I.iw[7] ,
    \top_I.branch[11].block[12].um_I.iw[6] ,
    \top_I.branch[11].block[12].um_I.iw[5] ,
    \top_I.branch[11].block[12].um_I.iw[4] ,
    \top_I.branch[11].block[12].um_I.iw[3] ,
    \top_I.branch[11].block[12].um_I.iw[2] ,
    \top_I.branch[11].block[12].um_I.iw[1] ,
    \top_I.branch[11].block[12].um_I.clk ,
    \top_I.branch[11].block[11].um_I.iw[17] ,
    \top_I.branch[11].block[11].um_I.iw[16] ,
    \top_I.branch[11].block[11].um_I.iw[15] ,
    \top_I.branch[11].block[11].um_I.iw[14] ,
    \top_I.branch[11].block[11].um_I.iw[13] ,
    \top_I.branch[11].block[11].um_I.iw[12] ,
    \top_I.branch[11].block[11].um_I.iw[11] ,
    \top_I.branch[11].block[11].um_I.iw[10] ,
    \top_I.branch[11].block[11].um_I.iw[9] ,
    \top_I.branch[11].block[11].um_I.iw[8] ,
    \top_I.branch[11].block[11].um_I.iw[7] ,
    \top_I.branch[11].block[11].um_I.iw[6] ,
    \top_I.branch[11].block[11].um_I.iw[5] ,
    \top_I.branch[11].block[11].um_I.iw[4] ,
    \top_I.branch[11].block[11].um_I.iw[3] ,
    \top_I.branch[11].block[11].um_I.iw[2] ,
    \top_I.branch[11].block[11].um_I.iw[1] ,
    \top_I.branch[11].block[11].um_I.clk ,
    \top_I.branch[11].block[10].um_I.iw[17] ,
    \top_I.branch[11].block[10].um_I.iw[16] ,
    \top_I.branch[11].block[10].um_I.iw[15] ,
    \top_I.branch[11].block[10].um_I.iw[14] ,
    \top_I.branch[11].block[10].um_I.iw[13] ,
    \top_I.branch[11].block[10].um_I.iw[12] ,
    \top_I.branch[11].block[10].um_I.iw[11] ,
    \top_I.branch[11].block[10].um_I.iw[10] ,
    \top_I.branch[11].block[10].um_I.iw[9] ,
    \top_I.branch[11].block[10].um_I.iw[8] ,
    \top_I.branch[11].block[10].um_I.iw[7] ,
    \top_I.branch[11].block[10].um_I.iw[6] ,
    \top_I.branch[11].block[10].um_I.iw[5] ,
    \top_I.branch[11].block[10].um_I.iw[4] ,
    \top_I.branch[11].block[10].um_I.iw[3] ,
    \top_I.branch[11].block[10].um_I.iw[2] ,
    \top_I.branch[11].block[10].um_I.iw[1] ,
    \top_I.branch[11].block[10].um_I.clk ,
    \top_I.branch[11].block[9].um_I.iw[17] ,
    \top_I.branch[11].block[9].um_I.iw[16] ,
    \top_I.branch[11].block[9].um_I.iw[15] ,
    \top_I.branch[11].block[9].um_I.iw[14] ,
    \top_I.branch[11].block[9].um_I.iw[13] ,
    \top_I.branch[11].block[9].um_I.iw[12] ,
    \top_I.branch[11].block[9].um_I.iw[11] ,
    \top_I.branch[11].block[9].um_I.iw[10] ,
    \top_I.branch[11].block[9].um_I.iw[9] ,
    \top_I.branch[11].block[9].um_I.iw[8] ,
    \top_I.branch[11].block[9].um_I.iw[7] ,
    \top_I.branch[11].block[9].um_I.iw[6] ,
    \top_I.branch[11].block[9].um_I.iw[5] ,
    \top_I.branch[11].block[9].um_I.iw[4] ,
    \top_I.branch[11].block[9].um_I.iw[3] ,
    \top_I.branch[11].block[9].um_I.iw[2] ,
    \top_I.branch[11].block[9].um_I.iw[1] ,
    \top_I.branch[11].block[9].um_I.clk ,
    \top_I.branch[11].block[8].um_I.iw[17] ,
    \top_I.branch[11].block[8].um_I.iw[16] ,
    \top_I.branch[11].block[8].um_I.iw[15] ,
    \top_I.branch[11].block[8].um_I.iw[14] ,
    \top_I.branch[11].block[8].um_I.iw[13] ,
    \top_I.branch[11].block[8].um_I.iw[12] ,
    \top_I.branch[11].block[8].um_I.iw[11] ,
    \top_I.branch[11].block[8].um_I.iw[10] ,
    \top_I.branch[11].block[8].um_I.iw[9] ,
    \top_I.branch[11].block[8].um_I.iw[8] ,
    \top_I.branch[11].block[8].um_I.iw[7] ,
    \top_I.branch[11].block[8].um_I.iw[6] ,
    \top_I.branch[11].block[8].um_I.iw[5] ,
    \top_I.branch[11].block[8].um_I.iw[4] ,
    \top_I.branch[11].block[8].um_I.iw[3] ,
    \top_I.branch[11].block[8].um_I.iw[2] ,
    \top_I.branch[11].block[8].um_I.iw[1] ,
    \top_I.branch[11].block[8].um_I.clk ,
    \top_I.branch[11].block[7].um_I.iw[17] ,
    \top_I.branch[11].block[7].um_I.iw[16] ,
    \top_I.branch[11].block[7].um_I.iw[15] ,
    \top_I.branch[11].block[7].um_I.iw[14] ,
    \top_I.branch[11].block[7].um_I.iw[13] ,
    \top_I.branch[11].block[7].um_I.iw[12] ,
    \top_I.branch[11].block[7].um_I.iw[11] ,
    \top_I.branch[11].block[7].um_I.iw[10] ,
    \top_I.branch[11].block[7].um_I.iw[9] ,
    \top_I.branch[11].block[7].um_I.iw[8] ,
    \top_I.branch[11].block[7].um_I.iw[7] ,
    \top_I.branch[11].block[7].um_I.iw[6] ,
    \top_I.branch[11].block[7].um_I.iw[5] ,
    \top_I.branch[11].block[7].um_I.iw[4] ,
    \top_I.branch[11].block[7].um_I.iw[3] ,
    \top_I.branch[11].block[7].um_I.iw[2] ,
    \top_I.branch[11].block[7].um_I.iw[1] ,
    \top_I.branch[11].block[7].um_I.clk ,
    \top_I.branch[11].block[6].um_I.iw[17] ,
    \top_I.branch[11].block[6].um_I.iw[16] ,
    \top_I.branch[11].block[6].um_I.iw[15] ,
    \top_I.branch[11].block[6].um_I.iw[14] ,
    \top_I.branch[11].block[6].um_I.iw[13] ,
    \top_I.branch[11].block[6].um_I.iw[12] ,
    \top_I.branch[11].block[6].um_I.iw[11] ,
    \top_I.branch[11].block[6].um_I.iw[10] ,
    \top_I.branch[11].block[6].um_I.iw[9] ,
    \top_I.branch[11].block[6].um_I.iw[8] ,
    \top_I.branch[11].block[6].um_I.iw[7] ,
    \top_I.branch[11].block[6].um_I.iw[6] ,
    \top_I.branch[11].block[6].um_I.iw[5] ,
    \top_I.branch[11].block[6].um_I.iw[4] ,
    \top_I.branch[11].block[6].um_I.iw[3] ,
    \top_I.branch[11].block[6].um_I.iw[2] ,
    \top_I.branch[11].block[6].um_I.iw[1] ,
    \top_I.branch[11].block[6].um_I.clk ,
    \top_I.branch[11].block[5].um_I.iw[17] ,
    \top_I.branch[11].block[5].um_I.iw[16] ,
    \top_I.branch[11].block[5].um_I.iw[15] ,
    \top_I.branch[11].block[5].um_I.iw[14] ,
    \top_I.branch[11].block[5].um_I.iw[13] ,
    \top_I.branch[11].block[5].um_I.iw[12] ,
    \top_I.branch[11].block[5].um_I.iw[11] ,
    \top_I.branch[11].block[5].um_I.iw[10] ,
    \top_I.branch[11].block[5].um_I.iw[9] ,
    \top_I.branch[11].block[5].um_I.iw[8] ,
    \top_I.branch[11].block[5].um_I.iw[7] ,
    \top_I.branch[11].block[5].um_I.iw[6] ,
    \top_I.branch[11].block[5].um_I.iw[5] ,
    \top_I.branch[11].block[5].um_I.iw[4] ,
    \top_I.branch[11].block[5].um_I.iw[3] ,
    \top_I.branch[11].block[5].um_I.iw[2] ,
    \top_I.branch[11].block[5].um_I.iw[1] ,
    \top_I.branch[11].block[5].um_I.clk ,
    \top_I.branch[11].block[4].um_I.iw[17] ,
    \top_I.branch[11].block[4].um_I.iw[16] ,
    \top_I.branch[11].block[4].um_I.iw[15] ,
    \top_I.branch[11].block[4].um_I.iw[14] ,
    \top_I.branch[11].block[4].um_I.iw[13] ,
    \top_I.branch[11].block[4].um_I.iw[12] ,
    \top_I.branch[11].block[4].um_I.iw[11] ,
    \top_I.branch[11].block[4].um_I.iw[10] ,
    \top_I.branch[11].block[4].um_I.iw[9] ,
    \top_I.branch[11].block[4].um_I.iw[8] ,
    \top_I.branch[11].block[4].um_I.iw[7] ,
    \top_I.branch[11].block[4].um_I.iw[6] ,
    \top_I.branch[11].block[4].um_I.iw[5] ,
    \top_I.branch[11].block[4].um_I.iw[4] ,
    \top_I.branch[11].block[4].um_I.iw[3] ,
    \top_I.branch[11].block[4].um_I.iw[2] ,
    \top_I.branch[11].block[4].um_I.iw[1] ,
    \top_I.branch[11].block[4].um_I.clk ,
    \top_I.branch[11].block[3].um_I.iw[17] ,
    \top_I.branch[11].block[3].um_I.iw[16] ,
    \top_I.branch[11].block[3].um_I.iw[15] ,
    \top_I.branch[11].block[3].um_I.iw[14] ,
    \top_I.branch[11].block[3].um_I.iw[13] ,
    \top_I.branch[11].block[3].um_I.iw[12] ,
    \top_I.branch[11].block[3].um_I.iw[11] ,
    \top_I.branch[11].block[3].um_I.iw[10] ,
    \top_I.branch[11].block[3].um_I.iw[9] ,
    \top_I.branch[11].block[3].um_I.iw[8] ,
    \top_I.branch[11].block[3].um_I.iw[7] ,
    \top_I.branch[11].block[3].um_I.iw[6] ,
    \top_I.branch[11].block[3].um_I.iw[5] ,
    \top_I.branch[11].block[3].um_I.iw[4] ,
    \top_I.branch[11].block[3].um_I.iw[3] ,
    \top_I.branch[11].block[3].um_I.iw[2] ,
    \top_I.branch[11].block[3].um_I.iw[1] ,
    \top_I.branch[11].block[3].um_I.clk ,
    \top_I.branch[11].block[2].um_I.iw[17] ,
    \top_I.branch[11].block[2].um_I.iw[16] ,
    \top_I.branch[11].block[2].um_I.iw[15] ,
    \top_I.branch[11].block[2].um_I.iw[14] ,
    \top_I.branch[11].block[2].um_I.iw[13] ,
    \top_I.branch[11].block[2].um_I.iw[12] ,
    \top_I.branch[11].block[2].um_I.iw[11] ,
    \top_I.branch[11].block[2].um_I.iw[10] ,
    \top_I.branch[11].block[2].um_I.iw[9] ,
    \top_I.branch[11].block[2].um_I.iw[8] ,
    \top_I.branch[11].block[2].um_I.iw[7] ,
    \top_I.branch[11].block[2].um_I.iw[6] ,
    \top_I.branch[11].block[2].um_I.iw[5] ,
    \top_I.branch[11].block[2].um_I.iw[4] ,
    \top_I.branch[11].block[2].um_I.iw[3] ,
    \top_I.branch[11].block[2].um_I.iw[2] ,
    \top_I.branch[11].block[2].um_I.iw[1] ,
    \top_I.branch[11].block[2].um_I.clk ,
    \top_I.branch[11].block[1].um_I.iw[17] ,
    \top_I.branch[11].block[1].um_I.iw[16] ,
    \top_I.branch[11].block[1].um_I.iw[15] ,
    \top_I.branch[11].block[1].um_I.iw[14] ,
    \top_I.branch[11].block[1].um_I.iw[13] ,
    \top_I.branch[11].block[1].um_I.iw[12] ,
    \top_I.branch[11].block[1].um_I.iw[11] ,
    \top_I.branch[11].block[1].um_I.iw[10] ,
    \top_I.branch[11].block[1].um_I.iw[9] ,
    \top_I.branch[11].block[1].um_I.iw[8] ,
    \top_I.branch[11].block[1].um_I.iw[7] ,
    \top_I.branch[11].block[1].um_I.iw[6] ,
    \top_I.branch[11].block[1].um_I.iw[5] ,
    \top_I.branch[11].block[1].um_I.iw[4] ,
    \top_I.branch[11].block[1].um_I.iw[3] ,
    \top_I.branch[11].block[1].um_I.iw[2] ,
    \top_I.branch[11].block[1].um_I.iw[1] ,
    \top_I.branch[11].block[1].um_I.clk ,
    \top_I.branch[11].block[0].um_I.iw[17] ,
    \top_I.branch[11].block[0].um_I.iw[16] ,
    \top_I.branch[11].block[0].um_I.iw[15] ,
    \top_I.branch[11].block[0].um_I.iw[14] ,
    \top_I.branch[11].block[0].um_I.iw[13] ,
    \top_I.branch[11].block[0].um_I.iw[12] ,
    \top_I.branch[11].block[0].um_I.iw[11] ,
    \top_I.branch[11].block[0].um_I.iw[10] ,
    \top_I.branch[11].block[0].um_I.iw[9] ,
    \top_I.branch[11].block[0].um_I.iw[8] ,
    \top_I.branch[11].block[0].um_I.iw[7] ,
    \top_I.branch[11].block[0].um_I.iw[6] ,
    \top_I.branch[11].block[0].um_I.iw[5] ,
    \top_I.branch[11].block[0].um_I.iw[4] ,
    \top_I.branch[11].block[0].um_I.iw[3] ,
    \top_I.branch[11].block[0].um_I.iw[2] ,
    \top_I.branch[11].block[0].um_I.iw[1] ,
    \top_I.branch[11].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[15].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[14].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[13].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[12].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[11].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[10].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[9].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[8].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[7].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[6].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[5].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[4].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[3].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[2].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[1].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero ,
    \top_I.branch[11].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[11].block[15].um_I.pg_vdd ,
    \top_I.branch[11].block[14].um_I.pg_vdd ,
    \top_I.branch[11].block[13].um_I.pg_vdd ,
    \top_I.branch[11].block[12].um_I.pg_vdd ,
    \top_I.branch[11].block[11].um_I.pg_vdd ,
    \top_I.branch[11].block[10].um_I.pg_vdd ,
    \top_I.branch[11].block[9].um_I.pg_vdd ,
    \top_I.branch[11].block[8].um_I.pg_vdd ,
    \top_I.branch[11].block[7].um_I.pg_vdd ,
    \top_I.branch[11].block[6].um_I.pg_vdd ,
    \top_I.branch[11].block[5].um_I.pg_vdd ,
    \top_I.branch[11].block[4].um_I.pg_vdd ,
    \top_I.branch[11].block[3].um_I.pg_vdd ,
    \top_I.branch[11].block[2].um_I.pg_vdd ,
    \top_I.branch[11].block[1].um_I.pg_vdd ,
    \top_I.branch[11].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[12].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[12].l_addr[1] ),
    .k_zero(\top_I.branch[12].l_addr[0] ),
    .addr({\top_I.branch[12].l_addr[0] ,
    \top_I.branch[12].l_addr[1] ,
    \top_I.branch[12].l_addr[1] ,
    \top_I.branch[12].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[12].block[15].um_I.ena ,
    \top_I.branch[12].block[14].um_I.ena ,
    \top_I.branch[12].block[13].um_I.ena ,
    \top_I.branch[12].block[12].um_I.ena ,
    \top_I.branch[12].block[11].um_I.ena ,
    \top_I.branch[12].block[10].um_I.ena ,
    \top_I.branch[12].block[9].um_I.ena ,
    \top_I.branch[12].block[8].um_I.ena ,
    \top_I.branch[12].block[7].um_I.ena ,
    \top_I.branch[12].block[6].um_I.ena ,
    \top_I.branch[12].block[5].um_I.ena ,
    \top_I.branch[12].block[4].um_I.ena ,
    \top_I.branch[12].block[3].um_I.ena ,
    \top_I.branch[12].block[2].um_I.ena ,
    \top_I.branch[12].block[1].um_I.ena ,
    \top_I.branch[12].block[0].um_I.ena }),
    .um_iw({\top_I.branch[12].block[15].um_I.iw[17] ,
    \top_I.branch[12].block[15].um_I.iw[16] ,
    \top_I.branch[12].block[15].um_I.iw[15] ,
    \top_I.branch[12].block[15].um_I.iw[14] ,
    \top_I.branch[12].block[15].um_I.iw[13] ,
    \top_I.branch[12].block[15].um_I.iw[12] ,
    \top_I.branch[12].block[15].um_I.iw[11] ,
    \top_I.branch[12].block[15].um_I.iw[10] ,
    \top_I.branch[12].block[15].um_I.iw[9] ,
    \top_I.branch[12].block[15].um_I.iw[8] ,
    \top_I.branch[12].block[15].um_I.iw[7] ,
    \top_I.branch[12].block[15].um_I.iw[6] ,
    \top_I.branch[12].block[15].um_I.iw[5] ,
    \top_I.branch[12].block[15].um_I.iw[4] ,
    \top_I.branch[12].block[15].um_I.iw[3] ,
    \top_I.branch[12].block[15].um_I.iw[2] ,
    \top_I.branch[12].block[15].um_I.iw[1] ,
    \top_I.branch[12].block[15].um_I.clk ,
    \top_I.branch[12].block[14].um_I.iw[17] ,
    \top_I.branch[12].block[14].um_I.iw[16] ,
    \top_I.branch[12].block[14].um_I.iw[15] ,
    \top_I.branch[12].block[14].um_I.iw[14] ,
    \top_I.branch[12].block[14].um_I.iw[13] ,
    \top_I.branch[12].block[14].um_I.iw[12] ,
    \top_I.branch[12].block[14].um_I.iw[11] ,
    \top_I.branch[12].block[14].um_I.iw[10] ,
    \top_I.branch[12].block[14].um_I.iw[9] ,
    \top_I.branch[12].block[14].um_I.iw[8] ,
    \top_I.branch[12].block[14].um_I.iw[7] ,
    \top_I.branch[12].block[14].um_I.iw[6] ,
    \top_I.branch[12].block[14].um_I.iw[5] ,
    \top_I.branch[12].block[14].um_I.iw[4] ,
    \top_I.branch[12].block[14].um_I.iw[3] ,
    \top_I.branch[12].block[14].um_I.iw[2] ,
    \top_I.branch[12].block[14].um_I.iw[1] ,
    \top_I.branch[12].block[14].um_I.clk ,
    \top_I.branch[12].block[13].um_I.iw[17] ,
    \top_I.branch[12].block[13].um_I.iw[16] ,
    \top_I.branch[12].block[13].um_I.iw[15] ,
    \top_I.branch[12].block[13].um_I.iw[14] ,
    \top_I.branch[12].block[13].um_I.iw[13] ,
    \top_I.branch[12].block[13].um_I.iw[12] ,
    \top_I.branch[12].block[13].um_I.iw[11] ,
    \top_I.branch[12].block[13].um_I.iw[10] ,
    \top_I.branch[12].block[13].um_I.iw[9] ,
    \top_I.branch[12].block[13].um_I.iw[8] ,
    \top_I.branch[12].block[13].um_I.iw[7] ,
    \top_I.branch[12].block[13].um_I.iw[6] ,
    \top_I.branch[12].block[13].um_I.iw[5] ,
    \top_I.branch[12].block[13].um_I.iw[4] ,
    \top_I.branch[12].block[13].um_I.iw[3] ,
    \top_I.branch[12].block[13].um_I.iw[2] ,
    \top_I.branch[12].block[13].um_I.iw[1] ,
    \top_I.branch[12].block[13].um_I.clk ,
    \top_I.branch[12].block[12].um_I.iw[17] ,
    \top_I.branch[12].block[12].um_I.iw[16] ,
    \top_I.branch[12].block[12].um_I.iw[15] ,
    \top_I.branch[12].block[12].um_I.iw[14] ,
    \top_I.branch[12].block[12].um_I.iw[13] ,
    \top_I.branch[12].block[12].um_I.iw[12] ,
    \top_I.branch[12].block[12].um_I.iw[11] ,
    \top_I.branch[12].block[12].um_I.iw[10] ,
    \top_I.branch[12].block[12].um_I.iw[9] ,
    \top_I.branch[12].block[12].um_I.iw[8] ,
    \top_I.branch[12].block[12].um_I.iw[7] ,
    \top_I.branch[12].block[12].um_I.iw[6] ,
    \top_I.branch[12].block[12].um_I.iw[5] ,
    \top_I.branch[12].block[12].um_I.iw[4] ,
    \top_I.branch[12].block[12].um_I.iw[3] ,
    \top_I.branch[12].block[12].um_I.iw[2] ,
    \top_I.branch[12].block[12].um_I.iw[1] ,
    \top_I.branch[12].block[12].um_I.clk ,
    \top_I.branch[12].block[11].um_I.iw[17] ,
    \top_I.branch[12].block[11].um_I.iw[16] ,
    \top_I.branch[12].block[11].um_I.iw[15] ,
    \top_I.branch[12].block[11].um_I.iw[14] ,
    \top_I.branch[12].block[11].um_I.iw[13] ,
    \top_I.branch[12].block[11].um_I.iw[12] ,
    \top_I.branch[12].block[11].um_I.iw[11] ,
    \top_I.branch[12].block[11].um_I.iw[10] ,
    \top_I.branch[12].block[11].um_I.iw[9] ,
    \top_I.branch[12].block[11].um_I.iw[8] ,
    \top_I.branch[12].block[11].um_I.iw[7] ,
    \top_I.branch[12].block[11].um_I.iw[6] ,
    \top_I.branch[12].block[11].um_I.iw[5] ,
    \top_I.branch[12].block[11].um_I.iw[4] ,
    \top_I.branch[12].block[11].um_I.iw[3] ,
    \top_I.branch[12].block[11].um_I.iw[2] ,
    \top_I.branch[12].block[11].um_I.iw[1] ,
    \top_I.branch[12].block[11].um_I.clk ,
    \top_I.branch[12].block[10].um_I.iw[17] ,
    \top_I.branch[12].block[10].um_I.iw[16] ,
    \top_I.branch[12].block[10].um_I.iw[15] ,
    \top_I.branch[12].block[10].um_I.iw[14] ,
    \top_I.branch[12].block[10].um_I.iw[13] ,
    \top_I.branch[12].block[10].um_I.iw[12] ,
    \top_I.branch[12].block[10].um_I.iw[11] ,
    \top_I.branch[12].block[10].um_I.iw[10] ,
    \top_I.branch[12].block[10].um_I.iw[9] ,
    \top_I.branch[12].block[10].um_I.iw[8] ,
    \top_I.branch[12].block[10].um_I.iw[7] ,
    \top_I.branch[12].block[10].um_I.iw[6] ,
    \top_I.branch[12].block[10].um_I.iw[5] ,
    \top_I.branch[12].block[10].um_I.iw[4] ,
    \top_I.branch[12].block[10].um_I.iw[3] ,
    \top_I.branch[12].block[10].um_I.iw[2] ,
    \top_I.branch[12].block[10].um_I.iw[1] ,
    \top_I.branch[12].block[10].um_I.clk ,
    \top_I.branch[12].block[9].um_I.iw[17] ,
    \top_I.branch[12].block[9].um_I.iw[16] ,
    \top_I.branch[12].block[9].um_I.iw[15] ,
    \top_I.branch[12].block[9].um_I.iw[14] ,
    \top_I.branch[12].block[9].um_I.iw[13] ,
    \top_I.branch[12].block[9].um_I.iw[12] ,
    \top_I.branch[12].block[9].um_I.iw[11] ,
    \top_I.branch[12].block[9].um_I.iw[10] ,
    \top_I.branch[12].block[9].um_I.iw[9] ,
    \top_I.branch[12].block[9].um_I.iw[8] ,
    \top_I.branch[12].block[9].um_I.iw[7] ,
    \top_I.branch[12].block[9].um_I.iw[6] ,
    \top_I.branch[12].block[9].um_I.iw[5] ,
    \top_I.branch[12].block[9].um_I.iw[4] ,
    \top_I.branch[12].block[9].um_I.iw[3] ,
    \top_I.branch[12].block[9].um_I.iw[2] ,
    \top_I.branch[12].block[9].um_I.iw[1] ,
    \top_I.branch[12].block[9].um_I.clk ,
    \top_I.branch[12].block[8].um_I.iw[17] ,
    \top_I.branch[12].block[8].um_I.iw[16] ,
    \top_I.branch[12].block[8].um_I.iw[15] ,
    \top_I.branch[12].block[8].um_I.iw[14] ,
    \top_I.branch[12].block[8].um_I.iw[13] ,
    \top_I.branch[12].block[8].um_I.iw[12] ,
    \top_I.branch[12].block[8].um_I.iw[11] ,
    \top_I.branch[12].block[8].um_I.iw[10] ,
    \top_I.branch[12].block[8].um_I.iw[9] ,
    \top_I.branch[12].block[8].um_I.iw[8] ,
    \top_I.branch[12].block[8].um_I.iw[7] ,
    \top_I.branch[12].block[8].um_I.iw[6] ,
    \top_I.branch[12].block[8].um_I.iw[5] ,
    \top_I.branch[12].block[8].um_I.iw[4] ,
    \top_I.branch[12].block[8].um_I.iw[3] ,
    \top_I.branch[12].block[8].um_I.iw[2] ,
    \top_I.branch[12].block[8].um_I.iw[1] ,
    \top_I.branch[12].block[8].um_I.clk ,
    \top_I.branch[12].block[7].um_I.iw[17] ,
    \top_I.branch[12].block[7].um_I.iw[16] ,
    \top_I.branch[12].block[7].um_I.iw[15] ,
    \top_I.branch[12].block[7].um_I.iw[14] ,
    \top_I.branch[12].block[7].um_I.iw[13] ,
    \top_I.branch[12].block[7].um_I.iw[12] ,
    \top_I.branch[12].block[7].um_I.iw[11] ,
    \top_I.branch[12].block[7].um_I.iw[10] ,
    \top_I.branch[12].block[7].um_I.iw[9] ,
    \top_I.branch[12].block[7].um_I.iw[8] ,
    \top_I.branch[12].block[7].um_I.iw[7] ,
    \top_I.branch[12].block[7].um_I.iw[6] ,
    \top_I.branch[12].block[7].um_I.iw[5] ,
    \top_I.branch[12].block[7].um_I.iw[4] ,
    \top_I.branch[12].block[7].um_I.iw[3] ,
    \top_I.branch[12].block[7].um_I.iw[2] ,
    \top_I.branch[12].block[7].um_I.iw[1] ,
    \top_I.branch[12].block[7].um_I.clk ,
    \top_I.branch[12].block[6].um_I.iw[17] ,
    \top_I.branch[12].block[6].um_I.iw[16] ,
    \top_I.branch[12].block[6].um_I.iw[15] ,
    \top_I.branch[12].block[6].um_I.iw[14] ,
    \top_I.branch[12].block[6].um_I.iw[13] ,
    \top_I.branch[12].block[6].um_I.iw[12] ,
    \top_I.branch[12].block[6].um_I.iw[11] ,
    \top_I.branch[12].block[6].um_I.iw[10] ,
    \top_I.branch[12].block[6].um_I.iw[9] ,
    \top_I.branch[12].block[6].um_I.iw[8] ,
    \top_I.branch[12].block[6].um_I.iw[7] ,
    \top_I.branch[12].block[6].um_I.iw[6] ,
    \top_I.branch[12].block[6].um_I.iw[5] ,
    \top_I.branch[12].block[6].um_I.iw[4] ,
    \top_I.branch[12].block[6].um_I.iw[3] ,
    \top_I.branch[12].block[6].um_I.iw[2] ,
    \top_I.branch[12].block[6].um_I.iw[1] ,
    \top_I.branch[12].block[6].um_I.clk ,
    \top_I.branch[12].block[5].um_I.iw[17] ,
    \top_I.branch[12].block[5].um_I.iw[16] ,
    \top_I.branch[12].block[5].um_I.iw[15] ,
    \top_I.branch[12].block[5].um_I.iw[14] ,
    \top_I.branch[12].block[5].um_I.iw[13] ,
    \top_I.branch[12].block[5].um_I.iw[12] ,
    \top_I.branch[12].block[5].um_I.iw[11] ,
    \top_I.branch[12].block[5].um_I.iw[10] ,
    \top_I.branch[12].block[5].um_I.iw[9] ,
    \top_I.branch[12].block[5].um_I.iw[8] ,
    \top_I.branch[12].block[5].um_I.iw[7] ,
    \top_I.branch[12].block[5].um_I.iw[6] ,
    \top_I.branch[12].block[5].um_I.iw[5] ,
    \top_I.branch[12].block[5].um_I.iw[4] ,
    \top_I.branch[12].block[5].um_I.iw[3] ,
    \top_I.branch[12].block[5].um_I.iw[2] ,
    \top_I.branch[12].block[5].um_I.iw[1] ,
    \top_I.branch[12].block[5].um_I.clk ,
    \top_I.branch[12].block[4].um_I.iw[17] ,
    \top_I.branch[12].block[4].um_I.iw[16] ,
    \top_I.branch[12].block[4].um_I.iw[15] ,
    \top_I.branch[12].block[4].um_I.iw[14] ,
    \top_I.branch[12].block[4].um_I.iw[13] ,
    \top_I.branch[12].block[4].um_I.iw[12] ,
    \top_I.branch[12].block[4].um_I.iw[11] ,
    \top_I.branch[12].block[4].um_I.iw[10] ,
    \top_I.branch[12].block[4].um_I.iw[9] ,
    \top_I.branch[12].block[4].um_I.iw[8] ,
    \top_I.branch[12].block[4].um_I.iw[7] ,
    \top_I.branch[12].block[4].um_I.iw[6] ,
    \top_I.branch[12].block[4].um_I.iw[5] ,
    \top_I.branch[12].block[4].um_I.iw[4] ,
    \top_I.branch[12].block[4].um_I.iw[3] ,
    \top_I.branch[12].block[4].um_I.iw[2] ,
    \top_I.branch[12].block[4].um_I.iw[1] ,
    \top_I.branch[12].block[4].um_I.clk ,
    \top_I.branch[12].block[3].um_I.iw[17] ,
    \top_I.branch[12].block[3].um_I.iw[16] ,
    \top_I.branch[12].block[3].um_I.iw[15] ,
    \top_I.branch[12].block[3].um_I.iw[14] ,
    \top_I.branch[12].block[3].um_I.iw[13] ,
    \top_I.branch[12].block[3].um_I.iw[12] ,
    \top_I.branch[12].block[3].um_I.iw[11] ,
    \top_I.branch[12].block[3].um_I.iw[10] ,
    \top_I.branch[12].block[3].um_I.iw[9] ,
    \top_I.branch[12].block[3].um_I.iw[8] ,
    \top_I.branch[12].block[3].um_I.iw[7] ,
    \top_I.branch[12].block[3].um_I.iw[6] ,
    \top_I.branch[12].block[3].um_I.iw[5] ,
    \top_I.branch[12].block[3].um_I.iw[4] ,
    \top_I.branch[12].block[3].um_I.iw[3] ,
    \top_I.branch[12].block[3].um_I.iw[2] ,
    \top_I.branch[12].block[3].um_I.iw[1] ,
    \top_I.branch[12].block[3].um_I.clk ,
    \top_I.branch[12].block[2].um_I.iw[17] ,
    \top_I.branch[12].block[2].um_I.iw[16] ,
    \top_I.branch[12].block[2].um_I.iw[15] ,
    \top_I.branch[12].block[2].um_I.iw[14] ,
    \top_I.branch[12].block[2].um_I.iw[13] ,
    \top_I.branch[12].block[2].um_I.iw[12] ,
    \top_I.branch[12].block[2].um_I.iw[11] ,
    \top_I.branch[12].block[2].um_I.iw[10] ,
    \top_I.branch[12].block[2].um_I.iw[9] ,
    \top_I.branch[12].block[2].um_I.iw[8] ,
    \top_I.branch[12].block[2].um_I.iw[7] ,
    \top_I.branch[12].block[2].um_I.iw[6] ,
    \top_I.branch[12].block[2].um_I.iw[5] ,
    \top_I.branch[12].block[2].um_I.iw[4] ,
    \top_I.branch[12].block[2].um_I.iw[3] ,
    \top_I.branch[12].block[2].um_I.iw[2] ,
    \top_I.branch[12].block[2].um_I.iw[1] ,
    \top_I.branch[12].block[2].um_I.clk ,
    \top_I.branch[12].block[1].um_I.iw[17] ,
    \top_I.branch[12].block[1].um_I.iw[16] ,
    \top_I.branch[12].block[1].um_I.iw[15] ,
    \top_I.branch[12].block[1].um_I.iw[14] ,
    \top_I.branch[12].block[1].um_I.iw[13] ,
    \top_I.branch[12].block[1].um_I.iw[12] ,
    \top_I.branch[12].block[1].um_I.iw[11] ,
    \top_I.branch[12].block[1].um_I.iw[10] ,
    \top_I.branch[12].block[1].um_I.iw[9] ,
    \top_I.branch[12].block[1].um_I.iw[8] ,
    \top_I.branch[12].block[1].um_I.iw[7] ,
    \top_I.branch[12].block[1].um_I.iw[6] ,
    \top_I.branch[12].block[1].um_I.iw[5] ,
    \top_I.branch[12].block[1].um_I.iw[4] ,
    \top_I.branch[12].block[1].um_I.iw[3] ,
    \top_I.branch[12].block[1].um_I.iw[2] ,
    \top_I.branch[12].block[1].um_I.iw[1] ,
    \top_I.branch[12].block[1].um_I.clk ,
    \top_I.branch[12].block[0].um_I.iw[17] ,
    \top_I.branch[12].block[0].um_I.iw[16] ,
    \top_I.branch[12].block[0].um_I.iw[15] ,
    \top_I.branch[12].block[0].um_I.iw[14] ,
    \top_I.branch[12].block[0].um_I.iw[13] ,
    \top_I.branch[12].block[0].um_I.iw[12] ,
    \top_I.branch[12].block[0].um_I.iw[11] ,
    \top_I.branch[12].block[0].um_I.iw[10] ,
    \top_I.branch[12].block[0].um_I.iw[9] ,
    \top_I.branch[12].block[0].um_I.iw[8] ,
    \top_I.branch[12].block[0].um_I.iw[7] ,
    \top_I.branch[12].block[0].um_I.iw[6] ,
    \top_I.branch[12].block[0].um_I.iw[5] ,
    \top_I.branch[12].block[0].um_I.iw[4] ,
    \top_I.branch[12].block[0].um_I.iw[3] ,
    \top_I.branch[12].block[0].um_I.iw[2] ,
    \top_I.branch[12].block[0].um_I.iw[1] ,
    \top_I.branch[12].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[15].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[14].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[13].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[12].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[11].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[10].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[9].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[8].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[7].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[6].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[5].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[4].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[3].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[2].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[1].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero ,
    \top_I.branch[12].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[12].block[15].um_I.pg_vdd ,
    \top_I.branch[12].block[14].um_I.pg_vdd ,
    \top_I.branch[12].block[13].um_I.pg_vdd ,
    \top_I.branch[12].block[12].um_I.pg_vdd ,
    \top_I.branch[12].block[11].um_I.pg_vdd ,
    \top_I.branch[12].block[10].um_I.pg_vdd ,
    \top_I.branch[12].block[9].um_I.pg_vdd ,
    \top_I.branch[12].block[8].um_I.pg_vdd ,
    \top_I.branch[12].block[7].um_I.pg_vdd ,
    \top_I.branch[12].block[6].um_I.pg_vdd ,
    \top_I.branch[12].block[5].um_I.pg_vdd ,
    \top_I.branch[12].block[4].um_I.pg_vdd ,
    \top_I.branch[12].block[3].um_I.pg_vdd ,
    \top_I.branch[12].block[2].um_I.pg_vdd ,
    \top_I.branch[12].block[1].um_I.pg_vdd ,
    \top_I.branch[12].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[13].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[13].l_addr[1] ),
    .k_zero(\top_I.branch[13].l_addr[0] ),
    .addr({\top_I.branch[13].l_addr[0] ,
    \top_I.branch[13].l_addr[1] ,
    \top_I.branch[13].l_addr[1] ,
    \top_I.branch[13].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[13].block[15].um_I.ena ,
    \top_I.branch[13].block[14].um_I.ena ,
    \top_I.branch[13].block[13].um_I.ena ,
    \top_I.branch[13].block[12].um_I.ena ,
    \top_I.branch[13].block[11].um_I.ena ,
    \top_I.branch[13].block[10].um_I.ena ,
    \top_I.branch[13].block[9].um_I.ena ,
    \top_I.branch[13].block[8].um_I.ena ,
    \top_I.branch[13].block[7].um_I.ena ,
    \top_I.branch[13].block[6].um_I.ena ,
    \top_I.branch[13].block[5].um_I.ena ,
    \top_I.branch[13].block[4].um_I.ena ,
    \top_I.branch[13].block[3].um_I.ena ,
    \top_I.branch[13].block[2].um_I.ena ,
    \top_I.branch[13].block[1].um_I.ena ,
    \top_I.branch[13].block[0].um_I.ena }),
    .um_iw({\top_I.branch[13].block[15].um_I.iw[17] ,
    \top_I.branch[13].block[15].um_I.iw[16] ,
    \top_I.branch[13].block[15].um_I.iw[15] ,
    \top_I.branch[13].block[15].um_I.iw[14] ,
    \top_I.branch[13].block[15].um_I.iw[13] ,
    \top_I.branch[13].block[15].um_I.iw[12] ,
    \top_I.branch[13].block[15].um_I.iw[11] ,
    \top_I.branch[13].block[15].um_I.iw[10] ,
    \top_I.branch[13].block[15].um_I.iw[9] ,
    \top_I.branch[13].block[15].um_I.iw[8] ,
    \top_I.branch[13].block[15].um_I.iw[7] ,
    \top_I.branch[13].block[15].um_I.iw[6] ,
    \top_I.branch[13].block[15].um_I.iw[5] ,
    \top_I.branch[13].block[15].um_I.iw[4] ,
    \top_I.branch[13].block[15].um_I.iw[3] ,
    \top_I.branch[13].block[15].um_I.iw[2] ,
    \top_I.branch[13].block[15].um_I.iw[1] ,
    \top_I.branch[13].block[15].um_I.clk ,
    \top_I.branch[13].block[14].um_I.iw[17] ,
    \top_I.branch[13].block[14].um_I.iw[16] ,
    \top_I.branch[13].block[14].um_I.iw[15] ,
    \top_I.branch[13].block[14].um_I.iw[14] ,
    \top_I.branch[13].block[14].um_I.iw[13] ,
    \top_I.branch[13].block[14].um_I.iw[12] ,
    \top_I.branch[13].block[14].um_I.iw[11] ,
    \top_I.branch[13].block[14].um_I.iw[10] ,
    \top_I.branch[13].block[14].um_I.iw[9] ,
    \top_I.branch[13].block[14].um_I.iw[8] ,
    \top_I.branch[13].block[14].um_I.iw[7] ,
    \top_I.branch[13].block[14].um_I.iw[6] ,
    \top_I.branch[13].block[14].um_I.iw[5] ,
    \top_I.branch[13].block[14].um_I.iw[4] ,
    \top_I.branch[13].block[14].um_I.iw[3] ,
    \top_I.branch[13].block[14].um_I.iw[2] ,
    \top_I.branch[13].block[14].um_I.iw[1] ,
    \top_I.branch[13].block[14].um_I.clk ,
    \top_I.branch[13].block[13].um_I.iw[17] ,
    \top_I.branch[13].block[13].um_I.iw[16] ,
    \top_I.branch[13].block[13].um_I.iw[15] ,
    \top_I.branch[13].block[13].um_I.iw[14] ,
    \top_I.branch[13].block[13].um_I.iw[13] ,
    \top_I.branch[13].block[13].um_I.iw[12] ,
    \top_I.branch[13].block[13].um_I.iw[11] ,
    \top_I.branch[13].block[13].um_I.iw[10] ,
    \top_I.branch[13].block[13].um_I.iw[9] ,
    \top_I.branch[13].block[13].um_I.iw[8] ,
    \top_I.branch[13].block[13].um_I.iw[7] ,
    \top_I.branch[13].block[13].um_I.iw[6] ,
    \top_I.branch[13].block[13].um_I.iw[5] ,
    \top_I.branch[13].block[13].um_I.iw[4] ,
    \top_I.branch[13].block[13].um_I.iw[3] ,
    \top_I.branch[13].block[13].um_I.iw[2] ,
    \top_I.branch[13].block[13].um_I.iw[1] ,
    \top_I.branch[13].block[13].um_I.clk ,
    \top_I.branch[13].block[12].um_I.iw[17] ,
    \top_I.branch[13].block[12].um_I.iw[16] ,
    \top_I.branch[13].block[12].um_I.iw[15] ,
    \top_I.branch[13].block[12].um_I.iw[14] ,
    \top_I.branch[13].block[12].um_I.iw[13] ,
    \top_I.branch[13].block[12].um_I.iw[12] ,
    \top_I.branch[13].block[12].um_I.iw[11] ,
    \top_I.branch[13].block[12].um_I.iw[10] ,
    \top_I.branch[13].block[12].um_I.iw[9] ,
    \top_I.branch[13].block[12].um_I.iw[8] ,
    \top_I.branch[13].block[12].um_I.iw[7] ,
    \top_I.branch[13].block[12].um_I.iw[6] ,
    \top_I.branch[13].block[12].um_I.iw[5] ,
    \top_I.branch[13].block[12].um_I.iw[4] ,
    \top_I.branch[13].block[12].um_I.iw[3] ,
    \top_I.branch[13].block[12].um_I.iw[2] ,
    \top_I.branch[13].block[12].um_I.iw[1] ,
    \top_I.branch[13].block[12].um_I.clk ,
    \top_I.branch[13].block[11].um_I.iw[17] ,
    \top_I.branch[13].block[11].um_I.iw[16] ,
    \top_I.branch[13].block[11].um_I.iw[15] ,
    \top_I.branch[13].block[11].um_I.iw[14] ,
    \top_I.branch[13].block[11].um_I.iw[13] ,
    \top_I.branch[13].block[11].um_I.iw[12] ,
    \top_I.branch[13].block[11].um_I.iw[11] ,
    \top_I.branch[13].block[11].um_I.iw[10] ,
    \top_I.branch[13].block[11].um_I.iw[9] ,
    \top_I.branch[13].block[11].um_I.iw[8] ,
    \top_I.branch[13].block[11].um_I.iw[7] ,
    \top_I.branch[13].block[11].um_I.iw[6] ,
    \top_I.branch[13].block[11].um_I.iw[5] ,
    \top_I.branch[13].block[11].um_I.iw[4] ,
    \top_I.branch[13].block[11].um_I.iw[3] ,
    \top_I.branch[13].block[11].um_I.iw[2] ,
    \top_I.branch[13].block[11].um_I.iw[1] ,
    \top_I.branch[13].block[11].um_I.clk ,
    \top_I.branch[13].block[10].um_I.iw[17] ,
    \top_I.branch[13].block[10].um_I.iw[16] ,
    \top_I.branch[13].block[10].um_I.iw[15] ,
    \top_I.branch[13].block[10].um_I.iw[14] ,
    \top_I.branch[13].block[10].um_I.iw[13] ,
    \top_I.branch[13].block[10].um_I.iw[12] ,
    \top_I.branch[13].block[10].um_I.iw[11] ,
    \top_I.branch[13].block[10].um_I.iw[10] ,
    \top_I.branch[13].block[10].um_I.iw[9] ,
    \top_I.branch[13].block[10].um_I.iw[8] ,
    \top_I.branch[13].block[10].um_I.iw[7] ,
    \top_I.branch[13].block[10].um_I.iw[6] ,
    \top_I.branch[13].block[10].um_I.iw[5] ,
    \top_I.branch[13].block[10].um_I.iw[4] ,
    \top_I.branch[13].block[10].um_I.iw[3] ,
    \top_I.branch[13].block[10].um_I.iw[2] ,
    \top_I.branch[13].block[10].um_I.iw[1] ,
    \top_I.branch[13].block[10].um_I.clk ,
    \top_I.branch[13].block[9].um_I.iw[17] ,
    \top_I.branch[13].block[9].um_I.iw[16] ,
    \top_I.branch[13].block[9].um_I.iw[15] ,
    \top_I.branch[13].block[9].um_I.iw[14] ,
    \top_I.branch[13].block[9].um_I.iw[13] ,
    \top_I.branch[13].block[9].um_I.iw[12] ,
    \top_I.branch[13].block[9].um_I.iw[11] ,
    \top_I.branch[13].block[9].um_I.iw[10] ,
    \top_I.branch[13].block[9].um_I.iw[9] ,
    \top_I.branch[13].block[9].um_I.iw[8] ,
    \top_I.branch[13].block[9].um_I.iw[7] ,
    \top_I.branch[13].block[9].um_I.iw[6] ,
    \top_I.branch[13].block[9].um_I.iw[5] ,
    \top_I.branch[13].block[9].um_I.iw[4] ,
    \top_I.branch[13].block[9].um_I.iw[3] ,
    \top_I.branch[13].block[9].um_I.iw[2] ,
    \top_I.branch[13].block[9].um_I.iw[1] ,
    \top_I.branch[13].block[9].um_I.clk ,
    \top_I.branch[13].block[8].um_I.iw[17] ,
    \top_I.branch[13].block[8].um_I.iw[16] ,
    \top_I.branch[13].block[8].um_I.iw[15] ,
    \top_I.branch[13].block[8].um_I.iw[14] ,
    \top_I.branch[13].block[8].um_I.iw[13] ,
    \top_I.branch[13].block[8].um_I.iw[12] ,
    \top_I.branch[13].block[8].um_I.iw[11] ,
    \top_I.branch[13].block[8].um_I.iw[10] ,
    \top_I.branch[13].block[8].um_I.iw[9] ,
    \top_I.branch[13].block[8].um_I.iw[8] ,
    \top_I.branch[13].block[8].um_I.iw[7] ,
    \top_I.branch[13].block[8].um_I.iw[6] ,
    \top_I.branch[13].block[8].um_I.iw[5] ,
    \top_I.branch[13].block[8].um_I.iw[4] ,
    \top_I.branch[13].block[8].um_I.iw[3] ,
    \top_I.branch[13].block[8].um_I.iw[2] ,
    \top_I.branch[13].block[8].um_I.iw[1] ,
    \top_I.branch[13].block[8].um_I.clk ,
    \top_I.branch[13].block[7].um_I.iw[17] ,
    \top_I.branch[13].block[7].um_I.iw[16] ,
    \top_I.branch[13].block[7].um_I.iw[15] ,
    \top_I.branch[13].block[7].um_I.iw[14] ,
    \top_I.branch[13].block[7].um_I.iw[13] ,
    \top_I.branch[13].block[7].um_I.iw[12] ,
    \top_I.branch[13].block[7].um_I.iw[11] ,
    \top_I.branch[13].block[7].um_I.iw[10] ,
    \top_I.branch[13].block[7].um_I.iw[9] ,
    \top_I.branch[13].block[7].um_I.iw[8] ,
    \top_I.branch[13].block[7].um_I.iw[7] ,
    \top_I.branch[13].block[7].um_I.iw[6] ,
    \top_I.branch[13].block[7].um_I.iw[5] ,
    \top_I.branch[13].block[7].um_I.iw[4] ,
    \top_I.branch[13].block[7].um_I.iw[3] ,
    \top_I.branch[13].block[7].um_I.iw[2] ,
    \top_I.branch[13].block[7].um_I.iw[1] ,
    \top_I.branch[13].block[7].um_I.clk ,
    \top_I.branch[13].block[6].um_I.iw[17] ,
    \top_I.branch[13].block[6].um_I.iw[16] ,
    \top_I.branch[13].block[6].um_I.iw[15] ,
    \top_I.branch[13].block[6].um_I.iw[14] ,
    \top_I.branch[13].block[6].um_I.iw[13] ,
    \top_I.branch[13].block[6].um_I.iw[12] ,
    \top_I.branch[13].block[6].um_I.iw[11] ,
    \top_I.branch[13].block[6].um_I.iw[10] ,
    \top_I.branch[13].block[6].um_I.iw[9] ,
    \top_I.branch[13].block[6].um_I.iw[8] ,
    \top_I.branch[13].block[6].um_I.iw[7] ,
    \top_I.branch[13].block[6].um_I.iw[6] ,
    \top_I.branch[13].block[6].um_I.iw[5] ,
    \top_I.branch[13].block[6].um_I.iw[4] ,
    \top_I.branch[13].block[6].um_I.iw[3] ,
    \top_I.branch[13].block[6].um_I.iw[2] ,
    \top_I.branch[13].block[6].um_I.iw[1] ,
    \top_I.branch[13].block[6].um_I.clk ,
    \top_I.branch[13].block[5].um_I.iw[17] ,
    \top_I.branch[13].block[5].um_I.iw[16] ,
    \top_I.branch[13].block[5].um_I.iw[15] ,
    \top_I.branch[13].block[5].um_I.iw[14] ,
    \top_I.branch[13].block[5].um_I.iw[13] ,
    \top_I.branch[13].block[5].um_I.iw[12] ,
    \top_I.branch[13].block[5].um_I.iw[11] ,
    \top_I.branch[13].block[5].um_I.iw[10] ,
    \top_I.branch[13].block[5].um_I.iw[9] ,
    \top_I.branch[13].block[5].um_I.iw[8] ,
    \top_I.branch[13].block[5].um_I.iw[7] ,
    \top_I.branch[13].block[5].um_I.iw[6] ,
    \top_I.branch[13].block[5].um_I.iw[5] ,
    \top_I.branch[13].block[5].um_I.iw[4] ,
    \top_I.branch[13].block[5].um_I.iw[3] ,
    \top_I.branch[13].block[5].um_I.iw[2] ,
    \top_I.branch[13].block[5].um_I.iw[1] ,
    \top_I.branch[13].block[5].um_I.clk ,
    \top_I.branch[13].block[4].um_I.iw[17] ,
    \top_I.branch[13].block[4].um_I.iw[16] ,
    \top_I.branch[13].block[4].um_I.iw[15] ,
    \top_I.branch[13].block[4].um_I.iw[14] ,
    \top_I.branch[13].block[4].um_I.iw[13] ,
    \top_I.branch[13].block[4].um_I.iw[12] ,
    \top_I.branch[13].block[4].um_I.iw[11] ,
    \top_I.branch[13].block[4].um_I.iw[10] ,
    \top_I.branch[13].block[4].um_I.iw[9] ,
    \top_I.branch[13].block[4].um_I.iw[8] ,
    \top_I.branch[13].block[4].um_I.iw[7] ,
    \top_I.branch[13].block[4].um_I.iw[6] ,
    \top_I.branch[13].block[4].um_I.iw[5] ,
    \top_I.branch[13].block[4].um_I.iw[4] ,
    \top_I.branch[13].block[4].um_I.iw[3] ,
    \top_I.branch[13].block[4].um_I.iw[2] ,
    \top_I.branch[13].block[4].um_I.iw[1] ,
    \top_I.branch[13].block[4].um_I.clk ,
    \top_I.branch[13].block[3].um_I.iw[17] ,
    \top_I.branch[13].block[3].um_I.iw[16] ,
    \top_I.branch[13].block[3].um_I.iw[15] ,
    \top_I.branch[13].block[3].um_I.iw[14] ,
    \top_I.branch[13].block[3].um_I.iw[13] ,
    \top_I.branch[13].block[3].um_I.iw[12] ,
    \top_I.branch[13].block[3].um_I.iw[11] ,
    \top_I.branch[13].block[3].um_I.iw[10] ,
    \top_I.branch[13].block[3].um_I.iw[9] ,
    \top_I.branch[13].block[3].um_I.iw[8] ,
    \top_I.branch[13].block[3].um_I.iw[7] ,
    \top_I.branch[13].block[3].um_I.iw[6] ,
    \top_I.branch[13].block[3].um_I.iw[5] ,
    \top_I.branch[13].block[3].um_I.iw[4] ,
    \top_I.branch[13].block[3].um_I.iw[3] ,
    \top_I.branch[13].block[3].um_I.iw[2] ,
    \top_I.branch[13].block[3].um_I.iw[1] ,
    \top_I.branch[13].block[3].um_I.clk ,
    \top_I.branch[13].block[2].um_I.iw[17] ,
    \top_I.branch[13].block[2].um_I.iw[16] ,
    \top_I.branch[13].block[2].um_I.iw[15] ,
    \top_I.branch[13].block[2].um_I.iw[14] ,
    \top_I.branch[13].block[2].um_I.iw[13] ,
    \top_I.branch[13].block[2].um_I.iw[12] ,
    \top_I.branch[13].block[2].um_I.iw[11] ,
    \top_I.branch[13].block[2].um_I.iw[10] ,
    \top_I.branch[13].block[2].um_I.iw[9] ,
    \top_I.branch[13].block[2].um_I.iw[8] ,
    \top_I.branch[13].block[2].um_I.iw[7] ,
    \top_I.branch[13].block[2].um_I.iw[6] ,
    \top_I.branch[13].block[2].um_I.iw[5] ,
    \top_I.branch[13].block[2].um_I.iw[4] ,
    \top_I.branch[13].block[2].um_I.iw[3] ,
    \top_I.branch[13].block[2].um_I.iw[2] ,
    \top_I.branch[13].block[2].um_I.iw[1] ,
    \top_I.branch[13].block[2].um_I.clk ,
    \top_I.branch[13].block[1].um_I.iw[17] ,
    \top_I.branch[13].block[1].um_I.iw[16] ,
    \top_I.branch[13].block[1].um_I.iw[15] ,
    \top_I.branch[13].block[1].um_I.iw[14] ,
    \top_I.branch[13].block[1].um_I.iw[13] ,
    \top_I.branch[13].block[1].um_I.iw[12] ,
    \top_I.branch[13].block[1].um_I.iw[11] ,
    \top_I.branch[13].block[1].um_I.iw[10] ,
    \top_I.branch[13].block[1].um_I.iw[9] ,
    \top_I.branch[13].block[1].um_I.iw[8] ,
    \top_I.branch[13].block[1].um_I.iw[7] ,
    \top_I.branch[13].block[1].um_I.iw[6] ,
    \top_I.branch[13].block[1].um_I.iw[5] ,
    \top_I.branch[13].block[1].um_I.iw[4] ,
    \top_I.branch[13].block[1].um_I.iw[3] ,
    \top_I.branch[13].block[1].um_I.iw[2] ,
    \top_I.branch[13].block[1].um_I.iw[1] ,
    \top_I.branch[13].block[1].um_I.clk ,
    \top_I.branch[13].block[0].um_I.iw[17] ,
    \top_I.branch[13].block[0].um_I.iw[16] ,
    \top_I.branch[13].block[0].um_I.iw[15] ,
    \top_I.branch[13].block[0].um_I.iw[14] ,
    \top_I.branch[13].block[0].um_I.iw[13] ,
    \top_I.branch[13].block[0].um_I.iw[12] ,
    \top_I.branch[13].block[0].um_I.iw[11] ,
    \top_I.branch[13].block[0].um_I.iw[10] ,
    \top_I.branch[13].block[0].um_I.iw[9] ,
    \top_I.branch[13].block[0].um_I.iw[8] ,
    \top_I.branch[13].block[0].um_I.iw[7] ,
    \top_I.branch[13].block[0].um_I.iw[6] ,
    \top_I.branch[13].block[0].um_I.iw[5] ,
    \top_I.branch[13].block[0].um_I.iw[4] ,
    \top_I.branch[13].block[0].um_I.iw[3] ,
    \top_I.branch[13].block[0].um_I.iw[2] ,
    \top_I.branch[13].block[0].um_I.iw[1] ,
    \top_I.branch[13].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[15].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[14].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[13].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[12].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[11].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[10].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[9].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[8].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[7].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[6].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[5].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[4].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[3].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[2].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[1].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero ,
    \top_I.branch[13].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[13].block[15].um_I.pg_vdd ,
    \top_I.branch[13].block[14].um_I.pg_vdd ,
    \top_I.branch[13].block[13].um_I.pg_vdd ,
    \top_I.branch[13].block[12].um_I.pg_vdd ,
    \top_I.branch[13].block[11].um_I.pg_vdd ,
    \top_I.branch[13].block[10].um_I.pg_vdd ,
    \top_I.branch[13].block[9].um_I.pg_vdd ,
    \top_I.branch[13].block[8].um_I.pg_vdd ,
    \top_I.branch[13].block[7].um_I.pg_vdd ,
    \top_I.branch[13].block[6].um_I.pg_vdd ,
    \top_I.branch[13].block[5].um_I.pg_vdd ,
    \top_I.branch[13].block[4].um_I.pg_vdd ,
    \top_I.branch[13].block[3].um_I.pg_vdd ,
    \top_I.branch[13].block[2].um_I.pg_vdd ,
    \top_I.branch[13].block[1].um_I.pg_vdd ,
    \top_I.branch[13].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[14].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[14].l_addr[0] ),
    .k_zero(\top_I.branch[14].l_addr[3] ),
    .addr({\top_I.branch[14].l_addr[3] ,
    \top_I.branch[14].l_addr[0] ,
    \top_I.branch[14].l_addr[0] ,
    \top_I.branch[14].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[14].block[15].um_I.ena ,
    \top_I.branch[14].block[14].um_I.ena ,
    \top_I.branch[14].block[13].um_I.ena ,
    \top_I.branch[14].block[12].um_I.ena ,
    \top_I.branch[14].block[11].um_I.ena ,
    \top_I.branch[14].block[10].um_I.ena ,
    \top_I.branch[14].block[9].um_I.ena ,
    \top_I.branch[14].block[8].um_I.ena ,
    \top_I.branch[14].block[7].um_I.ena ,
    \top_I.branch[14].block[6].um_I.ena ,
    \top_I.branch[14].block[5].um_I.ena ,
    \top_I.branch[14].block[4].um_I.ena ,
    \top_I.branch[14].block[3].um_I.ena ,
    \top_I.branch[14].block[2].um_I.ena ,
    \top_I.branch[14].block[1].um_I.ena ,
    \top_I.branch[14].block[0].um_I.ena }),
    .um_iw({\top_I.branch[14].block[15].um_I.iw[17] ,
    \top_I.branch[14].block[15].um_I.iw[16] ,
    \top_I.branch[14].block[15].um_I.iw[15] ,
    \top_I.branch[14].block[15].um_I.iw[14] ,
    \top_I.branch[14].block[15].um_I.iw[13] ,
    \top_I.branch[14].block[15].um_I.iw[12] ,
    \top_I.branch[14].block[15].um_I.iw[11] ,
    \top_I.branch[14].block[15].um_I.iw[10] ,
    \top_I.branch[14].block[15].um_I.iw[9] ,
    \top_I.branch[14].block[15].um_I.iw[8] ,
    \top_I.branch[14].block[15].um_I.iw[7] ,
    \top_I.branch[14].block[15].um_I.iw[6] ,
    \top_I.branch[14].block[15].um_I.iw[5] ,
    \top_I.branch[14].block[15].um_I.iw[4] ,
    \top_I.branch[14].block[15].um_I.iw[3] ,
    \top_I.branch[14].block[15].um_I.iw[2] ,
    \top_I.branch[14].block[15].um_I.iw[1] ,
    \top_I.branch[14].block[15].um_I.clk ,
    \top_I.branch[14].block[14].um_I.iw[17] ,
    \top_I.branch[14].block[14].um_I.iw[16] ,
    \top_I.branch[14].block[14].um_I.iw[15] ,
    \top_I.branch[14].block[14].um_I.iw[14] ,
    \top_I.branch[14].block[14].um_I.iw[13] ,
    \top_I.branch[14].block[14].um_I.iw[12] ,
    \top_I.branch[14].block[14].um_I.iw[11] ,
    \top_I.branch[14].block[14].um_I.iw[10] ,
    \top_I.branch[14].block[14].um_I.iw[9] ,
    \top_I.branch[14].block[14].um_I.iw[8] ,
    \top_I.branch[14].block[14].um_I.iw[7] ,
    \top_I.branch[14].block[14].um_I.iw[6] ,
    \top_I.branch[14].block[14].um_I.iw[5] ,
    \top_I.branch[14].block[14].um_I.iw[4] ,
    \top_I.branch[14].block[14].um_I.iw[3] ,
    \top_I.branch[14].block[14].um_I.iw[2] ,
    \top_I.branch[14].block[14].um_I.iw[1] ,
    \top_I.branch[14].block[14].um_I.clk ,
    \top_I.branch[14].block[13].um_I.iw[17] ,
    \top_I.branch[14].block[13].um_I.iw[16] ,
    \top_I.branch[14].block[13].um_I.iw[15] ,
    \top_I.branch[14].block[13].um_I.iw[14] ,
    \top_I.branch[14].block[13].um_I.iw[13] ,
    \top_I.branch[14].block[13].um_I.iw[12] ,
    \top_I.branch[14].block[13].um_I.iw[11] ,
    \top_I.branch[14].block[13].um_I.iw[10] ,
    \top_I.branch[14].block[13].um_I.iw[9] ,
    \top_I.branch[14].block[13].um_I.iw[8] ,
    \top_I.branch[14].block[13].um_I.iw[7] ,
    \top_I.branch[14].block[13].um_I.iw[6] ,
    \top_I.branch[14].block[13].um_I.iw[5] ,
    \top_I.branch[14].block[13].um_I.iw[4] ,
    \top_I.branch[14].block[13].um_I.iw[3] ,
    \top_I.branch[14].block[13].um_I.iw[2] ,
    \top_I.branch[14].block[13].um_I.iw[1] ,
    \top_I.branch[14].block[13].um_I.clk ,
    \top_I.branch[14].block[12].um_I.iw[17] ,
    \top_I.branch[14].block[12].um_I.iw[16] ,
    \top_I.branch[14].block[12].um_I.iw[15] ,
    \top_I.branch[14].block[12].um_I.iw[14] ,
    \top_I.branch[14].block[12].um_I.iw[13] ,
    \top_I.branch[14].block[12].um_I.iw[12] ,
    \top_I.branch[14].block[12].um_I.iw[11] ,
    \top_I.branch[14].block[12].um_I.iw[10] ,
    \top_I.branch[14].block[12].um_I.iw[9] ,
    \top_I.branch[14].block[12].um_I.iw[8] ,
    \top_I.branch[14].block[12].um_I.iw[7] ,
    \top_I.branch[14].block[12].um_I.iw[6] ,
    \top_I.branch[14].block[12].um_I.iw[5] ,
    \top_I.branch[14].block[12].um_I.iw[4] ,
    \top_I.branch[14].block[12].um_I.iw[3] ,
    \top_I.branch[14].block[12].um_I.iw[2] ,
    \top_I.branch[14].block[12].um_I.iw[1] ,
    \top_I.branch[14].block[12].um_I.clk ,
    \top_I.branch[14].block[11].um_I.iw[17] ,
    \top_I.branch[14].block[11].um_I.iw[16] ,
    \top_I.branch[14].block[11].um_I.iw[15] ,
    \top_I.branch[14].block[11].um_I.iw[14] ,
    \top_I.branch[14].block[11].um_I.iw[13] ,
    \top_I.branch[14].block[11].um_I.iw[12] ,
    \top_I.branch[14].block[11].um_I.iw[11] ,
    \top_I.branch[14].block[11].um_I.iw[10] ,
    \top_I.branch[14].block[11].um_I.iw[9] ,
    \top_I.branch[14].block[11].um_I.iw[8] ,
    \top_I.branch[14].block[11].um_I.iw[7] ,
    \top_I.branch[14].block[11].um_I.iw[6] ,
    \top_I.branch[14].block[11].um_I.iw[5] ,
    \top_I.branch[14].block[11].um_I.iw[4] ,
    \top_I.branch[14].block[11].um_I.iw[3] ,
    \top_I.branch[14].block[11].um_I.iw[2] ,
    \top_I.branch[14].block[11].um_I.iw[1] ,
    \top_I.branch[14].block[11].um_I.clk ,
    \top_I.branch[14].block[10].um_I.iw[17] ,
    \top_I.branch[14].block[10].um_I.iw[16] ,
    \top_I.branch[14].block[10].um_I.iw[15] ,
    \top_I.branch[14].block[10].um_I.iw[14] ,
    \top_I.branch[14].block[10].um_I.iw[13] ,
    \top_I.branch[14].block[10].um_I.iw[12] ,
    \top_I.branch[14].block[10].um_I.iw[11] ,
    \top_I.branch[14].block[10].um_I.iw[10] ,
    \top_I.branch[14].block[10].um_I.iw[9] ,
    \top_I.branch[14].block[10].um_I.iw[8] ,
    \top_I.branch[14].block[10].um_I.iw[7] ,
    \top_I.branch[14].block[10].um_I.iw[6] ,
    \top_I.branch[14].block[10].um_I.iw[5] ,
    \top_I.branch[14].block[10].um_I.iw[4] ,
    \top_I.branch[14].block[10].um_I.iw[3] ,
    \top_I.branch[14].block[10].um_I.iw[2] ,
    \top_I.branch[14].block[10].um_I.iw[1] ,
    \top_I.branch[14].block[10].um_I.clk ,
    \top_I.branch[14].block[9].um_I.iw[17] ,
    \top_I.branch[14].block[9].um_I.iw[16] ,
    \top_I.branch[14].block[9].um_I.iw[15] ,
    \top_I.branch[14].block[9].um_I.iw[14] ,
    \top_I.branch[14].block[9].um_I.iw[13] ,
    \top_I.branch[14].block[9].um_I.iw[12] ,
    \top_I.branch[14].block[9].um_I.iw[11] ,
    \top_I.branch[14].block[9].um_I.iw[10] ,
    \top_I.branch[14].block[9].um_I.iw[9] ,
    \top_I.branch[14].block[9].um_I.iw[8] ,
    \top_I.branch[14].block[9].um_I.iw[7] ,
    \top_I.branch[14].block[9].um_I.iw[6] ,
    \top_I.branch[14].block[9].um_I.iw[5] ,
    \top_I.branch[14].block[9].um_I.iw[4] ,
    \top_I.branch[14].block[9].um_I.iw[3] ,
    \top_I.branch[14].block[9].um_I.iw[2] ,
    \top_I.branch[14].block[9].um_I.iw[1] ,
    \top_I.branch[14].block[9].um_I.clk ,
    \top_I.branch[14].block[8].um_I.iw[17] ,
    \top_I.branch[14].block[8].um_I.iw[16] ,
    \top_I.branch[14].block[8].um_I.iw[15] ,
    \top_I.branch[14].block[8].um_I.iw[14] ,
    \top_I.branch[14].block[8].um_I.iw[13] ,
    \top_I.branch[14].block[8].um_I.iw[12] ,
    \top_I.branch[14].block[8].um_I.iw[11] ,
    \top_I.branch[14].block[8].um_I.iw[10] ,
    \top_I.branch[14].block[8].um_I.iw[9] ,
    \top_I.branch[14].block[8].um_I.iw[8] ,
    \top_I.branch[14].block[8].um_I.iw[7] ,
    \top_I.branch[14].block[8].um_I.iw[6] ,
    \top_I.branch[14].block[8].um_I.iw[5] ,
    \top_I.branch[14].block[8].um_I.iw[4] ,
    \top_I.branch[14].block[8].um_I.iw[3] ,
    \top_I.branch[14].block[8].um_I.iw[2] ,
    \top_I.branch[14].block[8].um_I.iw[1] ,
    \top_I.branch[14].block[8].um_I.clk ,
    \top_I.branch[14].block[7].um_I.iw[17] ,
    \top_I.branch[14].block[7].um_I.iw[16] ,
    \top_I.branch[14].block[7].um_I.iw[15] ,
    \top_I.branch[14].block[7].um_I.iw[14] ,
    \top_I.branch[14].block[7].um_I.iw[13] ,
    \top_I.branch[14].block[7].um_I.iw[12] ,
    \top_I.branch[14].block[7].um_I.iw[11] ,
    \top_I.branch[14].block[7].um_I.iw[10] ,
    \top_I.branch[14].block[7].um_I.iw[9] ,
    \top_I.branch[14].block[7].um_I.iw[8] ,
    \top_I.branch[14].block[7].um_I.iw[7] ,
    \top_I.branch[14].block[7].um_I.iw[6] ,
    \top_I.branch[14].block[7].um_I.iw[5] ,
    \top_I.branch[14].block[7].um_I.iw[4] ,
    \top_I.branch[14].block[7].um_I.iw[3] ,
    \top_I.branch[14].block[7].um_I.iw[2] ,
    \top_I.branch[14].block[7].um_I.iw[1] ,
    \top_I.branch[14].block[7].um_I.clk ,
    \top_I.branch[14].block[6].um_I.iw[17] ,
    \top_I.branch[14].block[6].um_I.iw[16] ,
    \top_I.branch[14].block[6].um_I.iw[15] ,
    \top_I.branch[14].block[6].um_I.iw[14] ,
    \top_I.branch[14].block[6].um_I.iw[13] ,
    \top_I.branch[14].block[6].um_I.iw[12] ,
    \top_I.branch[14].block[6].um_I.iw[11] ,
    \top_I.branch[14].block[6].um_I.iw[10] ,
    \top_I.branch[14].block[6].um_I.iw[9] ,
    \top_I.branch[14].block[6].um_I.iw[8] ,
    \top_I.branch[14].block[6].um_I.iw[7] ,
    \top_I.branch[14].block[6].um_I.iw[6] ,
    \top_I.branch[14].block[6].um_I.iw[5] ,
    \top_I.branch[14].block[6].um_I.iw[4] ,
    \top_I.branch[14].block[6].um_I.iw[3] ,
    \top_I.branch[14].block[6].um_I.iw[2] ,
    \top_I.branch[14].block[6].um_I.iw[1] ,
    \top_I.branch[14].block[6].um_I.clk ,
    \top_I.branch[14].block[5].um_I.iw[17] ,
    \top_I.branch[14].block[5].um_I.iw[16] ,
    \top_I.branch[14].block[5].um_I.iw[15] ,
    \top_I.branch[14].block[5].um_I.iw[14] ,
    \top_I.branch[14].block[5].um_I.iw[13] ,
    \top_I.branch[14].block[5].um_I.iw[12] ,
    \top_I.branch[14].block[5].um_I.iw[11] ,
    \top_I.branch[14].block[5].um_I.iw[10] ,
    \top_I.branch[14].block[5].um_I.iw[9] ,
    \top_I.branch[14].block[5].um_I.iw[8] ,
    \top_I.branch[14].block[5].um_I.iw[7] ,
    \top_I.branch[14].block[5].um_I.iw[6] ,
    \top_I.branch[14].block[5].um_I.iw[5] ,
    \top_I.branch[14].block[5].um_I.iw[4] ,
    \top_I.branch[14].block[5].um_I.iw[3] ,
    \top_I.branch[14].block[5].um_I.iw[2] ,
    \top_I.branch[14].block[5].um_I.iw[1] ,
    \top_I.branch[14].block[5].um_I.clk ,
    \top_I.branch[14].block[4].um_I.iw[17] ,
    \top_I.branch[14].block[4].um_I.iw[16] ,
    \top_I.branch[14].block[4].um_I.iw[15] ,
    \top_I.branch[14].block[4].um_I.iw[14] ,
    \top_I.branch[14].block[4].um_I.iw[13] ,
    \top_I.branch[14].block[4].um_I.iw[12] ,
    \top_I.branch[14].block[4].um_I.iw[11] ,
    \top_I.branch[14].block[4].um_I.iw[10] ,
    \top_I.branch[14].block[4].um_I.iw[9] ,
    \top_I.branch[14].block[4].um_I.iw[8] ,
    \top_I.branch[14].block[4].um_I.iw[7] ,
    \top_I.branch[14].block[4].um_I.iw[6] ,
    \top_I.branch[14].block[4].um_I.iw[5] ,
    \top_I.branch[14].block[4].um_I.iw[4] ,
    \top_I.branch[14].block[4].um_I.iw[3] ,
    \top_I.branch[14].block[4].um_I.iw[2] ,
    \top_I.branch[14].block[4].um_I.iw[1] ,
    \top_I.branch[14].block[4].um_I.clk ,
    \top_I.branch[14].block[3].um_I.iw[17] ,
    \top_I.branch[14].block[3].um_I.iw[16] ,
    \top_I.branch[14].block[3].um_I.iw[15] ,
    \top_I.branch[14].block[3].um_I.iw[14] ,
    \top_I.branch[14].block[3].um_I.iw[13] ,
    \top_I.branch[14].block[3].um_I.iw[12] ,
    \top_I.branch[14].block[3].um_I.iw[11] ,
    \top_I.branch[14].block[3].um_I.iw[10] ,
    \top_I.branch[14].block[3].um_I.iw[9] ,
    \top_I.branch[14].block[3].um_I.iw[8] ,
    \top_I.branch[14].block[3].um_I.iw[7] ,
    \top_I.branch[14].block[3].um_I.iw[6] ,
    \top_I.branch[14].block[3].um_I.iw[5] ,
    \top_I.branch[14].block[3].um_I.iw[4] ,
    \top_I.branch[14].block[3].um_I.iw[3] ,
    \top_I.branch[14].block[3].um_I.iw[2] ,
    \top_I.branch[14].block[3].um_I.iw[1] ,
    \top_I.branch[14].block[3].um_I.clk ,
    \top_I.branch[14].block[2].um_I.iw[17] ,
    \top_I.branch[14].block[2].um_I.iw[16] ,
    \top_I.branch[14].block[2].um_I.iw[15] ,
    \top_I.branch[14].block[2].um_I.iw[14] ,
    \top_I.branch[14].block[2].um_I.iw[13] ,
    \top_I.branch[14].block[2].um_I.iw[12] ,
    \top_I.branch[14].block[2].um_I.iw[11] ,
    \top_I.branch[14].block[2].um_I.iw[10] ,
    \top_I.branch[14].block[2].um_I.iw[9] ,
    \top_I.branch[14].block[2].um_I.iw[8] ,
    \top_I.branch[14].block[2].um_I.iw[7] ,
    \top_I.branch[14].block[2].um_I.iw[6] ,
    \top_I.branch[14].block[2].um_I.iw[5] ,
    \top_I.branch[14].block[2].um_I.iw[4] ,
    \top_I.branch[14].block[2].um_I.iw[3] ,
    \top_I.branch[14].block[2].um_I.iw[2] ,
    \top_I.branch[14].block[2].um_I.iw[1] ,
    \top_I.branch[14].block[2].um_I.clk ,
    \top_I.branch[14].block[1].um_I.iw[17] ,
    \top_I.branch[14].block[1].um_I.iw[16] ,
    \top_I.branch[14].block[1].um_I.iw[15] ,
    \top_I.branch[14].block[1].um_I.iw[14] ,
    \top_I.branch[14].block[1].um_I.iw[13] ,
    \top_I.branch[14].block[1].um_I.iw[12] ,
    \top_I.branch[14].block[1].um_I.iw[11] ,
    \top_I.branch[14].block[1].um_I.iw[10] ,
    \top_I.branch[14].block[1].um_I.iw[9] ,
    \top_I.branch[14].block[1].um_I.iw[8] ,
    \top_I.branch[14].block[1].um_I.iw[7] ,
    \top_I.branch[14].block[1].um_I.iw[6] ,
    \top_I.branch[14].block[1].um_I.iw[5] ,
    \top_I.branch[14].block[1].um_I.iw[4] ,
    \top_I.branch[14].block[1].um_I.iw[3] ,
    \top_I.branch[14].block[1].um_I.iw[2] ,
    \top_I.branch[14].block[1].um_I.iw[1] ,
    \top_I.branch[14].block[1].um_I.clk ,
    \top_I.branch[14].block[0].um_I.iw[17] ,
    \top_I.branch[14].block[0].um_I.iw[16] ,
    \top_I.branch[14].block[0].um_I.iw[15] ,
    \top_I.branch[14].block[0].um_I.iw[14] ,
    \top_I.branch[14].block[0].um_I.iw[13] ,
    \top_I.branch[14].block[0].um_I.iw[12] ,
    \top_I.branch[14].block[0].um_I.iw[11] ,
    \top_I.branch[14].block[0].um_I.iw[10] ,
    \top_I.branch[14].block[0].um_I.iw[9] ,
    \top_I.branch[14].block[0].um_I.iw[8] ,
    \top_I.branch[14].block[0].um_I.iw[7] ,
    \top_I.branch[14].block[0].um_I.iw[6] ,
    \top_I.branch[14].block[0].um_I.iw[5] ,
    \top_I.branch[14].block[0].um_I.iw[4] ,
    \top_I.branch[14].block[0].um_I.iw[3] ,
    \top_I.branch[14].block[0].um_I.iw[2] ,
    \top_I.branch[14].block[0].um_I.iw[1] ,
    \top_I.branch[14].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[15].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[14].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[13].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[12].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[11].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[10].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[9].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[8].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[7].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[6].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[5].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[4].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[3].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[2].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[1].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero ,
    \top_I.branch[14].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[14].block[15].um_I.pg_vdd ,
    \top_I.branch[14].block[14].um_I.pg_vdd ,
    \top_I.branch[14].block[13].um_I.pg_vdd ,
    \top_I.branch[14].block[12].um_I.pg_vdd ,
    \top_I.branch[14].block[11].um_I.pg_vdd ,
    \top_I.branch[14].block[10].um_I.pg_vdd ,
    \top_I.branch[14].block[9].um_I.pg_vdd ,
    \top_I.branch[14].block[8].um_I.pg_vdd ,
    \top_I.branch[14].block[7].um_I.pg_vdd ,
    \top_I.branch[14].block[6].um_I.pg_vdd ,
    \top_I.branch[14].block[5].um_I.pg_vdd ,
    \top_I.branch[14].block[4].um_I.pg_vdd ,
    \top_I.branch[14].block[3].um_I.pg_vdd ,
    \top_I.branch[14].block[2].um_I.pg_vdd ,
    \top_I.branch[14].block[1].um_I.pg_vdd ,
    \top_I.branch[14].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[15].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[15].l_addr[0] ),
    .k_zero(\top_I.branch[15].l_addr[3] ),
    .addr({\top_I.branch[15].l_addr[3] ,
    \top_I.branch[15].l_addr[0] ,
    \top_I.branch[15].l_addr[0] ,
    \top_I.branch[15].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[15].block[15].um_I.ena ,
    \top_I.branch[15].block[14].um_I.ena ,
    \top_I.branch[15].block[13].um_I.ena ,
    \top_I.branch[15].block[12].um_I.ena ,
    \top_I.branch[15].block[11].um_I.ena ,
    \top_I.branch[15].block[10].um_I.ena ,
    \top_I.branch[15].block[9].um_I.ena ,
    \top_I.branch[15].block[8].um_I.ena ,
    \top_I.branch[15].block[7].um_I.ena ,
    \top_I.branch[15].block[6].um_I.ena ,
    \top_I.branch[15].block[5].um_I.ena ,
    \top_I.branch[15].block[4].um_I.ena ,
    \top_I.branch[15].block[3].um_I.ena ,
    \top_I.branch[15].block[2].um_I.ena ,
    \top_I.branch[15].block[1].um_I.ena ,
    \top_I.branch[15].block[0].um_I.ena }),
    .um_iw({\top_I.branch[15].block[15].um_I.iw[17] ,
    \top_I.branch[15].block[15].um_I.iw[16] ,
    \top_I.branch[15].block[15].um_I.iw[15] ,
    \top_I.branch[15].block[15].um_I.iw[14] ,
    \top_I.branch[15].block[15].um_I.iw[13] ,
    \top_I.branch[15].block[15].um_I.iw[12] ,
    \top_I.branch[15].block[15].um_I.iw[11] ,
    \top_I.branch[15].block[15].um_I.iw[10] ,
    \top_I.branch[15].block[15].um_I.iw[9] ,
    \top_I.branch[15].block[15].um_I.iw[8] ,
    \top_I.branch[15].block[15].um_I.iw[7] ,
    \top_I.branch[15].block[15].um_I.iw[6] ,
    \top_I.branch[15].block[15].um_I.iw[5] ,
    \top_I.branch[15].block[15].um_I.iw[4] ,
    \top_I.branch[15].block[15].um_I.iw[3] ,
    \top_I.branch[15].block[15].um_I.iw[2] ,
    \top_I.branch[15].block[15].um_I.iw[1] ,
    \top_I.branch[15].block[15].um_I.clk ,
    \top_I.branch[15].block[14].um_I.iw[17] ,
    \top_I.branch[15].block[14].um_I.iw[16] ,
    \top_I.branch[15].block[14].um_I.iw[15] ,
    \top_I.branch[15].block[14].um_I.iw[14] ,
    \top_I.branch[15].block[14].um_I.iw[13] ,
    \top_I.branch[15].block[14].um_I.iw[12] ,
    \top_I.branch[15].block[14].um_I.iw[11] ,
    \top_I.branch[15].block[14].um_I.iw[10] ,
    \top_I.branch[15].block[14].um_I.iw[9] ,
    \top_I.branch[15].block[14].um_I.iw[8] ,
    \top_I.branch[15].block[14].um_I.iw[7] ,
    \top_I.branch[15].block[14].um_I.iw[6] ,
    \top_I.branch[15].block[14].um_I.iw[5] ,
    \top_I.branch[15].block[14].um_I.iw[4] ,
    \top_I.branch[15].block[14].um_I.iw[3] ,
    \top_I.branch[15].block[14].um_I.iw[2] ,
    \top_I.branch[15].block[14].um_I.iw[1] ,
    \top_I.branch[15].block[14].um_I.clk ,
    \top_I.branch[15].block[13].um_I.iw[17] ,
    \top_I.branch[15].block[13].um_I.iw[16] ,
    \top_I.branch[15].block[13].um_I.iw[15] ,
    \top_I.branch[15].block[13].um_I.iw[14] ,
    \top_I.branch[15].block[13].um_I.iw[13] ,
    \top_I.branch[15].block[13].um_I.iw[12] ,
    \top_I.branch[15].block[13].um_I.iw[11] ,
    \top_I.branch[15].block[13].um_I.iw[10] ,
    \top_I.branch[15].block[13].um_I.iw[9] ,
    \top_I.branch[15].block[13].um_I.iw[8] ,
    \top_I.branch[15].block[13].um_I.iw[7] ,
    \top_I.branch[15].block[13].um_I.iw[6] ,
    \top_I.branch[15].block[13].um_I.iw[5] ,
    \top_I.branch[15].block[13].um_I.iw[4] ,
    \top_I.branch[15].block[13].um_I.iw[3] ,
    \top_I.branch[15].block[13].um_I.iw[2] ,
    \top_I.branch[15].block[13].um_I.iw[1] ,
    \top_I.branch[15].block[13].um_I.clk ,
    \top_I.branch[15].block[12].um_I.iw[17] ,
    \top_I.branch[15].block[12].um_I.iw[16] ,
    \top_I.branch[15].block[12].um_I.iw[15] ,
    \top_I.branch[15].block[12].um_I.iw[14] ,
    \top_I.branch[15].block[12].um_I.iw[13] ,
    \top_I.branch[15].block[12].um_I.iw[12] ,
    \top_I.branch[15].block[12].um_I.iw[11] ,
    \top_I.branch[15].block[12].um_I.iw[10] ,
    \top_I.branch[15].block[12].um_I.iw[9] ,
    \top_I.branch[15].block[12].um_I.iw[8] ,
    \top_I.branch[15].block[12].um_I.iw[7] ,
    \top_I.branch[15].block[12].um_I.iw[6] ,
    \top_I.branch[15].block[12].um_I.iw[5] ,
    \top_I.branch[15].block[12].um_I.iw[4] ,
    \top_I.branch[15].block[12].um_I.iw[3] ,
    \top_I.branch[15].block[12].um_I.iw[2] ,
    \top_I.branch[15].block[12].um_I.iw[1] ,
    \top_I.branch[15].block[12].um_I.clk ,
    \top_I.branch[15].block[11].um_I.iw[17] ,
    \top_I.branch[15].block[11].um_I.iw[16] ,
    \top_I.branch[15].block[11].um_I.iw[15] ,
    \top_I.branch[15].block[11].um_I.iw[14] ,
    \top_I.branch[15].block[11].um_I.iw[13] ,
    \top_I.branch[15].block[11].um_I.iw[12] ,
    \top_I.branch[15].block[11].um_I.iw[11] ,
    \top_I.branch[15].block[11].um_I.iw[10] ,
    \top_I.branch[15].block[11].um_I.iw[9] ,
    \top_I.branch[15].block[11].um_I.iw[8] ,
    \top_I.branch[15].block[11].um_I.iw[7] ,
    \top_I.branch[15].block[11].um_I.iw[6] ,
    \top_I.branch[15].block[11].um_I.iw[5] ,
    \top_I.branch[15].block[11].um_I.iw[4] ,
    \top_I.branch[15].block[11].um_I.iw[3] ,
    \top_I.branch[15].block[11].um_I.iw[2] ,
    \top_I.branch[15].block[11].um_I.iw[1] ,
    \top_I.branch[15].block[11].um_I.clk ,
    \top_I.branch[15].block[10].um_I.iw[17] ,
    \top_I.branch[15].block[10].um_I.iw[16] ,
    \top_I.branch[15].block[10].um_I.iw[15] ,
    \top_I.branch[15].block[10].um_I.iw[14] ,
    \top_I.branch[15].block[10].um_I.iw[13] ,
    \top_I.branch[15].block[10].um_I.iw[12] ,
    \top_I.branch[15].block[10].um_I.iw[11] ,
    \top_I.branch[15].block[10].um_I.iw[10] ,
    \top_I.branch[15].block[10].um_I.iw[9] ,
    \top_I.branch[15].block[10].um_I.iw[8] ,
    \top_I.branch[15].block[10].um_I.iw[7] ,
    \top_I.branch[15].block[10].um_I.iw[6] ,
    \top_I.branch[15].block[10].um_I.iw[5] ,
    \top_I.branch[15].block[10].um_I.iw[4] ,
    \top_I.branch[15].block[10].um_I.iw[3] ,
    \top_I.branch[15].block[10].um_I.iw[2] ,
    \top_I.branch[15].block[10].um_I.iw[1] ,
    \top_I.branch[15].block[10].um_I.clk ,
    \top_I.branch[15].block[9].um_I.iw[17] ,
    \top_I.branch[15].block[9].um_I.iw[16] ,
    \top_I.branch[15].block[9].um_I.iw[15] ,
    \top_I.branch[15].block[9].um_I.iw[14] ,
    \top_I.branch[15].block[9].um_I.iw[13] ,
    \top_I.branch[15].block[9].um_I.iw[12] ,
    \top_I.branch[15].block[9].um_I.iw[11] ,
    \top_I.branch[15].block[9].um_I.iw[10] ,
    \top_I.branch[15].block[9].um_I.iw[9] ,
    \top_I.branch[15].block[9].um_I.iw[8] ,
    \top_I.branch[15].block[9].um_I.iw[7] ,
    \top_I.branch[15].block[9].um_I.iw[6] ,
    \top_I.branch[15].block[9].um_I.iw[5] ,
    \top_I.branch[15].block[9].um_I.iw[4] ,
    \top_I.branch[15].block[9].um_I.iw[3] ,
    \top_I.branch[15].block[9].um_I.iw[2] ,
    \top_I.branch[15].block[9].um_I.iw[1] ,
    \top_I.branch[15].block[9].um_I.clk ,
    \top_I.branch[15].block[8].um_I.iw[17] ,
    \top_I.branch[15].block[8].um_I.iw[16] ,
    \top_I.branch[15].block[8].um_I.iw[15] ,
    \top_I.branch[15].block[8].um_I.iw[14] ,
    \top_I.branch[15].block[8].um_I.iw[13] ,
    \top_I.branch[15].block[8].um_I.iw[12] ,
    \top_I.branch[15].block[8].um_I.iw[11] ,
    \top_I.branch[15].block[8].um_I.iw[10] ,
    \top_I.branch[15].block[8].um_I.iw[9] ,
    \top_I.branch[15].block[8].um_I.iw[8] ,
    \top_I.branch[15].block[8].um_I.iw[7] ,
    \top_I.branch[15].block[8].um_I.iw[6] ,
    \top_I.branch[15].block[8].um_I.iw[5] ,
    \top_I.branch[15].block[8].um_I.iw[4] ,
    \top_I.branch[15].block[8].um_I.iw[3] ,
    \top_I.branch[15].block[8].um_I.iw[2] ,
    \top_I.branch[15].block[8].um_I.iw[1] ,
    \top_I.branch[15].block[8].um_I.clk ,
    \top_I.branch[15].block[7].um_I.iw[17] ,
    \top_I.branch[15].block[7].um_I.iw[16] ,
    \top_I.branch[15].block[7].um_I.iw[15] ,
    \top_I.branch[15].block[7].um_I.iw[14] ,
    \top_I.branch[15].block[7].um_I.iw[13] ,
    \top_I.branch[15].block[7].um_I.iw[12] ,
    \top_I.branch[15].block[7].um_I.iw[11] ,
    \top_I.branch[15].block[7].um_I.iw[10] ,
    \top_I.branch[15].block[7].um_I.iw[9] ,
    \top_I.branch[15].block[7].um_I.iw[8] ,
    \top_I.branch[15].block[7].um_I.iw[7] ,
    \top_I.branch[15].block[7].um_I.iw[6] ,
    \top_I.branch[15].block[7].um_I.iw[5] ,
    \top_I.branch[15].block[7].um_I.iw[4] ,
    \top_I.branch[15].block[7].um_I.iw[3] ,
    \top_I.branch[15].block[7].um_I.iw[2] ,
    \top_I.branch[15].block[7].um_I.iw[1] ,
    \top_I.branch[15].block[7].um_I.clk ,
    \top_I.branch[15].block[6].um_I.iw[17] ,
    \top_I.branch[15].block[6].um_I.iw[16] ,
    \top_I.branch[15].block[6].um_I.iw[15] ,
    \top_I.branch[15].block[6].um_I.iw[14] ,
    \top_I.branch[15].block[6].um_I.iw[13] ,
    \top_I.branch[15].block[6].um_I.iw[12] ,
    \top_I.branch[15].block[6].um_I.iw[11] ,
    \top_I.branch[15].block[6].um_I.iw[10] ,
    \top_I.branch[15].block[6].um_I.iw[9] ,
    \top_I.branch[15].block[6].um_I.iw[8] ,
    \top_I.branch[15].block[6].um_I.iw[7] ,
    \top_I.branch[15].block[6].um_I.iw[6] ,
    \top_I.branch[15].block[6].um_I.iw[5] ,
    \top_I.branch[15].block[6].um_I.iw[4] ,
    \top_I.branch[15].block[6].um_I.iw[3] ,
    \top_I.branch[15].block[6].um_I.iw[2] ,
    \top_I.branch[15].block[6].um_I.iw[1] ,
    \top_I.branch[15].block[6].um_I.clk ,
    \top_I.branch[15].block[5].um_I.iw[17] ,
    \top_I.branch[15].block[5].um_I.iw[16] ,
    \top_I.branch[15].block[5].um_I.iw[15] ,
    \top_I.branch[15].block[5].um_I.iw[14] ,
    \top_I.branch[15].block[5].um_I.iw[13] ,
    \top_I.branch[15].block[5].um_I.iw[12] ,
    \top_I.branch[15].block[5].um_I.iw[11] ,
    \top_I.branch[15].block[5].um_I.iw[10] ,
    \top_I.branch[15].block[5].um_I.iw[9] ,
    \top_I.branch[15].block[5].um_I.iw[8] ,
    \top_I.branch[15].block[5].um_I.iw[7] ,
    \top_I.branch[15].block[5].um_I.iw[6] ,
    \top_I.branch[15].block[5].um_I.iw[5] ,
    \top_I.branch[15].block[5].um_I.iw[4] ,
    \top_I.branch[15].block[5].um_I.iw[3] ,
    \top_I.branch[15].block[5].um_I.iw[2] ,
    \top_I.branch[15].block[5].um_I.iw[1] ,
    \top_I.branch[15].block[5].um_I.clk ,
    \top_I.branch[15].block[4].um_I.iw[17] ,
    \top_I.branch[15].block[4].um_I.iw[16] ,
    \top_I.branch[15].block[4].um_I.iw[15] ,
    \top_I.branch[15].block[4].um_I.iw[14] ,
    \top_I.branch[15].block[4].um_I.iw[13] ,
    \top_I.branch[15].block[4].um_I.iw[12] ,
    \top_I.branch[15].block[4].um_I.iw[11] ,
    \top_I.branch[15].block[4].um_I.iw[10] ,
    \top_I.branch[15].block[4].um_I.iw[9] ,
    \top_I.branch[15].block[4].um_I.iw[8] ,
    \top_I.branch[15].block[4].um_I.iw[7] ,
    \top_I.branch[15].block[4].um_I.iw[6] ,
    \top_I.branch[15].block[4].um_I.iw[5] ,
    \top_I.branch[15].block[4].um_I.iw[4] ,
    \top_I.branch[15].block[4].um_I.iw[3] ,
    \top_I.branch[15].block[4].um_I.iw[2] ,
    \top_I.branch[15].block[4].um_I.iw[1] ,
    \top_I.branch[15].block[4].um_I.clk ,
    \top_I.branch[15].block[3].um_I.iw[17] ,
    \top_I.branch[15].block[3].um_I.iw[16] ,
    \top_I.branch[15].block[3].um_I.iw[15] ,
    \top_I.branch[15].block[3].um_I.iw[14] ,
    \top_I.branch[15].block[3].um_I.iw[13] ,
    \top_I.branch[15].block[3].um_I.iw[12] ,
    \top_I.branch[15].block[3].um_I.iw[11] ,
    \top_I.branch[15].block[3].um_I.iw[10] ,
    \top_I.branch[15].block[3].um_I.iw[9] ,
    \top_I.branch[15].block[3].um_I.iw[8] ,
    \top_I.branch[15].block[3].um_I.iw[7] ,
    \top_I.branch[15].block[3].um_I.iw[6] ,
    \top_I.branch[15].block[3].um_I.iw[5] ,
    \top_I.branch[15].block[3].um_I.iw[4] ,
    \top_I.branch[15].block[3].um_I.iw[3] ,
    \top_I.branch[15].block[3].um_I.iw[2] ,
    \top_I.branch[15].block[3].um_I.iw[1] ,
    \top_I.branch[15].block[3].um_I.clk ,
    \top_I.branch[15].block[2].um_I.iw[17] ,
    \top_I.branch[15].block[2].um_I.iw[16] ,
    \top_I.branch[15].block[2].um_I.iw[15] ,
    \top_I.branch[15].block[2].um_I.iw[14] ,
    \top_I.branch[15].block[2].um_I.iw[13] ,
    \top_I.branch[15].block[2].um_I.iw[12] ,
    \top_I.branch[15].block[2].um_I.iw[11] ,
    \top_I.branch[15].block[2].um_I.iw[10] ,
    \top_I.branch[15].block[2].um_I.iw[9] ,
    \top_I.branch[15].block[2].um_I.iw[8] ,
    \top_I.branch[15].block[2].um_I.iw[7] ,
    \top_I.branch[15].block[2].um_I.iw[6] ,
    \top_I.branch[15].block[2].um_I.iw[5] ,
    \top_I.branch[15].block[2].um_I.iw[4] ,
    \top_I.branch[15].block[2].um_I.iw[3] ,
    \top_I.branch[15].block[2].um_I.iw[2] ,
    \top_I.branch[15].block[2].um_I.iw[1] ,
    \top_I.branch[15].block[2].um_I.clk ,
    \top_I.branch[15].block[1].um_I.iw[17] ,
    \top_I.branch[15].block[1].um_I.iw[16] ,
    \top_I.branch[15].block[1].um_I.iw[15] ,
    \top_I.branch[15].block[1].um_I.iw[14] ,
    \top_I.branch[15].block[1].um_I.iw[13] ,
    \top_I.branch[15].block[1].um_I.iw[12] ,
    \top_I.branch[15].block[1].um_I.iw[11] ,
    \top_I.branch[15].block[1].um_I.iw[10] ,
    \top_I.branch[15].block[1].um_I.iw[9] ,
    \top_I.branch[15].block[1].um_I.iw[8] ,
    \top_I.branch[15].block[1].um_I.iw[7] ,
    \top_I.branch[15].block[1].um_I.iw[6] ,
    \top_I.branch[15].block[1].um_I.iw[5] ,
    \top_I.branch[15].block[1].um_I.iw[4] ,
    \top_I.branch[15].block[1].um_I.iw[3] ,
    \top_I.branch[15].block[1].um_I.iw[2] ,
    \top_I.branch[15].block[1].um_I.iw[1] ,
    \top_I.branch[15].block[1].um_I.clk ,
    \top_I.branch[15].block[0].um_I.iw[17] ,
    \top_I.branch[15].block[0].um_I.iw[16] ,
    \top_I.branch[15].block[0].um_I.iw[15] ,
    \top_I.branch[15].block[0].um_I.iw[14] ,
    \top_I.branch[15].block[0].um_I.iw[13] ,
    \top_I.branch[15].block[0].um_I.iw[12] ,
    \top_I.branch[15].block[0].um_I.iw[11] ,
    \top_I.branch[15].block[0].um_I.iw[10] ,
    \top_I.branch[15].block[0].um_I.iw[9] ,
    \top_I.branch[15].block[0].um_I.iw[8] ,
    \top_I.branch[15].block[0].um_I.iw[7] ,
    \top_I.branch[15].block[0].um_I.iw[6] ,
    \top_I.branch[15].block[0].um_I.iw[5] ,
    \top_I.branch[15].block[0].um_I.iw[4] ,
    \top_I.branch[15].block[0].um_I.iw[3] ,
    \top_I.branch[15].block[0].um_I.iw[2] ,
    \top_I.branch[15].block[0].um_I.iw[1] ,
    \top_I.branch[15].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[15].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[14].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[13].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[12].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[11].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[10].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[9].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[8].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[7].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[6].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[5].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[4].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[3].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[2].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[1].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero ,
    \top_I.branch[15].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[15].block[15].um_I.pg_vdd ,
    \top_I.branch[15].block[14].um_I.pg_vdd ,
    \top_I.branch[15].block[13].um_I.pg_vdd ,
    \top_I.branch[15].block[12].um_I.pg_vdd ,
    \top_I.branch[15].block[11].um_I.pg_vdd ,
    \top_I.branch[15].block[10].um_I.pg_vdd ,
    \top_I.branch[15].block[9].um_I.pg_vdd ,
    \top_I.branch[15].block[8].um_I.pg_vdd ,
    \top_I.branch[15].block[7].um_I.pg_vdd ,
    \top_I.branch[15].block[6].um_I.pg_vdd ,
    \top_I.branch[15].block[5].um_I.pg_vdd ,
    \top_I.branch[15].block[4].um_I.pg_vdd ,
    \top_I.branch[15].block[3].um_I.pg_vdd ,
    \top_I.branch[15].block[2].um_I.pg_vdd ,
    \top_I.branch[15].block[1].um_I.pg_vdd ,
    \top_I.branch[15].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[16].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[16].l_addr[3] ),
    .k_zero(\top_I.branch[16].l_addr[0] ),
    .addr({\top_I.branch[16].l_addr[3] ,
    \top_I.branch[16].l_addr[0] ,
    \top_I.branch[16].l_addr[0] ,
    \top_I.branch[16].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[16].block[15].um_I.ena ,
    \top_I.branch[16].block[14].um_I.ena ,
    \top_I.branch[16].block[13].um_I.ena ,
    \top_I.branch[16].block[12].um_I.ena ,
    \top_I.branch[16].block[11].um_I.ena ,
    \top_I.branch[16].block[10].um_I.ena ,
    \top_I.branch[16].block[9].um_I.ena ,
    \top_I.branch[16].block[8].um_I.ena ,
    \top_I.branch[16].block[7].um_I.ena ,
    \top_I.branch[16].block[6].um_I.ena ,
    \top_I.branch[16].block[5].um_I.ena ,
    \top_I.branch[16].block[4].um_I.ena ,
    \top_I.branch[16].block[3].um_I.ena ,
    \top_I.branch[16].block[2].um_I.ena ,
    \top_I.branch[16].block[1].um_I.ena ,
    \top_I.branch[16].block[0].um_I.ena }),
    .um_iw({\top_I.branch[16].block[15].um_I.iw[17] ,
    \top_I.branch[16].block[15].um_I.iw[16] ,
    \top_I.branch[16].block[15].um_I.iw[15] ,
    \top_I.branch[16].block[15].um_I.iw[14] ,
    \top_I.branch[16].block[15].um_I.iw[13] ,
    \top_I.branch[16].block[15].um_I.iw[12] ,
    \top_I.branch[16].block[15].um_I.iw[11] ,
    \top_I.branch[16].block[15].um_I.iw[10] ,
    \top_I.branch[16].block[15].um_I.iw[9] ,
    \top_I.branch[16].block[15].um_I.iw[8] ,
    \top_I.branch[16].block[15].um_I.iw[7] ,
    \top_I.branch[16].block[15].um_I.iw[6] ,
    \top_I.branch[16].block[15].um_I.iw[5] ,
    \top_I.branch[16].block[15].um_I.iw[4] ,
    \top_I.branch[16].block[15].um_I.iw[3] ,
    \top_I.branch[16].block[15].um_I.iw[2] ,
    \top_I.branch[16].block[15].um_I.iw[1] ,
    \top_I.branch[16].block[15].um_I.clk ,
    \top_I.branch[16].block[14].um_I.iw[17] ,
    \top_I.branch[16].block[14].um_I.iw[16] ,
    \top_I.branch[16].block[14].um_I.iw[15] ,
    \top_I.branch[16].block[14].um_I.iw[14] ,
    \top_I.branch[16].block[14].um_I.iw[13] ,
    \top_I.branch[16].block[14].um_I.iw[12] ,
    \top_I.branch[16].block[14].um_I.iw[11] ,
    \top_I.branch[16].block[14].um_I.iw[10] ,
    \top_I.branch[16].block[14].um_I.iw[9] ,
    \top_I.branch[16].block[14].um_I.iw[8] ,
    \top_I.branch[16].block[14].um_I.iw[7] ,
    \top_I.branch[16].block[14].um_I.iw[6] ,
    \top_I.branch[16].block[14].um_I.iw[5] ,
    \top_I.branch[16].block[14].um_I.iw[4] ,
    \top_I.branch[16].block[14].um_I.iw[3] ,
    \top_I.branch[16].block[14].um_I.iw[2] ,
    \top_I.branch[16].block[14].um_I.iw[1] ,
    \top_I.branch[16].block[14].um_I.clk ,
    \top_I.branch[16].block[13].um_I.iw[17] ,
    \top_I.branch[16].block[13].um_I.iw[16] ,
    \top_I.branch[16].block[13].um_I.iw[15] ,
    \top_I.branch[16].block[13].um_I.iw[14] ,
    \top_I.branch[16].block[13].um_I.iw[13] ,
    \top_I.branch[16].block[13].um_I.iw[12] ,
    \top_I.branch[16].block[13].um_I.iw[11] ,
    \top_I.branch[16].block[13].um_I.iw[10] ,
    \top_I.branch[16].block[13].um_I.iw[9] ,
    \top_I.branch[16].block[13].um_I.iw[8] ,
    \top_I.branch[16].block[13].um_I.iw[7] ,
    \top_I.branch[16].block[13].um_I.iw[6] ,
    \top_I.branch[16].block[13].um_I.iw[5] ,
    \top_I.branch[16].block[13].um_I.iw[4] ,
    \top_I.branch[16].block[13].um_I.iw[3] ,
    \top_I.branch[16].block[13].um_I.iw[2] ,
    \top_I.branch[16].block[13].um_I.iw[1] ,
    \top_I.branch[16].block[13].um_I.clk ,
    \top_I.branch[16].block[12].um_I.iw[17] ,
    \top_I.branch[16].block[12].um_I.iw[16] ,
    \top_I.branch[16].block[12].um_I.iw[15] ,
    \top_I.branch[16].block[12].um_I.iw[14] ,
    \top_I.branch[16].block[12].um_I.iw[13] ,
    \top_I.branch[16].block[12].um_I.iw[12] ,
    \top_I.branch[16].block[12].um_I.iw[11] ,
    \top_I.branch[16].block[12].um_I.iw[10] ,
    \top_I.branch[16].block[12].um_I.iw[9] ,
    \top_I.branch[16].block[12].um_I.iw[8] ,
    \top_I.branch[16].block[12].um_I.iw[7] ,
    \top_I.branch[16].block[12].um_I.iw[6] ,
    \top_I.branch[16].block[12].um_I.iw[5] ,
    \top_I.branch[16].block[12].um_I.iw[4] ,
    \top_I.branch[16].block[12].um_I.iw[3] ,
    \top_I.branch[16].block[12].um_I.iw[2] ,
    \top_I.branch[16].block[12].um_I.iw[1] ,
    \top_I.branch[16].block[12].um_I.clk ,
    \top_I.branch[16].block[11].um_I.iw[17] ,
    \top_I.branch[16].block[11].um_I.iw[16] ,
    \top_I.branch[16].block[11].um_I.iw[15] ,
    \top_I.branch[16].block[11].um_I.iw[14] ,
    \top_I.branch[16].block[11].um_I.iw[13] ,
    \top_I.branch[16].block[11].um_I.iw[12] ,
    \top_I.branch[16].block[11].um_I.iw[11] ,
    \top_I.branch[16].block[11].um_I.iw[10] ,
    \top_I.branch[16].block[11].um_I.iw[9] ,
    \top_I.branch[16].block[11].um_I.iw[8] ,
    \top_I.branch[16].block[11].um_I.iw[7] ,
    \top_I.branch[16].block[11].um_I.iw[6] ,
    \top_I.branch[16].block[11].um_I.iw[5] ,
    \top_I.branch[16].block[11].um_I.iw[4] ,
    \top_I.branch[16].block[11].um_I.iw[3] ,
    \top_I.branch[16].block[11].um_I.iw[2] ,
    \top_I.branch[16].block[11].um_I.iw[1] ,
    \top_I.branch[16].block[11].um_I.clk ,
    \top_I.branch[16].block[10].um_I.iw[17] ,
    \top_I.branch[16].block[10].um_I.iw[16] ,
    \top_I.branch[16].block[10].um_I.iw[15] ,
    \top_I.branch[16].block[10].um_I.iw[14] ,
    \top_I.branch[16].block[10].um_I.iw[13] ,
    \top_I.branch[16].block[10].um_I.iw[12] ,
    \top_I.branch[16].block[10].um_I.iw[11] ,
    \top_I.branch[16].block[10].um_I.iw[10] ,
    \top_I.branch[16].block[10].um_I.iw[9] ,
    \top_I.branch[16].block[10].um_I.iw[8] ,
    \top_I.branch[16].block[10].um_I.iw[7] ,
    \top_I.branch[16].block[10].um_I.iw[6] ,
    \top_I.branch[16].block[10].um_I.iw[5] ,
    \top_I.branch[16].block[10].um_I.iw[4] ,
    \top_I.branch[16].block[10].um_I.iw[3] ,
    \top_I.branch[16].block[10].um_I.iw[2] ,
    \top_I.branch[16].block[10].um_I.iw[1] ,
    \top_I.branch[16].block[10].um_I.clk ,
    \top_I.branch[16].block[9].um_I.iw[17] ,
    \top_I.branch[16].block[9].um_I.iw[16] ,
    \top_I.branch[16].block[9].um_I.iw[15] ,
    \top_I.branch[16].block[9].um_I.iw[14] ,
    \top_I.branch[16].block[9].um_I.iw[13] ,
    \top_I.branch[16].block[9].um_I.iw[12] ,
    \top_I.branch[16].block[9].um_I.iw[11] ,
    \top_I.branch[16].block[9].um_I.iw[10] ,
    \top_I.branch[16].block[9].um_I.iw[9] ,
    \top_I.branch[16].block[9].um_I.iw[8] ,
    \top_I.branch[16].block[9].um_I.iw[7] ,
    \top_I.branch[16].block[9].um_I.iw[6] ,
    \top_I.branch[16].block[9].um_I.iw[5] ,
    \top_I.branch[16].block[9].um_I.iw[4] ,
    \top_I.branch[16].block[9].um_I.iw[3] ,
    \top_I.branch[16].block[9].um_I.iw[2] ,
    \top_I.branch[16].block[9].um_I.iw[1] ,
    \top_I.branch[16].block[9].um_I.clk ,
    \top_I.branch[16].block[8].um_I.iw[17] ,
    \top_I.branch[16].block[8].um_I.iw[16] ,
    \top_I.branch[16].block[8].um_I.iw[15] ,
    \top_I.branch[16].block[8].um_I.iw[14] ,
    \top_I.branch[16].block[8].um_I.iw[13] ,
    \top_I.branch[16].block[8].um_I.iw[12] ,
    \top_I.branch[16].block[8].um_I.iw[11] ,
    \top_I.branch[16].block[8].um_I.iw[10] ,
    \top_I.branch[16].block[8].um_I.iw[9] ,
    \top_I.branch[16].block[8].um_I.iw[8] ,
    \top_I.branch[16].block[8].um_I.iw[7] ,
    \top_I.branch[16].block[8].um_I.iw[6] ,
    \top_I.branch[16].block[8].um_I.iw[5] ,
    \top_I.branch[16].block[8].um_I.iw[4] ,
    \top_I.branch[16].block[8].um_I.iw[3] ,
    \top_I.branch[16].block[8].um_I.iw[2] ,
    \top_I.branch[16].block[8].um_I.iw[1] ,
    \top_I.branch[16].block[8].um_I.clk ,
    \top_I.branch[16].block[7].um_I.iw[17] ,
    \top_I.branch[16].block[7].um_I.iw[16] ,
    \top_I.branch[16].block[7].um_I.iw[15] ,
    \top_I.branch[16].block[7].um_I.iw[14] ,
    \top_I.branch[16].block[7].um_I.iw[13] ,
    \top_I.branch[16].block[7].um_I.iw[12] ,
    \top_I.branch[16].block[7].um_I.iw[11] ,
    \top_I.branch[16].block[7].um_I.iw[10] ,
    \top_I.branch[16].block[7].um_I.iw[9] ,
    \top_I.branch[16].block[7].um_I.iw[8] ,
    \top_I.branch[16].block[7].um_I.iw[7] ,
    \top_I.branch[16].block[7].um_I.iw[6] ,
    \top_I.branch[16].block[7].um_I.iw[5] ,
    \top_I.branch[16].block[7].um_I.iw[4] ,
    \top_I.branch[16].block[7].um_I.iw[3] ,
    \top_I.branch[16].block[7].um_I.iw[2] ,
    \top_I.branch[16].block[7].um_I.iw[1] ,
    \top_I.branch[16].block[7].um_I.clk ,
    \top_I.branch[16].block[6].um_I.iw[17] ,
    \top_I.branch[16].block[6].um_I.iw[16] ,
    \top_I.branch[16].block[6].um_I.iw[15] ,
    \top_I.branch[16].block[6].um_I.iw[14] ,
    \top_I.branch[16].block[6].um_I.iw[13] ,
    \top_I.branch[16].block[6].um_I.iw[12] ,
    \top_I.branch[16].block[6].um_I.iw[11] ,
    \top_I.branch[16].block[6].um_I.iw[10] ,
    \top_I.branch[16].block[6].um_I.iw[9] ,
    \top_I.branch[16].block[6].um_I.iw[8] ,
    \top_I.branch[16].block[6].um_I.iw[7] ,
    \top_I.branch[16].block[6].um_I.iw[6] ,
    \top_I.branch[16].block[6].um_I.iw[5] ,
    \top_I.branch[16].block[6].um_I.iw[4] ,
    \top_I.branch[16].block[6].um_I.iw[3] ,
    \top_I.branch[16].block[6].um_I.iw[2] ,
    \top_I.branch[16].block[6].um_I.iw[1] ,
    \top_I.branch[16].block[6].um_I.clk ,
    \top_I.branch[16].block[5].um_I.iw[17] ,
    \top_I.branch[16].block[5].um_I.iw[16] ,
    \top_I.branch[16].block[5].um_I.iw[15] ,
    \top_I.branch[16].block[5].um_I.iw[14] ,
    \top_I.branch[16].block[5].um_I.iw[13] ,
    \top_I.branch[16].block[5].um_I.iw[12] ,
    \top_I.branch[16].block[5].um_I.iw[11] ,
    \top_I.branch[16].block[5].um_I.iw[10] ,
    \top_I.branch[16].block[5].um_I.iw[9] ,
    \top_I.branch[16].block[5].um_I.iw[8] ,
    \top_I.branch[16].block[5].um_I.iw[7] ,
    \top_I.branch[16].block[5].um_I.iw[6] ,
    \top_I.branch[16].block[5].um_I.iw[5] ,
    \top_I.branch[16].block[5].um_I.iw[4] ,
    \top_I.branch[16].block[5].um_I.iw[3] ,
    \top_I.branch[16].block[5].um_I.iw[2] ,
    \top_I.branch[16].block[5].um_I.iw[1] ,
    \top_I.branch[16].block[5].um_I.clk ,
    \top_I.branch[16].block[4].um_I.iw[17] ,
    \top_I.branch[16].block[4].um_I.iw[16] ,
    \top_I.branch[16].block[4].um_I.iw[15] ,
    \top_I.branch[16].block[4].um_I.iw[14] ,
    \top_I.branch[16].block[4].um_I.iw[13] ,
    \top_I.branch[16].block[4].um_I.iw[12] ,
    \top_I.branch[16].block[4].um_I.iw[11] ,
    \top_I.branch[16].block[4].um_I.iw[10] ,
    \top_I.branch[16].block[4].um_I.iw[9] ,
    \top_I.branch[16].block[4].um_I.iw[8] ,
    \top_I.branch[16].block[4].um_I.iw[7] ,
    \top_I.branch[16].block[4].um_I.iw[6] ,
    \top_I.branch[16].block[4].um_I.iw[5] ,
    \top_I.branch[16].block[4].um_I.iw[4] ,
    \top_I.branch[16].block[4].um_I.iw[3] ,
    \top_I.branch[16].block[4].um_I.iw[2] ,
    \top_I.branch[16].block[4].um_I.iw[1] ,
    \top_I.branch[16].block[4].um_I.clk ,
    \top_I.branch[16].block[3].um_I.iw[17] ,
    \top_I.branch[16].block[3].um_I.iw[16] ,
    \top_I.branch[16].block[3].um_I.iw[15] ,
    \top_I.branch[16].block[3].um_I.iw[14] ,
    \top_I.branch[16].block[3].um_I.iw[13] ,
    \top_I.branch[16].block[3].um_I.iw[12] ,
    \top_I.branch[16].block[3].um_I.iw[11] ,
    \top_I.branch[16].block[3].um_I.iw[10] ,
    \top_I.branch[16].block[3].um_I.iw[9] ,
    \top_I.branch[16].block[3].um_I.iw[8] ,
    \top_I.branch[16].block[3].um_I.iw[7] ,
    \top_I.branch[16].block[3].um_I.iw[6] ,
    \top_I.branch[16].block[3].um_I.iw[5] ,
    \top_I.branch[16].block[3].um_I.iw[4] ,
    \top_I.branch[16].block[3].um_I.iw[3] ,
    \top_I.branch[16].block[3].um_I.iw[2] ,
    \top_I.branch[16].block[3].um_I.iw[1] ,
    \top_I.branch[16].block[3].um_I.clk ,
    \top_I.branch[16].block[2].um_I.iw[17] ,
    \top_I.branch[16].block[2].um_I.iw[16] ,
    \top_I.branch[16].block[2].um_I.iw[15] ,
    \top_I.branch[16].block[2].um_I.iw[14] ,
    \top_I.branch[16].block[2].um_I.iw[13] ,
    \top_I.branch[16].block[2].um_I.iw[12] ,
    \top_I.branch[16].block[2].um_I.iw[11] ,
    \top_I.branch[16].block[2].um_I.iw[10] ,
    \top_I.branch[16].block[2].um_I.iw[9] ,
    \top_I.branch[16].block[2].um_I.iw[8] ,
    \top_I.branch[16].block[2].um_I.iw[7] ,
    \top_I.branch[16].block[2].um_I.iw[6] ,
    \top_I.branch[16].block[2].um_I.iw[5] ,
    \top_I.branch[16].block[2].um_I.iw[4] ,
    \top_I.branch[16].block[2].um_I.iw[3] ,
    \top_I.branch[16].block[2].um_I.iw[2] ,
    \top_I.branch[16].block[2].um_I.iw[1] ,
    \top_I.branch[16].block[2].um_I.clk ,
    \top_I.branch[16].block[1].um_I.iw[17] ,
    \top_I.branch[16].block[1].um_I.iw[16] ,
    \top_I.branch[16].block[1].um_I.iw[15] ,
    \top_I.branch[16].block[1].um_I.iw[14] ,
    \top_I.branch[16].block[1].um_I.iw[13] ,
    \top_I.branch[16].block[1].um_I.iw[12] ,
    \top_I.branch[16].block[1].um_I.iw[11] ,
    \top_I.branch[16].block[1].um_I.iw[10] ,
    \top_I.branch[16].block[1].um_I.iw[9] ,
    \top_I.branch[16].block[1].um_I.iw[8] ,
    \top_I.branch[16].block[1].um_I.iw[7] ,
    \top_I.branch[16].block[1].um_I.iw[6] ,
    \top_I.branch[16].block[1].um_I.iw[5] ,
    \top_I.branch[16].block[1].um_I.iw[4] ,
    \top_I.branch[16].block[1].um_I.iw[3] ,
    \top_I.branch[16].block[1].um_I.iw[2] ,
    \top_I.branch[16].block[1].um_I.iw[1] ,
    \top_I.branch[16].block[1].um_I.clk ,
    \top_I.branch[16].block[0].um_I.iw[17] ,
    \top_I.branch[16].block[0].um_I.iw[16] ,
    \top_I.branch[16].block[0].um_I.iw[15] ,
    \top_I.branch[16].block[0].um_I.iw[14] ,
    \top_I.branch[16].block[0].um_I.iw[13] ,
    \top_I.branch[16].block[0].um_I.iw[12] ,
    \top_I.branch[16].block[0].um_I.iw[11] ,
    \top_I.branch[16].block[0].um_I.iw[10] ,
    \top_I.branch[16].block[0].um_I.iw[9] ,
    \top_I.branch[16].block[0].um_I.iw[8] ,
    \top_I.branch[16].block[0].um_I.iw[7] ,
    \top_I.branch[16].block[0].um_I.iw[6] ,
    \top_I.branch[16].block[0].um_I.iw[5] ,
    \top_I.branch[16].block[0].um_I.iw[4] ,
    \top_I.branch[16].block[0].um_I.iw[3] ,
    \top_I.branch[16].block[0].um_I.iw[2] ,
    \top_I.branch[16].block[0].um_I.iw[1] ,
    \top_I.branch[16].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[15].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[14].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[13].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[12].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[11].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[10].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[9].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[8].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[7].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[6].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[5].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[4].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[3].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[2].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[1].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero ,
    \top_I.branch[16].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[16].block[15].um_I.pg_vdd ,
    \top_I.branch[16].block[14].um_I.pg_vdd ,
    \top_I.branch[16].block[13].um_I.pg_vdd ,
    \top_I.branch[16].block[12].um_I.pg_vdd ,
    \top_I.branch[16].block[11].um_I.pg_vdd ,
    \top_I.branch[16].block[10].um_I.pg_vdd ,
    \top_I.branch[16].block[9].um_I.pg_vdd ,
    \top_I.branch[16].block[8].um_I.pg_vdd ,
    \top_I.branch[16].block[7].um_I.pg_vdd ,
    \top_I.branch[16].block[6].um_I.pg_vdd ,
    \top_I.branch[16].block[5].um_I.pg_vdd ,
    \top_I.branch[16].block[4].um_I.pg_vdd ,
    \top_I.branch[16].block[3].um_I.pg_vdd ,
    \top_I.branch[16].block[2].um_I.pg_vdd ,
    \top_I.branch[16].block[1].um_I.pg_vdd ,
    \top_I.branch[16].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[17].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[17].l_addr[3] ),
    .k_zero(\top_I.branch[17].l_addr[0] ),
    .addr({\top_I.branch[17].l_addr[3] ,
    \top_I.branch[17].l_addr[0] ,
    \top_I.branch[17].l_addr[0] ,
    \top_I.branch[17].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[17].block[15].um_I.ena ,
    \top_I.branch[17].block[14].um_I.ena ,
    \top_I.branch[17].block[13].um_I.ena ,
    \top_I.branch[17].block[12].um_I.ena ,
    \top_I.branch[17].block[11].um_I.ena ,
    \top_I.branch[17].block[10].um_I.ena ,
    \top_I.branch[17].block[9].um_I.ena ,
    \top_I.branch[17].block[8].um_I.ena ,
    \top_I.branch[17].block[7].um_I.ena ,
    \top_I.branch[17].block[6].um_I.ena ,
    \top_I.branch[17].block[5].um_I.ena ,
    \top_I.branch[17].block[4].um_I.ena ,
    \top_I.branch[17].block[3].um_I.ena ,
    \top_I.branch[17].block[2].um_I.ena ,
    \top_I.branch[17].block[1].um_I.ena ,
    \top_I.branch[17].block[0].um_I.ena }),
    .um_iw({\top_I.branch[17].block[15].um_I.iw[17] ,
    \top_I.branch[17].block[15].um_I.iw[16] ,
    \top_I.branch[17].block[15].um_I.iw[15] ,
    \top_I.branch[17].block[15].um_I.iw[14] ,
    \top_I.branch[17].block[15].um_I.iw[13] ,
    \top_I.branch[17].block[15].um_I.iw[12] ,
    \top_I.branch[17].block[15].um_I.iw[11] ,
    \top_I.branch[17].block[15].um_I.iw[10] ,
    \top_I.branch[17].block[15].um_I.iw[9] ,
    \top_I.branch[17].block[15].um_I.iw[8] ,
    \top_I.branch[17].block[15].um_I.iw[7] ,
    \top_I.branch[17].block[15].um_I.iw[6] ,
    \top_I.branch[17].block[15].um_I.iw[5] ,
    \top_I.branch[17].block[15].um_I.iw[4] ,
    \top_I.branch[17].block[15].um_I.iw[3] ,
    \top_I.branch[17].block[15].um_I.iw[2] ,
    \top_I.branch[17].block[15].um_I.iw[1] ,
    \top_I.branch[17].block[15].um_I.clk ,
    \top_I.branch[17].block[14].um_I.iw[17] ,
    \top_I.branch[17].block[14].um_I.iw[16] ,
    \top_I.branch[17].block[14].um_I.iw[15] ,
    \top_I.branch[17].block[14].um_I.iw[14] ,
    \top_I.branch[17].block[14].um_I.iw[13] ,
    \top_I.branch[17].block[14].um_I.iw[12] ,
    \top_I.branch[17].block[14].um_I.iw[11] ,
    \top_I.branch[17].block[14].um_I.iw[10] ,
    \top_I.branch[17].block[14].um_I.iw[9] ,
    \top_I.branch[17].block[14].um_I.iw[8] ,
    \top_I.branch[17].block[14].um_I.iw[7] ,
    \top_I.branch[17].block[14].um_I.iw[6] ,
    \top_I.branch[17].block[14].um_I.iw[5] ,
    \top_I.branch[17].block[14].um_I.iw[4] ,
    \top_I.branch[17].block[14].um_I.iw[3] ,
    \top_I.branch[17].block[14].um_I.iw[2] ,
    \top_I.branch[17].block[14].um_I.iw[1] ,
    \top_I.branch[17].block[14].um_I.clk ,
    \top_I.branch[17].block[13].um_I.iw[17] ,
    \top_I.branch[17].block[13].um_I.iw[16] ,
    \top_I.branch[17].block[13].um_I.iw[15] ,
    \top_I.branch[17].block[13].um_I.iw[14] ,
    \top_I.branch[17].block[13].um_I.iw[13] ,
    \top_I.branch[17].block[13].um_I.iw[12] ,
    \top_I.branch[17].block[13].um_I.iw[11] ,
    \top_I.branch[17].block[13].um_I.iw[10] ,
    \top_I.branch[17].block[13].um_I.iw[9] ,
    \top_I.branch[17].block[13].um_I.iw[8] ,
    \top_I.branch[17].block[13].um_I.iw[7] ,
    \top_I.branch[17].block[13].um_I.iw[6] ,
    \top_I.branch[17].block[13].um_I.iw[5] ,
    \top_I.branch[17].block[13].um_I.iw[4] ,
    \top_I.branch[17].block[13].um_I.iw[3] ,
    \top_I.branch[17].block[13].um_I.iw[2] ,
    \top_I.branch[17].block[13].um_I.iw[1] ,
    \top_I.branch[17].block[13].um_I.clk ,
    \top_I.branch[17].block[12].um_I.iw[17] ,
    \top_I.branch[17].block[12].um_I.iw[16] ,
    \top_I.branch[17].block[12].um_I.iw[15] ,
    \top_I.branch[17].block[12].um_I.iw[14] ,
    \top_I.branch[17].block[12].um_I.iw[13] ,
    \top_I.branch[17].block[12].um_I.iw[12] ,
    \top_I.branch[17].block[12].um_I.iw[11] ,
    \top_I.branch[17].block[12].um_I.iw[10] ,
    \top_I.branch[17].block[12].um_I.iw[9] ,
    \top_I.branch[17].block[12].um_I.iw[8] ,
    \top_I.branch[17].block[12].um_I.iw[7] ,
    \top_I.branch[17].block[12].um_I.iw[6] ,
    \top_I.branch[17].block[12].um_I.iw[5] ,
    \top_I.branch[17].block[12].um_I.iw[4] ,
    \top_I.branch[17].block[12].um_I.iw[3] ,
    \top_I.branch[17].block[12].um_I.iw[2] ,
    \top_I.branch[17].block[12].um_I.iw[1] ,
    \top_I.branch[17].block[12].um_I.clk ,
    \top_I.branch[17].block[11].um_I.iw[17] ,
    \top_I.branch[17].block[11].um_I.iw[16] ,
    \top_I.branch[17].block[11].um_I.iw[15] ,
    \top_I.branch[17].block[11].um_I.iw[14] ,
    \top_I.branch[17].block[11].um_I.iw[13] ,
    \top_I.branch[17].block[11].um_I.iw[12] ,
    \top_I.branch[17].block[11].um_I.iw[11] ,
    \top_I.branch[17].block[11].um_I.iw[10] ,
    \top_I.branch[17].block[11].um_I.iw[9] ,
    \top_I.branch[17].block[11].um_I.iw[8] ,
    \top_I.branch[17].block[11].um_I.iw[7] ,
    \top_I.branch[17].block[11].um_I.iw[6] ,
    \top_I.branch[17].block[11].um_I.iw[5] ,
    \top_I.branch[17].block[11].um_I.iw[4] ,
    \top_I.branch[17].block[11].um_I.iw[3] ,
    \top_I.branch[17].block[11].um_I.iw[2] ,
    \top_I.branch[17].block[11].um_I.iw[1] ,
    \top_I.branch[17].block[11].um_I.clk ,
    \top_I.branch[17].block[10].um_I.iw[17] ,
    \top_I.branch[17].block[10].um_I.iw[16] ,
    \top_I.branch[17].block[10].um_I.iw[15] ,
    \top_I.branch[17].block[10].um_I.iw[14] ,
    \top_I.branch[17].block[10].um_I.iw[13] ,
    \top_I.branch[17].block[10].um_I.iw[12] ,
    \top_I.branch[17].block[10].um_I.iw[11] ,
    \top_I.branch[17].block[10].um_I.iw[10] ,
    \top_I.branch[17].block[10].um_I.iw[9] ,
    \top_I.branch[17].block[10].um_I.iw[8] ,
    \top_I.branch[17].block[10].um_I.iw[7] ,
    \top_I.branch[17].block[10].um_I.iw[6] ,
    \top_I.branch[17].block[10].um_I.iw[5] ,
    \top_I.branch[17].block[10].um_I.iw[4] ,
    \top_I.branch[17].block[10].um_I.iw[3] ,
    \top_I.branch[17].block[10].um_I.iw[2] ,
    \top_I.branch[17].block[10].um_I.iw[1] ,
    \top_I.branch[17].block[10].um_I.clk ,
    \top_I.branch[17].block[9].um_I.iw[17] ,
    \top_I.branch[17].block[9].um_I.iw[16] ,
    \top_I.branch[17].block[9].um_I.iw[15] ,
    \top_I.branch[17].block[9].um_I.iw[14] ,
    \top_I.branch[17].block[9].um_I.iw[13] ,
    \top_I.branch[17].block[9].um_I.iw[12] ,
    \top_I.branch[17].block[9].um_I.iw[11] ,
    \top_I.branch[17].block[9].um_I.iw[10] ,
    \top_I.branch[17].block[9].um_I.iw[9] ,
    \top_I.branch[17].block[9].um_I.iw[8] ,
    \top_I.branch[17].block[9].um_I.iw[7] ,
    \top_I.branch[17].block[9].um_I.iw[6] ,
    \top_I.branch[17].block[9].um_I.iw[5] ,
    \top_I.branch[17].block[9].um_I.iw[4] ,
    \top_I.branch[17].block[9].um_I.iw[3] ,
    \top_I.branch[17].block[9].um_I.iw[2] ,
    \top_I.branch[17].block[9].um_I.iw[1] ,
    \top_I.branch[17].block[9].um_I.clk ,
    \top_I.branch[17].block[8].um_I.iw[17] ,
    \top_I.branch[17].block[8].um_I.iw[16] ,
    \top_I.branch[17].block[8].um_I.iw[15] ,
    \top_I.branch[17].block[8].um_I.iw[14] ,
    \top_I.branch[17].block[8].um_I.iw[13] ,
    \top_I.branch[17].block[8].um_I.iw[12] ,
    \top_I.branch[17].block[8].um_I.iw[11] ,
    \top_I.branch[17].block[8].um_I.iw[10] ,
    \top_I.branch[17].block[8].um_I.iw[9] ,
    \top_I.branch[17].block[8].um_I.iw[8] ,
    \top_I.branch[17].block[8].um_I.iw[7] ,
    \top_I.branch[17].block[8].um_I.iw[6] ,
    \top_I.branch[17].block[8].um_I.iw[5] ,
    \top_I.branch[17].block[8].um_I.iw[4] ,
    \top_I.branch[17].block[8].um_I.iw[3] ,
    \top_I.branch[17].block[8].um_I.iw[2] ,
    \top_I.branch[17].block[8].um_I.iw[1] ,
    \top_I.branch[17].block[8].um_I.clk ,
    \top_I.branch[17].block[7].um_I.iw[17] ,
    \top_I.branch[17].block[7].um_I.iw[16] ,
    \top_I.branch[17].block[7].um_I.iw[15] ,
    \top_I.branch[17].block[7].um_I.iw[14] ,
    \top_I.branch[17].block[7].um_I.iw[13] ,
    \top_I.branch[17].block[7].um_I.iw[12] ,
    \top_I.branch[17].block[7].um_I.iw[11] ,
    \top_I.branch[17].block[7].um_I.iw[10] ,
    \top_I.branch[17].block[7].um_I.iw[9] ,
    \top_I.branch[17].block[7].um_I.iw[8] ,
    \top_I.branch[17].block[7].um_I.iw[7] ,
    \top_I.branch[17].block[7].um_I.iw[6] ,
    \top_I.branch[17].block[7].um_I.iw[5] ,
    \top_I.branch[17].block[7].um_I.iw[4] ,
    \top_I.branch[17].block[7].um_I.iw[3] ,
    \top_I.branch[17].block[7].um_I.iw[2] ,
    \top_I.branch[17].block[7].um_I.iw[1] ,
    \top_I.branch[17].block[7].um_I.clk ,
    \top_I.branch[17].block[6].um_I.iw[17] ,
    \top_I.branch[17].block[6].um_I.iw[16] ,
    \top_I.branch[17].block[6].um_I.iw[15] ,
    \top_I.branch[17].block[6].um_I.iw[14] ,
    \top_I.branch[17].block[6].um_I.iw[13] ,
    \top_I.branch[17].block[6].um_I.iw[12] ,
    \top_I.branch[17].block[6].um_I.iw[11] ,
    \top_I.branch[17].block[6].um_I.iw[10] ,
    \top_I.branch[17].block[6].um_I.iw[9] ,
    \top_I.branch[17].block[6].um_I.iw[8] ,
    \top_I.branch[17].block[6].um_I.iw[7] ,
    \top_I.branch[17].block[6].um_I.iw[6] ,
    \top_I.branch[17].block[6].um_I.iw[5] ,
    \top_I.branch[17].block[6].um_I.iw[4] ,
    \top_I.branch[17].block[6].um_I.iw[3] ,
    \top_I.branch[17].block[6].um_I.iw[2] ,
    \top_I.branch[17].block[6].um_I.iw[1] ,
    \top_I.branch[17].block[6].um_I.clk ,
    \top_I.branch[17].block[5].um_I.iw[17] ,
    \top_I.branch[17].block[5].um_I.iw[16] ,
    \top_I.branch[17].block[5].um_I.iw[15] ,
    \top_I.branch[17].block[5].um_I.iw[14] ,
    \top_I.branch[17].block[5].um_I.iw[13] ,
    \top_I.branch[17].block[5].um_I.iw[12] ,
    \top_I.branch[17].block[5].um_I.iw[11] ,
    \top_I.branch[17].block[5].um_I.iw[10] ,
    \top_I.branch[17].block[5].um_I.iw[9] ,
    \top_I.branch[17].block[5].um_I.iw[8] ,
    \top_I.branch[17].block[5].um_I.iw[7] ,
    \top_I.branch[17].block[5].um_I.iw[6] ,
    \top_I.branch[17].block[5].um_I.iw[5] ,
    \top_I.branch[17].block[5].um_I.iw[4] ,
    \top_I.branch[17].block[5].um_I.iw[3] ,
    \top_I.branch[17].block[5].um_I.iw[2] ,
    \top_I.branch[17].block[5].um_I.iw[1] ,
    \top_I.branch[17].block[5].um_I.clk ,
    \top_I.branch[17].block[4].um_I.iw[17] ,
    \top_I.branch[17].block[4].um_I.iw[16] ,
    \top_I.branch[17].block[4].um_I.iw[15] ,
    \top_I.branch[17].block[4].um_I.iw[14] ,
    \top_I.branch[17].block[4].um_I.iw[13] ,
    \top_I.branch[17].block[4].um_I.iw[12] ,
    \top_I.branch[17].block[4].um_I.iw[11] ,
    \top_I.branch[17].block[4].um_I.iw[10] ,
    \top_I.branch[17].block[4].um_I.iw[9] ,
    \top_I.branch[17].block[4].um_I.iw[8] ,
    \top_I.branch[17].block[4].um_I.iw[7] ,
    \top_I.branch[17].block[4].um_I.iw[6] ,
    \top_I.branch[17].block[4].um_I.iw[5] ,
    \top_I.branch[17].block[4].um_I.iw[4] ,
    \top_I.branch[17].block[4].um_I.iw[3] ,
    \top_I.branch[17].block[4].um_I.iw[2] ,
    \top_I.branch[17].block[4].um_I.iw[1] ,
    \top_I.branch[17].block[4].um_I.clk ,
    \top_I.branch[17].block[3].um_I.iw[17] ,
    \top_I.branch[17].block[3].um_I.iw[16] ,
    \top_I.branch[17].block[3].um_I.iw[15] ,
    \top_I.branch[17].block[3].um_I.iw[14] ,
    \top_I.branch[17].block[3].um_I.iw[13] ,
    \top_I.branch[17].block[3].um_I.iw[12] ,
    \top_I.branch[17].block[3].um_I.iw[11] ,
    \top_I.branch[17].block[3].um_I.iw[10] ,
    \top_I.branch[17].block[3].um_I.iw[9] ,
    \top_I.branch[17].block[3].um_I.iw[8] ,
    \top_I.branch[17].block[3].um_I.iw[7] ,
    \top_I.branch[17].block[3].um_I.iw[6] ,
    \top_I.branch[17].block[3].um_I.iw[5] ,
    \top_I.branch[17].block[3].um_I.iw[4] ,
    \top_I.branch[17].block[3].um_I.iw[3] ,
    \top_I.branch[17].block[3].um_I.iw[2] ,
    \top_I.branch[17].block[3].um_I.iw[1] ,
    \top_I.branch[17].block[3].um_I.clk ,
    \top_I.branch[17].block[2].um_I.iw[17] ,
    \top_I.branch[17].block[2].um_I.iw[16] ,
    \top_I.branch[17].block[2].um_I.iw[15] ,
    \top_I.branch[17].block[2].um_I.iw[14] ,
    \top_I.branch[17].block[2].um_I.iw[13] ,
    \top_I.branch[17].block[2].um_I.iw[12] ,
    \top_I.branch[17].block[2].um_I.iw[11] ,
    \top_I.branch[17].block[2].um_I.iw[10] ,
    \top_I.branch[17].block[2].um_I.iw[9] ,
    \top_I.branch[17].block[2].um_I.iw[8] ,
    \top_I.branch[17].block[2].um_I.iw[7] ,
    \top_I.branch[17].block[2].um_I.iw[6] ,
    \top_I.branch[17].block[2].um_I.iw[5] ,
    \top_I.branch[17].block[2].um_I.iw[4] ,
    \top_I.branch[17].block[2].um_I.iw[3] ,
    \top_I.branch[17].block[2].um_I.iw[2] ,
    \top_I.branch[17].block[2].um_I.iw[1] ,
    \top_I.branch[17].block[2].um_I.clk ,
    \top_I.branch[17].block[1].um_I.iw[17] ,
    \top_I.branch[17].block[1].um_I.iw[16] ,
    \top_I.branch[17].block[1].um_I.iw[15] ,
    \top_I.branch[17].block[1].um_I.iw[14] ,
    \top_I.branch[17].block[1].um_I.iw[13] ,
    \top_I.branch[17].block[1].um_I.iw[12] ,
    \top_I.branch[17].block[1].um_I.iw[11] ,
    \top_I.branch[17].block[1].um_I.iw[10] ,
    \top_I.branch[17].block[1].um_I.iw[9] ,
    \top_I.branch[17].block[1].um_I.iw[8] ,
    \top_I.branch[17].block[1].um_I.iw[7] ,
    \top_I.branch[17].block[1].um_I.iw[6] ,
    \top_I.branch[17].block[1].um_I.iw[5] ,
    \top_I.branch[17].block[1].um_I.iw[4] ,
    \top_I.branch[17].block[1].um_I.iw[3] ,
    \top_I.branch[17].block[1].um_I.iw[2] ,
    \top_I.branch[17].block[1].um_I.iw[1] ,
    \top_I.branch[17].block[1].um_I.clk ,
    \top_I.branch[17].block[0].um_I.iw[17] ,
    \top_I.branch[17].block[0].um_I.iw[16] ,
    \top_I.branch[17].block[0].um_I.iw[15] ,
    \top_I.branch[17].block[0].um_I.iw[14] ,
    \top_I.branch[17].block[0].um_I.iw[13] ,
    \top_I.branch[17].block[0].um_I.iw[12] ,
    \top_I.branch[17].block[0].um_I.iw[11] ,
    \top_I.branch[17].block[0].um_I.iw[10] ,
    \top_I.branch[17].block[0].um_I.iw[9] ,
    \top_I.branch[17].block[0].um_I.iw[8] ,
    \top_I.branch[17].block[0].um_I.iw[7] ,
    \top_I.branch[17].block[0].um_I.iw[6] ,
    \top_I.branch[17].block[0].um_I.iw[5] ,
    \top_I.branch[17].block[0].um_I.iw[4] ,
    \top_I.branch[17].block[0].um_I.iw[3] ,
    \top_I.branch[17].block[0].um_I.iw[2] ,
    \top_I.branch[17].block[0].um_I.iw[1] ,
    \top_I.branch[17].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[15].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[14].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[13].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[12].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[11].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[10].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[9].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[8].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[7].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[6].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[5].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[4].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[3].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[2].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[1].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero ,
    \top_I.branch[17].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[17].block[15].um_I.pg_vdd ,
    \top_I.branch[17].block[14].um_I.pg_vdd ,
    \top_I.branch[17].block[13].um_I.pg_vdd ,
    \top_I.branch[17].block[12].um_I.pg_vdd ,
    \top_I.branch[17].block[11].um_I.pg_vdd ,
    \top_I.branch[17].block[10].um_I.pg_vdd ,
    \top_I.branch[17].block[9].um_I.pg_vdd ,
    \top_I.branch[17].block[8].um_I.pg_vdd ,
    \top_I.branch[17].block[7].um_I.pg_vdd ,
    \top_I.branch[17].block[6].um_I.pg_vdd ,
    \top_I.branch[17].block[5].um_I.pg_vdd ,
    \top_I.branch[17].block[4].um_I.pg_vdd ,
    \top_I.branch[17].block[3].um_I.pg_vdd ,
    \top_I.branch[17].block[2].um_I.pg_vdd ,
    \top_I.branch[17].block[1].um_I.pg_vdd ,
    \top_I.branch[17].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[18].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[18].l_addr[0] ),
    .k_zero(\top_I.branch[18].l_addr[1] ),
    .addr({\top_I.branch[18].l_addr[0] ,
    \top_I.branch[18].l_addr[1] ,
    \top_I.branch[18].l_addr[1] ,
    \top_I.branch[18].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[18].block[15].um_I.ena ,
    \top_I.branch[18].block[14].um_I.ena ,
    \top_I.branch[18].block[13].um_I.ena ,
    \top_I.branch[18].block[12].um_I.ena ,
    \top_I.branch[18].block[11].um_I.ena ,
    \top_I.branch[18].block[10].um_I.ena ,
    \top_I.branch[18].block[9].um_I.ena ,
    \top_I.branch[18].block[8].um_I.ena ,
    \top_I.branch[18].block[7].um_I.ena ,
    \top_I.branch[18].block[6].um_I.ena ,
    \top_I.branch[18].block[5].um_I.ena ,
    \top_I.branch[18].block[4].um_I.ena ,
    \top_I.branch[18].block[3].um_I.ena ,
    \top_I.branch[18].block[2].um_I.ena ,
    \top_I.branch[18].block[1].um_I.ena ,
    \top_I.branch[18].block[0].um_I.ena }),
    .um_iw({\top_I.branch[18].block[15].um_I.iw[17] ,
    \top_I.branch[18].block[15].um_I.iw[16] ,
    \top_I.branch[18].block[15].um_I.iw[15] ,
    \top_I.branch[18].block[15].um_I.iw[14] ,
    \top_I.branch[18].block[15].um_I.iw[13] ,
    \top_I.branch[18].block[15].um_I.iw[12] ,
    \top_I.branch[18].block[15].um_I.iw[11] ,
    \top_I.branch[18].block[15].um_I.iw[10] ,
    \top_I.branch[18].block[15].um_I.iw[9] ,
    \top_I.branch[18].block[15].um_I.iw[8] ,
    \top_I.branch[18].block[15].um_I.iw[7] ,
    \top_I.branch[18].block[15].um_I.iw[6] ,
    \top_I.branch[18].block[15].um_I.iw[5] ,
    \top_I.branch[18].block[15].um_I.iw[4] ,
    \top_I.branch[18].block[15].um_I.iw[3] ,
    \top_I.branch[18].block[15].um_I.iw[2] ,
    \top_I.branch[18].block[15].um_I.iw[1] ,
    \top_I.branch[18].block[15].um_I.clk ,
    \top_I.branch[18].block[14].um_I.iw[17] ,
    \top_I.branch[18].block[14].um_I.iw[16] ,
    \top_I.branch[18].block[14].um_I.iw[15] ,
    \top_I.branch[18].block[14].um_I.iw[14] ,
    \top_I.branch[18].block[14].um_I.iw[13] ,
    \top_I.branch[18].block[14].um_I.iw[12] ,
    \top_I.branch[18].block[14].um_I.iw[11] ,
    \top_I.branch[18].block[14].um_I.iw[10] ,
    \top_I.branch[18].block[14].um_I.iw[9] ,
    \top_I.branch[18].block[14].um_I.iw[8] ,
    \top_I.branch[18].block[14].um_I.iw[7] ,
    \top_I.branch[18].block[14].um_I.iw[6] ,
    \top_I.branch[18].block[14].um_I.iw[5] ,
    \top_I.branch[18].block[14].um_I.iw[4] ,
    \top_I.branch[18].block[14].um_I.iw[3] ,
    \top_I.branch[18].block[14].um_I.iw[2] ,
    \top_I.branch[18].block[14].um_I.iw[1] ,
    \top_I.branch[18].block[14].um_I.clk ,
    \top_I.branch[18].block[13].um_I.iw[17] ,
    \top_I.branch[18].block[13].um_I.iw[16] ,
    \top_I.branch[18].block[13].um_I.iw[15] ,
    \top_I.branch[18].block[13].um_I.iw[14] ,
    \top_I.branch[18].block[13].um_I.iw[13] ,
    \top_I.branch[18].block[13].um_I.iw[12] ,
    \top_I.branch[18].block[13].um_I.iw[11] ,
    \top_I.branch[18].block[13].um_I.iw[10] ,
    \top_I.branch[18].block[13].um_I.iw[9] ,
    \top_I.branch[18].block[13].um_I.iw[8] ,
    \top_I.branch[18].block[13].um_I.iw[7] ,
    \top_I.branch[18].block[13].um_I.iw[6] ,
    \top_I.branch[18].block[13].um_I.iw[5] ,
    \top_I.branch[18].block[13].um_I.iw[4] ,
    \top_I.branch[18].block[13].um_I.iw[3] ,
    \top_I.branch[18].block[13].um_I.iw[2] ,
    \top_I.branch[18].block[13].um_I.iw[1] ,
    \top_I.branch[18].block[13].um_I.clk ,
    \top_I.branch[18].block[12].um_I.iw[17] ,
    \top_I.branch[18].block[12].um_I.iw[16] ,
    \top_I.branch[18].block[12].um_I.iw[15] ,
    \top_I.branch[18].block[12].um_I.iw[14] ,
    \top_I.branch[18].block[12].um_I.iw[13] ,
    \top_I.branch[18].block[12].um_I.iw[12] ,
    \top_I.branch[18].block[12].um_I.iw[11] ,
    \top_I.branch[18].block[12].um_I.iw[10] ,
    \top_I.branch[18].block[12].um_I.iw[9] ,
    \top_I.branch[18].block[12].um_I.iw[8] ,
    \top_I.branch[18].block[12].um_I.iw[7] ,
    \top_I.branch[18].block[12].um_I.iw[6] ,
    \top_I.branch[18].block[12].um_I.iw[5] ,
    \top_I.branch[18].block[12].um_I.iw[4] ,
    \top_I.branch[18].block[12].um_I.iw[3] ,
    \top_I.branch[18].block[12].um_I.iw[2] ,
    \top_I.branch[18].block[12].um_I.iw[1] ,
    \top_I.branch[18].block[12].um_I.clk ,
    \top_I.branch[18].block[11].um_I.iw[17] ,
    \top_I.branch[18].block[11].um_I.iw[16] ,
    \top_I.branch[18].block[11].um_I.iw[15] ,
    \top_I.branch[18].block[11].um_I.iw[14] ,
    \top_I.branch[18].block[11].um_I.iw[13] ,
    \top_I.branch[18].block[11].um_I.iw[12] ,
    \top_I.branch[18].block[11].um_I.iw[11] ,
    \top_I.branch[18].block[11].um_I.iw[10] ,
    \top_I.branch[18].block[11].um_I.iw[9] ,
    \top_I.branch[18].block[11].um_I.iw[8] ,
    \top_I.branch[18].block[11].um_I.iw[7] ,
    \top_I.branch[18].block[11].um_I.iw[6] ,
    \top_I.branch[18].block[11].um_I.iw[5] ,
    \top_I.branch[18].block[11].um_I.iw[4] ,
    \top_I.branch[18].block[11].um_I.iw[3] ,
    \top_I.branch[18].block[11].um_I.iw[2] ,
    \top_I.branch[18].block[11].um_I.iw[1] ,
    \top_I.branch[18].block[11].um_I.clk ,
    \top_I.branch[18].block[10].um_I.iw[17] ,
    \top_I.branch[18].block[10].um_I.iw[16] ,
    \top_I.branch[18].block[10].um_I.iw[15] ,
    \top_I.branch[18].block[10].um_I.iw[14] ,
    \top_I.branch[18].block[10].um_I.iw[13] ,
    \top_I.branch[18].block[10].um_I.iw[12] ,
    \top_I.branch[18].block[10].um_I.iw[11] ,
    \top_I.branch[18].block[10].um_I.iw[10] ,
    \top_I.branch[18].block[10].um_I.iw[9] ,
    \top_I.branch[18].block[10].um_I.iw[8] ,
    \top_I.branch[18].block[10].um_I.iw[7] ,
    \top_I.branch[18].block[10].um_I.iw[6] ,
    \top_I.branch[18].block[10].um_I.iw[5] ,
    \top_I.branch[18].block[10].um_I.iw[4] ,
    \top_I.branch[18].block[10].um_I.iw[3] ,
    \top_I.branch[18].block[10].um_I.iw[2] ,
    \top_I.branch[18].block[10].um_I.iw[1] ,
    \top_I.branch[18].block[10].um_I.clk ,
    \top_I.branch[18].block[9].um_I.iw[17] ,
    \top_I.branch[18].block[9].um_I.iw[16] ,
    \top_I.branch[18].block[9].um_I.iw[15] ,
    \top_I.branch[18].block[9].um_I.iw[14] ,
    \top_I.branch[18].block[9].um_I.iw[13] ,
    \top_I.branch[18].block[9].um_I.iw[12] ,
    \top_I.branch[18].block[9].um_I.iw[11] ,
    \top_I.branch[18].block[9].um_I.iw[10] ,
    \top_I.branch[18].block[9].um_I.iw[9] ,
    \top_I.branch[18].block[9].um_I.iw[8] ,
    \top_I.branch[18].block[9].um_I.iw[7] ,
    \top_I.branch[18].block[9].um_I.iw[6] ,
    \top_I.branch[18].block[9].um_I.iw[5] ,
    \top_I.branch[18].block[9].um_I.iw[4] ,
    \top_I.branch[18].block[9].um_I.iw[3] ,
    \top_I.branch[18].block[9].um_I.iw[2] ,
    \top_I.branch[18].block[9].um_I.iw[1] ,
    \top_I.branch[18].block[9].um_I.clk ,
    \top_I.branch[18].block[8].um_I.iw[17] ,
    \top_I.branch[18].block[8].um_I.iw[16] ,
    \top_I.branch[18].block[8].um_I.iw[15] ,
    \top_I.branch[18].block[8].um_I.iw[14] ,
    \top_I.branch[18].block[8].um_I.iw[13] ,
    \top_I.branch[18].block[8].um_I.iw[12] ,
    \top_I.branch[18].block[8].um_I.iw[11] ,
    \top_I.branch[18].block[8].um_I.iw[10] ,
    \top_I.branch[18].block[8].um_I.iw[9] ,
    \top_I.branch[18].block[8].um_I.iw[8] ,
    \top_I.branch[18].block[8].um_I.iw[7] ,
    \top_I.branch[18].block[8].um_I.iw[6] ,
    \top_I.branch[18].block[8].um_I.iw[5] ,
    \top_I.branch[18].block[8].um_I.iw[4] ,
    \top_I.branch[18].block[8].um_I.iw[3] ,
    \top_I.branch[18].block[8].um_I.iw[2] ,
    \top_I.branch[18].block[8].um_I.iw[1] ,
    \top_I.branch[18].block[8].um_I.clk ,
    \top_I.branch[18].block[7].um_I.iw[17] ,
    \top_I.branch[18].block[7].um_I.iw[16] ,
    \top_I.branch[18].block[7].um_I.iw[15] ,
    \top_I.branch[18].block[7].um_I.iw[14] ,
    \top_I.branch[18].block[7].um_I.iw[13] ,
    \top_I.branch[18].block[7].um_I.iw[12] ,
    \top_I.branch[18].block[7].um_I.iw[11] ,
    \top_I.branch[18].block[7].um_I.iw[10] ,
    \top_I.branch[18].block[7].um_I.iw[9] ,
    \top_I.branch[18].block[7].um_I.iw[8] ,
    \top_I.branch[18].block[7].um_I.iw[7] ,
    \top_I.branch[18].block[7].um_I.iw[6] ,
    \top_I.branch[18].block[7].um_I.iw[5] ,
    \top_I.branch[18].block[7].um_I.iw[4] ,
    \top_I.branch[18].block[7].um_I.iw[3] ,
    \top_I.branch[18].block[7].um_I.iw[2] ,
    \top_I.branch[18].block[7].um_I.iw[1] ,
    \top_I.branch[18].block[7].um_I.clk ,
    \top_I.branch[18].block[6].um_I.iw[17] ,
    \top_I.branch[18].block[6].um_I.iw[16] ,
    \top_I.branch[18].block[6].um_I.iw[15] ,
    \top_I.branch[18].block[6].um_I.iw[14] ,
    \top_I.branch[18].block[6].um_I.iw[13] ,
    \top_I.branch[18].block[6].um_I.iw[12] ,
    \top_I.branch[18].block[6].um_I.iw[11] ,
    \top_I.branch[18].block[6].um_I.iw[10] ,
    \top_I.branch[18].block[6].um_I.iw[9] ,
    \top_I.branch[18].block[6].um_I.iw[8] ,
    \top_I.branch[18].block[6].um_I.iw[7] ,
    \top_I.branch[18].block[6].um_I.iw[6] ,
    \top_I.branch[18].block[6].um_I.iw[5] ,
    \top_I.branch[18].block[6].um_I.iw[4] ,
    \top_I.branch[18].block[6].um_I.iw[3] ,
    \top_I.branch[18].block[6].um_I.iw[2] ,
    \top_I.branch[18].block[6].um_I.iw[1] ,
    \top_I.branch[18].block[6].um_I.clk ,
    \top_I.branch[18].block[5].um_I.iw[17] ,
    \top_I.branch[18].block[5].um_I.iw[16] ,
    \top_I.branch[18].block[5].um_I.iw[15] ,
    \top_I.branch[18].block[5].um_I.iw[14] ,
    \top_I.branch[18].block[5].um_I.iw[13] ,
    \top_I.branch[18].block[5].um_I.iw[12] ,
    \top_I.branch[18].block[5].um_I.iw[11] ,
    \top_I.branch[18].block[5].um_I.iw[10] ,
    \top_I.branch[18].block[5].um_I.iw[9] ,
    \top_I.branch[18].block[5].um_I.iw[8] ,
    \top_I.branch[18].block[5].um_I.iw[7] ,
    \top_I.branch[18].block[5].um_I.iw[6] ,
    \top_I.branch[18].block[5].um_I.iw[5] ,
    \top_I.branch[18].block[5].um_I.iw[4] ,
    \top_I.branch[18].block[5].um_I.iw[3] ,
    \top_I.branch[18].block[5].um_I.iw[2] ,
    \top_I.branch[18].block[5].um_I.iw[1] ,
    \top_I.branch[18].block[5].um_I.clk ,
    \top_I.branch[18].block[4].um_I.iw[17] ,
    \top_I.branch[18].block[4].um_I.iw[16] ,
    \top_I.branch[18].block[4].um_I.iw[15] ,
    \top_I.branch[18].block[4].um_I.iw[14] ,
    \top_I.branch[18].block[4].um_I.iw[13] ,
    \top_I.branch[18].block[4].um_I.iw[12] ,
    \top_I.branch[18].block[4].um_I.iw[11] ,
    \top_I.branch[18].block[4].um_I.iw[10] ,
    \top_I.branch[18].block[4].um_I.iw[9] ,
    \top_I.branch[18].block[4].um_I.iw[8] ,
    \top_I.branch[18].block[4].um_I.iw[7] ,
    \top_I.branch[18].block[4].um_I.iw[6] ,
    \top_I.branch[18].block[4].um_I.iw[5] ,
    \top_I.branch[18].block[4].um_I.iw[4] ,
    \top_I.branch[18].block[4].um_I.iw[3] ,
    \top_I.branch[18].block[4].um_I.iw[2] ,
    \top_I.branch[18].block[4].um_I.iw[1] ,
    \top_I.branch[18].block[4].um_I.clk ,
    \top_I.branch[18].block[3].um_I.iw[17] ,
    \top_I.branch[18].block[3].um_I.iw[16] ,
    \top_I.branch[18].block[3].um_I.iw[15] ,
    \top_I.branch[18].block[3].um_I.iw[14] ,
    \top_I.branch[18].block[3].um_I.iw[13] ,
    \top_I.branch[18].block[3].um_I.iw[12] ,
    \top_I.branch[18].block[3].um_I.iw[11] ,
    \top_I.branch[18].block[3].um_I.iw[10] ,
    \top_I.branch[18].block[3].um_I.iw[9] ,
    \top_I.branch[18].block[3].um_I.iw[8] ,
    \top_I.branch[18].block[3].um_I.iw[7] ,
    \top_I.branch[18].block[3].um_I.iw[6] ,
    \top_I.branch[18].block[3].um_I.iw[5] ,
    \top_I.branch[18].block[3].um_I.iw[4] ,
    \top_I.branch[18].block[3].um_I.iw[3] ,
    \top_I.branch[18].block[3].um_I.iw[2] ,
    \top_I.branch[18].block[3].um_I.iw[1] ,
    \top_I.branch[18].block[3].um_I.clk ,
    \top_I.branch[18].block[2].um_I.iw[17] ,
    \top_I.branch[18].block[2].um_I.iw[16] ,
    \top_I.branch[18].block[2].um_I.iw[15] ,
    \top_I.branch[18].block[2].um_I.iw[14] ,
    \top_I.branch[18].block[2].um_I.iw[13] ,
    \top_I.branch[18].block[2].um_I.iw[12] ,
    \top_I.branch[18].block[2].um_I.iw[11] ,
    \top_I.branch[18].block[2].um_I.iw[10] ,
    \top_I.branch[18].block[2].um_I.iw[9] ,
    \top_I.branch[18].block[2].um_I.iw[8] ,
    \top_I.branch[18].block[2].um_I.iw[7] ,
    \top_I.branch[18].block[2].um_I.iw[6] ,
    \top_I.branch[18].block[2].um_I.iw[5] ,
    \top_I.branch[18].block[2].um_I.iw[4] ,
    \top_I.branch[18].block[2].um_I.iw[3] ,
    \top_I.branch[18].block[2].um_I.iw[2] ,
    \top_I.branch[18].block[2].um_I.iw[1] ,
    \top_I.branch[18].block[2].um_I.clk ,
    \top_I.branch[18].block[1].um_I.iw[17] ,
    \top_I.branch[18].block[1].um_I.iw[16] ,
    \top_I.branch[18].block[1].um_I.iw[15] ,
    \top_I.branch[18].block[1].um_I.iw[14] ,
    \top_I.branch[18].block[1].um_I.iw[13] ,
    \top_I.branch[18].block[1].um_I.iw[12] ,
    \top_I.branch[18].block[1].um_I.iw[11] ,
    \top_I.branch[18].block[1].um_I.iw[10] ,
    \top_I.branch[18].block[1].um_I.iw[9] ,
    \top_I.branch[18].block[1].um_I.iw[8] ,
    \top_I.branch[18].block[1].um_I.iw[7] ,
    \top_I.branch[18].block[1].um_I.iw[6] ,
    \top_I.branch[18].block[1].um_I.iw[5] ,
    \top_I.branch[18].block[1].um_I.iw[4] ,
    \top_I.branch[18].block[1].um_I.iw[3] ,
    \top_I.branch[18].block[1].um_I.iw[2] ,
    \top_I.branch[18].block[1].um_I.iw[1] ,
    \top_I.branch[18].block[1].um_I.clk ,
    \top_I.branch[18].block[0].um_I.iw[17] ,
    \top_I.branch[18].block[0].um_I.iw[16] ,
    \top_I.branch[18].block[0].um_I.iw[15] ,
    \top_I.branch[18].block[0].um_I.iw[14] ,
    \top_I.branch[18].block[0].um_I.iw[13] ,
    \top_I.branch[18].block[0].um_I.iw[12] ,
    \top_I.branch[18].block[0].um_I.iw[11] ,
    \top_I.branch[18].block[0].um_I.iw[10] ,
    \top_I.branch[18].block[0].um_I.iw[9] ,
    \top_I.branch[18].block[0].um_I.iw[8] ,
    \top_I.branch[18].block[0].um_I.iw[7] ,
    \top_I.branch[18].block[0].um_I.iw[6] ,
    \top_I.branch[18].block[0].um_I.iw[5] ,
    \top_I.branch[18].block[0].um_I.iw[4] ,
    \top_I.branch[18].block[0].um_I.iw[3] ,
    \top_I.branch[18].block[0].um_I.iw[2] ,
    \top_I.branch[18].block[0].um_I.iw[1] ,
    \top_I.branch[18].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[15].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[14].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[13].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[12].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[11].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[10].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[9].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[8].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[7].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[6].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[5].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[4].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[3].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[2].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[1].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero ,
    \top_I.branch[18].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[18].block[15].um_I.pg_vdd ,
    \top_I.branch[18].block[14].um_I.pg_vdd ,
    \top_I.branch[18].block[13].um_I.pg_vdd ,
    \top_I.branch[18].block[12].um_I.pg_vdd ,
    \top_I.branch[18].block[11].um_I.pg_vdd ,
    \top_I.branch[18].block[10].um_I.pg_vdd ,
    \top_I.branch[18].block[9].um_I.pg_vdd ,
    \top_I.branch[18].block[8].um_I.pg_vdd ,
    \top_I.branch[18].block[7].um_I.pg_vdd ,
    \top_I.branch[18].block[6].um_I.pg_vdd ,
    \top_I.branch[18].block[5].um_I.pg_vdd ,
    \top_I.branch[18].block[4].um_I.pg_vdd ,
    \top_I.branch[18].block[3].um_I.pg_vdd ,
    \top_I.branch[18].block[2].um_I.pg_vdd ,
    \top_I.branch[18].block[1].um_I.pg_vdd ,
    \top_I.branch[18].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[19].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[19].l_addr[0] ),
    .k_zero(\top_I.branch[19].l_addr[1] ),
    .addr({\top_I.branch[19].l_addr[0] ,
    \top_I.branch[19].l_addr[1] ,
    \top_I.branch[19].l_addr[1] ,
    \top_I.branch[19].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[19].block[15].um_I.ena ,
    \top_I.branch[19].block[14].um_I.ena ,
    \top_I.branch[19].block[13].um_I.ena ,
    \top_I.branch[19].block[12].um_I.ena ,
    \top_I.branch[19].block[11].um_I.ena ,
    \top_I.branch[19].block[10].um_I.ena ,
    \top_I.branch[19].block[9].um_I.ena ,
    \top_I.branch[19].block[8].um_I.ena ,
    \top_I.branch[19].block[7].um_I.ena ,
    \top_I.branch[19].block[6].um_I.ena ,
    \top_I.branch[19].block[5].um_I.ena ,
    \top_I.branch[19].block[4].um_I.ena ,
    \top_I.branch[19].block[3].um_I.ena ,
    \top_I.branch[19].block[2].um_I.ena ,
    \top_I.branch[19].block[1].um_I.ena ,
    \top_I.branch[19].block[0].um_I.ena }),
    .um_iw({\top_I.branch[19].block[15].um_I.iw[17] ,
    \top_I.branch[19].block[15].um_I.iw[16] ,
    \top_I.branch[19].block[15].um_I.iw[15] ,
    \top_I.branch[19].block[15].um_I.iw[14] ,
    \top_I.branch[19].block[15].um_I.iw[13] ,
    \top_I.branch[19].block[15].um_I.iw[12] ,
    \top_I.branch[19].block[15].um_I.iw[11] ,
    \top_I.branch[19].block[15].um_I.iw[10] ,
    \top_I.branch[19].block[15].um_I.iw[9] ,
    \top_I.branch[19].block[15].um_I.iw[8] ,
    \top_I.branch[19].block[15].um_I.iw[7] ,
    \top_I.branch[19].block[15].um_I.iw[6] ,
    \top_I.branch[19].block[15].um_I.iw[5] ,
    \top_I.branch[19].block[15].um_I.iw[4] ,
    \top_I.branch[19].block[15].um_I.iw[3] ,
    \top_I.branch[19].block[15].um_I.iw[2] ,
    \top_I.branch[19].block[15].um_I.iw[1] ,
    \top_I.branch[19].block[15].um_I.clk ,
    \top_I.branch[19].block[14].um_I.iw[17] ,
    \top_I.branch[19].block[14].um_I.iw[16] ,
    \top_I.branch[19].block[14].um_I.iw[15] ,
    \top_I.branch[19].block[14].um_I.iw[14] ,
    \top_I.branch[19].block[14].um_I.iw[13] ,
    \top_I.branch[19].block[14].um_I.iw[12] ,
    \top_I.branch[19].block[14].um_I.iw[11] ,
    \top_I.branch[19].block[14].um_I.iw[10] ,
    \top_I.branch[19].block[14].um_I.iw[9] ,
    \top_I.branch[19].block[14].um_I.iw[8] ,
    \top_I.branch[19].block[14].um_I.iw[7] ,
    \top_I.branch[19].block[14].um_I.iw[6] ,
    \top_I.branch[19].block[14].um_I.iw[5] ,
    \top_I.branch[19].block[14].um_I.iw[4] ,
    \top_I.branch[19].block[14].um_I.iw[3] ,
    \top_I.branch[19].block[14].um_I.iw[2] ,
    \top_I.branch[19].block[14].um_I.iw[1] ,
    \top_I.branch[19].block[14].um_I.clk ,
    \top_I.branch[19].block[13].um_I.iw[17] ,
    \top_I.branch[19].block[13].um_I.iw[16] ,
    \top_I.branch[19].block[13].um_I.iw[15] ,
    \top_I.branch[19].block[13].um_I.iw[14] ,
    \top_I.branch[19].block[13].um_I.iw[13] ,
    \top_I.branch[19].block[13].um_I.iw[12] ,
    \top_I.branch[19].block[13].um_I.iw[11] ,
    \top_I.branch[19].block[13].um_I.iw[10] ,
    \top_I.branch[19].block[13].um_I.iw[9] ,
    \top_I.branch[19].block[13].um_I.iw[8] ,
    \top_I.branch[19].block[13].um_I.iw[7] ,
    \top_I.branch[19].block[13].um_I.iw[6] ,
    \top_I.branch[19].block[13].um_I.iw[5] ,
    \top_I.branch[19].block[13].um_I.iw[4] ,
    \top_I.branch[19].block[13].um_I.iw[3] ,
    \top_I.branch[19].block[13].um_I.iw[2] ,
    \top_I.branch[19].block[13].um_I.iw[1] ,
    \top_I.branch[19].block[13].um_I.clk ,
    \top_I.branch[19].block[12].um_I.iw[17] ,
    \top_I.branch[19].block[12].um_I.iw[16] ,
    \top_I.branch[19].block[12].um_I.iw[15] ,
    \top_I.branch[19].block[12].um_I.iw[14] ,
    \top_I.branch[19].block[12].um_I.iw[13] ,
    \top_I.branch[19].block[12].um_I.iw[12] ,
    \top_I.branch[19].block[12].um_I.iw[11] ,
    \top_I.branch[19].block[12].um_I.iw[10] ,
    \top_I.branch[19].block[12].um_I.iw[9] ,
    \top_I.branch[19].block[12].um_I.iw[8] ,
    \top_I.branch[19].block[12].um_I.iw[7] ,
    \top_I.branch[19].block[12].um_I.iw[6] ,
    \top_I.branch[19].block[12].um_I.iw[5] ,
    \top_I.branch[19].block[12].um_I.iw[4] ,
    \top_I.branch[19].block[12].um_I.iw[3] ,
    \top_I.branch[19].block[12].um_I.iw[2] ,
    \top_I.branch[19].block[12].um_I.iw[1] ,
    \top_I.branch[19].block[12].um_I.clk ,
    \top_I.branch[19].block[11].um_I.iw[17] ,
    \top_I.branch[19].block[11].um_I.iw[16] ,
    \top_I.branch[19].block[11].um_I.iw[15] ,
    \top_I.branch[19].block[11].um_I.iw[14] ,
    \top_I.branch[19].block[11].um_I.iw[13] ,
    \top_I.branch[19].block[11].um_I.iw[12] ,
    \top_I.branch[19].block[11].um_I.iw[11] ,
    \top_I.branch[19].block[11].um_I.iw[10] ,
    \top_I.branch[19].block[11].um_I.iw[9] ,
    \top_I.branch[19].block[11].um_I.iw[8] ,
    \top_I.branch[19].block[11].um_I.iw[7] ,
    \top_I.branch[19].block[11].um_I.iw[6] ,
    \top_I.branch[19].block[11].um_I.iw[5] ,
    \top_I.branch[19].block[11].um_I.iw[4] ,
    \top_I.branch[19].block[11].um_I.iw[3] ,
    \top_I.branch[19].block[11].um_I.iw[2] ,
    \top_I.branch[19].block[11].um_I.iw[1] ,
    \top_I.branch[19].block[11].um_I.clk ,
    \top_I.branch[19].block[10].um_I.iw[17] ,
    \top_I.branch[19].block[10].um_I.iw[16] ,
    \top_I.branch[19].block[10].um_I.iw[15] ,
    \top_I.branch[19].block[10].um_I.iw[14] ,
    \top_I.branch[19].block[10].um_I.iw[13] ,
    \top_I.branch[19].block[10].um_I.iw[12] ,
    \top_I.branch[19].block[10].um_I.iw[11] ,
    \top_I.branch[19].block[10].um_I.iw[10] ,
    \top_I.branch[19].block[10].um_I.iw[9] ,
    \top_I.branch[19].block[10].um_I.iw[8] ,
    \top_I.branch[19].block[10].um_I.iw[7] ,
    \top_I.branch[19].block[10].um_I.iw[6] ,
    \top_I.branch[19].block[10].um_I.iw[5] ,
    \top_I.branch[19].block[10].um_I.iw[4] ,
    \top_I.branch[19].block[10].um_I.iw[3] ,
    \top_I.branch[19].block[10].um_I.iw[2] ,
    \top_I.branch[19].block[10].um_I.iw[1] ,
    \top_I.branch[19].block[10].um_I.clk ,
    \top_I.branch[19].block[9].um_I.iw[17] ,
    \top_I.branch[19].block[9].um_I.iw[16] ,
    \top_I.branch[19].block[9].um_I.iw[15] ,
    \top_I.branch[19].block[9].um_I.iw[14] ,
    \top_I.branch[19].block[9].um_I.iw[13] ,
    \top_I.branch[19].block[9].um_I.iw[12] ,
    \top_I.branch[19].block[9].um_I.iw[11] ,
    \top_I.branch[19].block[9].um_I.iw[10] ,
    \top_I.branch[19].block[9].um_I.iw[9] ,
    \top_I.branch[19].block[9].um_I.iw[8] ,
    \top_I.branch[19].block[9].um_I.iw[7] ,
    \top_I.branch[19].block[9].um_I.iw[6] ,
    \top_I.branch[19].block[9].um_I.iw[5] ,
    \top_I.branch[19].block[9].um_I.iw[4] ,
    \top_I.branch[19].block[9].um_I.iw[3] ,
    \top_I.branch[19].block[9].um_I.iw[2] ,
    \top_I.branch[19].block[9].um_I.iw[1] ,
    \top_I.branch[19].block[9].um_I.clk ,
    \top_I.branch[19].block[8].um_I.iw[17] ,
    \top_I.branch[19].block[8].um_I.iw[16] ,
    \top_I.branch[19].block[8].um_I.iw[15] ,
    \top_I.branch[19].block[8].um_I.iw[14] ,
    \top_I.branch[19].block[8].um_I.iw[13] ,
    \top_I.branch[19].block[8].um_I.iw[12] ,
    \top_I.branch[19].block[8].um_I.iw[11] ,
    \top_I.branch[19].block[8].um_I.iw[10] ,
    \top_I.branch[19].block[8].um_I.iw[9] ,
    \top_I.branch[19].block[8].um_I.iw[8] ,
    \top_I.branch[19].block[8].um_I.iw[7] ,
    \top_I.branch[19].block[8].um_I.iw[6] ,
    \top_I.branch[19].block[8].um_I.iw[5] ,
    \top_I.branch[19].block[8].um_I.iw[4] ,
    \top_I.branch[19].block[8].um_I.iw[3] ,
    \top_I.branch[19].block[8].um_I.iw[2] ,
    \top_I.branch[19].block[8].um_I.iw[1] ,
    \top_I.branch[19].block[8].um_I.clk ,
    \top_I.branch[19].block[7].um_I.iw[17] ,
    \top_I.branch[19].block[7].um_I.iw[16] ,
    \top_I.branch[19].block[7].um_I.iw[15] ,
    \top_I.branch[19].block[7].um_I.iw[14] ,
    \top_I.branch[19].block[7].um_I.iw[13] ,
    \top_I.branch[19].block[7].um_I.iw[12] ,
    \top_I.branch[19].block[7].um_I.iw[11] ,
    \top_I.branch[19].block[7].um_I.iw[10] ,
    \top_I.branch[19].block[7].um_I.iw[9] ,
    \top_I.branch[19].block[7].um_I.iw[8] ,
    \top_I.branch[19].block[7].um_I.iw[7] ,
    \top_I.branch[19].block[7].um_I.iw[6] ,
    \top_I.branch[19].block[7].um_I.iw[5] ,
    \top_I.branch[19].block[7].um_I.iw[4] ,
    \top_I.branch[19].block[7].um_I.iw[3] ,
    \top_I.branch[19].block[7].um_I.iw[2] ,
    \top_I.branch[19].block[7].um_I.iw[1] ,
    \top_I.branch[19].block[7].um_I.clk ,
    \top_I.branch[19].block[6].um_I.iw[17] ,
    \top_I.branch[19].block[6].um_I.iw[16] ,
    \top_I.branch[19].block[6].um_I.iw[15] ,
    \top_I.branch[19].block[6].um_I.iw[14] ,
    \top_I.branch[19].block[6].um_I.iw[13] ,
    \top_I.branch[19].block[6].um_I.iw[12] ,
    \top_I.branch[19].block[6].um_I.iw[11] ,
    \top_I.branch[19].block[6].um_I.iw[10] ,
    \top_I.branch[19].block[6].um_I.iw[9] ,
    \top_I.branch[19].block[6].um_I.iw[8] ,
    \top_I.branch[19].block[6].um_I.iw[7] ,
    \top_I.branch[19].block[6].um_I.iw[6] ,
    \top_I.branch[19].block[6].um_I.iw[5] ,
    \top_I.branch[19].block[6].um_I.iw[4] ,
    \top_I.branch[19].block[6].um_I.iw[3] ,
    \top_I.branch[19].block[6].um_I.iw[2] ,
    \top_I.branch[19].block[6].um_I.iw[1] ,
    \top_I.branch[19].block[6].um_I.clk ,
    \top_I.branch[19].block[5].um_I.iw[17] ,
    \top_I.branch[19].block[5].um_I.iw[16] ,
    \top_I.branch[19].block[5].um_I.iw[15] ,
    \top_I.branch[19].block[5].um_I.iw[14] ,
    \top_I.branch[19].block[5].um_I.iw[13] ,
    \top_I.branch[19].block[5].um_I.iw[12] ,
    \top_I.branch[19].block[5].um_I.iw[11] ,
    \top_I.branch[19].block[5].um_I.iw[10] ,
    \top_I.branch[19].block[5].um_I.iw[9] ,
    \top_I.branch[19].block[5].um_I.iw[8] ,
    \top_I.branch[19].block[5].um_I.iw[7] ,
    \top_I.branch[19].block[5].um_I.iw[6] ,
    \top_I.branch[19].block[5].um_I.iw[5] ,
    \top_I.branch[19].block[5].um_I.iw[4] ,
    \top_I.branch[19].block[5].um_I.iw[3] ,
    \top_I.branch[19].block[5].um_I.iw[2] ,
    \top_I.branch[19].block[5].um_I.iw[1] ,
    \top_I.branch[19].block[5].um_I.clk ,
    \top_I.branch[19].block[4].um_I.iw[17] ,
    \top_I.branch[19].block[4].um_I.iw[16] ,
    \top_I.branch[19].block[4].um_I.iw[15] ,
    \top_I.branch[19].block[4].um_I.iw[14] ,
    \top_I.branch[19].block[4].um_I.iw[13] ,
    \top_I.branch[19].block[4].um_I.iw[12] ,
    \top_I.branch[19].block[4].um_I.iw[11] ,
    \top_I.branch[19].block[4].um_I.iw[10] ,
    \top_I.branch[19].block[4].um_I.iw[9] ,
    \top_I.branch[19].block[4].um_I.iw[8] ,
    \top_I.branch[19].block[4].um_I.iw[7] ,
    \top_I.branch[19].block[4].um_I.iw[6] ,
    \top_I.branch[19].block[4].um_I.iw[5] ,
    \top_I.branch[19].block[4].um_I.iw[4] ,
    \top_I.branch[19].block[4].um_I.iw[3] ,
    \top_I.branch[19].block[4].um_I.iw[2] ,
    \top_I.branch[19].block[4].um_I.iw[1] ,
    \top_I.branch[19].block[4].um_I.clk ,
    \top_I.branch[19].block[3].um_I.iw[17] ,
    \top_I.branch[19].block[3].um_I.iw[16] ,
    \top_I.branch[19].block[3].um_I.iw[15] ,
    \top_I.branch[19].block[3].um_I.iw[14] ,
    \top_I.branch[19].block[3].um_I.iw[13] ,
    \top_I.branch[19].block[3].um_I.iw[12] ,
    \top_I.branch[19].block[3].um_I.iw[11] ,
    \top_I.branch[19].block[3].um_I.iw[10] ,
    \top_I.branch[19].block[3].um_I.iw[9] ,
    \top_I.branch[19].block[3].um_I.iw[8] ,
    \top_I.branch[19].block[3].um_I.iw[7] ,
    \top_I.branch[19].block[3].um_I.iw[6] ,
    \top_I.branch[19].block[3].um_I.iw[5] ,
    \top_I.branch[19].block[3].um_I.iw[4] ,
    \top_I.branch[19].block[3].um_I.iw[3] ,
    \top_I.branch[19].block[3].um_I.iw[2] ,
    \top_I.branch[19].block[3].um_I.iw[1] ,
    \top_I.branch[19].block[3].um_I.clk ,
    \top_I.branch[19].block[2].um_I.iw[17] ,
    \top_I.branch[19].block[2].um_I.iw[16] ,
    \top_I.branch[19].block[2].um_I.iw[15] ,
    \top_I.branch[19].block[2].um_I.iw[14] ,
    \top_I.branch[19].block[2].um_I.iw[13] ,
    \top_I.branch[19].block[2].um_I.iw[12] ,
    \top_I.branch[19].block[2].um_I.iw[11] ,
    \top_I.branch[19].block[2].um_I.iw[10] ,
    \top_I.branch[19].block[2].um_I.iw[9] ,
    \top_I.branch[19].block[2].um_I.iw[8] ,
    \top_I.branch[19].block[2].um_I.iw[7] ,
    \top_I.branch[19].block[2].um_I.iw[6] ,
    \top_I.branch[19].block[2].um_I.iw[5] ,
    \top_I.branch[19].block[2].um_I.iw[4] ,
    \top_I.branch[19].block[2].um_I.iw[3] ,
    \top_I.branch[19].block[2].um_I.iw[2] ,
    \top_I.branch[19].block[2].um_I.iw[1] ,
    \top_I.branch[19].block[2].um_I.clk ,
    \top_I.branch[19].block[1].um_I.iw[17] ,
    \top_I.branch[19].block[1].um_I.iw[16] ,
    \top_I.branch[19].block[1].um_I.iw[15] ,
    \top_I.branch[19].block[1].um_I.iw[14] ,
    \top_I.branch[19].block[1].um_I.iw[13] ,
    \top_I.branch[19].block[1].um_I.iw[12] ,
    \top_I.branch[19].block[1].um_I.iw[11] ,
    \top_I.branch[19].block[1].um_I.iw[10] ,
    \top_I.branch[19].block[1].um_I.iw[9] ,
    \top_I.branch[19].block[1].um_I.iw[8] ,
    \top_I.branch[19].block[1].um_I.iw[7] ,
    \top_I.branch[19].block[1].um_I.iw[6] ,
    \top_I.branch[19].block[1].um_I.iw[5] ,
    \top_I.branch[19].block[1].um_I.iw[4] ,
    \top_I.branch[19].block[1].um_I.iw[3] ,
    \top_I.branch[19].block[1].um_I.iw[2] ,
    \top_I.branch[19].block[1].um_I.iw[1] ,
    \top_I.branch[19].block[1].um_I.clk ,
    \top_I.branch[19].block[0].um_I.iw[17] ,
    \top_I.branch[19].block[0].um_I.iw[16] ,
    \top_I.branch[19].block[0].um_I.iw[15] ,
    \top_I.branch[19].block[0].um_I.iw[14] ,
    \top_I.branch[19].block[0].um_I.iw[13] ,
    \top_I.branch[19].block[0].um_I.iw[12] ,
    \top_I.branch[19].block[0].um_I.iw[11] ,
    \top_I.branch[19].block[0].um_I.iw[10] ,
    \top_I.branch[19].block[0].um_I.iw[9] ,
    \top_I.branch[19].block[0].um_I.iw[8] ,
    \top_I.branch[19].block[0].um_I.iw[7] ,
    \top_I.branch[19].block[0].um_I.iw[6] ,
    \top_I.branch[19].block[0].um_I.iw[5] ,
    \top_I.branch[19].block[0].um_I.iw[4] ,
    \top_I.branch[19].block[0].um_I.iw[3] ,
    \top_I.branch[19].block[0].um_I.iw[2] ,
    \top_I.branch[19].block[0].um_I.iw[1] ,
    \top_I.branch[19].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[15].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[14].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[13].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[12].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[11].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[10].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[9].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[8].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[7].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[6].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[5].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[4].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[3].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[2].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[1].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero ,
    \top_I.branch[19].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[19].block[15].um_I.pg_vdd ,
    \top_I.branch[19].block[14].um_I.pg_vdd ,
    \top_I.branch[19].block[13].um_I.pg_vdd ,
    \top_I.branch[19].block[12].um_I.pg_vdd ,
    \top_I.branch[19].block[11].um_I.pg_vdd ,
    \top_I.branch[19].block[10].um_I.pg_vdd ,
    \top_I.branch[19].block[9].um_I.pg_vdd ,
    \top_I.branch[19].block[8].um_I.pg_vdd ,
    \top_I.branch[19].block[7].um_I.pg_vdd ,
    \top_I.branch[19].block[6].um_I.pg_vdd ,
    \top_I.branch[19].block[5].um_I.pg_vdd ,
    \top_I.branch[19].block[4].um_I.pg_vdd ,
    \top_I.branch[19].block[3].um_I.pg_vdd ,
    \top_I.branch[19].block[2].um_I.pg_vdd ,
    \top_I.branch[19].block[1].um_I.pg_vdd ,
    \top_I.branch[19].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[1].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[1].l_k_one ),
    .k_zero(\top_I.branch[1].l_addr[0] ),
    .addr({\top_I.branch[1].l_addr[0] ,
    \top_I.branch[1].l_addr[0] ,
    \top_I.branch[1].l_addr[0] ,
    \top_I.branch[1].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[1].block[15].um_I.ena ,
    \top_I.branch[1].block[14].um_I.ena ,
    \top_I.branch[1].block[13].um_I.ena ,
    \top_I.branch[1].block[12].um_I.ena ,
    \top_I.branch[1].block[11].um_I.ena ,
    \top_I.branch[1].block[10].um_I.ena ,
    \top_I.branch[1].block[9].um_I.ena ,
    \top_I.branch[1].block[8].um_I.ena ,
    \top_I.branch[1].block[7].um_I.ena ,
    \top_I.branch[1].block[6].um_I.ena ,
    \top_I.branch[1].block[5].um_I.ena ,
    \top_I.branch[1].block[4].um_I.ena ,
    \top_I.branch[1].block[3].um_I.ena ,
    \top_I.branch[1].block[2].um_I.ena ,
    \top_I.branch[1].block[1].um_I.ena ,
    \top_I.branch[1].block[0].um_I.ena }),
    .um_iw({\top_I.branch[1].block[15].um_I.iw[17] ,
    \top_I.branch[1].block[15].um_I.iw[16] ,
    \top_I.branch[1].block[15].um_I.iw[15] ,
    \top_I.branch[1].block[15].um_I.iw[14] ,
    \top_I.branch[1].block[15].um_I.iw[13] ,
    \top_I.branch[1].block[15].um_I.iw[12] ,
    \top_I.branch[1].block[15].um_I.iw[11] ,
    \top_I.branch[1].block[15].um_I.iw[10] ,
    \top_I.branch[1].block[15].um_I.iw[9] ,
    \top_I.branch[1].block[15].um_I.iw[8] ,
    \top_I.branch[1].block[15].um_I.iw[7] ,
    \top_I.branch[1].block[15].um_I.iw[6] ,
    \top_I.branch[1].block[15].um_I.iw[5] ,
    \top_I.branch[1].block[15].um_I.iw[4] ,
    \top_I.branch[1].block[15].um_I.iw[3] ,
    \top_I.branch[1].block[15].um_I.iw[2] ,
    \top_I.branch[1].block[15].um_I.iw[1] ,
    \top_I.branch[1].block[15].um_I.clk ,
    \top_I.branch[1].block[14].um_I.iw[17] ,
    \top_I.branch[1].block[14].um_I.iw[16] ,
    \top_I.branch[1].block[14].um_I.iw[15] ,
    \top_I.branch[1].block[14].um_I.iw[14] ,
    \top_I.branch[1].block[14].um_I.iw[13] ,
    \top_I.branch[1].block[14].um_I.iw[12] ,
    \top_I.branch[1].block[14].um_I.iw[11] ,
    \top_I.branch[1].block[14].um_I.iw[10] ,
    \top_I.branch[1].block[14].um_I.iw[9] ,
    \top_I.branch[1].block[14].um_I.iw[8] ,
    \top_I.branch[1].block[14].um_I.iw[7] ,
    \top_I.branch[1].block[14].um_I.iw[6] ,
    \top_I.branch[1].block[14].um_I.iw[5] ,
    \top_I.branch[1].block[14].um_I.iw[4] ,
    \top_I.branch[1].block[14].um_I.iw[3] ,
    \top_I.branch[1].block[14].um_I.iw[2] ,
    \top_I.branch[1].block[14].um_I.iw[1] ,
    \top_I.branch[1].block[14].um_I.clk ,
    \top_I.branch[1].block[13].um_I.iw[17] ,
    \top_I.branch[1].block[13].um_I.iw[16] ,
    \top_I.branch[1].block[13].um_I.iw[15] ,
    \top_I.branch[1].block[13].um_I.iw[14] ,
    \top_I.branch[1].block[13].um_I.iw[13] ,
    \top_I.branch[1].block[13].um_I.iw[12] ,
    \top_I.branch[1].block[13].um_I.iw[11] ,
    \top_I.branch[1].block[13].um_I.iw[10] ,
    \top_I.branch[1].block[13].um_I.iw[9] ,
    \top_I.branch[1].block[13].um_I.iw[8] ,
    \top_I.branch[1].block[13].um_I.iw[7] ,
    \top_I.branch[1].block[13].um_I.iw[6] ,
    \top_I.branch[1].block[13].um_I.iw[5] ,
    \top_I.branch[1].block[13].um_I.iw[4] ,
    \top_I.branch[1].block[13].um_I.iw[3] ,
    \top_I.branch[1].block[13].um_I.iw[2] ,
    \top_I.branch[1].block[13].um_I.iw[1] ,
    \top_I.branch[1].block[13].um_I.clk ,
    \top_I.branch[1].block[12].um_I.iw[17] ,
    \top_I.branch[1].block[12].um_I.iw[16] ,
    \top_I.branch[1].block[12].um_I.iw[15] ,
    \top_I.branch[1].block[12].um_I.iw[14] ,
    \top_I.branch[1].block[12].um_I.iw[13] ,
    \top_I.branch[1].block[12].um_I.iw[12] ,
    \top_I.branch[1].block[12].um_I.iw[11] ,
    \top_I.branch[1].block[12].um_I.iw[10] ,
    \top_I.branch[1].block[12].um_I.iw[9] ,
    \top_I.branch[1].block[12].um_I.iw[8] ,
    \top_I.branch[1].block[12].um_I.iw[7] ,
    \top_I.branch[1].block[12].um_I.iw[6] ,
    \top_I.branch[1].block[12].um_I.iw[5] ,
    \top_I.branch[1].block[12].um_I.iw[4] ,
    \top_I.branch[1].block[12].um_I.iw[3] ,
    \top_I.branch[1].block[12].um_I.iw[2] ,
    \top_I.branch[1].block[12].um_I.iw[1] ,
    \top_I.branch[1].block[12].um_I.clk ,
    \top_I.branch[1].block[11].um_I.iw[17] ,
    \top_I.branch[1].block[11].um_I.iw[16] ,
    \top_I.branch[1].block[11].um_I.iw[15] ,
    \top_I.branch[1].block[11].um_I.iw[14] ,
    \top_I.branch[1].block[11].um_I.iw[13] ,
    \top_I.branch[1].block[11].um_I.iw[12] ,
    \top_I.branch[1].block[11].um_I.iw[11] ,
    \top_I.branch[1].block[11].um_I.iw[10] ,
    \top_I.branch[1].block[11].um_I.iw[9] ,
    \top_I.branch[1].block[11].um_I.iw[8] ,
    \top_I.branch[1].block[11].um_I.iw[7] ,
    \top_I.branch[1].block[11].um_I.iw[6] ,
    \top_I.branch[1].block[11].um_I.iw[5] ,
    \top_I.branch[1].block[11].um_I.iw[4] ,
    \top_I.branch[1].block[11].um_I.iw[3] ,
    \top_I.branch[1].block[11].um_I.iw[2] ,
    \top_I.branch[1].block[11].um_I.iw[1] ,
    \top_I.branch[1].block[11].um_I.clk ,
    \top_I.branch[1].block[10].um_I.iw[17] ,
    \top_I.branch[1].block[10].um_I.iw[16] ,
    \top_I.branch[1].block[10].um_I.iw[15] ,
    \top_I.branch[1].block[10].um_I.iw[14] ,
    \top_I.branch[1].block[10].um_I.iw[13] ,
    \top_I.branch[1].block[10].um_I.iw[12] ,
    \top_I.branch[1].block[10].um_I.iw[11] ,
    \top_I.branch[1].block[10].um_I.iw[10] ,
    \top_I.branch[1].block[10].um_I.iw[9] ,
    \top_I.branch[1].block[10].um_I.iw[8] ,
    \top_I.branch[1].block[10].um_I.iw[7] ,
    \top_I.branch[1].block[10].um_I.iw[6] ,
    \top_I.branch[1].block[10].um_I.iw[5] ,
    \top_I.branch[1].block[10].um_I.iw[4] ,
    \top_I.branch[1].block[10].um_I.iw[3] ,
    \top_I.branch[1].block[10].um_I.iw[2] ,
    \top_I.branch[1].block[10].um_I.iw[1] ,
    \top_I.branch[1].block[10].um_I.clk ,
    \top_I.branch[1].block[9].um_I.iw[17] ,
    \top_I.branch[1].block[9].um_I.iw[16] ,
    \top_I.branch[1].block[9].um_I.iw[15] ,
    \top_I.branch[1].block[9].um_I.iw[14] ,
    \top_I.branch[1].block[9].um_I.iw[13] ,
    \top_I.branch[1].block[9].um_I.iw[12] ,
    \top_I.branch[1].block[9].um_I.iw[11] ,
    \top_I.branch[1].block[9].um_I.iw[10] ,
    \top_I.branch[1].block[9].um_I.iw[9] ,
    \top_I.branch[1].block[9].um_I.iw[8] ,
    \top_I.branch[1].block[9].um_I.iw[7] ,
    \top_I.branch[1].block[9].um_I.iw[6] ,
    \top_I.branch[1].block[9].um_I.iw[5] ,
    \top_I.branch[1].block[9].um_I.iw[4] ,
    \top_I.branch[1].block[9].um_I.iw[3] ,
    \top_I.branch[1].block[9].um_I.iw[2] ,
    \top_I.branch[1].block[9].um_I.iw[1] ,
    \top_I.branch[1].block[9].um_I.clk ,
    \top_I.branch[1].block[8].um_I.iw[17] ,
    \top_I.branch[1].block[8].um_I.iw[16] ,
    \top_I.branch[1].block[8].um_I.iw[15] ,
    \top_I.branch[1].block[8].um_I.iw[14] ,
    \top_I.branch[1].block[8].um_I.iw[13] ,
    \top_I.branch[1].block[8].um_I.iw[12] ,
    \top_I.branch[1].block[8].um_I.iw[11] ,
    \top_I.branch[1].block[8].um_I.iw[10] ,
    \top_I.branch[1].block[8].um_I.iw[9] ,
    \top_I.branch[1].block[8].um_I.iw[8] ,
    \top_I.branch[1].block[8].um_I.iw[7] ,
    \top_I.branch[1].block[8].um_I.iw[6] ,
    \top_I.branch[1].block[8].um_I.iw[5] ,
    \top_I.branch[1].block[8].um_I.iw[4] ,
    \top_I.branch[1].block[8].um_I.iw[3] ,
    \top_I.branch[1].block[8].um_I.iw[2] ,
    \top_I.branch[1].block[8].um_I.iw[1] ,
    \top_I.branch[1].block[8].um_I.clk ,
    \top_I.branch[1].block[7].um_I.iw[17] ,
    \top_I.branch[1].block[7].um_I.iw[16] ,
    \top_I.branch[1].block[7].um_I.iw[15] ,
    \top_I.branch[1].block[7].um_I.iw[14] ,
    \top_I.branch[1].block[7].um_I.iw[13] ,
    \top_I.branch[1].block[7].um_I.iw[12] ,
    \top_I.branch[1].block[7].um_I.iw[11] ,
    \top_I.branch[1].block[7].um_I.iw[10] ,
    \top_I.branch[1].block[7].um_I.iw[9] ,
    \top_I.branch[1].block[7].um_I.iw[8] ,
    \top_I.branch[1].block[7].um_I.iw[7] ,
    \top_I.branch[1].block[7].um_I.iw[6] ,
    \top_I.branch[1].block[7].um_I.iw[5] ,
    \top_I.branch[1].block[7].um_I.iw[4] ,
    \top_I.branch[1].block[7].um_I.iw[3] ,
    \top_I.branch[1].block[7].um_I.iw[2] ,
    \top_I.branch[1].block[7].um_I.iw[1] ,
    \top_I.branch[1].block[7].um_I.clk ,
    \top_I.branch[1].block[6].um_I.iw[17] ,
    \top_I.branch[1].block[6].um_I.iw[16] ,
    \top_I.branch[1].block[6].um_I.iw[15] ,
    \top_I.branch[1].block[6].um_I.iw[14] ,
    \top_I.branch[1].block[6].um_I.iw[13] ,
    \top_I.branch[1].block[6].um_I.iw[12] ,
    \top_I.branch[1].block[6].um_I.iw[11] ,
    \top_I.branch[1].block[6].um_I.iw[10] ,
    \top_I.branch[1].block[6].um_I.iw[9] ,
    \top_I.branch[1].block[6].um_I.iw[8] ,
    \top_I.branch[1].block[6].um_I.iw[7] ,
    \top_I.branch[1].block[6].um_I.iw[6] ,
    \top_I.branch[1].block[6].um_I.iw[5] ,
    \top_I.branch[1].block[6].um_I.iw[4] ,
    \top_I.branch[1].block[6].um_I.iw[3] ,
    \top_I.branch[1].block[6].um_I.iw[2] ,
    \top_I.branch[1].block[6].um_I.iw[1] ,
    \top_I.branch[1].block[6].um_I.clk ,
    \top_I.branch[1].block[5].um_I.iw[17] ,
    \top_I.branch[1].block[5].um_I.iw[16] ,
    \top_I.branch[1].block[5].um_I.iw[15] ,
    \top_I.branch[1].block[5].um_I.iw[14] ,
    \top_I.branch[1].block[5].um_I.iw[13] ,
    \top_I.branch[1].block[5].um_I.iw[12] ,
    \top_I.branch[1].block[5].um_I.iw[11] ,
    \top_I.branch[1].block[5].um_I.iw[10] ,
    \top_I.branch[1].block[5].um_I.iw[9] ,
    \top_I.branch[1].block[5].um_I.iw[8] ,
    \top_I.branch[1].block[5].um_I.iw[7] ,
    \top_I.branch[1].block[5].um_I.iw[6] ,
    \top_I.branch[1].block[5].um_I.iw[5] ,
    \top_I.branch[1].block[5].um_I.iw[4] ,
    \top_I.branch[1].block[5].um_I.iw[3] ,
    \top_I.branch[1].block[5].um_I.iw[2] ,
    \top_I.branch[1].block[5].um_I.iw[1] ,
    \top_I.branch[1].block[5].um_I.clk ,
    \top_I.branch[1].block[4].um_I.iw[17] ,
    \top_I.branch[1].block[4].um_I.iw[16] ,
    \top_I.branch[1].block[4].um_I.iw[15] ,
    \top_I.branch[1].block[4].um_I.iw[14] ,
    \top_I.branch[1].block[4].um_I.iw[13] ,
    \top_I.branch[1].block[4].um_I.iw[12] ,
    \top_I.branch[1].block[4].um_I.iw[11] ,
    \top_I.branch[1].block[4].um_I.iw[10] ,
    \top_I.branch[1].block[4].um_I.iw[9] ,
    \top_I.branch[1].block[4].um_I.iw[8] ,
    \top_I.branch[1].block[4].um_I.iw[7] ,
    \top_I.branch[1].block[4].um_I.iw[6] ,
    \top_I.branch[1].block[4].um_I.iw[5] ,
    \top_I.branch[1].block[4].um_I.iw[4] ,
    \top_I.branch[1].block[4].um_I.iw[3] ,
    \top_I.branch[1].block[4].um_I.iw[2] ,
    \top_I.branch[1].block[4].um_I.iw[1] ,
    \top_I.branch[1].block[4].um_I.clk ,
    \top_I.branch[1].block[3].um_I.iw[17] ,
    \top_I.branch[1].block[3].um_I.iw[16] ,
    \top_I.branch[1].block[3].um_I.iw[15] ,
    \top_I.branch[1].block[3].um_I.iw[14] ,
    \top_I.branch[1].block[3].um_I.iw[13] ,
    \top_I.branch[1].block[3].um_I.iw[12] ,
    \top_I.branch[1].block[3].um_I.iw[11] ,
    \top_I.branch[1].block[3].um_I.iw[10] ,
    \top_I.branch[1].block[3].um_I.iw[9] ,
    \top_I.branch[1].block[3].um_I.iw[8] ,
    \top_I.branch[1].block[3].um_I.iw[7] ,
    \top_I.branch[1].block[3].um_I.iw[6] ,
    \top_I.branch[1].block[3].um_I.iw[5] ,
    \top_I.branch[1].block[3].um_I.iw[4] ,
    \top_I.branch[1].block[3].um_I.iw[3] ,
    \top_I.branch[1].block[3].um_I.iw[2] ,
    \top_I.branch[1].block[3].um_I.iw[1] ,
    \top_I.branch[1].block[3].um_I.clk ,
    \top_I.branch[1].block[2].um_I.iw[17] ,
    \top_I.branch[1].block[2].um_I.iw[16] ,
    \top_I.branch[1].block[2].um_I.iw[15] ,
    \top_I.branch[1].block[2].um_I.iw[14] ,
    \top_I.branch[1].block[2].um_I.iw[13] ,
    \top_I.branch[1].block[2].um_I.iw[12] ,
    \top_I.branch[1].block[2].um_I.iw[11] ,
    \top_I.branch[1].block[2].um_I.iw[10] ,
    \top_I.branch[1].block[2].um_I.iw[9] ,
    \top_I.branch[1].block[2].um_I.iw[8] ,
    \top_I.branch[1].block[2].um_I.iw[7] ,
    \top_I.branch[1].block[2].um_I.iw[6] ,
    \top_I.branch[1].block[2].um_I.iw[5] ,
    \top_I.branch[1].block[2].um_I.iw[4] ,
    \top_I.branch[1].block[2].um_I.iw[3] ,
    \top_I.branch[1].block[2].um_I.iw[2] ,
    \top_I.branch[1].block[2].um_I.iw[1] ,
    \top_I.branch[1].block[2].um_I.clk ,
    \top_I.branch[1].block[1].um_I.iw[17] ,
    \top_I.branch[1].block[1].um_I.iw[16] ,
    \top_I.branch[1].block[1].um_I.iw[15] ,
    \top_I.branch[1].block[1].um_I.iw[14] ,
    \top_I.branch[1].block[1].um_I.iw[13] ,
    \top_I.branch[1].block[1].um_I.iw[12] ,
    \top_I.branch[1].block[1].um_I.iw[11] ,
    \top_I.branch[1].block[1].um_I.iw[10] ,
    \top_I.branch[1].block[1].um_I.iw[9] ,
    \top_I.branch[1].block[1].um_I.iw[8] ,
    \top_I.branch[1].block[1].um_I.iw[7] ,
    \top_I.branch[1].block[1].um_I.iw[6] ,
    \top_I.branch[1].block[1].um_I.iw[5] ,
    \top_I.branch[1].block[1].um_I.iw[4] ,
    \top_I.branch[1].block[1].um_I.iw[3] ,
    \top_I.branch[1].block[1].um_I.iw[2] ,
    \top_I.branch[1].block[1].um_I.iw[1] ,
    \top_I.branch[1].block[1].um_I.clk ,
    \top_I.branch[1].block[0].um_I.iw[17] ,
    \top_I.branch[1].block[0].um_I.iw[16] ,
    \top_I.branch[1].block[0].um_I.iw[15] ,
    \top_I.branch[1].block[0].um_I.iw[14] ,
    \top_I.branch[1].block[0].um_I.iw[13] ,
    \top_I.branch[1].block[0].um_I.iw[12] ,
    \top_I.branch[1].block[0].um_I.iw[11] ,
    \top_I.branch[1].block[0].um_I.iw[10] ,
    \top_I.branch[1].block[0].um_I.iw[9] ,
    \top_I.branch[1].block[0].um_I.iw[8] ,
    \top_I.branch[1].block[0].um_I.iw[7] ,
    \top_I.branch[1].block[0].um_I.iw[6] ,
    \top_I.branch[1].block[0].um_I.iw[5] ,
    \top_I.branch[1].block[0].um_I.iw[4] ,
    \top_I.branch[1].block[0].um_I.iw[3] ,
    \top_I.branch[1].block[0].um_I.iw[2] ,
    \top_I.branch[1].block[0].um_I.iw[1] ,
    \top_I.branch[1].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[15].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[14].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[13].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[12].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[11].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[10].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[9].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[8].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[7].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[6].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[5].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[4].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[3].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[2].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[1].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero ,
    \top_I.branch[1].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[1].block[15].um_I.pg_vdd ,
    \top_I.branch[1].block[14].um_I.pg_vdd ,
    \top_I.branch[1].block[13].um_I.pg_vdd ,
    \top_I.branch[1].block[12].um_I.pg_vdd ,
    \top_I.branch[1].block[11].um_I.pg_vdd ,
    \top_I.branch[1].block[10].um_I.pg_vdd ,
    \top_I.branch[1].block[9].um_I.pg_vdd ,
    \top_I.branch[1].block[8].um_I.pg_vdd ,
    \top_I.branch[1].block[7].um_I.pg_vdd ,
    \top_I.branch[1].block[6].um_I.pg_vdd ,
    \top_I.branch[1].block[5].um_I.pg_vdd ,
    \top_I.branch[1].block[4].um_I.pg_vdd ,
    \top_I.branch[1].block[3].um_I.pg_vdd ,
    \top_I.branch[1].block[2].um_I.pg_vdd ,
    \top_I.branch[1].block[1].um_I.pg_vdd ,
    \top_I.branch[1].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[20].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[20].l_addr[1] ),
    .k_zero(\top_I.branch[20].l_addr[0] ),
    .addr({\top_I.branch[20].l_addr[1] ,
    \top_I.branch[20].l_addr[0] ,
    \top_I.branch[20].l_addr[1] ,
    \top_I.branch[20].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[20].block[15].um_I.ena ,
    \top_I.branch[20].block[14].um_I.ena ,
    \top_I.branch[20].block[13].um_I.ena ,
    \top_I.branch[20].block[12].um_I.ena ,
    \top_I.branch[20].block[11].um_I.ena ,
    \top_I.branch[20].block[10].um_I.ena ,
    \top_I.branch[20].block[9].um_I.ena ,
    \top_I.branch[20].block[8].um_I.ena ,
    \top_I.branch[20].block[7].um_I.ena ,
    \top_I.branch[20].block[6].um_I.ena ,
    \top_I.branch[20].block[5].um_I.ena ,
    \top_I.branch[20].block[4].um_I.ena ,
    \top_I.branch[20].block[3].um_I.ena ,
    \top_I.branch[20].block[2].um_I.ena ,
    \top_I.branch[20].block[1].um_I.ena ,
    \top_I.branch[20].block[0].um_I.ena }),
    .um_iw({\top_I.branch[20].block[15].um_I.iw[17] ,
    \top_I.branch[20].block[15].um_I.iw[16] ,
    \top_I.branch[20].block[15].um_I.iw[15] ,
    \top_I.branch[20].block[15].um_I.iw[14] ,
    \top_I.branch[20].block[15].um_I.iw[13] ,
    \top_I.branch[20].block[15].um_I.iw[12] ,
    \top_I.branch[20].block[15].um_I.iw[11] ,
    \top_I.branch[20].block[15].um_I.iw[10] ,
    \top_I.branch[20].block[15].um_I.iw[9] ,
    \top_I.branch[20].block[15].um_I.iw[8] ,
    \top_I.branch[20].block[15].um_I.iw[7] ,
    \top_I.branch[20].block[15].um_I.iw[6] ,
    \top_I.branch[20].block[15].um_I.iw[5] ,
    \top_I.branch[20].block[15].um_I.iw[4] ,
    \top_I.branch[20].block[15].um_I.iw[3] ,
    \top_I.branch[20].block[15].um_I.iw[2] ,
    \top_I.branch[20].block[15].um_I.iw[1] ,
    \top_I.branch[20].block[15].um_I.clk ,
    \top_I.branch[20].block[14].um_I.iw[17] ,
    \top_I.branch[20].block[14].um_I.iw[16] ,
    \top_I.branch[20].block[14].um_I.iw[15] ,
    \top_I.branch[20].block[14].um_I.iw[14] ,
    \top_I.branch[20].block[14].um_I.iw[13] ,
    \top_I.branch[20].block[14].um_I.iw[12] ,
    \top_I.branch[20].block[14].um_I.iw[11] ,
    \top_I.branch[20].block[14].um_I.iw[10] ,
    \top_I.branch[20].block[14].um_I.iw[9] ,
    \top_I.branch[20].block[14].um_I.iw[8] ,
    \top_I.branch[20].block[14].um_I.iw[7] ,
    \top_I.branch[20].block[14].um_I.iw[6] ,
    \top_I.branch[20].block[14].um_I.iw[5] ,
    \top_I.branch[20].block[14].um_I.iw[4] ,
    \top_I.branch[20].block[14].um_I.iw[3] ,
    \top_I.branch[20].block[14].um_I.iw[2] ,
    \top_I.branch[20].block[14].um_I.iw[1] ,
    \top_I.branch[20].block[14].um_I.clk ,
    \top_I.branch[20].block[13].um_I.iw[17] ,
    \top_I.branch[20].block[13].um_I.iw[16] ,
    \top_I.branch[20].block[13].um_I.iw[15] ,
    \top_I.branch[20].block[13].um_I.iw[14] ,
    \top_I.branch[20].block[13].um_I.iw[13] ,
    \top_I.branch[20].block[13].um_I.iw[12] ,
    \top_I.branch[20].block[13].um_I.iw[11] ,
    \top_I.branch[20].block[13].um_I.iw[10] ,
    \top_I.branch[20].block[13].um_I.iw[9] ,
    \top_I.branch[20].block[13].um_I.iw[8] ,
    \top_I.branch[20].block[13].um_I.iw[7] ,
    \top_I.branch[20].block[13].um_I.iw[6] ,
    \top_I.branch[20].block[13].um_I.iw[5] ,
    \top_I.branch[20].block[13].um_I.iw[4] ,
    \top_I.branch[20].block[13].um_I.iw[3] ,
    \top_I.branch[20].block[13].um_I.iw[2] ,
    \top_I.branch[20].block[13].um_I.iw[1] ,
    \top_I.branch[20].block[13].um_I.clk ,
    \top_I.branch[20].block[12].um_I.iw[17] ,
    \top_I.branch[20].block[12].um_I.iw[16] ,
    \top_I.branch[20].block[12].um_I.iw[15] ,
    \top_I.branch[20].block[12].um_I.iw[14] ,
    \top_I.branch[20].block[12].um_I.iw[13] ,
    \top_I.branch[20].block[12].um_I.iw[12] ,
    \top_I.branch[20].block[12].um_I.iw[11] ,
    \top_I.branch[20].block[12].um_I.iw[10] ,
    \top_I.branch[20].block[12].um_I.iw[9] ,
    \top_I.branch[20].block[12].um_I.iw[8] ,
    \top_I.branch[20].block[12].um_I.iw[7] ,
    \top_I.branch[20].block[12].um_I.iw[6] ,
    \top_I.branch[20].block[12].um_I.iw[5] ,
    \top_I.branch[20].block[12].um_I.iw[4] ,
    \top_I.branch[20].block[12].um_I.iw[3] ,
    \top_I.branch[20].block[12].um_I.iw[2] ,
    \top_I.branch[20].block[12].um_I.iw[1] ,
    \top_I.branch[20].block[12].um_I.clk ,
    \top_I.branch[20].block[11].um_I.iw[17] ,
    \top_I.branch[20].block[11].um_I.iw[16] ,
    \top_I.branch[20].block[11].um_I.iw[15] ,
    \top_I.branch[20].block[11].um_I.iw[14] ,
    \top_I.branch[20].block[11].um_I.iw[13] ,
    \top_I.branch[20].block[11].um_I.iw[12] ,
    \top_I.branch[20].block[11].um_I.iw[11] ,
    \top_I.branch[20].block[11].um_I.iw[10] ,
    \top_I.branch[20].block[11].um_I.iw[9] ,
    \top_I.branch[20].block[11].um_I.iw[8] ,
    \top_I.branch[20].block[11].um_I.iw[7] ,
    \top_I.branch[20].block[11].um_I.iw[6] ,
    \top_I.branch[20].block[11].um_I.iw[5] ,
    \top_I.branch[20].block[11].um_I.iw[4] ,
    \top_I.branch[20].block[11].um_I.iw[3] ,
    \top_I.branch[20].block[11].um_I.iw[2] ,
    \top_I.branch[20].block[11].um_I.iw[1] ,
    \top_I.branch[20].block[11].um_I.clk ,
    \top_I.branch[20].block[10].um_I.iw[17] ,
    \top_I.branch[20].block[10].um_I.iw[16] ,
    \top_I.branch[20].block[10].um_I.iw[15] ,
    \top_I.branch[20].block[10].um_I.iw[14] ,
    \top_I.branch[20].block[10].um_I.iw[13] ,
    \top_I.branch[20].block[10].um_I.iw[12] ,
    \top_I.branch[20].block[10].um_I.iw[11] ,
    \top_I.branch[20].block[10].um_I.iw[10] ,
    \top_I.branch[20].block[10].um_I.iw[9] ,
    \top_I.branch[20].block[10].um_I.iw[8] ,
    \top_I.branch[20].block[10].um_I.iw[7] ,
    \top_I.branch[20].block[10].um_I.iw[6] ,
    \top_I.branch[20].block[10].um_I.iw[5] ,
    \top_I.branch[20].block[10].um_I.iw[4] ,
    \top_I.branch[20].block[10].um_I.iw[3] ,
    \top_I.branch[20].block[10].um_I.iw[2] ,
    \top_I.branch[20].block[10].um_I.iw[1] ,
    \top_I.branch[20].block[10].um_I.clk ,
    \top_I.branch[20].block[9].um_I.iw[17] ,
    \top_I.branch[20].block[9].um_I.iw[16] ,
    \top_I.branch[20].block[9].um_I.iw[15] ,
    \top_I.branch[20].block[9].um_I.iw[14] ,
    \top_I.branch[20].block[9].um_I.iw[13] ,
    \top_I.branch[20].block[9].um_I.iw[12] ,
    \top_I.branch[20].block[9].um_I.iw[11] ,
    \top_I.branch[20].block[9].um_I.iw[10] ,
    \top_I.branch[20].block[9].um_I.iw[9] ,
    \top_I.branch[20].block[9].um_I.iw[8] ,
    \top_I.branch[20].block[9].um_I.iw[7] ,
    \top_I.branch[20].block[9].um_I.iw[6] ,
    \top_I.branch[20].block[9].um_I.iw[5] ,
    \top_I.branch[20].block[9].um_I.iw[4] ,
    \top_I.branch[20].block[9].um_I.iw[3] ,
    \top_I.branch[20].block[9].um_I.iw[2] ,
    \top_I.branch[20].block[9].um_I.iw[1] ,
    \top_I.branch[20].block[9].um_I.clk ,
    \top_I.branch[20].block[8].um_I.iw[17] ,
    \top_I.branch[20].block[8].um_I.iw[16] ,
    \top_I.branch[20].block[8].um_I.iw[15] ,
    \top_I.branch[20].block[8].um_I.iw[14] ,
    \top_I.branch[20].block[8].um_I.iw[13] ,
    \top_I.branch[20].block[8].um_I.iw[12] ,
    \top_I.branch[20].block[8].um_I.iw[11] ,
    \top_I.branch[20].block[8].um_I.iw[10] ,
    \top_I.branch[20].block[8].um_I.iw[9] ,
    \top_I.branch[20].block[8].um_I.iw[8] ,
    \top_I.branch[20].block[8].um_I.iw[7] ,
    \top_I.branch[20].block[8].um_I.iw[6] ,
    \top_I.branch[20].block[8].um_I.iw[5] ,
    \top_I.branch[20].block[8].um_I.iw[4] ,
    \top_I.branch[20].block[8].um_I.iw[3] ,
    \top_I.branch[20].block[8].um_I.iw[2] ,
    \top_I.branch[20].block[8].um_I.iw[1] ,
    \top_I.branch[20].block[8].um_I.clk ,
    \top_I.branch[20].block[7].um_I.iw[17] ,
    \top_I.branch[20].block[7].um_I.iw[16] ,
    \top_I.branch[20].block[7].um_I.iw[15] ,
    \top_I.branch[20].block[7].um_I.iw[14] ,
    \top_I.branch[20].block[7].um_I.iw[13] ,
    \top_I.branch[20].block[7].um_I.iw[12] ,
    \top_I.branch[20].block[7].um_I.iw[11] ,
    \top_I.branch[20].block[7].um_I.iw[10] ,
    \top_I.branch[20].block[7].um_I.iw[9] ,
    \top_I.branch[20].block[7].um_I.iw[8] ,
    \top_I.branch[20].block[7].um_I.iw[7] ,
    \top_I.branch[20].block[7].um_I.iw[6] ,
    \top_I.branch[20].block[7].um_I.iw[5] ,
    \top_I.branch[20].block[7].um_I.iw[4] ,
    \top_I.branch[20].block[7].um_I.iw[3] ,
    \top_I.branch[20].block[7].um_I.iw[2] ,
    \top_I.branch[20].block[7].um_I.iw[1] ,
    \top_I.branch[20].block[7].um_I.clk ,
    \top_I.branch[20].block[6].um_I.iw[17] ,
    \top_I.branch[20].block[6].um_I.iw[16] ,
    \top_I.branch[20].block[6].um_I.iw[15] ,
    \top_I.branch[20].block[6].um_I.iw[14] ,
    \top_I.branch[20].block[6].um_I.iw[13] ,
    \top_I.branch[20].block[6].um_I.iw[12] ,
    \top_I.branch[20].block[6].um_I.iw[11] ,
    \top_I.branch[20].block[6].um_I.iw[10] ,
    \top_I.branch[20].block[6].um_I.iw[9] ,
    \top_I.branch[20].block[6].um_I.iw[8] ,
    \top_I.branch[20].block[6].um_I.iw[7] ,
    \top_I.branch[20].block[6].um_I.iw[6] ,
    \top_I.branch[20].block[6].um_I.iw[5] ,
    \top_I.branch[20].block[6].um_I.iw[4] ,
    \top_I.branch[20].block[6].um_I.iw[3] ,
    \top_I.branch[20].block[6].um_I.iw[2] ,
    \top_I.branch[20].block[6].um_I.iw[1] ,
    \top_I.branch[20].block[6].um_I.clk ,
    \top_I.branch[20].block[5].um_I.iw[17] ,
    \top_I.branch[20].block[5].um_I.iw[16] ,
    \top_I.branch[20].block[5].um_I.iw[15] ,
    \top_I.branch[20].block[5].um_I.iw[14] ,
    \top_I.branch[20].block[5].um_I.iw[13] ,
    \top_I.branch[20].block[5].um_I.iw[12] ,
    \top_I.branch[20].block[5].um_I.iw[11] ,
    \top_I.branch[20].block[5].um_I.iw[10] ,
    \top_I.branch[20].block[5].um_I.iw[9] ,
    \top_I.branch[20].block[5].um_I.iw[8] ,
    \top_I.branch[20].block[5].um_I.iw[7] ,
    \top_I.branch[20].block[5].um_I.iw[6] ,
    \top_I.branch[20].block[5].um_I.iw[5] ,
    \top_I.branch[20].block[5].um_I.iw[4] ,
    \top_I.branch[20].block[5].um_I.iw[3] ,
    \top_I.branch[20].block[5].um_I.iw[2] ,
    \top_I.branch[20].block[5].um_I.iw[1] ,
    \top_I.branch[20].block[5].um_I.clk ,
    \top_I.branch[20].block[4].um_I.iw[17] ,
    \top_I.branch[20].block[4].um_I.iw[16] ,
    \top_I.branch[20].block[4].um_I.iw[15] ,
    \top_I.branch[20].block[4].um_I.iw[14] ,
    \top_I.branch[20].block[4].um_I.iw[13] ,
    \top_I.branch[20].block[4].um_I.iw[12] ,
    \top_I.branch[20].block[4].um_I.iw[11] ,
    \top_I.branch[20].block[4].um_I.iw[10] ,
    \top_I.branch[20].block[4].um_I.iw[9] ,
    \top_I.branch[20].block[4].um_I.iw[8] ,
    \top_I.branch[20].block[4].um_I.iw[7] ,
    \top_I.branch[20].block[4].um_I.iw[6] ,
    \top_I.branch[20].block[4].um_I.iw[5] ,
    \top_I.branch[20].block[4].um_I.iw[4] ,
    \top_I.branch[20].block[4].um_I.iw[3] ,
    \top_I.branch[20].block[4].um_I.iw[2] ,
    \top_I.branch[20].block[4].um_I.iw[1] ,
    \top_I.branch[20].block[4].um_I.clk ,
    \top_I.branch[20].block[3].um_I.iw[17] ,
    \top_I.branch[20].block[3].um_I.iw[16] ,
    \top_I.branch[20].block[3].um_I.iw[15] ,
    \top_I.branch[20].block[3].um_I.iw[14] ,
    \top_I.branch[20].block[3].um_I.iw[13] ,
    \top_I.branch[20].block[3].um_I.iw[12] ,
    \top_I.branch[20].block[3].um_I.iw[11] ,
    \top_I.branch[20].block[3].um_I.iw[10] ,
    \top_I.branch[20].block[3].um_I.iw[9] ,
    \top_I.branch[20].block[3].um_I.iw[8] ,
    \top_I.branch[20].block[3].um_I.iw[7] ,
    \top_I.branch[20].block[3].um_I.iw[6] ,
    \top_I.branch[20].block[3].um_I.iw[5] ,
    \top_I.branch[20].block[3].um_I.iw[4] ,
    \top_I.branch[20].block[3].um_I.iw[3] ,
    \top_I.branch[20].block[3].um_I.iw[2] ,
    \top_I.branch[20].block[3].um_I.iw[1] ,
    \top_I.branch[20].block[3].um_I.clk ,
    \top_I.branch[20].block[2].um_I.iw[17] ,
    \top_I.branch[20].block[2].um_I.iw[16] ,
    \top_I.branch[20].block[2].um_I.iw[15] ,
    \top_I.branch[20].block[2].um_I.iw[14] ,
    \top_I.branch[20].block[2].um_I.iw[13] ,
    \top_I.branch[20].block[2].um_I.iw[12] ,
    \top_I.branch[20].block[2].um_I.iw[11] ,
    \top_I.branch[20].block[2].um_I.iw[10] ,
    \top_I.branch[20].block[2].um_I.iw[9] ,
    \top_I.branch[20].block[2].um_I.iw[8] ,
    \top_I.branch[20].block[2].um_I.iw[7] ,
    \top_I.branch[20].block[2].um_I.iw[6] ,
    \top_I.branch[20].block[2].um_I.iw[5] ,
    \top_I.branch[20].block[2].um_I.iw[4] ,
    \top_I.branch[20].block[2].um_I.iw[3] ,
    \top_I.branch[20].block[2].um_I.iw[2] ,
    \top_I.branch[20].block[2].um_I.iw[1] ,
    \top_I.branch[20].block[2].um_I.clk ,
    \top_I.branch[20].block[1].um_I.iw[17] ,
    \top_I.branch[20].block[1].um_I.iw[16] ,
    \top_I.branch[20].block[1].um_I.iw[15] ,
    \top_I.branch[20].block[1].um_I.iw[14] ,
    \top_I.branch[20].block[1].um_I.iw[13] ,
    \top_I.branch[20].block[1].um_I.iw[12] ,
    \top_I.branch[20].block[1].um_I.iw[11] ,
    \top_I.branch[20].block[1].um_I.iw[10] ,
    \top_I.branch[20].block[1].um_I.iw[9] ,
    \top_I.branch[20].block[1].um_I.iw[8] ,
    \top_I.branch[20].block[1].um_I.iw[7] ,
    \top_I.branch[20].block[1].um_I.iw[6] ,
    \top_I.branch[20].block[1].um_I.iw[5] ,
    \top_I.branch[20].block[1].um_I.iw[4] ,
    \top_I.branch[20].block[1].um_I.iw[3] ,
    \top_I.branch[20].block[1].um_I.iw[2] ,
    \top_I.branch[20].block[1].um_I.iw[1] ,
    \top_I.branch[20].block[1].um_I.clk ,
    \top_I.branch[20].block[0].um_I.iw[17] ,
    \top_I.branch[20].block[0].um_I.iw[16] ,
    \top_I.branch[20].block[0].um_I.iw[15] ,
    \top_I.branch[20].block[0].um_I.iw[14] ,
    \top_I.branch[20].block[0].um_I.iw[13] ,
    \top_I.branch[20].block[0].um_I.iw[12] ,
    \top_I.branch[20].block[0].um_I.iw[11] ,
    \top_I.branch[20].block[0].um_I.iw[10] ,
    \top_I.branch[20].block[0].um_I.iw[9] ,
    \top_I.branch[20].block[0].um_I.iw[8] ,
    \top_I.branch[20].block[0].um_I.iw[7] ,
    \top_I.branch[20].block[0].um_I.iw[6] ,
    \top_I.branch[20].block[0].um_I.iw[5] ,
    \top_I.branch[20].block[0].um_I.iw[4] ,
    \top_I.branch[20].block[0].um_I.iw[3] ,
    \top_I.branch[20].block[0].um_I.iw[2] ,
    \top_I.branch[20].block[0].um_I.iw[1] ,
    \top_I.branch[20].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[15].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[14].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[13].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[12].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[11].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[10].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[9].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[8].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[7].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[6].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[5].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[4].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[3].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[2].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[1].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero ,
    \top_I.branch[20].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[20].block[15].um_I.pg_vdd ,
    \top_I.branch[20].block[14].um_I.pg_vdd ,
    \top_I.branch[20].block[13].um_I.pg_vdd ,
    \top_I.branch[20].block[12].um_I.pg_vdd ,
    \top_I.branch[20].block[11].um_I.pg_vdd ,
    \top_I.branch[20].block[10].um_I.pg_vdd ,
    \top_I.branch[20].block[9].um_I.pg_vdd ,
    \top_I.branch[20].block[8].um_I.pg_vdd ,
    \top_I.branch[20].block[7].um_I.pg_vdd ,
    \top_I.branch[20].block[6].um_I.pg_vdd ,
    \top_I.branch[20].block[5].um_I.pg_vdd ,
    \top_I.branch[20].block[4].um_I.pg_vdd ,
    \top_I.branch[20].block[3].um_I.pg_vdd ,
    \top_I.branch[20].block[2].um_I.pg_vdd ,
    \top_I.branch[20].block[1].um_I.pg_vdd ,
    \top_I.branch[20].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[21].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[21].l_addr[1] ),
    .k_zero(\top_I.branch[21].l_addr[0] ),
    .addr({\top_I.branch[21].l_addr[1] ,
    \top_I.branch[21].l_addr[0] ,
    \top_I.branch[21].l_addr[1] ,
    \top_I.branch[21].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[21].block[15].um_I.ena ,
    \top_I.branch[21].block[14].um_I.ena ,
    \top_I.branch[21].block[13].um_I.ena ,
    \top_I.branch[21].block[12].um_I.ena ,
    \top_I.branch[21].block[11].um_I.ena ,
    \top_I.branch[21].block[10].um_I.ena ,
    \top_I.branch[21].block[9].um_I.ena ,
    \top_I.branch[21].block[8].um_I.ena ,
    \top_I.branch[21].block[7].um_I.ena ,
    \top_I.branch[21].block[6].um_I.ena ,
    \top_I.branch[21].block[5].um_I.ena ,
    \top_I.branch[21].block[4].um_I.ena ,
    \top_I.branch[21].block[3].um_I.ena ,
    \top_I.branch[21].block[2].um_I.ena ,
    \top_I.branch[21].block[1].um_I.ena ,
    \top_I.branch[21].block[0].um_I.ena }),
    .um_iw({\top_I.branch[21].block[15].um_I.iw[17] ,
    \top_I.branch[21].block[15].um_I.iw[16] ,
    \top_I.branch[21].block[15].um_I.iw[15] ,
    \top_I.branch[21].block[15].um_I.iw[14] ,
    \top_I.branch[21].block[15].um_I.iw[13] ,
    \top_I.branch[21].block[15].um_I.iw[12] ,
    \top_I.branch[21].block[15].um_I.iw[11] ,
    \top_I.branch[21].block[15].um_I.iw[10] ,
    \top_I.branch[21].block[15].um_I.iw[9] ,
    \top_I.branch[21].block[15].um_I.iw[8] ,
    \top_I.branch[21].block[15].um_I.iw[7] ,
    \top_I.branch[21].block[15].um_I.iw[6] ,
    \top_I.branch[21].block[15].um_I.iw[5] ,
    \top_I.branch[21].block[15].um_I.iw[4] ,
    \top_I.branch[21].block[15].um_I.iw[3] ,
    \top_I.branch[21].block[15].um_I.iw[2] ,
    \top_I.branch[21].block[15].um_I.iw[1] ,
    \top_I.branch[21].block[15].um_I.clk ,
    \top_I.branch[21].block[14].um_I.iw[17] ,
    \top_I.branch[21].block[14].um_I.iw[16] ,
    \top_I.branch[21].block[14].um_I.iw[15] ,
    \top_I.branch[21].block[14].um_I.iw[14] ,
    \top_I.branch[21].block[14].um_I.iw[13] ,
    \top_I.branch[21].block[14].um_I.iw[12] ,
    \top_I.branch[21].block[14].um_I.iw[11] ,
    \top_I.branch[21].block[14].um_I.iw[10] ,
    \top_I.branch[21].block[14].um_I.iw[9] ,
    \top_I.branch[21].block[14].um_I.iw[8] ,
    \top_I.branch[21].block[14].um_I.iw[7] ,
    \top_I.branch[21].block[14].um_I.iw[6] ,
    \top_I.branch[21].block[14].um_I.iw[5] ,
    \top_I.branch[21].block[14].um_I.iw[4] ,
    \top_I.branch[21].block[14].um_I.iw[3] ,
    \top_I.branch[21].block[14].um_I.iw[2] ,
    \top_I.branch[21].block[14].um_I.iw[1] ,
    \top_I.branch[21].block[14].um_I.clk ,
    \top_I.branch[21].block[13].um_I.iw[17] ,
    \top_I.branch[21].block[13].um_I.iw[16] ,
    \top_I.branch[21].block[13].um_I.iw[15] ,
    \top_I.branch[21].block[13].um_I.iw[14] ,
    \top_I.branch[21].block[13].um_I.iw[13] ,
    \top_I.branch[21].block[13].um_I.iw[12] ,
    \top_I.branch[21].block[13].um_I.iw[11] ,
    \top_I.branch[21].block[13].um_I.iw[10] ,
    \top_I.branch[21].block[13].um_I.iw[9] ,
    \top_I.branch[21].block[13].um_I.iw[8] ,
    \top_I.branch[21].block[13].um_I.iw[7] ,
    \top_I.branch[21].block[13].um_I.iw[6] ,
    \top_I.branch[21].block[13].um_I.iw[5] ,
    \top_I.branch[21].block[13].um_I.iw[4] ,
    \top_I.branch[21].block[13].um_I.iw[3] ,
    \top_I.branch[21].block[13].um_I.iw[2] ,
    \top_I.branch[21].block[13].um_I.iw[1] ,
    \top_I.branch[21].block[13].um_I.clk ,
    \top_I.branch[21].block[12].um_I.iw[17] ,
    \top_I.branch[21].block[12].um_I.iw[16] ,
    \top_I.branch[21].block[12].um_I.iw[15] ,
    \top_I.branch[21].block[12].um_I.iw[14] ,
    \top_I.branch[21].block[12].um_I.iw[13] ,
    \top_I.branch[21].block[12].um_I.iw[12] ,
    \top_I.branch[21].block[12].um_I.iw[11] ,
    \top_I.branch[21].block[12].um_I.iw[10] ,
    \top_I.branch[21].block[12].um_I.iw[9] ,
    \top_I.branch[21].block[12].um_I.iw[8] ,
    \top_I.branch[21].block[12].um_I.iw[7] ,
    \top_I.branch[21].block[12].um_I.iw[6] ,
    \top_I.branch[21].block[12].um_I.iw[5] ,
    \top_I.branch[21].block[12].um_I.iw[4] ,
    \top_I.branch[21].block[12].um_I.iw[3] ,
    \top_I.branch[21].block[12].um_I.iw[2] ,
    \top_I.branch[21].block[12].um_I.iw[1] ,
    \top_I.branch[21].block[12].um_I.clk ,
    \top_I.branch[21].block[11].um_I.iw[17] ,
    \top_I.branch[21].block[11].um_I.iw[16] ,
    \top_I.branch[21].block[11].um_I.iw[15] ,
    \top_I.branch[21].block[11].um_I.iw[14] ,
    \top_I.branch[21].block[11].um_I.iw[13] ,
    \top_I.branch[21].block[11].um_I.iw[12] ,
    \top_I.branch[21].block[11].um_I.iw[11] ,
    \top_I.branch[21].block[11].um_I.iw[10] ,
    \top_I.branch[21].block[11].um_I.iw[9] ,
    \top_I.branch[21].block[11].um_I.iw[8] ,
    \top_I.branch[21].block[11].um_I.iw[7] ,
    \top_I.branch[21].block[11].um_I.iw[6] ,
    \top_I.branch[21].block[11].um_I.iw[5] ,
    \top_I.branch[21].block[11].um_I.iw[4] ,
    \top_I.branch[21].block[11].um_I.iw[3] ,
    \top_I.branch[21].block[11].um_I.iw[2] ,
    \top_I.branch[21].block[11].um_I.iw[1] ,
    \top_I.branch[21].block[11].um_I.clk ,
    \top_I.branch[21].block[10].um_I.iw[17] ,
    \top_I.branch[21].block[10].um_I.iw[16] ,
    \top_I.branch[21].block[10].um_I.iw[15] ,
    \top_I.branch[21].block[10].um_I.iw[14] ,
    \top_I.branch[21].block[10].um_I.iw[13] ,
    \top_I.branch[21].block[10].um_I.iw[12] ,
    \top_I.branch[21].block[10].um_I.iw[11] ,
    \top_I.branch[21].block[10].um_I.iw[10] ,
    \top_I.branch[21].block[10].um_I.iw[9] ,
    \top_I.branch[21].block[10].um_I.iw[8] ,
    \top_I.branch[21].block[10].um_I.iw[7] ,
    \top_I.branch[21].block[10].um_I.iw[6] ,
    \top_I.branch[21].block[10].um_I.iw[5] ,
    \top_I.branch[21].block[10].um_I.iw[4] ,
    \top_I.branch[21].block[10].um_I.iw[3] ,
    \top_I.branch[21].block[10].um_I.iw[2] ,
    \top_I.branch[21].block[10].um_I.iw[1] ,
    \top_I.branch[21].block[10].um_I.clk ,
    \top_I.branch[21].block[9].um_I.iw[17] ,
    \top_I.branch[21].block[9].um_I.iw[16] ,
    \top_I.branch[21].block[9].um_I.iw[15] ,
    \top_I.branch[21].block[9].um_I.iw[14] ,
    \top_I.branch[21].block[9].um_I.iw[13] ,
    \top_I.branch[21].block[9].um_I.iw[12] ,
    \top_I.branch[21].block[9].um_I.iw[11] ,
    \top_I.branch[21].block[9].um_I.iw[10] ,
    \top_I.branch[21].block[9].um_I.iw[9] ,
    \top_I.branch[21].block[9].um_I.iw[8] ,
    \top_I.branch[21].block[9].um_I.iw[7] ,
    \top_I.branch[21].block[9].um_I.iw[6] ,
    \top_I.branch[21].block[9].um_I.iw[5] ,
    \top_I.branch[21].block[9].um_I.iw[4] ,
    \top_I.branch[21].block[9].um_I.iw[3] ,
    \top_I.branch[21].block[9].um_I.iw[2] ,
    \top_I.branch[21].block[9].um_I.iw[1] ,
    \top_I.branch[21].block[9].um_I.clk ,
    \top_I.branch[21].block[8].um_I.iw[17] ,
    \top_I.branch[21].block[8].um_I.iw[16] ,
    \top_I.branch[21].block[8].um_I.iw[15] ,
    \top_I.branch[21].block[8].um_I.iw[14] ,
    \top_I.branch[21].block[8].um_I.iw[13] ,
    \top_I.branch[21].block[8].um_I.iw[12] ,
    \top_I.branch[21].block[8].um_I.iw[11] ,
    \top_I.branch[21].block[8].um_I.iw[10] ,
    \top_I.branch[21].block[8].um_I.iw[9] ,
    \top_I.branch[21].block[8].um_I.iw[8] ,
    \top_I.branch[21].block[8].um_I.iw[7] ,
    \top_I.branch[21].block[8].um_I.iw[6] ,
    \top_I.branch[21].block[8].um_I.iw[5] ,
    \top_I.branch[21].block[8].um_I.iw[4] ,
    \top_I.branch[21].block[8].um_I.iw[3] ,
    \top_I.branch[21].block[8].um_I.iw[2] ,
    \top_I.branch[21].block[8].um_I.iw[1] ,
    \top_I.branch[21].block[8].um_I.clk ,
    \top_I.branch[21].block[7].um_I.iw[17] ,
    \top_I.branch[21].block[7].um_I.iw[16] ,
    \top_I.branch[21].block[7].um_I.iw[15] ,
    \top_I.branch[21].block[7].um_I.iw[14] ,
    \top_I.branch[21].block[7].um_I.iw[13] ,
    \top_I.branch[21].block[7].um_I.iw[12] ,
    \top_I.branch[21].block[7].um_I.iw[11] ,
    \top_I.branch[21].block[7].um_I.iw[10] ,
    \top_I.branch[21].block[7].um_I.iw[9] ,
    \top_I.branch[21].block[7].um_I.iw[8] ,
    \top_I.branch[21].block[7].um_I.iw[7] ,
    \top_I.branch[21].block[7].um_I.iw[6] ,
    \top_I.branch[21].block[7].um_I.iw[5] ,
    \top_I.branch[21].block[7].um_I.iw[4] ,
    \top_I.branch[21].block[7].um_I.iw[3] ,
    \top_I.branch[21].block[7].um_I.iw[2] ,
    \top_I.branch[21].block[7].um_I.iw[1] ,
    \top_I.branch[21].block[7].um_I.clk ,
    \top_I.branch[21].block[6].um_I.iw[17] ,
    \top_I.branch[21].block[6].um_I.iw[16] ,
    \top_I.branch[21].block[6].um_I.iw[15] ,
    \top_I.branch[21].block[6].um_I.iw[14] ,
    \top_I.branch[21].block[6].um_I.iw[13] ,
    \top_I.branch[21].block[6].um_I.iw[12] ,
    \top_I.branch[21].block[6].um_I.iw[11] ,
    \top_I.branch[21].block[6].um_I.iw[10] ,
    \top_I.branch[21].block[6].um_I.iw[9] ,
    \top_I.branch[21].block[6].um_I.iw[8] ,
    \top_I.branch[21].block[6].um_I.iw[7] ,
    \top_I.branch[21].block[6].um_I.iw[6] ,
    \top_I.branch[21].block[6].um_I.iw[5] ,
    \top_I.branch[21].block[6].um_I.iw[4] ,
    \top_I.branch[21].block[6].um_I.iw[3] ,
    \top_I.branch[21].block[6].um_I.iw[2] ,
    \top_I.branch[21].block[6].um_I.iw[1] ,
    \top_I.branch[21].block[6].um_I.clk ,
    \top_I.branch[21].block[5].um_I.iw[17] ,
    \top_I.branch[21].block[5].um_I.iw[16] ,
    \top_I.branch[21].block[5].um_I.iw[15] ,
    \top_I.branch[21].block[5].um_I.iw[14] ,
    \top_I.branch[21].block[5].um_I.iw[13] ,
    \top_I.branch[21].block[5].um_I.iw[12] ,
    \top_I.branch[21].block[5].um_I.iw[11] ,
    \top_I.branch[21].block[5].um_I.iw[10] ,
    \top_I.branch[21].block[5].um_I.iw[9] ,
    \top_I.branch[21].block[5].um_I.iw[8] ,
    \top_I.branch[21].block[5].um_I.iw[7] ,
    \top_I.branch[21].block[5].um_I.iw[6] ,
    \top_I.branch[21].block[5].um_I.iw[5] ,
    \top_I.branch[21].block[5].um_I.iw[4] ,
    \top_I.branch[21].block[5].um_I.iw[3] ,
    \top_I.branch[21].block[5].um_I.iw[2] ,
    \top_I.branch[21].block[5].um_I.iw[1] ,
    \top_I.branch[21].block[5].um_I.clk ,
    \top_I.branch[21].block[4].um_I.iw[17] ,
    \top_I.branch[21].block[4].um_I.iw[16] ,
    \top_I.branch[21].block[4].um_I.iw[15] ,
    \top_I.branch[21].block[4].um_I.iw[14] ,
    \top_I.branch[21].block[4].um_I.iw[13] ,
    \top_I.branch[21].block[4].um_I.iw[12] ,
    \top_I.branch[21].block[4].um_I.iw[11] ,
    \top_I.branch[21].block[4].um_I.iw[10] ,
    \top_I.branch[21].block[4].um_I.iw[9] ,
    \top_I.branch[21].block[4].um_I.iw[8] ,
    \top_I.branch[21].block[4].um_I.iw[7] ,
    \top_I.branch[21].block[4].um_I.iw[6] ,
    \top_I.branch[21].block[4].um_I.iw[5] ,
    \top_I.branch[21].block[4].um_I.iw[4] ,
    \top_I.branch[21].block[4].um_I.iw[3] ,
    \top_I.branch[21].block[4].um_I.iw[2] ,
    \top_I.branch[21].block[4].um_I.iw[1] ,
    \top_I.branch[21].block[4].um_I.clk ,
    \top_I.branch[21].block[3].um_I.iw[17] ,
    \top_I.branch[21].block[3].um_I.iw[16] ,
    \top_I.branch[21].block[3].um_I.iw[15] ,
    \top_I.branch[21].block[3].um_I.iw[14] ,
    \top_I.branch[21].block[3].um_I.iw[13] ,
    \top_I.branch[21].block[3].um_I.iw[12] ,
    \top_I.branch[21].block[3].um_I.iw[11] ,
    \top_I.branch[21].block[3].um_I.iw[10] ,
    \top_I.branch[21].block[3].um_I.iw[9] ,
    \top_I.branch[21].block[3].um_I.iw[8] ,
    \top_I.branch[21].block[3].um_I.iw[7] ,
    \top_I.branch[21].block[3].um_I.iw[6] ,
    \top_I.branch[21].block[3].um_I.iw[5] ,
    \top_I.branch[21].block[3].um_I.iw[4] ,
    \top_I.branch[21].block[3].um_I.iw[3] ,
    \top_I.branch[21].block[3].um_I.iw[2] ,
    \top_I.branch[21].block[3].um_I.iw[1] ,
    \top_I.branch[21].block[3].um_I.clk ,
    \top_I.branch[21].block[2].um_I.iw[17] ,
    \top_I.branch[21].block[2].um_I.iw[16] ,
    \top_I.branch[21].block[2].um_I.iw[15] ,
    \top_I.branch[21].block[2].um_I.iw[14] ,
    \top_I.branch[21].block[2].um_I.iw[13] ,
    \top_I.branch[21].block[2].um_I.iw[12] ,
    \top_I.branch[21].block[2].um_I.iw[11] ,
    \top_I.branch[21].block[2].um_I.iw[10] ,
    \top_I.branch[21].block[2].um_I.iw[9] ,
    \top_I.branch[21].block[2].um_I.iw[8] ,
    \top_I.branch[21].block[2].um_I.iw[7] ,
    \top_I.branch[21].block[2].um_I.iw[6] ,
    \top_I.branch[21].block[2].um_I.iw[5] ,
    \top_I.branch[21].block[2].um_I.iw[4] ,
    \top_I.branch[21].block[2].um_I.iw[3] ,
    \top_I.branch[21].block[2].um_I.iw[2] ,
    \top_I.branch[21].block[2].um_I.iw[1] ,
    \top_I.branch[21].block[2].um_I.clk ,
    \top_I.branch[21].block[1].um_I.iw[17] ,
    \top_I.branch[21].block[1].um_I.iw[16] ,
    \top_I.branch[21].block[1].um_I.iw[15] ,
    \top_I.branch[21].block[1].um_I.iw[14] ,
    \top_I.branch[21].block[1].um_I.iw[13] ,
    \top_I.branch[21].block[1].um_I.iw[12] ,
    \top_I.branch[21].block[1].um_I.iw[11] ,
    \top_I.branch[21].block[1].um_I.iw[10] ,
    \top_I.branch[21].block[1].um_I.iw[9] ,
    \top_I.branch[21].block[1].um_I.iw[8] ,
    \top_I.branch[21].block[1].um_I.iw[7] ,
    \top_I.branch[21].block[1].um_I.iw[6] ,
    \top_I.branch[21].block[1].um_I.iw[5] ,
    \top_I.branch[21].block[1].um_I.iw[4] ,
    \top_I.branch[21].block[1].um_I.iw[3] ,
    \top_I.branch[21].block[1].um_I.iw[2] ,
    \top_I.branch[21].block[1].um_I.iw[1] ,
    \top_I.branch[21].block[1].um_I.clk ,
    \top_I.branch[21].block[0].um_I.iw[17] ,
    \top_I.branch[21].block[0].um_I.iw[16] ,
    \top_I.branch[21].block[0].um_I.iw[15] ,
    \top_I.branch[21].block[0].um_I.iw[14] ,
    \top_I.branch[21].block[0].um_I.iw[13] ,
    \top_I.branch[21].block[0].um_I.iw[12] ,
    \top_I.branch[21].block[0].um_I.iw[11] ,
    \top_I.branch[21].block[0].um_I.iw[10] ,
    \top_I.branch[21].block[0].um_I.iw[9] ,
    \top_I.branch[21].block[0].um_I.iw[8] ,
    \top_I.branch[21].block[0].um_I.iw[7] ,
    \top_I.branch[21].block[0].um_I.iw[6] ,
    \top_I.branch[21].block[0].um_I.iw[5] ,
    \top_I.branch[21].block[0].um_I.iw[4] ,
    \top_I.branch[21].block[0].um_I.iw[3] ,
    \top_I.branch[21].block[0].um_I.iw[2] ,
    \top_I.branch[21].block[0].um_I.iw[1] ,
    \top_I.branch[21].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[15].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[14].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[13].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[12].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[11].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[10].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[9].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[8].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[7].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[6].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[5].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[4].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[3].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[2].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[1].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero ,
    \top_I.branch[21].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[21].block[15].um_I.pg_vdd ,
    \top_I.branch[21].block[14].um_I.pg_vdd ,
    \top_I.branch[21].block[13].um_I.pg_vdd ,
    \top_I.branch[21].block[12].um_I.pg_vdd ,
    \top_I.branch[21].block[11].um_I.pg_vdd ,
    \top_I.branch[21].block[10].um_I.pg_vdd ,
    \top_I.branch[21].block[9].um_I.pg_vdd ,
    \top_I.branch[21].block[8].um_I.pg_vdd ,
    \top_I.branch[21].block[7].um_I.pg_vdd ,
    \top_I.branch[21].block[6].um_I.pg_vdd ,
    \top_I.branch[21].block[5].um_I.pg_vdd ,
    \top_I.branch[21].block[4].um_I.pg_vdd ,
    \top_I.branch[21].block[3].um_I.pg_vdd ,
    \top_I.branch[21].block[2].um_I.pg_vdd ,
    \top_I.branch[21].block[1].um_I.pg_vdd ,
    \top_I.branch[21].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[22].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[22].l_addr[0] ),
    .k_zero(\top_I.branch[22].l_addr[2] ),
    .addr({\top_I.branch[22].l_addr[0] ,
    \top_I.branch[22].l_addr[2] ,
    \top_I.branch[22].l_addr[0] ,
    \top_I.branch[22].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[22].block[15].um_I.ena ,
    \top_I.branch[22].block[14].um_I.ena ,
    \top_I.branch[22].block[13].um_I.ena ,
    \top_I.branch[22].block[12].um_I.ena ,
    \top_I.branch[22].block[11].um_I.ena ,
    \top_I.branch[22].block[10].um_I.ena ,
    \top_I.branch[22].block[9].um_I.ena ,
    \top_I.branch[22].block[8].um_I.ena ,
    \top_I.branch[22].block[7].um_I.ena ,
    \top_I.branch[22].block[6].um_I.ena ,
    \top_I.branch[22].block[5].um_I.ena ,
    \top_I.branch[22].block[4].um_I.ena ,
    \top_I.branch[22].block[3].um_I.ena ,
    \top_I.branch[22].block[2].um_I.ena ,
    \top_I.branch[22].block[1].um_I.ena ,
    \top_I.branch[22].block[0].um_I.ena }),
    .um_iw({\top_I.branch[22].block[15].um_I.iw[17] ,
    \top_I.branch[22].block[15].um_I.iw[16] ,
    \top_I.branch[22].block[15].um_I.iw[15] ,
    \top_I.branch[22].block[15].um_I.iw[14] ,
    \top_I.branch[22].block[15].um_I.iw[13] ,
    \top_I.branch[22].block[15].um_I.iw[12] ,
    \top_I.branch[22].block[15].um_I.iw[11] ,
    \top_I.branch[22].block[15].um_I.iw[10] ,
    \top_I.branch[22].block[15].um_I.iw[9] ,
    \top_I.branch[22].block[15].um_I.iw[8] ,
    \top_I.branch[22].block[15].um_I.iw[7] ,
    \top_I.branch[22].block[15].um_I.iw[6] ,
    \top_I.branch[22].block[15].um_I.iw[5] ,
    \top_I.branch[22].block[15].um_I.iw[4] ,
    \top_I.branch[22].block[15].um_I.iw[3] ,
    \top_I.branch[22].block[15].um_I.iw[2] ,
    \top_I.branch[22].block[15].um_I.iw[1] ,
    \top_I.branch[22].block[15].um_I.clk ,
    \top_I.branch[22].block[14].um_I.iw[17] ,
    \top_I.branch[22].block[14].um_I.iw[16] ,
    \top_I.branch[22].block[14].um_I.iw[15] ,
    \top_I.branch[22].block[14].um_I.iw[14] ,
    \top_I.branch[22].block[14].um_I.iw[13] ,
    \top_I.branch[22].block[14].um_I.iw[12] ,
    \top_I.branch[22].block[14].um_I.iw[11] ,
    \top_I.branch[22].block[14].um_I.iw[10] ,
    \top_I.branch[22].block[14].um_I.iw[9] ,
    \top_I.branch[22].block[14].um_I.iw[8] ,
    \top_I.branch[22].block[14].um_I.iw[7] ,
    \top_I.branch[22].block[14].um_I.iw[6] ,
    \top_I.branch[22].block[14].um_I.iw[5] ,
    \top_I.branch[22].block[14].um_I.iw[4] ,
    \top_I.branch[22].block[14].um_I.iw[3] ,
    \top_I.branch[22].block[14].um_I.iw[2] ,
    \top_I.branch[22].block[14].um_I.iw[1] ,
    \top_I.branch[22].block[14].um_I.clk ,
    \top_I.branch[22].block[13].um_I.iw[17] ,
    \top_I.branch[22].block[13].um_I.iw[16] ,
    \top_I.branch[22].block[13].um_I.iw[15] ,
    \top_I.branch[22].block[13].um_I.iw[14] ,
    \top_I.branch[22].block[13].um_I.iw[13] ,
    \top_I.branch[22].block[13].um_I.iw[12] ,
    \top_I.branch[22].block[13].um_I.iw[11] ,
    \top_I.branch[22].block[13].um_I.iw[10] ,
    \top_I.branch[22].block[13].um_I.iw[9] ,
    \top_I.branch[22].block[13].um_I.iw[8] ,
    \top_I.branch[22].block[13].um_I.iw[7] ,
    \top_I.branch[22].block[13].um_I.iw[6] ,
    \top_I.branch[22].block[13].um_I.iw[5] ,
    \top_I.branch[22].block[13].um_I.iw[4] ,
    \top_I.branch[22].block[13].um_I.iw[3] ,
    \top_I.branch[22].block[13].um_I.iw[2] ,
    \top_I.branch[22].block[13].um_I.iw[1] ,
    \top_I.branch[22].block[13].um_I.clk ,
    \top_I.branch[22].block[12].um_I.iw[17] ,
    \top_I.branch[22].block[12].um_I.iw[16] ,
    \top_I.branch[22].block[12].um_I.iw[15] ,
    \top_I.branch[22].block[12].um_I.iw[14] ,
    \top_I.branch[22].block[12].um_I.iw[13] ,
    \top_I.branch[22].block[12].um_I.iw[12] ,
    \top_I.branch[22].block[12].um_I.iw[11] ,
    \top_I.branch[22].block[12].um_I.iw[10] ,
    \top_I.branch[22].block[12].um_I.iw[9] ,
    \top_I.branch[22].block[12].um_I.iw[8] ,
    \top_I.branch[22].block[12].um_I.iw[7] ,
    \top_I.branch[22].block[12].um_I.iw[6] ,
    \top_I.branch[22].block[12].um_I.iw[5] ,
    \top_I.branch[22].block[12].um_I.iw[4] ,
    \top_I.branch[22].block[12].um_I.iw[3] ,
    \top_I.branch[22].block[12].um_I.iw[2] ,
    \top_I.branch[22].block[12].um_I.iw[1] ,
    \top_I.branch[22].block[12].um_I.clk ,
    \top_I.branch[22].block[11].um_I.iw[17] ,
    \top_I.branch[22].block[11].um_I.iw[16] ,
    \top_I.branch[22].block[11].um_I.iw[15] ,
    \top_I.branch[22].block[11].um_I.iw[14] ,
    \top_I.branch[22].block[11].um_I.iw[13] ,
    \top_I.branch[22].block[11].um_I.iw[12] ,
    \top_I.branch[22].block[11].um_I.iw[11] ,
    \top_I.branch[22].block[11].um_I.iw[10] ,
    \top_I.branch[22].block[11].um_I.iw[9] ,
    \top_I.branch[22].block[11].um_I.iw[8] ,
    \top_I.branch[22].block[11].um_I.iw[7] ,
    \top_I.branch[22].block[11].um_I.iw[6] ,
    \top_I.branch[22].block[11].um_I.iw[5] ,
    \top_I.branch[22].block[11].um_I.iw[4] ,
    \top_I.branch[22].block[11].um_I.iw[3] ,
    \top_I.branch[22].block[11].um_I.iw[2] ,
    \top_I.branch[22].block[11].um_I.iw[1] ,
    \top_I.branch[22].block[11].um_I.clk ,
    \top_I.branch[22].block[10].um_I.iw[17] ,
    \top_I.branch[22].block[10].um_I.iw[16] ,
    \top_I.branch[22].block[10].um_I.iw[15] ,
    \top_I.branch[22].block[10].um_I.iw[14] ,
    \top_I.branch[22].block[10].um_I.iw[13] ,
    \top_I.branch[22].block[10].um_I.iw[12] ,
    \top_I.branch[22].block[10].um_I.iw[11] ,
    \top_I.branch[22].block[10].um_I.iw[10] ,
    \top_I.branch[22].block[10].um_I.iw[9] ,
    \top_I.branch[22].block[10].um_I.iw[8] ,
    \top_I.branch[22].block[10].um_I.iw[7] ,
    \top_I.branch[22].block[10].um_I.iw[6] ,
    \top_I.branch[22].block[10].um_I.iw[5] ,
    \top_I.branch[22].block[10].um_I.iw[4] ,
    \top_I.branch[22].block[10].um_I.iw[3] ,
    \top_I.branch[22].block[10].um_I.iw[2] ,
    \top_I.branch[22].block[10].um_I.iw[1] ,
    \top_I.branch[22].block[10].um_I.clk ,
    \top_I.branch[22].block[9].um_I.iw[17] ,
    \top_I.branch[22].block[9].um_I.iw[16] ,
    \top_I.branch[22].block[9].um_I.iw[15] ,
    \top_I.branch[22].block[9].um_I.iw[14] ,
    \top_I.branch[22].block[9].um_I.iw[13] ,
    \top_I.branch[22].block[9].um_I.iw[12] ,
    \top_I.branch[22].block[9].um_I.iw[11] ,
    \top_I.branch[22].block[9].um_I.iw[10] ,
    \top_I.branch[22].block[9].um_I.iw[9] ,
    \top_I.branch[22].block[9].um_I.iw[8] ,
    \top_I.branch[22].block[9].um_I.iw[7] ,
    \top_I.branch[22].block[9].um_I.iw[6] ,
    \top_I.branch[22].block[9].um_I.iw[5] ,
    \top_I.branch[22].block[9].um_I.iw[4] ,
    \top_I.branch[22].block[9].um_I.iw[3] ,
    \top_I.branch[22].block[9].um_I.iw[2] ,
    \top_I.branch[22].block[9].um_I.iw[1] ,
    \top_I.branch[22].block[9].um_I.clk ,
    \top_I.branch[22].block[8].um_I.iw[17] ,
    \top_I.branch[22].block[8].um_I.iw[16] ,
    \top_I.branch[22].block[8].um_I.iw[15] ,
    \top_I.branch[22].block[8].um_I.iw[14] ,
    \top_I.branch[22].block[8].um_I.iw[13] ,
    \top_I.branch[22].block[8].um_I.iw[12] ,
    \top_I.branch[22].block[8].um_I.iw[11] ,
    \top_I.branch[22].block[8].um_I.iw[10] ,
    \top_I.branch[22].block[8].um_I.iw[9] ,
    \top_I.branch[22].block[8].um_I.iw[8] ,
    \top_I.branch[22].block[8].um_I.iw[7] ,
    \top_I.branch[22].block[8].um_I.iw[6] ,
    \top_I.branch[22].block[8].um_I.iw[5] ,
    \top_I.branch[22].block[8].um_I.iw[4] ,
    \top_I.branch[22].block[8].um_I.iw[3] ,
    \top_I.branch[22].block[8].um_I.iw[2] ,
    \top_I.branch[22].block[8].um_I.iw[1] ,
    \top_I.branch[22].block[8].um_I.clk ,
    \top_I.branch[22].block[7].um_I.iw[17] ,
    \top_I.branch[22].block[7].um_I.iw[16] ,
    \top_I.branch[22].block[7].um_I.iw[15] ,
    \top_I.branch[22].block[7].um_I.iw[14] ,
    \top_I.branch[22].block[7].um_I.iw[13] ,
    \top_I.branch[22].block[7].um_I.iw[12] ,
    \top_I.branch[22].block[7].um_I.iw[11] ,
    \top_I.branch[22].block[7].um_I.iw[10] ,
    \top_I.branch[22].block[7].um_I.iw[9] ,
    \top_I.branch[22].block[7].um_I.iw[8] ,
    \top_I.branch[22].block[7].um_I.iw[7] ,
    \top_I.branch[22].block[7].um_I.iw[6] ,
    \top_I.branch[22].block[7].um_I.iw[5] ,
    \top_I.branch[22].block[7].um_I.iw[4] ,
    \top_I.branch[22].block[7].um_I.iw[3] ,
    \top_I.branch[22].block[7].um_I.iw[2] ,
    \top_I.branch[22].block[7].um_I.iw[1] ,
    \top_I.branch[22].block[7].um_I.clk ,
    \top_I.branch[22].block[6].um_I.iw[17] ,
    \top_I.branch[22].block[6].um_I.iw[16] ,
    \top_I.branch[22].block[6].um_I.iw[15] ,
    \top_I.branch[22].block[6].um_I.iw[14] ,
    \top_I.branch[22].block[6].um_I.iw[13] ,
    \top_I.branch[22].block[6].um_I.iw[12] ,
    \top_I.branch[22].block[6].um_I.iw[11] ,
    \top_I.branch[22].block[6].um_I.iw[10] ,
    \top_I.branch[22].block[6].um_I.iw[9] ,
    \top_I.branch[22].block[6].um_I.iw[8] ,
    \top_I.branch[22].block[6].um_I.iw[7] ,
    \top_I.branch[22].block[6].um_I.iw[6] ,
    \top_I.branch[22].block[6].um_I.iw[5] ,
    \top_I.branch[22].block[6].um_I.iw[4] ,
    \top_I.branch[22].block[6].um_I.iw[3] ,
    \top_I.branch[22].block[6].um_I.iw[2] ,
    \top_I.branch[22].block[6].um_I.iw[1] ,
    \top_I.branch[22].block[6].um_I.clk ,
    \top_I.branch[22].block[5].um_I.iw[17] ,
    \top_I.branch[22].block[5].um_I.iw[16] ,
    \top_I.branch[22].block[5].um_I.iw[15] ,
    \top_I.branch[22].block[5].um_I.iw[14] ,
    \top_I.branch[22].block[5].um_I.iw[13] ,
    \top_I.branch[22].block[5].um_I.iw[12] ,
    \top_I.branch[22].block[5].um_I.iw[11] ,
    \top_I.branch[22].block[5].um_I.iw[10] ,
    \top_I.branch[22].block[5].um_I.iw[9] ,
    \top_I.branch[22].block[5].um_I.iw[8] ,
    \top_I.branch[22].block[5].um_I.iw[7] ,
    \top_I.branch[22].block[5].um_I.iw[6] ,
    \top_I.branch[22].block[5].um_I.iw[5] ,
    \top_I.branch[22].block[5].um_I.iw[4] ,
    \top_I.branch[22].block[5].um_I.iw[3] ,
    \top_I.branch[22].block[5].um_I.iw[2] ,
    \top_I.branch[22].block[5].um_I.iw[1] ,
    \top_I.branch[22].block[5].um_I.clk ,
    \top_I.branch[22].block[4].um_I.iw[17] ,
    \top_I.branch[22].block[4].um_I.iw[16] ,
    \top_I.branch[22].block[4].um_I.iw[15] ,
    \top_I.branch[22].block[4].um_I.iw[14] ,
    \top_I.branch[22].block[4].um_I.iw[13] ,
    \top_I.branch[22].block[4].um_I.iw[12] ,
    \top_I.branch[22].block[4].um_I.iw[11] ,
    \top_I.branch[22].block[4].um_I.iw[10] ,
    \top_I.branch[22].block[4].um_I.iw[9] ,
    \top_I.branch[22].block[4].um_I.iw[8] ,
    \top_I.branch[22].block[4].um_I.iw[7] ,
    \top_I.branch[22].block[4].um_I.iw[6] ,
    \top_I.branch[22].block[4].um_I.iw[5] ,
    \top_I.branch[22].block[4].um_I.iw[4] ,
    \top_I.branch[22].block[4].um_I.iw[3] ,
    \top_I.branch[22].block[4].um_I.iw[2] ,
    \top_I.branch[22].block[4].um_I.iw[1] ,
    \top_I.branch[22].block[4].um_I.clk ,
    \top_I.branch[22].block[3].um_I.iw[17] ,
    \top_I.branch[22].block[3].um_I.iw[16] ,
    \top_I.branch[22].block[3].um_I.iw[15] ,
    \top_I.branch[22].block[3].um_I.iw[14] ,
    \top_I.branch[22].block[3].um_I.iw[13] ,
    \top_I.branch[22].block[3].um_I.iw[12] ,
    \top_I.branch[22].block[3].um_I.iw[11] ,
    \top_I.branch[22].block[3].um_I.iw[10] ,
    \top_I.branch[22].block[3].um_I.iw[9] ,
    \top_I.branch[22].block[3].um_I.iw[8] ,
    \top_I.branch[22].block[3].um_I.iw[7] ,
    \top_I.branch[22].block[3].um_I.iw[6] ,
    \top_I.branch[22].block[3].um_I.iw[5] ,
    \top_I.branch[22].block[3].um_I.iw[4] ,
    \top_I.branch[22].block[3].um_I.iw[3] ,
    \top_I.branch[22].block[3].um_I.iw[2] ,
    \top_I.branch[22].block[3].um_I.iw[1] ,
    \top_I.branch[22].block[3].um_I.clk ,
    \top_I.branch[22].block[2].um_I.iw[17] ,
    \top_I.branch[22].block[2].um_I.iw[16] ,
    \top_I.branch[22].block[2].um_I.iw[15] ,
    \top_I.branch[22].block[2].um_I.iw[14] ,
    \top_I.branch[22].block[2].um_I.iw[13] ,
    \top_I.branch[22].block[2].um_I.iw[12] ,
    \top_I.branch[22].block[2].um_I.iw[11] ,
    \top_I.branch[22].block[2].um_I.iw[10] ,
    \top_I.branch[22].block[2].um_I.iw[9] ,
    \top_I.branch[22].block[2].um_I.iw[8] ,
    \top_I.branch[22].block[2].um_I.iw[7] ,
    \top_I.branch[22].block[2].um_I.iw[6] ,
    \top_I.branch[22].block[2].um_I.iw[5] ,
    \top_I.branch[22].block[2].um_I.iw[4] ,
    \top_I.branch[22].block[2].um_I.iw[3] ,
    \top_I.branch[22].block[2].um_I.iw[2] ,
    \top_I.branch[22].block[2].um_I.iw[1] ,
    \top_I.branch[22].block[2].um_I.clk ,
    \top_I.branch[22].block[1].um_I.iw[17] ,
    \top_I.branch[22].block[1].um_I.iw[16] ,
    \top_I.branch[22].block[1].um_I.iw[15] ,
    \top_I.branch[22].block[1].um_I.iw[14] ,
    \top_I.branch[22].block[1].um_I.iw[13] ,
    \top_I.branch[22].block[1].um_I.iw[12] ,
    \top_I.branch[22].block[1].um_I.iw[11] ,
    \top_I.branch[22].block[1].um_I.iw[10] ,
    \top_I.branch[22].block[1].um_I.iw[9] ,
    \top_I.branch[22].block[1].um_I.iw[8] ,
    \top_I.branch[22].block[1].um_I.iw[7] ,
    \top_I.branch[22].block[1].um_I.iw[6] ,
    \top_I.branch[22].block[1].um_I.iw[5] ,
    \top_I.branch[22].block[1].um_I.iw[4] ,
    \top_I.branch[22].block[1].um_I.iw[3] ,
    \top_I.branch[22].block[1].um_I.iw[2] ,
    \top_I.branch[22].block[1].um_I.iw[1] ,
    \top_I.branch[22].block[1].um_I.clk ,
    \top_I.branch[22].block[0].um_I.iw[17] ,
    \top_I.branch[22].block[0].um_I.iw[16] ,
    \top_I.branch[22].block[0].um_I.iw[15] ,
    \top_I.branch[22].block[0].um_I.iw[14] ,
    \top_I.branch[22].block[0].um_I.iw[13] ,
    \top_I.branch[22].block[0].um_I.iw[12] ,
    \top_I.branch[22].block[0].um_I.iw[11] ,
    \top_I.branch[22].block[0].um_I.iw[10] ,
    \top_I.branch[22].block[0].um_I.iw[9] ,
    \top_I.branch[22].block[0].um_I.iw[8] ,
    \top_I.branch[22].block[0].um_I.iw[7] ,
    \top_I.branch[22].block[0].um_I.iw[6] ,
    \top_I.branch[22].block[0].um_I.iw[5] ,
    \top_I.branch[22].block[0].um_I.iw[4] ,
    \top_I.branch[22].block[0].um_I.iw[3] ,
    \top_I.branch[22].block[0].um_I.iw[2] ,
    \top_I.branch[22].block[0].um_I.iw[1] ,
    \top_I.branch[22].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[15].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[14].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[13].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[12].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[11].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[10].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[9].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[8].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[7].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[6].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[5].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[4].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[3].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[2].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[1].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero ,
    \top_I.branch[22].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[22].block[15].um_I.pg_vdd ,
    \top_I.branch[22].block[14].um_I.pg_vdd ,
    \top_I.branch[22].block[13].um_I.pg_vdd ,
    \top_I.branch[22].block[12].um_I.pg_vdd ,
    \top_I.branch[22].block[11].um_I.pg_vdd ,
    \top_I.branch[22].block[10].um_I.pg_vdd ,
    \top_I.branch[22].block[9].um_I.pg_vdd ,
    \top_I.branch[22].block[8].um_I.pg_vdd ,
    \top_I.branch[22].block[7].um_I.pg_vdd ,
    \top_I.branch[22].block[6].um_I.pg_vdd ,
    \top_I.branch[22].block[5].um_I.pg_vdd ,
    \top_I.branch[22].block[4].um_I.pg_vdd ,
    \top_I.branch[22].block[3].um_I.pg_vdd ,
    \top_I.branch[22].block[2].um_I.pg_vdd ,
    \top_I.branch[22].block[1].um_I.pg_vdd ,
    \top_I.branch[22].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[23].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[23].l_addr[0] ),
    .k_zero(\top_I.branch[23].l_addr[2] ),
    .addr({\top_I.branch[23].l_addr[0] ,
    \top_I.branch[23].l_addr[2] ,
    \top_I.branch[23].l_addr[0] ,
    \top_I.branch[23].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[23].block[15].um_I.ena ,
    \top_I.branch[23].block[14].um_I.ena ,
    \top_I.branch[23].block[13].um_I.ena ,
    \top_I.branch[23].block[12].um_I.ena ,
    \top_I.branch[23].block[11].um_I.ena ,
    \top_I.branch[23].block[10].um_I.ena ,
    \top_I.branch[23].block[9].um_I.ena ,
    \top_I.branch[23].block[8].um_I.ena ,
    \top_I.branch[23].block[7].um_I.ena ,
    \top_I.branch[23].block[6].um_I.ena ,
    \top_I.branch[23].block[5].um_I.ena ,
    \top_I.branch[23].block[4].um_I.ena ,
    \top_I.branch[23].block[3].um_I.ena ,
    \top_I.branch[23].block[2].um_I.ena ,
    \top_I.branch[23].block[1].um_I.ena ,
    \top_I.branch[23].block[0].um_I.ena }),
    .um_iw({\top_I.branch[23].block[15].um_I.iw[17] ,
    \top_I.branch[23].block[15].um_I.iw[16] ,
    \top_I.branch[23].block[15].um_I.iw[15] ,
    \top_I.branch[23].block[15].um_I.iw[14] ,
    \top_I.branch[23].block[15].um_I.iw[13] ,
    \top_I.branch[23].block[15].um_I.iw[12] ,
    \top_I.branch[23].block[15].um_I.iw[11] ,
    \top_I.branch[23].block[15].um_I.iw[10] ,
    \top_I.branch[23].block[15].um_I.iw[9] ,
    \top_I.branch[23].block[15].um_I.iw[8] ,
    \top_I.branch[23].block[15].um_I.iw[7] ,
    \top_I.branch[23].block[15].um_I.iw[6] ,
    \top_I.branch[23].block[15].um_I.iw[5] ,
    \top_I.branch[23].block[15].um_I.iw[4] ,
    \top_I.branch[23].block[15].um_I.iw[3] ,
    \top_I.branch[23].block[15].um_I.iw[2] ,
    \top_I.branch[23].block[15].um_I.iw[1] ,
    \top_I.branch[23].block[15].um_I.clk ,
    \top_I.branch[23].block[14].um_I.iw[17] ,
    \top_I.branch[23].block[14].um_I.iw[16] ,
    \top_I.branch[23].block[14].um_I.iw[15] ,
    \top_I.branch[23].block[14].um_I.iw[14] ,
    \top_I.branch[23].block[14].um_I.iw[13] ,
    \top_I.branch[23].block[14].um_I.iw[12] ,
    \top_I.branch[23].block[14].um_I.iw[11] ,
    \top_I.branch[23].block[14].um_I.iw[10] ,
    \top_I.branch[23].block[14].um_I.iw[9] ,
    \top_I.branch[23].block[14].um_I.iw[8] ,
    \top_I.branch[23].block[14].um_I.iw[7] ,
    \top_I.branch[23].block[14].um_I.iw[6] ,
    \top_I.branch[23].block[14].um_I.iw[5] ,
    \top_I.branch[23].block[14].um_I.iw[4] ,
    \top_I.branch[23].block[14].um_I.iw[3] ,
    \top_I.branch[23].block[14].um_I.iw[2] ,
    \top_I.branch[23].block[14].um_I.iw[1] ,
    \top_I.branch[23].block[14].um_I.clk ,
    \top_I.branch[23].block[13].um_I.iw[17] ,
    \top_I.branch[23].block[13].um_I.iw[16] ,
    \top_I.branch[23].block[13].um_I.iw[15] ,
    \top_I.branch[23].block[13].um_I.iw[14] ,
    \top_I.branch[23].block[13].um_I.iw[13] ,
    \top_I.branch[23].block[13].um_I.iw[12] ,
    \top_I.branch[23].block[13].um_I.iw[11] ,
    \top_I.branch[23].block[13].um_I.iw[10] ,
    \top_I.branch[23].block[13].um_I.iw[9] ,
    \top_I.branch[23].block[13].um_I.iw[8] ,
    \top_I.branch[23].block[13].um_I.iw[7] ,
    \top_I.branch[23].block[13].um_I.iw[6] ,
    \top_I.branch[23].block[13].um_I.iw[5] ,
    \top_I.branch[23].block[13].um_I.iw[4] ,
    \top_I.branch[23].block[13].um_I.iw[3] ,
    \top_I.branch[23].block[13].um_I.iw[2] ,
    \top_I.branch[23].block[13].um_I.iw[1] ,
    \top_I.branch[23].block[13].um_I.clk ,
    \top_I.branch[23].block[12].um_I.iw[17] ,
    \top_I.branch[23].block[12].um_I.iw[16] ,
    \top_I.branch[23].block[12].um_I.iw[15] ,
    \top_I.branch[23].block[12].um_I.iw[14] ,
    \top_I.branch[23].block[12].um_I.iw[13] ,
    \top_I.branch[23].block[12].um_I.iw[12] ,
    \top_I.branch[23].block[12].um_I.iw[11] ,
    \top_I.branch[23].block[12].um_I.iw[10] ,
    \top_I.branch[23].block[12].um_I.iw[9] ,
    \top_I.branch[23].block[12].um_I.iw[8] ,
    \top_I.branch[23].block[12].um_I.iw[7] ,
    \top_I.branch[23].block[12].um_I.iw[6] ,
    \top_I.branch[23].block[12].um_I.iw[5] ,
    \top_I.branch[23].block[12].um_I.iw[4] ,
    \top_I.branch[23].block[12].um_I.iw[3] ,
    \top_I.branch[23].block[12].um_I.iw[2] ,
    \top_I.branch[23].block[12].um_I.iw[1] ,
    \top_I.branch[23].block[12].um_I.clk ,
    \top_I.branch[23].block[11].um_I.iw[17] ,
    \top_I.branch[23].block[11].um_I.iw[16] ,
    \top_I.branch[23].block[11].um_I.iw[15] ,
    \top_I.branch[23].block[11].um_I.iw[14] ,
    \top_I.branch[23].block[11].um_I.iw[13] ,
    \top_I.branch[23].block[11].um_I.iw[12] ,
    \top_I.branch[23].block[11].um_I.iw[11] ,
    \top_I.branch[23].block[11].um_I.iw[10] ,
    \top_I.branch[23].block[11].um_I.iw[9] ,
    \top_I.branch[23].block[11].um_I.iw[8] ,
    \top_I.branch[23].block[11].um_I.iw[7] ,
    \top_I.branch[23].block[11].um_I.iw[6] ,
    \top_I.branch[23].block[11].um_I.iw[5] ,
    \top_I.branch[23].block[11].um_I.iw[4] ,
    \top_I.branch[23].block[11].um_I.iw[3] ,
    \top_I.branch[23].block[11].um_I.iw[2] ,
    \top_I.branch[23].block[11].um_I.iw[1] ,
    \top_I.branch[23].block[11].um_I.clk ,
    \top_I.branch[23].block[10].um_I.iw[17] ,
    \top_I.branch[23].block[10].um_I.iw[16] ,
    \top_I.branch[23].block[10].um_I.iw[15] ,
    \top_I.branch[23].block[10].um_I.iw[14] ,
    \top_I.branch[23].block[10].um_I.iw[13] ,
    \top_I.branch[23].block[10].um_I.iw[12] ,
    \top_I.branch[23].block[10].um_I.iw[11] ,
    \top_I.branch[23].block[10].um_I.iw[10] ,
    \top_I.branch[23].block[10].um_I.iw[9] ,
    \top_I.branch[23].block[10].um_I.iw[8] ,
    \top_I.branch[23].block[10].um_I.iw[7] ,
    \top_I.branch[23].block[10].um_I.iw[6] ,
    \top_I.branch[23].block[10].um_I.iw[5] ,
    \top_I.branch[23].block[10].um_I.iw[4] ,
    \top_I.branch[23].block[10].um_I.iw[3] ,
    \top_I.branch[23].block[10].um_I.iw[2] ,
    \top_I.branch[23].block[10].um_I.iw[1] ,
    \top_I.branch[23].block[10].um_I.clk ,
    \top_I.branch[23].block[9].um_I.iw[17] ,
    \top_I.branch[23].block[9].um_I.iw[16] ,
    \top_I.branch[23].block[9].um_I.iw[15] ,
    \top_I.branch[23].block[9].um_I.iw[14] ,
    \top_I.branch[23].block[9].um_I.iw[13] ,
    \top_I.branch[23].block[9].um_I.iw[12] ,
    \top_I.branch[23].block[9].um_I.iw[11] ,
    \top_I.branch[23].block[9].um_I.iw[10] ,
    \top_I.branch[23].block[9].um_I.iw[9] ,
    \top_I.branch[23].block[9].um_I.iw[8] ,
    \top_I.branch[23].block[9].um_I.iw[7] ,
    \top_I.branch[23].block[9].um_I.iw[6] ,
    \top_I.branch[23].block[9].um_I.iw[5] ,
    \top_I.branch[23].block[9].um_I.iw[4] ,
    \top_I.branch[23].block[9].um_I.iw[3] ,
    \top_I.branch[23].block[9].um_I.iw[2] ,
    \top_I.branch[23].block[9].um_I.iw[1] ,
    \top_I.branch[23].block[9].um_I.clk ,
    \top_I.branch[23].block[8].um_I.iw[17] ,
    \top_I.branch[23].block[8].um_I.iw[16] ,
    \top_I.branch[23].block[8].um_I.iw[15] ,
    \top_I.branch[23].block[8].um_I.iw[14] ,
    \top_I.branch[23].block[8].um_I.iw[13] ,
    \top_I.branch[23].block[8].um_I.iw[12] ,
    \top_I.branch[23].block[8].um_I.iw[11] ,
    \top_I.branch[23].block[8].um_I.iw[10] ,
    \top_I.branch[23].block[8].um_I.iw[9] ,
    \top_I.branch[23].block[8].um_I.iw[8] ,
    \top_I.branch[23].block[8].um_I.iw[7] ,
    \top_I.branch[23].block[8].um_I.iw[6] ,
    \top_I.branch[23].block[8].um_I.iw[5] ,
    \top_I.branch[23].block[8].um_I.iw[4] ,
    \top_I.branch[23].block[8].um_I.iw[3] ,
    \top_I.branch[23].block[8].um_I.iw[2] ,
    \top_I.branch[23].block[8].um_I.iw[1] ,
    \top_I.branch[23].block[8].um_I.clk ,
    \top_I.branch[23].block[7].um_I.iw[17] ,
    \top_I.branch[23].block[7].um_I.iw[16] ,
    \top_I.branch[23].block[7].um_I.iw[15] ,
    \top_I.branch[23].block[7].um_I.iw[14] ,
    \top_I.branch[23].block[7].um_I.iw[13] ,
    \top_I.branch[23].block[7].um_I.iw[12] ,
    \top_I.branch[23].block[7].um_I.iw[11] ,
    \top_I.branch[23].block[7].um_I.iw[10] ,
    \top_I.branch[23].block[7].um_I.iw[9] ,
    \top_I.branch[23].block[7].um_I.iw[8] ,
    \top_I.branch[23].block[7].um_I.iw[7] ,
    \top_I.branch[23].block[7].um_I.iw[6] ,
    \top_I.branch[23].block[7].um_I.iw[5] ,
    \top_I.branch[23].block[7].um_I.iw[4] ,
    \top_I.branch[23].block[7].um_I.iw[3] ,
    \top_I.branch[23].block[7].um_I.iw[2] ,
    \top_I.branch[23].block[7].um_I.iw[1] ,
    \top_I.branch[23].block[7].um_I.clk ,
    \top_I.branch[23].block[6].um_I.iw[17] ,
    \top_I.branch[23].block[6].um_I.iw[16] ,
    \top_I.branch[23].block[6].um_I.iw[15] ,
    \top_I.branch[23].block[6].um_I.iw[14] ,
    \top_I.branch[23].block[6].um_I.iw[13] ,
    \top_I.branch[23].block[6].um_I.iw[12] ,
    \top_I.branch[23].block[6].um_I.iw[11] ,
    \top_I.branch[23].block[6].um_I.iw[10] ,
    \top_I.branch[23].block[6].um_I.iw[9] ,
    \top_I.branch[23].block[6].um_I.iw[8] ,
    \top_I.branch[23].block[6].um_I.iw[7] ,
    \top_I.branch[23].block[6].um_I.iw[6] ,
    \top_I.branch[23].block[6].um_I.iw[5] ,
    \top_I.branch[23].block[6].um_I.iw[4] ,
    \top_I.branch[23].block[6].um_I.iw[3] ,
    \top_I.branch[23].block[6].um_I.iw[2] ,
    \top_I.branch[23].block[6].um_I.iw[1] ,
    \top_I.branch[23].block[6].um_I.clk ,
    \top_I.branch[23].block[5].um_I.iw[17] ,
    \top_I.branch[23].block[5].um_I.iw[16] ,
    \top_I.branch[23].block[5].um_I.iw[15] ,
    \top_I.branch[23].block[5].um_I.iw[14] ,
    \top_I.branch[23].block[5].um_I.iw[13] ,
    \top_I.branch[23].block[5].um_I.iw[12] ,
    \top_I.branch[23].block[5].um_I.iw[11] ,
    \top_I.branch[23].block[5].um_I.iw[10] ,
    \top_I.branch[23].block[5].um_I.iw[9] ,
    \top_I.branch[23].block[5].um_I.iw[8] ,
    \top_I.branch[23].block[5].um_I.iw[7] ,
    \top_I.branch[23].block[5].um_I.iw[6] ,
    \top_I.branch[23].block[5].um_I.iw[5] ,
    \top_I.branch[23].block[5].um_I.iw[4] ,
    \top_I.branch[23].block[5].um_I.iw[3] ,
    \top_I.branch[23].block[5].um_I.iw[2] ,
    \top_I.branch[23].block[5].um_I.iw[1] ,
    \top_I.branch[23].block[5].um_I.clk ,
    \top_I.branch[23].block[4].um_I.iw[17] ,
    \top_I.branch[23].block[4].um_I.iw[16] ,
    \top_I.branch[23].block[4].um_I.iw[15] ,
    \top_I.branch[23].block[4].um_I.iw[14] ,
    \top_I.branch[23].block[4].um_I.iw[13] ,
    \top_I.branch[23].block[4].um_I.iw[12] ,
    \top_I.branch[23].block[4].um_I.iw[11] ,
    \top_I.branch[23].block[4].um_I.iw[10] ,
    \top_I.branch[23].block[4].um_I.iw[9] ,
    \top_I.branch[23].block[4].um_I.iw[8] ,
    \top_I.branch[23].block[4].um_I.iw[7] ,
    \top_I.branch[23].block[4].um_I.iw[6] ,
    \top_I.branch[23].block[4].um_I.iw[5] ,
    \top_I.branch[23].block[4].um_I.iw[4] ,
    \top_I.branch[23].block[4].um_I.iw[3] ,
    \top_I.branch[23].block[4].um_I.iw[2] ,
    \top_I.branch[23].block[4].um_I.iw[1] ,
    \top_I.branch[23].block[4].um_I.clk ,
    \top_I.branch[23].block[3].um_I.iw[17] ,
    \top_I.branch[23].block[3].um_I.iw[16] ,
    \top_I.branch[23].block[3].um_I.iw[15] ,
    \top_I.branch[23].block[3].um_I.iw[14] ,
    \top_I.branch[23].block[3].um_I.iw[13] ,
    \top_I.branch[23].block[3].um_I.iw[12] ,
    \top_I.branch[23].block[3].um_I.iw[11] ,
    \top_I.branch[23].block[3].um_I.iw[10] ,
    \top_I.branch[23].block[3].um_I.iw[9] ,
    \top_I.branch[23].block[3].um_I.iw[8] ,
    \top_I.branch[23].block[3].um_I.iw[7] ,
    \top_I.branch[23].block[3].um_I.iw[6] ,
    \top_I.branch[23].block[3].um_I.iw[5] ,
    \top_I.branch[23].block[3].um_I.iw[4] ,
    \top_I.branch[23].block[3].um_I.iw[3] ,
    \top_I.branch[23].block[3].um_I.iw[2] ,
    \top_I.branch[23].block[3].um_I.iw[1] ,
    \top_I.branch[23].block[3].um_I.clk ,
    \top_I.branch[23].block[2].um_I.iw[17] ,
    \top_I.branch[23].block[2].um_I.iw[16] ,
    \top_I.branch[23].block[2].um_I.iw[15] ,
    \top_I.branch[23].block[2].um_I.iw[14] ,
    \top_I.branch[23].block[2].um_I.iw[13] ,
    \top_I.branch[23].block[2].um_I.iw[12] ,
    \top_I.branch[23].block[2].um_I.iw[11] ,
    \top_I.branch[23].block[2].um_I.iw[10] ,
    \top_I.branch[23].block[2].um_I.iw[9] ,
    \top_I.branch[23].block[2].um_I.iw[8] ,
    \top_I.branch[23].block[2].um_I.iw[7] ,
    \top_I.branch[23].block[2].um_I.iw[6] ,
    \top_I.branch[23].block[2].um_I.iw[5] ,
    \top_I.branch[23].block[2].um_I.iw[4] ,
    \top_I.branch[23].block[2].um_I.iw[3] ,
    \top_I.branch[23].block[2].um_I.iw[2] ,
    \top_I.branch[23].block[2].um_I.iw[1] ,
    \top_I.branch[23].block[2].um_I.clk ,
    \top_I.branch[23].block[1].um_I.iw[17] ,
    \top_I.branch[23].block[1].um_I.iw[16] ,
    \top_I.branch[23].block[1].um_I.iw[15] ,
    \top_I.branch[23].block[1].um_I.iw[14] ,
    \top_I.branch[23].block[1].um_I.iw[13] ,
    \top_I.branch[23].block[1].um_I.iw[12] ,
    \top_I.branch[23].block[1].um_I.iw[11] ,
    \top_I.branch[23].block[1].um_I.iw[10] ,
    \top_I.branch[23].block[1].um_I.iw[9] ,
    \top_I.branch[23].block[1].um_I.iw[8] ,
    \top_I.branch[23].block[1].um_I.iw[7] ,
    \top_I.branch[23].block[1].um_I.iw[6] ,
    \top_I.branch[23].block[1].um_I.iw[5] ,
    \top_I.branch[23].block[1].um_I.iw[4] ,
    \top_I.branch[23].block[1].um_I.iw[3] ,
    \top_I.branch[23].block[1].um_I.iw[2] ,
    \top_I.branch[23].block[1].um_I.iw[1] ,
    \top_I.branch[23].block[1].um_I.clk ,
    \top_I.branch[23].block[0].um_I.iw[17] ,
    \top_I.branch[23].block[0].um_I.iw[16] ,
    \top_I.branch[23].block[0].um_I.iw[15] ,
    \top_I.branch[23].block[0].um_I.iw[14] ,
    \top_I.branch[23].block[0].um_I.iw[13] ,
    \top_I.branch[23].block[0].um_I.iw[12] ,
    \top_I.branch[23].block[0].um_I.iw[11] ,
    \top_I.branch[23].block[0].um_I.iw[10] ,
    \top_I.branch[23].block[0].um_I.iw[9] ,
    \top_I.branch[23].block[0].um_I.iw[8] ,
    \top_I.branch[23].block[0].um_I.iw[7] ,
    \top_I.branch[23].block[0].um_I.iw[6] ,
    \top_I.branch[23].block[0].um_I.iw[5] ,
    \top_I.branch[23].block[0].um_I.iw[4] ,
    \top_I.branch[23].block[0].um_I.iw[3] ,
    \top_I.branch[23].block[0].um_I.iw[2] ,
    \top_I.branch[23].block[0].um_I.iw[1] ,
    \top_I.branch[23].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[15].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[14].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[13].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[12].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[11].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[10].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[9].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[8].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[7].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[6].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[5].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[4].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[3].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[2].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[1].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero ,
    \top_I.branch[23].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[23].block[15].um_I.pg_vdd ,
    \top_I.branch[23].block[14].um_I.pg_vdd ,
    \top_I.branch[23].block[13].um_I.pg_vdd ,
    \top_I.branch[23].block[12].um_I.pg_vdd ,
    \top_I.branch[23].block[11].um_I.pg_vdd ,
    \top_I.branch[23].block[10].um_I.pg_vdd ,
    \top_I.branch[23].block[9].um_I.pg_vdd ,
    \top_I.branch[23].block[8].um_I.pg_vdd ,
    \top_I.branch[23].block[7].um_I.pg_vdd ,
    \top_I.branch[23].block[6].um_I.pg_vdd ,
    \top_I.branch[23].block[5].um_I.pg_vdd ,
    \top_I.branch[23].block[4].um_I.pg_vdd ,
    \top_I.branch[23].block[3].um_I.pg_vdd ,
    \top_I.branch[23].block[2].um_I.pg_vdd ,
    \top_I.branch[23].block[1].um_I.pg_vdd ,
    \top_I.branch[23].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[24].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[24].l_addr[2] ),
    .k_zero(\top_I.branch[24].l_addr[0] ),
    .addr({\top_I.branch[24].l_addr[2] ,
    \top_I.branch[24].l_addr[2] ,
    \top_I.branch[24].l_addr[0] ,
    \top_I.branch[24].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[24].block[15].um_I.ena ,
    \top_I.branch[24].block[14].um_I.ena ,
    \top_I.branch[24].block[13].um_I.ena ,
    \top_I.branch[24].block[12].um_I.ena ,
    \top_I.branch[24].block[11].um_I.ena ,
    \top_I.branch[24].block[10].um_I.ena ,
    \top_I.branch[24].block[9].um_I.ena ,
    \top_I.branch[24].block[8].um_I.ena ,
    \top_I.branch[24].block[7].um_I.ena ,
    \top_I.branch[24].block[6].um_I.ena ,
    \top_I.branch[24].block[5].um_I.ena ,
    \top_I.branch[24].block[4].um_I.ena ,
    \top_I.branch[24].block[3].um_I.ena ,
    \top_I.branch[24].block[2].um_I.ena ,
    \top_I.branch[24].block[1].um_I.ena ,
    \top_I.branch[24].block[0].um_I.ena }),
    .um_iw({\top_I.branch[24].block[15].um_I.iw[17] ,
    \top_I.branch[24].block[15].um_I.iw[16] ,
    \top_I.branch[24].block[15].um_I.iw[15] ,
    \top_I.branch[24].block[15].um_I.iw[14] ,
    \top_I.branch[24].block[15].um_I.iw[13] ,
    \top_I.branch[24].block[15].um_I.iw[12] ,
    \top_I.branch[24].block[15].um_I.iw[11] ,
    \top_I.branch[24].block[15].um_I.iw[10] ,
    \top_I.branch[24].block[15].um_I.iw[9] ,
    \top_I.branch[24].block[15].um_I.iw[8] ,
    \top_I.branch[24].block[15].um_I.iw[7] ,
    \top_I.branch[24].block[15].um_I.iw[6] ,
    \top_I.branch[24].block[15].um_I.iw[5] ,
    \top_I.branch[24].block[15].um_I.iw[4] ,
    \top_I.branch[24].block[15].um_I.iw[3] ,
    \top_I.branch[24].block[15].um_I.iw[2] ,
    \top_I.branch[24].block[15].um_I.iw[1] ,
    \top_I.branch[24].block[15].um_I.clk ,
    \top_I.branch[24].block[14].um_I.iw[17] ,
    \top_I.branch[24].block[14].um_I.iw[16] ,
    \top_I.branch[24].block[14].um_I.iw[15] ,
    \top_I.branch[24].block[14].um_I.iw[14] ,
    \top_I.branch[24].block[14].um_I.iw[13] ,
    \top_I.branch[24].block[14].um_I.iw[12] ,
    \top_I.branch[24].block[14].um_I.iw[11] ,
    \top_I.branch[24].block[14].um_I.iw[10] ,
    \top_I.branch[24].block[14].um_I.iw[9] ,
    \top_I.branch[24].block[14].um_I.iw[8] ,
    \top_I.branch[24].block[14].um_I.iw[7] ,
    \top_I.branch[24].block[14].um_I.iw[6] ,
    \top_I.branch[24].block[14].um_I.iw[5] ,
    \top_I.branch[24].block[14].um_I.iw[4] ,
    \top_I.branch[24].block[14].um_I.iw[3] ,
    \top_I.branch[24].block[14].um_I.iw[2] ,
    \top_I.branch[24].block[14].um_I.iw[1] ,
    \top_I.branch[24].block[14].um_I.clk ,
    \top_I.branch[24].block[13].um_I.iw[17] ,
    \top_I.branch[24].block[13].um_I.iw[16] ,
    \top_I.branch[24].block[13].um_I.iw[15] ,
    \top_I.branch[24].block[13].um_I.iw[14] ,
    \top_I.branch[24].block[13].um_I.iw[13] ,
    \top_I.branch[24].block[13].um_I.iw[12] ,
    \top_I.branch[24].block[13].um_I.iw[11] ,
    \top_I.branch[24].block[13].um_I.iw[10] ,
    \top_I.branch[24].block[13].um_I.iw[9] ,
    \top_I.branch[24].block[13].um_I.iw[8] ,
    \top_I.branch[24].block[13].um_I.iw[7] ,
    \top_I.branch[24].block[13].um_I.iw[6] ,
    \top_I.branch[24].block[13].um_I.iw[5] ,
    \top_I.branch[24].block[13].um_I.iw[4] ,
    \top_I.branch[24].block[13].um_I.iw[3] ,
    \top_I.branch[24].block[13].um_I.iw[2] ,
    \top_I.branch[24].block[13].um_I.iw[1] ,
    \top_I.branch[24].block[13].um_I.clk ,
    \top_I.branch[24].block[12].um_I.iw[17] ,
    \top_I.branch[24].block[12].um_I.iw[16] ,
    \top_I.branch[24].block[12].um_I.iw[15] ,
    \top_I.branch[24].block[12].um_I.iw[14] ,
    \top_I.branch[24].block[12].um_I.iw[13] ,
    \top_I.branch[24].block[12].um_I.iw[12] ,
    \top_I.branch[24].block[12].um_I.iw[11] ,
    \top_I.branch[24].block[12].um_I.iw[10] ,
    \top_I.branch[24].block[12].um_I.iw[9] ,
    \top_I.branch[24].block[12].um_I.iw[8] ,
    \top_I.branch[24].block[12].um_I.iw[7] ,
    \top_I.branch[24].block[12].um_I.iw[6] ,
    \top_I.branch[24].block[12].um_I.iw[5] ,
    \top_I.branch[24].block[12].um_I.iw[4] ,
    \top_I.branch[24].block[12].um_I.iw[3] ,
    \top_I.branch[24].block[12].um_I.iw[2] ,
    \top_I.branch[24].block[12].um_I.iw[1] ,
    \top_I.branch[24].block[12].um_I.clk ,
    \top_I.branch[24].block[11].um_I.iw[17] ,
    \top_I.branch[24].block[11].um_I.iw[16] ,
    \top_I.branch[24].block[11].um_I.iw[15] ,
    \top_I.branch[24].block[11].um_I.iw[14] ,
    \top_I.branch[24].block[11].um_I.iw[13] ,
    \top_I.branch[24].block[11].um_I.iw[12] ,
    \top_I.branch[24].block[11].um_I.iw[11] ,
    \top_I.branch[24].block[11].um_I.iw[10] ,
    \top_I.branch[24].block[11].um_I.iw[9] ,
    \top_I.branch[24].block[11].um_I.iw[8] ,
    \top_I.branch[24].block[11].um_I.iw[7] ,
    \top_I.branch[24].block[11].um_I.iw[6] ,
    \top_I.branch[24].block[11].um_I.iw[5] ,
    \top_I.branch[24].block[11].um_I.iw[4] ,
    \top_I.branch[24].block[11].um_I.iw[3] ,
    \top_I.branch[24].block[11].um_I.iw[2] ,
    \top_I.branch[24].block[11].um_I.iw[1] ,
    \top_I.branch[24].block[11].um_I.clk ,
    \top_I.branch[24].block[10].um_I.iw[17] ,
    \top_I.branch[24].block[10].um_I.iw[16] ,
    \top_I.branch[24].block[10].um_I.iw[15] ,
    \top_I.branch[24].block[10].um_I.iw[14] ,
    \top_I.branch[24].block[10].um_I.iw[13] ,
    \top_I.branch[24].block[10].um_I.iw[12] ,
    \top_I.branch[24].block[10].um_I.iw[11] ,
    \top_I.branch[24].block[10].um_I.iw[10] ,
    \top_I.branch[24].block[10].um_I.iw[9] ,
    \top_I.branch[24].block[10].um_I.iw[8] ,
    \top_I.branch[24].block[10].um_I.iw[7] ,
    \top_I.branch[24].block[10].um_I.iw[6] ,
    \top_I.branch[24].block[10].um_I.iw[5] ,
    \top_I.branch[24].block[10].um_I.iw[4] ,
    \top_I.branch[24].block[10].um_I.iw[3] ,
    \top_I.branch[24].block[10].um_I.iw[2] ,
    \top_I.branch[24].block[10].um_I.iw[1] ,
    \top_I.branch[24].block[10].um_I.clk ,
    \top_I.branch[24].block[9].um_I.iw[17] ,
    \top_I.branch[24].block[9].um_I.iw[16] ,
    \top_I.branch[24].block[9].um_I.iw[15] ,
    \top_I.branch[24].block[9].um_I.iw[14] ,
    \top_I.branch[24].block[9].um_I.iw[13] ,
    \top_I.branch[24].block[9].um_I.iw[12] ,
    \top_I.branch[24].block[9].um_I.iw[11] ,
    \top_I.branch[24].block[9].um_I.iw[10] ,
    \top_I.branch[24].block[9].um_I.iw[9] ,
    \top_I.branch[24].block[9].um_I.iw[8] ,
    \top_I.branch[24].block[9].um_I.iw[7] ,
    \top_I.branch[24].block[9].um_I.iw[6] ,
    \top_I.branch[24].block[9].um_I.iw[5] ,
    \top_I.branch[24].block[9].um_I.iw[4] ,
    \top_I.branch[24].block[9].um_I.iw[3] ,
    \top_I.branch[24].block[9].um_I.iw[2] ,
    \top_I.branch[24].block[9].um_I.iw[1] ,
    \top_I.branch[24].block[9].um_I.clk ,
    \top_I.branch[24].block[8].um_I.iw[17] ,
    \top_I.branch[24].block[8].um_I.iw[16] ,
    \top_I.branch[24].block[8].um_I.iw[15] ,
    \top_I.branch[24].block[8].um_I.iw[14] ,
    \top_I.branch[24].block[8].um_I.iw[13] ,
    \top_I.branch[24].block[8].um_I.iw[12] ,
    \top_I.branch[24].block[8].um_I.iw[11] ,
    \top_I.branch[24].block[8].um_I.iw[10] ,
    \top_I.branch[24].block[8].um_I.iw[9] ,
    \top_I.branch[24].block[8].um_I.iw[8] ,
    \top_I.branch[24].block[8].um_I.iw[7] ,
    \top_I.branch[24].block[8].um_I.iw[6] ,
    \top_I.branch[24].block[8].um_I.iw[5] ,
    \top_I.branch[24].block[8].um_I.iw[4] ,
    \top_I.branch[24].block[8].um_I.iw[3] ,
    \top_I.branch[24].block[8].um_I.iw[2] ,
    \top_I.branch[24].block[8].um_I.iw[1] ,
    \top_I.branch[24].block[8].um_I.clk ,
    \top_I.branch[24].block[7].um_I.iw[17] ,
    \top_I.branch[24].block[7].um_I.iw[16] ,
    \top_I.branch[24].block[7].um_I.iw[15] ,
    \top_I.branch[24].block[7].um_I.iw[14] ,
    \top_I.branch[24].block[7].um_I.iw[13] ,
    \top_I.branch[24].block[7].um_I.iw[12] ,
    \top_I.branch[24].block[7].um_I.iw[11] ,
    \top_I.branch[24].block[7].um_I.iw[10] ,
    \top_I.branch[24].block[7].um_I.iw[9] ,
    \top_I.branch[24].block[7].um_I.iw[8] ,
    \top_I.branch[24].block[7].um_I.iw[7] ,
    \top_I.branch[24].block[7].um_I.iw[6] ,
    \top_I.branch[24].block[7].um_I.iw[5] ,
    \top_I.branch[24].block[7].um_I.iw[4] ,
    \top_I.branch[24].block[7].um_I.iw[3] ,
    \top_I.branch[24].block[7].um_I.iw[2] ,
    \top_I.branch[24].block[7].um_I.iw[1] ,
    \top_I.branch[24].block[7].um_I.clk ,
    \top_I.branch[24].block[6].um_I.iw[17] ,
    \top_I.branch[24].block[6].um_I.iw[16] ,
    \top_I.branch[24].block[6].um_I.iw[15] ,
    \top_I.branch[24].block[6].um_I.iw[14] ,
    \top_I.branch[24].block[6].um_I.iw[13] ,
    \top_I.branch[24].block[6].um_I.iw[12] ,
    \top_I.branch[24].block[6].um_I.iw[11] ,
    \top_I.branch[24].block[6].um_I.iw[10] ,
    \top_I.branch[24].block[6].um_I.iw[9] ,
    \top_I.branch[24].block[6].um_I.iw[8] ,
    \top_I.branch[24].block[6].um_I.iw[7] ,
    \top_I.branch[24].block[6].um_I.iw[6] ,
    \top_I.branch[24].block[6].um_I.iw[5] ,
    \top_I.branch[24].block[6].um_I.iw[4] ,
    \top_I.branch[24].block[6].um_I.iw[3] ,
    \top_I.branch[24].block[6].um_I.iw[2] ,
    \top_I.branch[24].block[6].um_I.iw[1] ,
    \top_I.branch[24].block[6].um_I.clk ,
    \top_I.branch[24].block[5].um_I.iw[17] ,
    \top_I.branch[24].block[5].um_I.iw[16] ,
    \top_I.branch[24].block[5].um_I.iw[15] ,
    \top_I.branch[24].block[5].um_I.iw[14] ,
    \top_I.branch[24].block[5].um_I.iw[13] ,
    \top_I.branch[24].block[5].um_I.iw[12] ,
    \top_I.branch[24].block[5].um_I.iw[11] ,
    \top_I.branch[24].block[5].um_I.iw[10] ,
    \top_I.branch[24].block[5].um_I.iw[9] ,
    \top_I.branch[24].block[5].um_I.iw[8] ,
    \top_I.branch[24].block[5].um_I.iw[7] ,
    \top_I.branch[24].block[5].um_I.iw[6] ,
    \top_I.branch[24].block[5].um_I.iw[5] ,
    \top_I.branch[24].block[5].um_I.iw[4] ,
    \top_I.branch[24].block[5].um_I.iw[3] ,
    \top_I.branch[24].block[5].um_I.iw[2] ,
    \top_I.branch[24].block[5].um_I.iw[1] ,
    \top_I.branch[24].block[5].um_I.clk ,
    \top_I.branch[24].block[4].um_I.iw[17] ,
    \top_I.branch[24].block[4].um_I.iw[16] ,
    \top_I.branch[24].block[4].um_I.iw[15] ,
    \top_I.branch[24].block[4].um_I.iw[14] ,
    \top_I.branch[24].block[4].um_I.iw[13] ,
    \top_I.branch[24].block[4].um_I.iw[12] ,
    \top_I.branch[24].block[4].um_I.iw[11] ,
    \top_I.branch[24].block[4].um_I.iw[10] ,
    \top_I.branch[24].block[4].um_I.iw[9] ,
    \top_I.branch[24].block[4].um_I.iw[8] ,
    \top_I.branch[24].block[4].um_I.iw[7] ,
    \top_I.branch[24].block[4].um_I.iw[6] ,
    \top_I.branch[24].block[4].um_I.iw[5] ,
    \top_I.branch[24].block[4].um_I.iw[4] ,
    \top_I.branch[24].block[4].um_I.iw[3] ,
    \top_I.branch[24].block[4].um_I.iw[2] ,
    \top_I.branch[24].block[4].um_I.iw[1] ,
    \top_I.branch[24].block[4].um_I.clk ,
    \top_I.branch[24].block[3].um_I.iw[17] ,
    \top_I.branch[24].block[3].um_I.iw[16] ,
    \top_I.branch[24].block[3].um_I.iw[15] ,
    \top_I.branch[24].block[3].um_I.iw[14] ,
    \top_I.branch[24].block[3].um_I.iw[13] ,
    \top_I.branch[24].block[3].um_I.iw[12] ,
    \top_I.branch[24].block[3].um_I.iw[11] ,
    \top_I.branch[24].block[3].um_I.iw[10] ,
    \top_I.branch[24].block[3].um_I.iw[9] ,
    \top_I.branch[24].block[3].um_I.iw[8] ,
    \top_I.branch[24].block[3].um_I.iw[7] ,
    \top_I.branch[24].block[3].um_I.iw[6] ,
    \top_I.branch[24].block[3].um_I.iw[5] ,
    \top_I.branch[24].block[3].um_I.iw[4] ,
    \top_I.branch[24].block[3].um_I.iw[3] ,
    \top_I.branch[24].block[3].um_I.iw[2] ,
    \top_I.branch[24].block[3].um_I.iw[1] ,
    \top_I.branch[24].block[3].um_I.clk ,
    \top_I.branch[24].block[2].um_I.iw[17] ,
    \top_I.branch[24].block[2].um_I.iw[16] ,
    \top_I.branch[24].block[2].um_I.iw[15] ,
    \top_I.branch[24].block[2].um_I.iw[14] ,
    \top_I.branch[24].block[2].um_I.iw[13] ,
    \top_I.branch[24].block[2].um_I.iw[12] ,
    \top_I.branch[24].block[2].um_I.iw[11] ,
    \top_I.branch[24].block[2].um_I.iw[10] ,
    \top_I.branch[24].block[2].um_I.iw[9] ,
    \top_I.branch[24].block[2].um_I.iw[8] ,
    \top_I.branch[24].block[2].um_I.iw[7] ,
    \top_I.branch[24].block[2].um_I.iw[6] ,
    \top_I.branch[24].block[2].um_I.iw[5] ,
    \top_I.branch[24].block[2].um_I.iw[4] ,
    \top_I.branch[24].block[2].um_I.iw[3] ,
    \top_I.branch[24].block[2].um_I.iw[2] ,
    \top_I.branch[24].block[2].um_I.iw[1] ,
    \top_I.branch[24].block[2].um_I.clk ,
    \top_I.branch[24].block[1].um_I.iw[17] ,
    \top_I.branch[24].block[1].um_I.iw[16] ,
    \top_I.branch[24].block[1].um_I.iw[15] ,
    \top_I.branch[24].block[1].um_I.iw[14] ,
    \top_I.branch[24].block[1].um_I.iw[13] ,
    \top_I.branch[24].block[1].um_I.iw[12] ,
    \top_I.branch[24].block[1].um_I.iw[11] ,
    \top_I.branch[24].block[1].um_I.iw[10] ,
    \top_I.branch[24].block[1].um_I.iw[9] ,
    \top_I.branch[24].block[1].um_I.iw[8] ,
    \top_I.branch[24].block[1].um_I.iw[7] ,
    \top_I.branch[24].block[1].um_I.iw[6] ,
    \top_I.branch[24].block[1].um_I.iw[5] ,
    \top_I.branch[24].block[1].um_I.iw[4] ,
    \top_I.branch[24].block[1].um_I.iw[3] ,
    \top_I.branch[24].block[1].um_I.iw[2] ,
    \top_I.branch[24].block[1].um_I.iw[1] ,
    \top_I.branch[24].block[1].um_I.clk ,
    \top_I.branch[24].block[0].um_I.iw[17] ,
    \top_I.branch[24].block[0].um_I.iw[16] ,
    \top_I.branch[24].block[0].um_I.iw[15] ,
    \top_I.branch[24].block[0].um_I.iw[14] ,
    \top_I.branch[24].block[0].um_I.iw[13] ,
    \top_I.branch[24].block[0].um_I.iw[12] ,
    \top_I.branch[24].block[0].um_I.iw[11] ,
    \top_I.branch[24].block[0].um_I.iw[10] ,
    \top_I.branch[24].block[0].um_I.iw[9] ,
    \top_I.branch[24].block[0].um_I.iw[8] ,
    \top_I.branch[24].block[0].um_I.iw[7] ,
    \top_I.branch[24].block[0].um_I.iw[6] ,
    \top_I.branch[24].block[0].um_I.iw[5] ,
    \top_I.branch[24].block[0].um_I.iw[4] ,
    \top_I.branch[24].block[0].um_I.iw[3] ,
    \top_I.branch[24].block[0].um_I.iw[2] ,
    \top_I.branch[24].block[0].um_I.iw[1] ,
    \top_I.branch[24].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[15].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[14].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[13].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[12].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[11].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[10].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[9].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[8].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[7].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[6].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[5].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[4].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[3].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[2].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[1].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero ,
    \top_I.branch[24].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[24].block[15].um_I.pg_vdd ,
    \top_I.branch[24].block[14].um_I.pg_vdd ,
    \top_I.branch[24].block[13].um_I.pg_vdd ,
    \top_I.branch[24].block[12].um_I.pg_vdd ,
    \top_I.branch[24].block[11].um_I.pg_vdd ,
    \top_I.branch[24].block[10].um_I.pg_vdd ,
    \top_I.branch[24].block[9].um_I.pg_vdd ,
    \top_I.branch[24].block[8].um_I.pg_vdd ,
    \top_I.branch[24].block[7].um_I.pg_vdd ,
    \top_I.branch[24].block[6].um_I.pg_vdd ,
    \top_I.branch[24].block[5].um_I.pg_vdd ,
    \top_I.branch[24].block[4].um_I.pg_vdd ,
    \top_I.branch[24].block[3].um_I.pg_vdd ,
    \top_I.branch[24].block[2].um_I.pg_vdd ,
    \top_I.branch[24].block[1].um_I.pg_vdd ,
    \top_I.branch[24].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[25].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[25].l_addr[2] ),
    .k_zero(\top_I.branch[25].l_addr[0] ),
    .addr({\top_I.branch[25].l_addr[2] ,
    \top_I.branch[25].l_addr[2] ,
    \top_I.branch[25].l_addr[0] ,
    \top_I.branch[25].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[25].block[15].um_I.ena ,
    \top_I.branch[25].block[14].um_I.ena ,
    \top_I.branch[25].block[13].um_I.ena ,
    \top_I.branch[25].block[12].um_I.ena ,
    \top_I.branch[25].block[11].um_I.ena ,
    \top_I.branch[25].block[10].um_I.ena ,
    \top_I.branch[25].block[9].um_I.ena ,
    \top_I.branch[25].block[8].um_I.ena ,
    \top_I.branch[25].block[7].um_I.ena ,
    \top_I.branch[25].block[6].um_I.ena ,
    \top_I.branch[25].block[5].um_I.ena ,
    \top_I.branch[25].block[4].um_I.ena ,
    \top_I.branch[25].block[3].um_I.ena ,
    \top_I.branch[25].block[2].um_I.ena ,
    \top_I.branch[25].block[1].um_I.ena ,
    \top_I.branch[25].block[0].um_I.ena }),
    .um_iw({\top_I.branch[25].block[15].um_I.iw[17] ,
    \top_I.branch[25].block[15].um_I.iw[16] ,
    \top_I.branch[25].block[15].um_I.iw[15] ,
    \top_I.branch[25].block[15].um_I.iw[14] ,
    \top_I.branch[25].block[15].um_I.iw[13] ,
    \top_I.branch[25].block[15].um_I.iw[12] ,
    \top_I.branch[25].block[15].um_I.iw[11] ,
    \top_I.branch[25].block[15].um_I.iw[10] ,
    \top_I.branch[25].block[15].um_I.iw[9] ,
    \top_I.branch[25].block[15].um_I.iw[8] ,
    \top_I.branch[25].block[15].um_I.iw[7] ,
    \top_I.branch[25].block[15].um_I.iw[6] ,
    \top_I.branch[25].block[15].um_I.iw[5] ,
    \top_I.branch[25].block[15].um_I.iw[4] ,
    \top_I.branch[25].block[15].um_I.iw[3] ,
    \top_I.branch[25].block[15].um_I.iw[2] ,
    \top_I.branch[25].block[15].um_I.iw[1] ,
    \top_I.branch[25].block[15].um_I.clk ,
    \top_I.branch[25].block[14].um_I.iw[17] ,
    \top_I.branch[25].block[14].um_I.iw[16] ,
    \top_I.branch[25].block[14].um_I.iw[15] ,
    \top_I.branch[25].block[14].um_I.iw[14] ,
    \top_I.branch[25].block[14].um_I.iw[13] ,
    \top_I.branch[25].block[14].um_I.iw[12] ,
    \top_I.branch[25].block[14].um_I.iw[11] ,
    \top_I.branch[25].block[14].um_I.iw[10] ,
    \top_I.branch[25].block[14].um_I.iw[9] ,
    \top_I.branch[25].block[14].um_I.iw[8] ,
    \top_I.branch[25].block[14].um_I.iw[7] ,
    \top_I.branch[25].block[14].um_I.iw[6] ,
    \top_I.branch[25].block[14].um_I.iw[5] ,
    \top_I.branch[25].block[14].um_I.iw[4] ,
    \top_I.branch[25].block[14].um_I.iw[3] ,
    \top_I.branch[25].block[14].um_I.iw[2] ,
    \top_I.branch[25].block[14].um_I.iw[1] ,
    \top_I.branch[25].block[14].um_I.clk ,
    \top_I.branch[25].block[13].um_I.iw[17] ,
    \top_I.branch[25].block[13].um_I.iw[16] ,
    \top_I.branch[25].block[13].um_I.iw[15] ,
    \top_I.branch[25].block[13].um_I.iw[14] ,
    \top_I.branch[25].block[13].um_I.iw[13] ,
    \top_I.branch[25].block[13].um_I.iw[12] ,
    \top_I.branch[25].block[13].um_I.iw[11] ,
    \top_I.branch[25].block[13].um_I.iw[10] ,
    \top_I.branch[25].block[13].um_I.iw[9] ,
    \top_I.branch[25].block[13].um_I.iw[8] ,
    \top_I.branch[25].block[13].um_I.iw[7] ,
    \top_I.branch[25].block[13].um_I.iw[6] ,
    \top_I.branch[25].block[13].um_I.iw[5] ,
    \top_I.branch[25].block[13].um_I.iw[4] ,
    \top_I.branch[25].block[13].um_I.iw[3] ,
    \top_I.branch[25].block[13].um_I.iw[2] ,
    \top_I.branch[25].block[13].um_I.iw[1] ,
    \top_I.branch[25].block[13].um_I.clk ,
    \top_I.branch[25].block[12].um_I.iw[17] ,
    \top_I.branch[25].block[12].um_I.iw[16] ,
    \top_I.branch[25].block[12].um_I.iw[15] ,
    \top_I.branch[25].block[12].um_I.iw[14] ,
    \top_I.branch[25].block[12].um_I.iw[13] ,
    \top_I.branch[25].block[12].um_I.iw[12] ,
    \top_I.branch[25].block[12].um_I.iw[11] ,
    \top_I.branch[25].block[12].um_I.iw[10] ,
    \top_I.branch[25].block[12].um_I.iw[9] ,
    \top_I.branch[25].block[12].um_I.iw[8] ,
    \top_I.branch[25].block[12].um_I.iw[7] ,
    \top_I.branch[25].block[12].um_I.iw[6] ,
    \top_I.branch[25].block[12].um_I.iw[5] ,
    \top_I.branch[25].block[12].um_I.iw[4] ,
    \top_I.branch[25].block[12].um_I.iw[3] ,
    \top_I.branch[25].block[12].um_I.iw[2] ,
    \top_I.branch[25].block[12].um_I.iw[1] ,
    \top_I.branch[25].block[12].um_I.clk ,
    \top_I.branch[25].block[11].um_I.iw[17] ,
    \top_I.branch[25].block[11].um_I.iw[16] ,
    \top_I.branch[25].block[11].um_I.iw[15] ,
    \top_I.branch[25].block[11].um_I.iw[14] ,
    \top_I.branch[25].block[11].um_I.iw[13] ,
    \top_I.branch[25].block[11].um_I.iw[12] ,
    \top_I.branch[25].block[11].um_I.iw[11] ,
    \top_I.branch[25].block[11].um_I.iw[10] ,
    \top_I.branch[25].block[11].um_I.iw[9] ,
    \top_I.branch[25].block[11].um_I.iw[8] ,
    \top_I.branch[25].block[11].um_I.iw[7] ,
    \top_I.branch[25].block[11].um_I.iw[6] ,
    \top_I.branch[25].block[11].um_I.iw[5] ,
    \top_I.branch[25].block[11].um_I.iw[4] ,
    \top_I.branch[25].block[11].um_I.iw[3] ,
    \top_I.branch[25].block[11].um_I.iw[2] ,
    \top_I.branch[25].block[11].um_I.iw[1] ,
    \top_I.branch[25].block[11].um_I.clk ,
    \top_I.branch[25].block[10].um_I.iw[17] ,
    \top_I.branch[25].block[10].um_I.iw[16] ,
    \top_I.branch[25].block[10].um_I.iw[15] ,
    \top_I.branch[25].block[10].um_I.iw[14] ,
    \top_I.branch[25].block[10].um_I.iw[13] ,
    \top_I.branch[25].block[10].um_I.iw[12] ,
    \top_I.branch[25].block[10].um_I.iw[11] ,
    \top_I.branch[25].block[10].um_I.iw[10] ,
    \top_I.branch[25].block[10].um_I.iw[9] ,
    \top_I.branch[25].block[10].um_I.iw[8] ,
    \top_I.branch[25].block[10].um_I.iw[7] ,
    \top_I.branch[25].block[10].um_I.iw[6] ,
    \top_I.branch[25].block[10].um_I.iw[5] ,
    \top_I.branch[25].block[10].um_I.iw[4] ,
    \top_I.branch[25].block[10].um_I.iw[3] ,
    \top_I.branch[25].block[10].um_I.iw[2] ,
    \top_I.branch[25].block[10].um_I.iw[1] ,
    \top_I.branch[25].block[10].um_I.clk ,
    \top_I.branch[25].block[9].um_I.iw[17] ,
    \top_I.branch[25].block[9].um_I.iw[16] ,
    \top_I.branch[25].block[9].um_I.iw[15] ,
    \top_I.branch[25].block[9].um_I.iw[14] ,
    \top_I.branch[25].block[9].um_I.iw[13] ,
    \top_I.branch[25].block[9].um_I.iw[12] ,
    \top_I.branch[25].block[9].um_I.iw[11] ,
    \top_I.branch[25].block[9].um_I.iw[10] ,
    \top_I.branch[25].block[9].um_I.iw[9] ,
    \top_I.branch[25].block[9].um_I.iw[8] ,
    \top_I.branch[25].block[9].um_I.iw[7] ,
    \top_I.branch[25].block[9].um_I.iw[6] ,
    \top_I.branch[25].block[9].um_I.iw[5] ,
    \top_I.branch[25].block[9].um_I.iw[4] ,
    \top_I.branch[25].block[9].um_I.iw[3] ,
    \top_I.branch[25].block[9].um_I.iw[2] ,
    \top_I.branch[25].block[9].um_I.iw[1] ,
    \top_I.branch[25].block[9].um_I.clk ,
    \top_I.branch[25].block[8].um_I.iw[17] ,
    \top_I.branch[25].block[8].um_I.iw[16] ,
    \top_I.branch[25].block[8].um_I.iw[15] ,
    \top_I.branch[25].block[8].um_I.iw[14] ,
    \top_I.branch[25].block[8].um_I.iw[13] ,
    \top_I.branch[25].block[8].um_I.iw[12] ,
    \top_I.branch[25].block[8].um_I.iw[11] ,
    \top_I.branch[25].block[8].um_I.iw[10] ,
    \top_I.branch[25].block[8].um_I.iw[9] ,
    \top_I.branch[25].block[8].um_I.iw[8] ,
    \top_I.branch[25].block[8].um_I.iw[7] ,
    \top_I.branch[25].block[8].um_I.iw[6] ,
    \top_I.branch[25].block[8].um_I.iw[5] ,
    \top_I.branch[25].block[8].um_I.iw[4] ,
    \top_I.branch[25].block[8].um_I.iw[3] ,
    \top_I.branch[25].block[8].um_I.iw[2] ,
    \top_I.branch[25].block[8].um_I.iw[1] ,
    \top_I.branch[25].block[8].um_I.clk ,
    \top_I.branch[25].block[7].um_I.iw[17] ,
    \top_I.branch[25].block[7].um_I.iw[16] ,
    \top_I.branch[25].block[7].um_I.iw[15] ,
    \top_I.branch[25].block[7].um_I.iw[14] ,
    \top_I.branch[25].block[7].um_I.iw[13] ,
    \top_I.branch[25].block[7].um_I.iw[12] ,
    \top_I.branch[25].block[7].um_I.iw[11] ,
    \top_I.branch[25].block[7].um_I.iw[10] ,
    \top_I.branch[25].block[7].um_I.iw[9] ,
    \top_I.branch[25].block[7].um_I.iw[8] ,
    \top_I.branch[25].block[7].um_I.iw[7] ,
    \top_I.branch[25].block[7].um_I.iw[6] ,
    \top_I.branch[25].block[7].um_I.iw[5] ,
    \top_I.branch[25].block[7].um_I.iw[4] ,
    \top_I.branch[25].block[7].um_I.iw[3] ,
    \top_I.branch[25].block[7].um_I.iw[2] ,
    \top_I.branch[25].block[7].um_I.iw[1] ,
    \top_I.branch[25].block[7].um_I.clk ,
    \top_I.branch[25].block[6].um_I.iw[17] ,
    \top_I.branch[25].block[6].um_I.iw[16] ,
    \top_I.branch[25].block[6].um_I.iw[15] ,
    \top_I.branch[25].block[6].um_I.iw[14] ,
    \top_I.branch[25].block[6].um_I.iw[13] ,
    \top_I.branch[25].block[6].um_I.iw[12] ,
    \top_I.branch[25].block[6].um_I.iw[11] ,
    \top_I.branch[25].block[6].um_I.iw[10] ,
    \top_I.branch[25].block[6].um_I.iw[9] ,
    \top_I.branch[25].block[6].um_I.iw[8] ,
    \top_I.branch[25].block[6].um_I.iw[7] ,
    \top_I.branch[25].block[6].um_I.iw[6] ,
    \top_I.branch[25].block[6].um_I.iw[5] ,
    \top_I.branch[25].block[6].um_I.iw[4] ,
    \top_I.branch[25].block[6].um_I.iw[3] ,
    \top_I.branch[25].block[6].um_I.iw[2] ,
    \top_I.branch[25].block[6].um_I.iw[1] ,
    \top_I.branch[25].block[6].um_I.clk ,
    \top_I.branch[25].block[5].um_I.iw[17] ,
    \top_I.branch[25].block[5].um_I.iw[16] ,
    \top_I.branch[25].block[5].um_I.iw[15] ,
    \top_I.branch[25].block[5].um_I.iw[14] ,
    \top_I.branch[25].block[5].um_I.iw[13] ,
    \top_I.branch[25].block[5].um_I.iw[12] ,
    \top_I.branch[25].block[5].um_I.iw[11] ,
    \top_I.branch[25].block[5].um_I.iw[10] ,
    \top_I.branch[25].block[5].um_I.iw[9] ,
    \top_I.branch[25].block[5].um_I.iw[8] ,
    \top_I.branch[25].block[5].um_I.iw[7] ,
    \top_I.branch[25].block[5].um_I.iw[6] ,
    \top_I.branch[25].block[5].um_I.iw[5] ,
    \top_I.branch[25].block[5].um_I.iw[4] ,
    \top_I.branch[25].block[5].um_I.iw[3] ,
    \top_I.branch[25].block[5].um_I.iw[2] ,
    \top_I.branch[25].block[5].um_I.iw[1] ,
    \top_I.branch[25].block[5].um_I.clk ,
    \top_I.branch[25].block[4].um_I.iw[17] ,
    \top_I.branch[25].block[4].um_I.iw[16] ,
    \top_I.branch[25].block[4].um_I.iw[15] ,
    \top_I.branch[25].block[4].um_I.iw[14] ,
    \top_I.branch[25].block[4].um_I.iw[13] ,
    \top_I.branch[25].block[4].um_I.iw[12] ,
    \top_I.branch[25].block[4].um_I.iw[11] ,
    \top_I.branch[25].block[4].um_I.iw[10] ,
    \top_I.branch[25].block[4].um_I.iw[9] ,
    \top_I.branch[25].block[4].um_I.iw[8] ,
    \top_I.branch[25].block[4].um_I.iw[7] ,
    \top_I.branch[25].block[4].um_I.iw[6] ,
    \top_I.branch[25].block[4].um_I.iw[5] ,
    \top_I.branch[25].block[4].um_I.iw[4] ,
    \top_I.branch[25].block[4].um_I.iw[3] ,
    \top_I.branch[25].block[4].um_I.iw[2] ,
    \top_I.branch[25].block[4].um_I.iw[1] ,
    \top_I.branch[25].block[4].um_I.clk ,
    \top_I.branch[25].block[3].um_I.iw[17] ,
    \top_I.branch[25].block[3].um_I.iw[16] ,
    \top_I.branch[25].block[3].um_I.iw[15] ,
    \top_I.branch[25].block[3].um_I.iw[14] ,
    \top_I.branch[25].block[3].um_I.iw[13] ,
    \top_I.branch[25].block[3].um_I.iw[12] ,
    \top_I.branch[25].block[3].um_I.iw[11] ,
    \top_I.branch[25].block[3].um_I.iw[10] ,
    \top_I.branch[25].block[3].um_I.iw[9] ,
    \top_I.branch[25].block[3].um_I.iw[8] ,
    \top_I.branch[25].block[3].um_I.iw[7] ,
    \top_I.branch[25].block[3].um_I.iw[6] ,
    \top_I.branch[25].block[3].um_I.iw[5] ,
    \top_I.branch[25].block[3].um_I.iw[4] ,
    \top_I.branch[25].block[3].um_I.iw[3] ,
    \top_I.branch[25].block[3].um_I.iw[2] ,
    \top_I.branch[25].block[3].um_I.iw[1] ,
    \top_I.branch[25].block[3].um_I.clk ,
    \top_I.branch[25].block[2].um_I.iw[17] ,
    \top_I.branch[25].block[2].um_I.iw[16] ,
    \top_I.branch[25].block[2].um_I.iw[15] ,
    \top_I.branch[25].block[2].um_I.iw[14] ,
    \top_I.branch[25].block[2].um_I.iw[13] ,
    \top_I.branch[25].block[2].um_I.iw[12] ,
    \top_I.branch[25].block[2].um_I.iw[11] ,
    \top_I.branch[25].block[2].um_I.iw[10] ,
    \top_I.branch[25].block[2].um_I.iw[9] ,
    \top_I.branch[25].block[2].um_I.iw[8] ,
    \top_I.branch[25].block[2].um_I.iw[7] ,
    \top_I.branch[25].block[2].um_I.iw[6] ,
    \top_I.branch[25].block[2].um_I.iw[5] ,
    \top_I.branch[25].block[2].um_I.iw[4] ,
    \top_I.branch[25].block[2].um_I.iw[3] ,
    \top_I.branch[25].block[2].um_I.iw[2] ,
    \top_I.branch[25].block[2].um_I.iw[1] ,
    \top_I.branch[25].block[2].um_I.clk ,
    \top_I.branch[25].block[1].um_I.iw[17] ,
    \top_I.branch[25].block[1].um_I.iw[16] ,
    \top_I.branch[25].block[1].um_I.iw[15] ,
    \top_I.branch[25].block[1].um_I.iw[14] ,
    \top_I.branch[25].block[1].um_I.iw[13] ,
    \top_I.branch[25].block[1].um_I.iw[12] ,
    \top_I.branch[25].block[1].um_I.iw[11] ,
    \top_I.branch[25].block[1].um_I.iw[10] ,
    \top_I.branch[25].block[1].um_I.iw[9] ,
    \top_I.branch[25].block[1].um_I.iw[8] ,
    \top_I.branch[25].block[1].um_I.iw[7] ,
    \top_I.branch[25].block[1].um_I.iw[6] ,
    \top_I.branch[25].block[1].um_I.iw[5] ,
    \top_I.branch[25].block[1].um_I.iw[4] ,
    \top_I.branch[25].block[1].um_I.iw[3] ,
    \top_I.branch[25].block[1].um_I.iw[2] ,
    \top_I.branch[25].block[1].um_I.iw[1] ,
    \top_I.branch[25].block[1].um_I.clk ,
    \top_I.branch[25].block[0].um_I.iw[17] ,
    \top_I.branch[25].block[0].um_I.iw[16] ,
    \top_I.branch[25].block[0].um_I.iw[15] ,
    \top_I.branch[25].block[0].um_I.iw[14] ,
    \top_I.branch[25].block[0].um_I.iw[13] ,
    \top_I.branch[25].block[0].um_I.iw[12] ,
    \top_I.branch[25].block[0].um_I.iw[11] ,
    \top_I.branch[25].block[0].um_I.iw[10] ,
    \top_I.branch[25].block[0].um_I.iw[9] ,
    \top_I.branch[25].block[0].um_I.iw[8] ,
    \top_I.branch[25].block[0].um_I.iw[7] ,
    \top_I.branch[25].block[0].um_I.iw[6] ,
    \top_I.branch[25].block[0].um_I.iw[5] ,
    \top_I.branch[25].block[0].um_I.iw[4] ,
    \top_I.branch[25].block[0].um_I.iw[3] ,
    \top_I.branch[25].block[0].um_I.iw[2] ,
    \top_I.branch[25].block[0].um_I.iw[1] ,
    \top_I.branch[25].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[15].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[14].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[13].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[12].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[11].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[10].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[9].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[8].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[7].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[6].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[5].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[4].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[3].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[2].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[1].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero ,
    \top_I.branch[25].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[25].block[15].um_I.pg_vdd ,
    \top_I.branch[25].block[14].um_I.pg_vdd ,
    \top_I.branch[25].block[13].um_I.pg_vdd ,
    \top_I.branch[25].block[12].um_I.pg_vdd ,
    \top_I.branch[25].block[11].um_I.pg_vdd ,
    \top_I.branch[25].block[10].um_I.pg_vdd ,
    \top_I.branch[25].block[9].um_I.pg_vdd ,
    \top_I.branch[25].block[8].um_I.pg_vdd ,
    \top_I.branch[25].block[7].um_I.pg_vdd ,
    \top_I.branch[25].block[6].um_I.pg_vdd ,
    \top_I.branch[25].block[5].um_I.pg_vdd ,
    \top_I.branch[25].block[4].um_I.pg_vdd ,
    \top_I.branch[25].block[3].um_I.pg_vdd ,
    \top_I.branch[25].block[2].um_I.pg_vdd ,
    \top_I.branch[25].block[1].um_I.pg_vdd ,
    \top_I.branch[25].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[26].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[26].l_addr[0] ),
    .k_zero(\top_I.branch[26].l_addr[1] ),
    .addr({\top_I.branch[26].l_addr[0] ,
    \top_I.branch[26].l_addr[0] ,
    \top_I.branch[26].l_addr[1] ,
    \top_I.branch[26].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[26].block[15].um_I.ena ,
    \top_I.branch[26].block[14].um_I.ena ,
    \top_I.branch[26].block[13].um_I.ena ,
    \top_I.branch[26].block[12].um_I.ena ,
    \top_I.branch[26].block[11].um_I.ena ,
    \top_I.branch[26].block[10].um_I.ena ,
    \top_I.branch[26].block[9].um_I.ena ,
    \top_I.branch[26].block[8].um_I.ena ,
    \top_I.branch[26].block[7].um_I.ena ,
    \top_I.branch[26].block[6].um_I.ena ,
    \top_I.branch[26].block[5].um_I.ena ,
    \top_I.branch[26].block[4].um_I.ena ,
    \top_I.branch[26].block[3].um_I.ena ,
    \top_I.branch[26].block[2].um_I.ena ,
    \top_I.branch[26].block[1].um_I.ena ,
    \top_I.branch[26].block[0].um_I.ena }),
    .um_iw({\top_I.branch[26].block[15].um_I.iw[17] ,
    \top_I.branch[26].block[15].um_I.iw[16] ,
    \top_I.branch[26].block[15].um_I.iw[15] ,
    \top_I.branch[26].block[15].um_I.iw[14] ,
    \top_I.branch[26].block[15].um_I.iw[13] ,
    \top_I.branch[26].block[15].um_I.iw[12] ,
    \top_I.branch[26].block[15].um_I.iw[11] ,
    \top_I.branch[26].block[15].um_I.iw[10] ,
    \top_I.branch[26].block[15].um_I.iw[9] ,
    \top_I.branch[26].block[15].um_I.iw[8] ,
    \top_I.branch[26].block[15].um_I.iw[7] ,
    \top_I.branch[26].block[15].um_I.iw[6] ,
    \top_I.branch[26].block[15].um_I.iw[5] ,
    \top_I.branch[26].block[15].um_I.iw[4] ,
    \top_I.branch[26].block[15].um_I.iw[3] ,
    \top_I.branch[26].block[15].um_I.iw[2] ,
    \top_I.branch[26].block[15].um_I.iw[1] ,
    \top_I.branch[26].block[15].um_I.clk ,
    \top_I.branch[26].block[14].um_I.iw[17] ,
    \top_I.branch[26].block[14].um_I.iw[16] ,
    \top_I.branch[26].block[14].um_I.iw[15] ,
    \top_I.branch[26].block[14].um_I.iw[14] ,
    \top_I.branch[26].block[14].um_I.iw[13] ,
    \top_I.branch[26].block[14].um_I.iw[12] ,
    \top_I.branch[26].block[14].um_I.iw[11] ,
    \top_I.branch[26].block[14].um_I.iw[10] ,
    \top_I.branch[26].block[14].um_I.iw[9] ,
    \top_I.branch[26].block[14].um_I.iw[8] ,
    \top_I.branch[26].block[14].um_I.iw[7] ,
    \top_I.branch[26].block[14].um_I.iw[6] ,
    \top_I.branch[26].block[14].um_I.iw[5] ,
    \top_I.branch[26].block[14].um_I.iw[4] ,
    \top_I.branch[26].block[14].um_I.iw[3] ,
    \top_I.branch[26].block[14].um_I.iw[2] ,
    \top_I.branch[26].block[14].um_I.iw[1] ,
    \top_I.branch[26].block[14].um_I.clk ,
    \top_I.branch[26].block[13].um_I.iw[17] ,
    \top_I.branch[26].block[13].um_I.iw[16] ,
    \top_I.branch[26].block[13].um_I.iw[15] ,
    \top_I.branch[26].block[13].um_I.iw[14] ,
    \top_I.branch[26].block[13].um_I.iw[13] ,
    \top_I.branch[26].block[13].um_I.iw[12] ,
    \top_I.branch[26].block[13].um_I.iw[11] ,
    \top_I.branch[26].block[13].um_I.iw[10] ,
    \top_I.branch[26].block[13].um_I.iw[9] ,
    \top_I.branch[26].block[13].um_I.iw[8] ,
    \top_I.branch[26].block[13].um_I.iw[7] ,
    \top_I.branch[26].block[13].um_I.iw[6] ,
    \top_I.branch[26].block[13].um_I.iw[5] ,
    \top_I.branch[26].block[13].um_I.iw[4] ,
    \top_I.branch[26].block[13].um_I.iw[3] ,
    \top_I.branch[26].block[13].um_I.iw[2] ,
    \top_I.branch[26].block[13].um_I.iw[1] ,
    \top_I.branch[26].block[13].um_I.clk ,
    \top_I.branch[26].block[12].um_I.iw[17] ,
    \top_I.branch[26].block[12].um_I.iw[16] ,
    \top_I.branch[26].block[12].um_I.iw[15] ,
    \top_I.branch[26].block[12].um_I.iw[14] ,
    \top_I.branch[26].block[12].um_I.iw[13] ,
    \top_I.branch[26].block[12].um_I.iw[12] ,
    \top_I.branch[26].block[12].um_I.iw[11] ,
    \top_I.branch[26].block[12].um_I.iw[10] ,
    \top_I.branch[26].block[12].um_I.iw[9] ,
    \top_I.branch[26].block[12].um_I.iw[8] ,
    \top_I.branch[26].block[12].um_I.iw[7] ,
    \top_I.branch[26].block[12].um_I.iw[6] ,
    \top_I.branch[26].block[12].um_I.iw[5] ,
    \top_I.branch[26].block[12].um_I.iw[4] ,
    \top_I.branch[26].block[12].um_I.iw[3] ,
    \top_I.branch[26].block[12].um_I.iw[2] ,
    \top_I.branch[26].block[12].um_I.iw[1] ,
    \top_I.branch[26].block[12].um_I.clk ,
    \top_I.branch[26].block[11].um_I.iw[17] ,
    \top_I.branch[26].block[11].um_I.iw[16] ,
    \top_I.branch[26].block[11].um_I.iw[15] ,
    \top_I.branch[26].block[11].um_I.iw[14] ,
    \top_I.branch[26].block[11].um_I.iw[13] ,
    \top_I.branch[26].block[11].um_I.iw[12] ,
    \top_I.branch[26].block[11].um_I.iw[11] ,
    \top_I.branch[26].block[11].um_I.iw[10] ,
    \top_I.branch[26].block[11].um_I.iw[9] ,
    \top_I.branch[26].block[11].um_I.iw[8] ,
    \top_I.branch[26].block[11].um_I.iw[7] ,
    \top_I.branch[26].block[11].um_I.iw[6] ,
    \top_I.branch[26].block[11].um_I.iw[5] ,
    \top_I.branch[26].block[11].um_I.iw[4] ,
    \top_I.branch[26].block[11].um_I.iw[3] ,
    \top_I.branch[26].block[11].um_I.iw[2] ,
    \top_I.branch[26].block[11].um_I.iw[1] ,
    \top_I.branch[26].block[11].um_I.clk ,
    \top_I.branch[26].block[10].um_I.iw[17] ,
    \top_I.branch[26].block[10].um_I.iw[16] ,
    \top_I.branch[26].block[10].um_I.iw[15] ,
    \top_I.branch[26].block[10].um_I.iw[14] ,
    \top_I.branch[26].block[10].um_I.iw[13] ,
    \top_I.branch[26].block[10].um_I.iw[12] ,
    \top_I.branch[26].block[10].um_I.iw[11] ,
    \top_I.branch[26].block[10].um_I.iw[10] ,
    \top_I.branch[26].block[10].um_I.iw[9] ,
    \top_I.branch[26].block[10].um_I.iw[8] ,
    \top_I.branch[26].block[10].um_I.iw[7] ,
    \top_I.branch[26].block[10].um_I.iw[6] ,
    \top_I.branch[26].block[10].um_I.iw[5] ,
    \top_I.branch[26].block[10].um_I.iw[4] ,
    \top_I.branch[26].block[10].um_I.iw[3] ,
    \top_I.branch[26].block[10].um_I.iw[2] ,
    \top_I.branch[26].block[10].um_I.iw[1] ,
    \top_I.branch[26].block[10].um_I.clk ,
    \top_I.branch[26].block[9].um_I.iw[17] ,
    \top_I.branch[26].block[9].um_I.iw[16] ,
    \top_I.branch[26].block[9].um_I.iw[15] ,
    \top_I.branch[26].block[9].um_I.iw[14] ,
    \top_I.branch[26].block[9].um_I.iw[13] ,
    \top_I.branch[26].block[9].um_I.iw[12] ,
    \top_I.branch[26].block[9].um_I.iw[11] ,
    \top_I.branch[26].block[9].um_I.iw[10] ,
    \top_I.branch[26].block[9].um_I.iw[9] ,
    \top_I.branch[26].block[9].um_I.iw[8] ,
    \top_I.branch[26].block[9].um_I.iw[7] ,
    \top_I.branch[26].block[9].um_I.iw[6] ,
    \top_I.branch[26].block[9].um_I.iw[5] ,
    \top_I.branch[26].block[9].um_I.iw[4] ,
    \top_I.branch[26].block[9].um_I.iw[3] ,
    \top_I.branch[26].block[9].um_I.iw[2] ,
    \top_I.branch[26].block[9].um_I.iw[1] ,
    \top_I.branch[26].block[9].um_I.clk ,
    \top_I.branch[26].block[8].um_I.iw[17] ,
    \top_I.branch[26].block[8].um_I.iw[16] ,
    \top_I.branch[26].block[8].um_I.iw[15] ,
    \top_I.branch[26].block[8].um_I.iw[14] ,
    \top_I.branch[26].block[8].um_I.iw[13] ,
    \top_I.branch[26].block[8].um_I.iw[12] ,
    \top_I.branch[26].block[8].um_I.iw[11] ,
    \top_I.branch[26].block[8].um_I.iw[10] ,
    \top_I.branch[26].block[8].um_I.iw[9] ,
    \top_I.branch[26].block[8].um_I.iw[8] ,
    \top_I.branch[26].block[8].um_I.iw[7] ,
    \top_I.branch[26].block[8].um_I.iw[6] ,
    \top_I.branch[26].block[8].um_I.iw[5] ,
    \top_I.branch[26].block[8].um_I.iw[4] ,
    \top_I.branch[26].block[8].um_I.iw[3] ,
    \top_I.branch[26].block[8].um_I.iw[2] ,
    \top_I.branch[26].block[8].um_I.iw[1] ,
    \top_I.branch[26].block[8].um_I.clk ,
    \top_I.branch[26].block[7].um_I.iw[17] ,
    \top_I.branch[26].block[7].um_I.iw[16] ,
    \top_I.branch[26].block[7].um_I.iw[15] ,
    \top_I.branch[26].block[7].um_I.iw[14] ,
    \top_I.branch[26].block[7].um_I.iw[13] ,
    \top_I.branch[26].block[7].um_I.iw[12] ,
    \top_I.branch[26].block[7].um_I.iw[11] ,
    \top_I.branch[26].block[7].um_I.iw[10] ,
    \top_I.branch[26].block[7].um_I.iw[9] ,
    \top_I.branch[26].block[7].um_I.iw[8] ,
    \top_I.branch[26].block[7].um_I.iw[7] ,
    \top_I.branch[26].block[7].um_I.iw[6] ,
    \top_I.branch[26].block[7].um_I.iw[5] ,
    \top_I.branch[26].block[7].um_I.iw[4] ,
    \top_I.branch[26].block[7].um_I.iw[3] ,
    \top_I.branch[26].block[7].um_I.iw[2] ,
    \top_I.branch[26].block[7].um_I.iw[1] ,
    \top_I.branch[26].block[7].um_I.clk ,
    \top_I.branch[26].block[6].um_I.iw[17] ,
    \top_I.branch[26].block[6].um_I.iw[16] ,
    \top_I.branch[26].block[6].um_I.iw[15] ,
    \top_I.branch[26].block[6].um_I.iw[14] ,
    \top_I.branch[26].block[6].um_I.iw[13] ,
    \top_I.branch[26].block[6].um_I.iw[12] ,
    \top_I.branch[26].block[6].um_I.iw[11] ,
    \top_I.branch[26].block[6].um_I.iw[10] ,
    \top_I.branch[26].block[6].um_I.iw[9] ,
    \top_I.branch[26].block[6].um_I.iw[8] ,
    \top_I.branch[26].block[6].um_I.iw[7] ,
    \top_I.branch[26].block[6].um_I.iw[6] ,
    \top_I.branch[26].block[6].um_I.iw[5] ,
    \top_I.branch[26].block[6].um_I.iw[4] ,
    \top_I.branch[26].block[6].um_I.iw[3] ,
    \top_I.branch[26].block[6].um_I.iw[2] ,
    \top_I.branch[26].block[6].um_I.iw[1] ,
    \top_I.branch[26].block[6].um_I.clk ,
    \top_I.branch[26].block[5].um_I.iw[17] ,
    \top_I.branch[26].block[5].um_I.iw[16] ,
    \top_I.branch[26].block[5].um_I.iw[15] ,
    \top_I.branch[26].block[5].um_I.iw[14] ,
    \top_I.branch[26].block[5].um_I.iw[13] ,
    \top_I.branch[26].block[5].um_I.iw[12] ,
    \top_I.branch[26].block[5].um_I.iw[11] ,
    \top_I.branch[26].block[5].um_I.iw[10] ,
    \top_I.branch[26].block[5].um_I.iw[9] ,
    \top_I.branch[26].block[5].um_I.iw[8] ,
    \top_I.branch[26].block[5].um_I.iw[7] ,
    \top_I.branch[26].block[5].um_I.iw[6] ,
    \top_I.branch[26].block[5].um_I.iw[5] ,
    \top_I.branch[26].block[5].um_I.iw[4] ,
    \top_I.branch[26].block[5].um_I.iw[3] ,
    \top_I.branch[26].block[5].um_I.iw[2] ,
    \top_I.branch[26].block[5].um_I.iw[1] ,
    \top_I.branch[26].block[5].um_I.clk ,
    \top_I.branch[26].block[4].um_I.iw[17] ,
    \top_I.branch[26].block[4].um_I.iw[16] ,
    \top_I.branch[26].block[4].um_I.iw[15] ,
    \top_I.branch[26].block[4].um_I.iw[14] ,
    \top_I.branch[26].block[4].um_I.iw[13] ,
    \top_I.branch[26].block[4].um_I.iw[12] ,
    \top_I.branch[26].block[4].um_I.iw[11] ,
    \top_I.branch[26].block[4].um_I.iw[10] ,
    \top_I.branch[26].block[4].um_I.iw[9] ,
    \top_I.branch[26].block[4].um_I.iw[8] ,
    \top_I.branch[26].block[4].um_I.iw[7] ,
    \top_I.branch[26].block[4].um_I.iw[6] ,
    \top_I.branch[26].block[4].um_I.iw[5] ,
    \top_I.branch[26].block[4].um_I.iw[4] ,
    \top_I.branch[26].block[4].um_I.iw[3] ,
    \top_I.branch[26].block[4].um_I.iw[2] ,
    \top_I.branch[26].block[4].um_I.iw[1] ,
    \top_I.branch[26].block[4].um_I.clk ,
    \top_I.branch[26].block[3].um_I.iw[17] ,
    \top_I.branch[26].block[3].um_I.iw[16] ,
    \top_I.branch[26].block[3].um_I.iw[15] ,
    \top_I.branch[26].block[3].um_I.iw[14] ,
    \top_I.branch[26].block[3].um_I.iw[13] ,
    \top_I.branch[26].block[3].um_I.iw[12] ,
    \top_I.branch[26].block[3].um_I.iw[11] ,
    \top_I.branch[26].block[3].um_I.iw[10] ,
    \top_I.branch[26].block[3].um_I.iw[9] ,
    \top_I.branch[26].block[3].um_I.iw[8] ,
    \top_I.branch[26].block[3].um_I.iw[7] ,
    \top_I.branch[26].block[3].um_I.iw[6] ,
    \top_I.branch[26].block[3].um_I.iw[5] ,
    \top_I.branch[26].block[3].um_I.iw[4] ,
    \top_I.branch[26].block[3].um_I.iw[3] ,
    \top_I.branch[26].block[3].um_I.iw[2] ,
    \top_I.branch[26].block[3].um_I.iw[1] ,
    \top_I.branch[26].block[3].um_I.clk ,
    \top_I.branch[26].block[2].um_I.iw[17] ,
    \top_I.branch[26].block[2].um_I.iw[16] ,
    \top_I.branch[26].block[2].um_I.iw[15] ,
    \top_I.branch[26].block[2].um_I.iw[14] ,
    \top_I.branch[26].block[2].um_I.iw[13] ,
    \top_I.branch[26].block[2].um_I.iw[12] ,
    \top_I.branch[26].block[2].um_I.iw[11] ,
    \top_I.branch[26].block[2].um_I.iw[10] ,
    \top_I.branch[26].block[2].um_I.iw[9] ,
    \top_I.branch[26].block[2].um_I.iw[8] ,
    \top_I.branch[26].block[2].um_I.iw[7] ,
    \top_I.branch[26].block[2].um_I.iw[6] ,
    \top_I.branch[26].block[2].um_I.iw[5] ,
    \top_I.branch[26].block[2].um_I.iw[4] ,
    \top_I.branch[26].block[2].um_I.iw[3] ,
    \top_I.branch[26].block[2].um_I.iw[2] ,
    \top_I.branch[26].block[2].um_I.iw[1] ,
    \top_I.branch[26].block[2].um_I.clk ,
    \top_I.branch[26].block[1].um_I.iw[17] ,
    \top_I.branch[26].block[1].um_I.iw[16] ,
    \top_I.branch[26].block[1].um_I.iw[15] ,
    \top_I.branch[26].block[1].um_I.iw[14] ,
    \top_I.branch[26].block[1].um_I.iw[13] ,
    \top_I.branch[26].block[1].um_I.iw[12] ,
    \top_I.branch[26].block[1].um_I.iw[11] ,
    \top_I.branch[26].block[1].um_I.iw[10] ,
    \top_I.branch[26].block[1].um_I.iw[9] ,
    \top_I.branch[26].block[1].um_I.iw[8] ,
    \top_I.branch[26].block[1].um_I.iw[7] ,
    \top_I.branch[26].block[1].um_I.iw[6] ,
    \top_I.branch[26].block[1].um_I.iw[5] ,
    \top_I.branch[26].block[1].um_I.iw[4] ,
    \top_I.branch[26].block[1].um_I.iw[3] ,
    \top_I.branch[26].block[1].um_I.iw[2] ,
    \top_I.branch[26].block[1].um_I.iw[1] ,
    \top_I.branch[26].block[1].um_I.clk ,
    \top_I.branch[26].block[0].um_I.iw[17] ,
    \top_I.branch[26].block[0].um_I.iw[16] ,
    \top_I.branch[26].block[0].um_I.iw[15] ,
    \top_I.branch[26].block[0].um_I.iw[14] ,
    \top_I.branch[26].block[0].um_I.iw[13] ,
    \top_I.branch[26].block[0].um_I.iw[12] ,
    \top_I.branch[26].block[0].um_I.iw[11] ,
    \top_I.branch[26].block[0].um_I.iw[10] ,
    \top_I.branch[26].block[0].um_I.iw[9] ,
    \top_I.branch[26].block[0].um_I.iw[8] ,
    \top_I.branch[26].block[0].um_I.iw[7] ,
    \top_I.branch[26].block[0].um_I.iw[6] ,
    \top_I.branch[26].block[0].um_I.iw[5] ,
    \top_I.branch[26].block[0].um_I.iw[4] ,
    \top_I.branch[26].block[0].um_I.iw[3] ,
    \top_I.branch[26].block[0].um_I.iw[2] ,
    \top_I.branch[26].block[0].um_I.iw[1] ,
    \top_I.branch[26].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[15].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[14].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[13].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[12].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[11].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[10].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[9].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[8].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[7].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[6].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[5].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[4].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[3].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[2].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[1].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero ,
    \top_I.branch[26].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[26].block[15].um_I.pg_vdd ,
    \top_I.branch[26].block[14].um_I.pg_vdd ,
    \top_I.branch[26].block[13].um_I.pg_vdd ,
    \top_I.branch[26].block[12].um_I.pg_vdd ,
    \top_I.branch[26].block[11].um_I.pg_vdd ,
    \top_I.branch[26].block[10].um_I.pg_vdd ,
    \top_I.branch[26].block[9].um_I.pg_vdd ,
    \top_I.branch[26].block[8].um_I.pg_vdd ,
    \top_I.branch[26].block[7].um_I.pg_vdd ,
    \top_I.branch[26].block[6].um_I.pg_vdd ,
    \top_I.branch[26].block[5].um_I.pg_vdd ,
    \top_I.branch[26].block[4].um_I.pg_vdd ,
    \top_I.branch[26].block[3].um_I.pg_vdd ,
    \top_I.branch[26].block[2].um_I.pg_vdd ,
    \top_I.branch[26].block[1].um_I.pg_vdd ,
    \top_I.branch[26].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[27].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[27].l_addr[0] ),
    .k_zero(\top_I.branch[27].l_addr[1] ),
    .addr({\top_I.branch[27].l_addr[0] ,
    \top_I.branch[27].l_addr[0] ,
    \top_I.branch[27].l_addr[1] ,
    \top_I.branch[27].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[27].block[15].um_I.ena ,
    \top_I.branch[27].block[14].um_I.ena ,
    \top_I.branch[27].block[13].um_I.ena ,
    \top_I.branch[27].block[12].um_I.ena ,
    \top_I.branch[27].block[11].um_I.ena ,
    \top_I.branch[27].block[10].um_I.ena ,
    \top_I.branch[27].block[9].um_I.ena ,
    \top_I.branch[27].block[8].um_I.ena ,
    \top_I.branch[27].block[7].um_I.ena ,
    \top_I.branch[27].block[6].um_I.ena ,
    \top_I.branch[27].block[5].um_I.ena ,
    \top_I.branch[27].block[4].um_I.ena ,
    \top_I.branch[27].block[3].um_I.ena ,
    \top_I.branch[27].block[2].um_I.ena ,
    \top_I.branch[27].block[1].um_I.ena ,
    \top_I.branch[27].block[0].um_I.ena }),
    .um_iw({\top_I.branch[27].block[15].um_I.iw[17] ,
    \top_I.branch[27].block[15].um_I.iw[16] ,
    \top_I.branch[27].block[15].um_I.iw[15] ,
    \top_I.branch[27].block[15].um_I.iw[14] ,
    \top_I.branch[27].block[15].um_I.iw[13] ,
    \top_I.branch[27].block[15].um_I.iw[12] ,
    \top_I.branch[27].block[15].um_I.iw[11] ,
    \top_I.branch[27].block[15].um_I.iw[10] ,
    \top_I.branch[27].block[15].um_I.iw[9] ,
    \top_I.branch[27].block[15].um_I.iw[8] ,
    \top_I.branch[27].block[15].um_I.iw[7] ,
    \top_I.branch[27].block[15].um_I.iw[6] ,
    \top_I.branch[27].block[15].um_I.iw[5] ,
    \top_I.branch[27].block[15].um_I.iw[4] ,
    \top_I.branch[27].block[15].um_I.iw[3] ,
    \top_I.branch[27].block[15].um_I.iw[2] ,
    \top_I.branch[27].block[15].um_I.iw[1] ,
    \top_I.branch[27].block[15].um_I.clk ,
    \top_I.branch[27].block[14].um_I.iw[17] ,
    \top_I.branch[27].block[14].um_I.iw[16] ,
    \top_I.branch[27].block[14].um_I.iw[15] ,
    \top_I.branch[27].block[14].um_I.iw[14] ,
    \top_I.branch[27].block[14].um_I.iw[13] ,
    \top_I.branch[27].block[14].um_I.iw[12] ,
    \top_I.branch[27].block[14].um_I.iw[11] ,
    \top_I.branch[27].block[14].um_I.iw[10] ,
    \top_I.branch[27].block[14].um_I.iw[9] ,
    \top_I.branch[27].block[14].um_I.iw[8] ,
    \top_I.branch[27].block[14].um_I.iw[7] ,
    \top_I.branch[27].block[14].um_I.iw[6] ,
    \top_I.branch[27].block[14].um_I.iw[5] ,
    \top_I.branch[27].block[14].um_I.iw[4] ,
    \top_I.branch[27].block[14].um_I.iw[3] ,
    \top_I.branch[27].block[14].um_I.iw[2] ,
    \top_I.branch[27].block[14].um_I.iw[1] ,
    \top_I.branch[27].block[14].um_I.clk ,
    \top_I.branch[27].block[13].um_I.iw[17] ,
    \top_I.branch[27].block[13].um_I.iw[16] ,
    \top_I.branch[27].block[13].um_I.iw[15] ,
    \top_I.branch[27].block[13].um_I.iw[14] ,
    \top_I.branch[27].block[13].um_I.iw[13] ,
    \top_I.branch[27].block[13].um_I.iw[12] ,
    \top_I.branch[27].block[13].um_I.iw[11] ,
    \top_I.branch[27].block[13].um_I.iw[10] ,
    \top_I.branch[27].block[13].um_I.iw[9] ,
    \top_I.branch[27].block[13].um_I.iw[8] ,
    \top_I.branch[27].block[13].um_I.iw[7] ,
    \top_I.branch[27].block[13].um_I.iw[6] ,
    \top_I.branch[27].block[13].um_I.iw[5] ,
    \top_I.branch[27].block[13].um_I.iw[4] ,
    \top_I.branch[27].block[13].um_I.iw[3] ,
    \top_I.branch[27].block[13].um_I.iw[2] ,
    \top_I.branch[27].block[13].um_I.iw[1] ,
    \top_I.branch[27].block[13].um_I.clk ,
    \top_I.branch[27].block[12].um_I.iw[17] ,
    \top_I.branch[27].block[12].um_I.iw[16] ,
    \top_I.branch[27].block[12].um_I.iw[15] ,
    \top_I.branch[27].block[12].um_I.iw[14] ,
    \top_I.branch[27].block[12].um_I.iw[13] ,
    \top_I.branch[27].block[12].um_I.iw[12] ,
    \top_I.branch[27].block[12].um_I.iw[11] ,
    \top_I.branch[27].block[12].um_I.iw[10] ,
    \top_I.branch[27].block[12].um_I.iw[9] ,
    \top_I.branch[27].block[12].um_I.iw[8] ,
    \top_I.branch[27].block[12].um_I.iw[7] ,
    \top_I.branch[27].block[12].um_I.iw[6] ,
    \top_I.branch[27].block[12].um_I.iw[5] ,
    \top_I.branch[27].block[12].um_I.iw[4] ,
    \top_I.branch[27].block[12].um_I.iw[3] ,
    \top_I.branch[27].block[12].um_I.iw[2] ,
    \top_I.branch[27].block[12].um_I.iw[1] ,
    \top_I.branch[27].block[12].um_I.clk ,
    \top_I.branch[27].block[11].um_I.iw[17] ,
    \top_I.branch[27].block[11].um_I.iw[16] ,
    \top_I.branch[27].block[11].um_I.iw[15] ,
    \top_I.branch[27].block[11].um_I.iw[14] ,
    \top_I.branch[27].block[11].um_I.iw[13] ,
    \top_I.branch[27].block[11].um_I.iw[12] ,
    \top_I.branch[27].block[11].um_I.iw[11] ,
    \top_I.branch[27].block[11].um_I.iw[10] ,
    \top_I.branch[27].block[11].um_I.iw[9] ,
    \top_I.branch[27].block[11].um_I.iw[8] ,
    \top_I.branch[27].block[11].um_I.iw[7] ,
    \top_I.branch[27].block[11].um_I.iw[6] ,
    \top_I.branch[27].block[11].um_I.iw[5] ,
    \top_I.branch[27].block[11].um_I.iw[4] ,
    \top_I.branch[27].block[11].um_I.iw[3] ,
    \top_I.branch[27].block[11].um_I.iw[2] ,
    \top_I.branch[27].block[11].um_I.iw[1] ,
    \top_I.branch[27].block[11].um_I.clk ,
    \top_I.branch[27].block[10].um_I.iw[17] ,
    \top_I.branch[27].block[10].um_I.iw[16] ,
    \top_I.branch[27].block[10].um_I.iw[15] ,
    \top_I.branch[27].block[10].um_I.iw[14] ,
    \top_I.branch[27].block[10].um_I.iw[13] ,
    \top_I.branch[27].block[10].um_I.iw[12] ,
    \top_I.branch[27].block[10].um_I.iw[11] ,
    \top_I.branch[27].block[10].um_I.iw[10] ,
    \top_I.branch[27].block[10].um_I.iw[9] ,
    \top_I.branch[27].block[10].um_I.iw[8] ,
    \top_I.branch[27].block[10].um_I.iw[7] ,
    \top_I.branch[27].block[10].um_I.iw[6] ,
    \top_I.branch[27].block[10].um_I.iw[5] ,
    \top_I.branch[27].block[10].um_I.iw[4] ,
    \top_I.branch[27].block[10].um_I.iw[3] ,
    \top_I.branch[27].block[10].um_I.iw[2] ,
    \top_I.branch[27].block[10].um_I.iw[1] ,
    \top_I.branch[27].block[10].um_I.clk ,
    \top_I.branch[27].block[9].um_I.iw[17] ,
    \top_I.branch[27].block[9].um_I.iw[16] ,
    \top_I.branch[27].block[9].um_I.iw[15] ,
    \top_I.branch[27].block[9].um_I.iw[14] ,
    \top_I.branch[27].block[9].um_I.iw[13] ,
    \top_I.branch[27].block[9].um_I.iw[12] ,
    \top_I.branch[27].block[9].um_I.iw[11] ,
    \top_I.branch[27].block[9].um_I.iw[10] ,
    \top_I.branch[27].block[9].um_I.iw[9] ,
    \top_I.branch[27].block[9].um_I.iw[8] ,
    \top_I.branch[27].block[9].um_I.iw[7] ,
    \top_I.branch[27].block[9].um_I.iw[6] ,
    \top_I.branch[27].block[9].um_I.iw[5] ,
    \top_I.branch[27].block[9].um_I.iw[4] ,
    \top_I.branch[27].block[9].um_I.iw[3] ,
    \top_I.branch[27].block[9].um_I.iw[2] ,
    \top_I.branch[27].block[9].um_I.iw[1] ,
    \top_I.branch[27].block[9].um_I.clk ,
    \top_I.branch[27].block[8].um_I.iw[17] ,
    \top_I.branch[27].block[8].um_I.iw[16] ,
    \top_I.branch[27].block[8].um_I.iw[15] ,
    \top_I.branch[27].block[8].um_I.iw[14] ,
    \top_I.branch[27].block[8].um_I.iw[13] ,
    \top_I.branch[27].block[8].um_I.iw[12] ,
    \top_I.branch[27].block[8].um_I.iw[11] ,
    \top_I.branch[27].block[8].um_I.iw[10] ,
    \top_I.branch[27].block[8].um_I.iw[9] ,
    \top_I.branch[27].block[8].um_I.iw[8] ,
    \top_I.branch[27].block[8].um_I.iw[7] ,
    \top_I.branch[27].block[8].um_I.iw[6] ,
    \top_I.branch[27].block[8].um_I.iw[5] ,
    \top_I.branch[27].block[8].um_I.iw[4] ,
    \top_I.branch[27].block[8].um_I.iw[3] ,
    \top_I.branch[27].block[8].um_I.iw[2] ,
    \top_I.branch[27].block[8].um_I.iw[1] ,
    \top_I.branch[27].block[8].um_I.clk ,
    \top_I.branch[27].block[7].um_I.iw[17] ,
    \top_I.branch[27].block[7].um_I.iw[16] ,
    \top_I.branch[27].block[7].um_I.iw[15] ,
    \top_I.branch[27].block[7].um_I.iw[14] ,
    \top_I.branch[27].block[7].um_I.iw[13] ,
    \top_I.branch[27].block[7].um_I.iw[12] ,
    \top_I.branch[27].block[7].um_I.iw[11] ,
    \top_I.branch[27].block[7].um_I.iw[10] ,
    \top_I.branch[27].block[7].um_I.iw[9] ,
    \top_I.branch[27].block[7].um_I.iw[8] ,
    \top_I.branch[27].block[7].um_I.iw[7] ,
    \top_I.branch[27].block[7].um_I.iw[6] ,
    \top_I.branch[27].block[7].um_I.iw[5] ,
    \top_I.branch[27].block[7].um_I.iw[4] ,
    \top_I.branch[27].block[7].um_I.iw[3] ,
    \top_I.branch[27].block[7].um_I.iw[2] ,
    \top_I.branch[27].block[7].um_I.iw[1] ,
    \top_I.branch[27].block[7].um_I.clk ,
    \top_I.branch[27].block[6].um_I.iw[17] ,
    \top_I.branch[27].block[6].um_I.iw[16] ,
    \top_I.branch[27].block[6].um_I.iw[15] ,
    \top_I.branch[27].block[6].um_I.iw[14] ,
    \top_I.branch[27].block[6].um_I.iw[13] ,
    \top_I.branch[27].block[6].um_I.iw[12] ,
    \top_I.branch[27].block[6].um_I.iw[11] ,
    \top_I.branch[27].block[6].um_I.iw[10] ,
    \top_I.branch[27].block[6].um_I.iw[9] ,
    \top_I.branch[27].block[6].um_I.iw[8] ,
    \top_I.branch[27].block[6].um_I.iw[7] ,
    \top_I.branch[27].block[6].um_I.iw[6] ,
    \top_I.branch[27].block[6].um_I.iw[5] ,
    \top_I.branch[27].block[6].um_I.iw[4] ,
    \top_I.branch[27].block[6].um_I.iw[3] ,
    \top_I.branch[27].block[6].um_I.iw[2] ,
    \top_I.branch[27].block[6].um_I.iw[1] ,
    \top_I.branch[27].block[6].um_I.clk ,
    \top_I.branch[27].block[5].um_I.iw[17] ,
    \top_I.branch[27].block[5].um_I.iw[16] ,
    \top_I.branch[27].block[5].um_I.iw[15] ,
    \top_I.branch[27].block[5].um_I.iw[14] ,
    \top_I.branch[27].block[5].um_I.iw[13] ,
    \top_I.branch[27].block[5].um_I.iw[12] ,
    \top_I.branch[27].block[5].um_I.iw[11] ,
    \top_I.branch[27].block[5].um_I.iw[10] ,
    \top_I.branch[27].block[5].um_I.iw[9] ,
    \top_I.branch[27].block[5].um_I.iw[8] ,
    \top_I.branch[27].block[5].um_I.iw[7] ,
    \top_I.branch[27].block[5].um_I.iw[6] ,
    \top_I.branch[27].block[5].um_I.iw[5] ,
    \top_I.branch[27].block[5].um_I.iw[4] ,
    \top_I.branch[27].block[5].um_I.iw[3] ,
    \top_I.branch[27].block[5].um_I.iw[2] ,
    \top_I.branch[27].block[5].um_I.iw[1] ,
    \top_I.branch[27].block[5].um_I.clk ,
    \top_I.branch[27].block[4].um_I.iw[17] ,
    \top_I.branch[27].block[4].um_I.iw[16] ,
    \top_I.branch[27].block[4].um_I.iw[15] ,
    \top_I.branch[27].block[4].um_I.iw[14] ,
    \top_I.branch[27].block[4].um_I.iw[13] ,
    \top_I.branch[27].block[4].um_I.iw[12] ,
    \top_I.branch[27].block[4].um_I.iw[11] ,
    \top_I.branch[27].block[4].um_I.iw[10] ,
    \top_I.branch[27].block[4].um_I.iw[9] ,
    \top_I.branch[27].block[4].um_I.iw[8] ,
    \top_I.branch[27].block[4].um_I.iw[7] ,
    \top_I.branch[27].block[4].um_I.iw[6] ,
    \top_I.branch[27].block[4].um_I.iw[5] ,
    \top_I.branch[27].block[4].um_I.iw[4] ,
    \top_I.branch[27].block[4].um_I.iw[3] ,
    \top_I.branch[27].block[4].um_I.iw[2] ,
    \top_I.branch[27].block[4].um_I.iw[1] ,
    \top_I.branch[27].block[4].um_I.clk ,
    \top_I.branch[27].block[3].um_I.iw[17] ,
    \top_I.branch[27].block[3].um_I.iw[16] ,
    \top_I.branch[27].block[3].um_I.iw[15] ,
    \top_I.branch[27].block[3].um_I.iw[14] ,
    \top_I.branch[27].block[3].um_I.iw[13] ,
    \top_I.branch[27].block[3].um_I.iw[12] ,
    \top_I.branch[27].block[3].um_I.iw[11] ,
    \top_I.branch[27].block[3].um_I.iw[10] ,
    \top_I.branch[27].block[3].um_I.iw[9] ,
    \top_I.branch[27].block[3].um_I.iw[8] ,
    \top_I.branch[27].block[3].um_I.iw[7] ,
    \top_I.branch[27].block[3].um_I.iw[6] ,
    \top_I.branch[27].block[3].um_I.iw[5] ,
    \top_I.branch[27].block[3].um_I.iw[4] ,
    \top_I.branch[27].block[3].um_I.iw[3] ,
    \top_I.branch[27].block[3].um_I.iw[2] ,
    \top_I.branch[27].block[3].um_I.iw[1] ,
    \top_I.branch[27].block[3].um_I.clk ,
    \top_I.branch[27].block[2].um_I.iw[17] ,
    \top_I.branch[27].block[2].um_I.iw[16] ,
    \top_I.branch[27].block[2].um_I.iw[15] ,
    \top_I.branch[27].block[2].um_I.iw[14] ,
    \top_I.branch[27].block[2].um_I.iw[13] ,
    \top_I.branch[27].block[2].um_I.iw[12] ,
    \top_I.branch[27].block[2].um_I.iw[11] ,
    \top_I.branch[27].block[2].um_I.iw[10] ,
    \top_I.branch[27].block[2].um_I.iw[9] ,
    \top_I.branch[27].block[2].um_I.iw[8] ,
    \top_I.branch[27].block[2].um_I.iw[7] ,
    \top_I.branch[27].block[2].um_I.iw[6] ,
    \top_I.branch[27].block[2].um_I.iw[5] ,
    \top_I.branch[27].block[2].um_I.iw[4] ,
    \top_I.branch[27].block[2].um_I.iw[3] ,
    \top_I.branch[27].block[2].um_I.iw[2] ,
    \top_I.branch[27].block[2].um_I.iw[1] ,
    \top_I.branch[27].block[2].um_I.clk ,
    \top_I.branch[27].block[1].um_I.iw[17] ,
    \top_I.branch[27].block[1].um_I.iw[16] ,
    \top_I.branch[27].block[1].um_I.iw[15] ,
    \top_I.branch[27].block[1].um_I.iw[14] ,
    \top_I.branch[27].block[1].um_I.iw[13] ,
    \top_I.branch[27].block[1].um_I.iw[12] ,
    \top_I.branch[27].block[1].um_I.iw[11] ,
    \top_I.branch[27].block[1].um_I.iw[10] ,
    \top_I.branch[27].block[1].um_I.iw[9] ,
    \top_I.branch[27].block[1].um_I.iw[8] ,
    \top_I.branch[27].block[1].um_I.iw[7] ,
    \top_I.branch[27].block[1].um_I.iw[6] ,
    \top_I.branch[27].block[1].um_I.iw[5] ,
    \top_I.branch[27].block[1].um_I.iw[4] ,
    \top_I.branch[27].block[1].um_I.iw[3] ,
    \top_I.branch[27].block[1].um_I.iw[2] ,
    \top_I.branch[27].block[1].um_I.iw[1] ,
    \top_I.branch[27].block[1].um_I.clk ,
    \top_I.branch[27].block[0].um_I.iw[17] ,
    \top_I.branch[27].block[0].um_I.iw[16] ,
    \top_I.branch[27].block[0].um_I.iw[15] ,
    \top_I.branch[27].block[0].um_I.iw[14] ,
    \top_I.branch[27].block[0].um_I.iw[13] ,
    \top_I.branch[27].block[0].um_I.iw[12] ,
    \top_I.branch[27].block[0].um_I.iw[11] ,
    \top_I.branch[27].block[0].um_I.iw[10] ,
    \top_I.branch[27].block[0].um_I.iw[9] ,
    \top_I.branch[27].block[0].um_I.iw[8] ,
    \top_I.branch[27].block[0].um_I.iw[7] ,
    \top_I.branch[27].block[0].um_I.iw[6] ,
    \top_I.branch[27].block[0].um_I.iw[5] ,
    \top_I.branch[27].block[0].um_I.iw[4] ,
    \top_I.branch[27].block[0].um_I.iw[3] ,
    \top_I.branch[27].block[0].um_I.iw[2] ,
    \top_I.branch[27].block[0].um_I.iw[1] ,
    \top_I.branch[27].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[15].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[14].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[13].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[12].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[11].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[10].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[9].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[8].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[7].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[6].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[5].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[4].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[3].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[2].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[1].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero ,
    \top_I.branch[27].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[27].block[15].um_I.pg_vdd ,
    \top_I.branch[27].block[14].um_I.pg_vdd ,
    \top_I.branch[27].block[13].um_I.pg_vdd ,
    \top_I.branch[27].block[12].um_I.pg_vdd ,
    \top_I.branch[27].block[11].um_I.pg_vdd ,
    \top_I.branch[27].block[10].um_I.pg_vdd ,
    \top_I.branch[27].block[9].um_I.pg_vdd ,
    \top_I.branch[27].block[8].um_I.pg_vdd ,
    \top_I.branch[27].block[7].um_I.pg_vdd ,
    \top_I.branch[27].block[6].um_I.pg_vdd ,
    \top_I.branch[27].block[5].um_I.pg_vdd ,
    \top_I.branch[27].block[4].um_I.pg_vdd ,
    \top_I.branch[27].block[3].um_I.pg_vdd ,
    \top_I.branch[27].block[2].um_I.pg_vdd ,
    \top_I.branch[27].block[1].um_I.pg_vdd ,
    \top_I.branch[27].block[0].um_I.pg_vdd }));
 tt_pg_vdd_1 \top_I.branch[28].block[0].um_I.block_28_0.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[0].um_I.block_28_0.vpwr ),
    .ctrl(\top_I.branch[28].block[0].um_I.pg_vdd ));
 tt_um_haeuslermarkus_fir_filter \top_I.branch[28].block[0].um_I.block_28_0.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[0].um_I.block_28_0.vpwr ),
    .clk(\top_I.branch[28].block[0].um_I.clk ),
    .ena(\top_I.branch[28].block[0].um_I.ena ),
    .rst_n(\top_I.branch[28].block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[0].um_I.iw[9] ,
    \top_I.branch[28].block[0].um_I.iw[8] ,
    \top_I.branch[28].block[0].um_I.iw[7] ,
    \top_I.branch[28].block[0].um_I.iw[6] ,
    \top_I.branch[28].block[0].um_I.iw[5] ,
    \top_I.branch[28].block[0].um_I.iw[4] ,
    \top_I.branch[28].block[0].um_I.iw[3] ,
    \top_I.branch[28].block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[0].um_I.iw[17] ,
    \top_I.branch[28].block[0].um_I.iw[16] ,
    \top_I.branch[28].block[0].um_I.iw[15] ,
    \top_I.branch[28].block[0].um_I.iw[14] ,
    \top_I.branch[28].block[0].um_I.iw[13] ,
    \top_I.branch[28].block[0].um_I.iw[12] ,
    \top_I.branch[28].block[0].um_I.iw[11] ,
    \top_I.branch[28].block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[0].um_I.ow[23] ,
    \top_I.branch[28].block[0].um_I.ow[22] ,
    \top_I.branch[28].block[0].um_I.ow[21] ,
    \top_I.branch[28].block[0].um_I.ow[20] ,
    \top_I.branch[28].block[0].um_I.ow[19] ,
    \top_I.branch[28].block[0].um_I.ow[18] ,
    \top_I.branch[28].block[0].um_I.ow[17] ,
    \top_I.branch[28].block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[0].um_I.ow[15] ,
    \top_I.branch[28].block[0].um_I.ow[14] ,
    \top_I.branch[28].block[0].um_I.ow[13] ,
    \top_I.branch[28].block[0].um_I.ow[12] ,
    \top_I.branch[28].block[0].um_I.ow[11] ,
    \top_I.branch[28].block[0].um_I.ow[10] ,
    \top_I.branch[28].block[0].um_I.ow[9] ,
    \top_I.branch[28].block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[0].um_I.ow[7] ,
    \top_I.branch[28].block[0].um_I.ow[6] ,
    \top_I.branch[28].block[0].um_I.ow[5] ,
    \top_I.branch[28].block[0].um_I.ow[4] ,
    \top_I.branch[28].block[0].um_I.ow[3] ,
    \top_I.branch[28].block[0].um_I.ow[2] ,
    \top_I.branch[28].block[0].um_I.ow[1] ,
    \top_I.branch[28].block[0].um_I.ow[0] }));
 tt_pg_vdd_2 \top_I.branch[28].block[10].um_I.block_28_10.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[10].um_I.block_28_10.vpwr ),
    .ctrl(\top_I.branch[28].block[10].um_I.pg_vdd ));
 tt_um_mattvenn_r2r_dac \top_I.branch[28].block[10].um_I.block_28_10.tt_um_I  (.clk(\top_I.branch[28].block[10].um_I.clk ),
    .ena(\top_I.branch[28].block[10].um_I.ena ),
    .rst_n(\top_I.branch[28].block[10].um_I.iw[1] ),
    .VPWR(\top_I.branch[28].block[10].um_I.block_28_10.vpwr ),
    .VGND(vssd1),
    .ua({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8}),
    .ui_in({\top_I.branch[28].block[10].um_I.iw[9] ,
    \top_I.branch[28].block[10].um_I.iw[8] ,
    \top_I.branch[28].block[10].um_I.iw[7] ,
    \top_I.branch[28].block[10].um_I.iw[6] ,
    \top_I.branch[28].block[10].um_I.iw[5] ,
    \top_I.branch[28].block[10].um_I.iw[4] ,
    \top_I.branch[28].block[10].um_I.iw[3] ,
    \top_I.branch[28].block[10].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[10].um_I.iw[17] ,
    \top_I.branch[28].block[10].um_I.iw[16] ,
    \top_I.branch[28].block[10].um_I.iw[15] ,
    \top_I.branch[28].block[10].um_I.iw[14] ,
    \top_I.branch[28].block[10].um_I.iw[13] ,
    \top_I.branch[28].block[10].um_I.iw[12] ,
    \top_I.branch[28].block[10].um_I.iw[11] ,
    \top_I.branch[28].block[10].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[10].um_I.ow[23] ,
    \top_I.branch[28].block[10].um_I.ow[22] ,
    \top_I.branch[28].block[10].um_I.ow[21] ,
    \top_I.branch[28].block[10].um_I.ow[20] ,
    \top_I.branch[28].block[10].um_I.ow[19] ,
    \top_I.branch[28].block[10].um_I.ow[18] ,
    \top_I.branch[28].block[10].um_I.ow[17] ,
    \top_I.branch[28].block[10].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[10].um_I.ow[15] ,
    \top_I.branch[28].block[10].um_I.ow[14] ,
    \top_I.branch[28].block[10].um_I.ow[13] ,
    \top_I.branch[28].block[10].um_I.ow[12] ,
    \top_I.branch[28].block[10].um_I.ow[11] ,
    \top_I.branch[28].block[10].um_I.ow[10] ,
    \top_I.branch[28].block[10].um_I.ow[9] ,
    \top_I.branch[28].block[10].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[10].um_I.ow[7] ,
    \top_I.branch[28].block[10].um_I.ow[6] ,
    \top_I.branch[28].block[10].um_I.ow[5] ,
    \top_I.branch[28].block[10].um_I.ow[4] ,
    \top_I.branch[28].block[10].um_I.ow[3] ,
    \top_I.branch[28].block[10].um_I.ow[2] ,
    \top_I.branch[28].block[10].um_I.ow[1] ,
    \top_I.branch[28].block[10].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[11].um_I.block_28_11.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[11].um_I.block_28_11.vpwr ),
    .ctrl(\top_I.branch[28].block[11].um_I.pg_vdd ));
 tt_um_iron_violet_simon \top_I.branch[28].block[11].um_I.block_28_11.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[11].um_I.block_28_11.vpwr ),
    .clk(\top_I.branch[28].block[11].um_I.clk ),
    .ena(\top_I.branch[28].block[11].um_I.ena ),
    .rst_n(\top_I.branch[28].block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[11].um_I.iw[9] ,
    \top_I.branch[28].block[11].um_I.iw[8] ,
    \top_I.branch[28].block[11].um_I.iw[7] ,
    \top_I.branch[28].block[11].um_I.iw[6] ,
    \top_I.branch[28].block[11].um_I.iw[5] ,
    \top_I.branch[28].block[11].um_I.iw[4] ,
    \top_I.branch[28].block[11].um_I.iw[3] ,
    \top_I.branch[28].block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[11].um_I.iw[17] ,
    \top_I.branch[28].block[11].um_I.iw[16] ,
    \top_I.branch[28].block[11].um_I.iw[15] ,
    \top_I.branch[28].block[11].um_I.iw[14] ,
    \top_I.branch[28].block[11].um_I.iw[13] ,
    \top_I.branch[28].block[11].um_I.iw[12] ,
    \top_I.branch[28].block[11].um_I.iw[11] ,
    \top_I.branch[28].block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[11].um_I.ow[23] ,
    \top_I.branch[28].block[11].um_I.ow[22] ,
    \top_I.branch[28].block[11].um_I.ow[21] ,
    \top_I.branch[28].block[11].um_I.ow[20] ,
    \top_I.branch[28].block[11].um_I.ow[19] ,
    \top_I.branch[28].block[11].um_I.ow[18] ,
    \top_I.branch[28].block[11].um_I.ow[17] ,
    \top_I.branch[28].block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[11].um_I.ow[15] ,
    \top_I.branch[28].block[11].um_I.ow[14] ,
    \top_I.branch[28].block[11].um_I.ow[13] ,
    \top_I.branch[28].block[11].um_I.ow[12] ,
    \top_I.branch[28].block[11].um_I.ow[11] ,
    \top_I.branch[28].block[11].um_I.ow[10] ,
    \top_I.branch[28].block[11].um_I.ow[9] ,
    \top_I.branch[28].block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[11].um_I.ow[7] ,
    \top_I.branch[28].block[11].um_I.ow[6] ,
    \top_I.branch[28].block[11].um_I.ow[5] ,
    \top_I.branch[28].block[11].um_I.ow[4] ,
    \top_I.branch[28].block[11].um_I.ow[3] ,
    \top_I.branch[28].block[11].um_I.ow[2] ,
    \top_I.branch[28].block[11].um_I.ow[1] ,
    \top_I.branch[28].block[11].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[13].um_I.block_28_13.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[13].um_I.block_28_13.vpwr ),
    .ctrl(\top_I.branch[28].block[13].um_I.pg_vdd ));
 tt_um_alexsegura_pong \top_I.branch[28].block[13].um_I.block_28_13.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[13].um_I.block_28_13.vpwr ),
    .clk(\top_I.branch[28].block[13].um_I.clk ),
    .ena(\top_I.branch[28].block[13].um_I.ena ),
    .rst_n(\top_I.branch[28].block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[13].um_I.iw[9] ,
    \top_I.branch[28].block[13].um_I.iw[8] ,
    \top_I.branch[28].block[13].um_I.iw[7] ,
    \top_I.branch[28].block[13].um_I.iw[6] ,
    \top_I.branch[28].block[13].um_I.iw[5] ,
    \top_I.branch[28].block[13].um_I.iw[4] ,
    \top_I.branch[28].block[13].um_I.iw[3] ,
    \top_I.branch[28].block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[13].um_I.iw[17] ,
    \top_I.branch[28].block[13].um_I.iw[16] ,
    \top_I.branch[28].block[13].um_I.iw[15] ,
    \top_I.branch[28].block[13].um_I.iw[14] ,
    \top_I.branch[28].block[13].um_I.iw[13] ,
    \top_I.branch[28].block[13].um_I.iw[12] ,
    \top_I.branch[28].block[13].um_I.iw[11] ,
    \top_I.branch[28].block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[13].um_I.ow[23] ,
    \top_I.branch[28].block[13].um_I.ow[22] ,
    \top_I.branch[28].block[13].um_I.ow[21] ,
    \top_I.branch[28].block[13].um_I.ow[20] ,
    \top_I.branch[28].block[13].um_I.ow[19] ,
    \top_I.branch[28].block[13].um_I.ow[18] ,
    \top_I.branch[28].block[13].um_I.ow[17] ,
    \top_I.branch[28].block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[13].um_I.ow[15] ,
    \top_I.branch[28].block[13].um_I.ow[14] ,
    \top_I.branch[28].block[13].um_I.ow[13] ,
    \top_I.branch[28].block[13].um_I.ow[12] ,
    \top_I.branch[28].block[13].um_I.ow[11] ,
    \top_I.branch[28].block[13].um_I.ow[10] ,
    \top_I.branch[28].block[13].um_I.ow[9] ,
    \top_I.branch[28].block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[13].um_I.ow[7] ,
    \top_I.branch[28].block[13].um_I.ow[6] ,
    \top_I.branch[28].block[13].um_I.ow[5] ,
    \top_I.branch[28].block[13].um_I.ow[4] ,
    \top_I.branch[28].block[13].um_I.ow[3] ,
    \top_I.branch[28].block[13].um_I.ow[2] ,
    \top_I.branch[28].block[13].um_I.ow[1] ,
    \top_I.branch[28].block[13].um_I.ow[0] }));
 tt_pg_vdd_2 \top_I.branch[28].block[14].um_I.block_28_14.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[14].um_I.block_28_14.vpwr ),
    .ctrl(\top_I.branch[28].block[14].um_I.pg_vdd ));
 tt_um_MichaelBell_tinyQV \top_I.branch[28].block[14].um_I.block_28_14.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[14].um_I.block_28_14.vpwr ),
    .clk(\top_I.branch[28].block[14].um_I.clk ),
    .ena(\top_I.branch[28].block[14].um_I.ena ),
    .rst_n(\top_I.branch[28].block[14].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[14].um_I.iw[9] ,
    \top_I.branch[28].block[14].um_I.iw[8] ,
    \top_I.branch[28].block[14].um_I.iw[7] ,
    \top_I.branch[28].block[14].um_I.iw[6] ,
    \top_I.branch[28].block[14].um_I.iw[5] ,
    \top_I.branch[28].block[14].um_I.iw[4] ,
    \top_I.branch[28].block[14].um_I.iw[3] ,
    \top_I.branch[28].block[14].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[14].um_I.iw[17] ,
    \top_I.branch[28].block[14].um_I.iw[16] ,
    \top_I.branch[28].block[14].um_I.iw[15] ,
    \top_I.branch[28].block[14].um_I.iw[14] ,
    \top_I.branch[28].block[14].um_I.iw[13] ,
    \top_I.branch[28].block[14].um_I.iw[12] ,
    \top_I.branch[28].block[14].um_I.iw[11] ,
    \top_I.branch[28].block[14].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[14].um_I.ow[23] ,
    \top_I.branch[28].block[14].um_I.ow[22] ,
    \top_I.branch[28].block[14].um_I.ow[21] ,
    \top_I.branch[28].block[14].um_I.ow[20] ,
    \top_I.branch[28].block[14].um_I.ow[19] ,
    \top_I.branch[28].block[14].um_I.ow[18] ,
    \top_I.branch[28].block[14].um_I.ow[17] ,
    \top_I.branch[28].block[14].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[14].um_I.ow[15] ,
    \top_I.branch[28].block[14].um_I.ow[14] ,
    \top_I.branch[28].block[14].um_I.ow[13] ,
    \top_I.branch[28].block[14].um_I.ow[12] ,
    \top_I.branch[28].block[14].um_I.ow[11] ,
    \top_I.branch[28].block[14].um_I.ow[10] ,
    \top_I.branch[28].block[14].um_I.ow[9] ,
    \top_I.branch[28].block[14].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[14].um_I.ow[7] ,
    \top_I.branch[28].block[14].um_I.ow[6] ,
    \top_I.branch[28].block[14].um_I.ow[5] ,
    \top_I.branch[28].block[14].um_I.ow[4] ,
    \top_I.branch[28].block[14].um_I.ow[3] ,
    \top_I.branch[28].block[14].um_I.ow[2] ,
    \top_I.branch[28].block[14].um_I.ow[1] ,
    \top_I.branch[28].block[14].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[15].um_I.block_28_15.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[15].um_I.block_28_15.vpwr ),
    .ctrl(\top_I.branch[28].block[15].um_I.pg_vdd ));
 tt_um_coloquinte_moosic \top_I.branch[28].block[15].um_I.block_28_15.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[15].um_I.block_28_15.vpwr ),
    .clk(\top_I.branch[28].block[15].um_I.clk ),
    .ena(\top_I.branch[28].block[15].um_I.ena ),
    .rst_n(\top_I.branch[28].block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[15].um_I.iw[9] ,
    \top_I.branch[28].block[15].um_I.iw[8] ,
    \top_I.branch[28].block[15].um_I.iw[7] ,
    \top_I.branch[28].block[15].um_I.iw[6] ,
    \top_I.branch[28].block[15].um_I.iw[5] ,
    \top_I.branch[28].block[15].um_I.iw[4] ,
    \top_I.branch[28].block[15].um_I.iw[3] ,
    \top_I.branch[28].block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[15].um_I.iw[17] ,
    \top_I.branch[28].block[15].um_I.iw[16] ,
    \top_I.branch[28].block[15].um_I.iw[15] ,
    \top_I.branch[28].block[15].um_I.iw[14] ,
    \top_I.branch[28].block[15].um_I.iw[13] ,
    \top_I.branch[28].block[15].um_I.iw[12] ,
    \top_I.branch[28].block[15].um_I.iw[11] ,
    \top_I.branch[28].block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[15].um_I.ow[23] ,
    \top_I.branch[28].block[15].um_I.ow[22] ,
    \top_I.branch[28].block[15].um_I.ow[21] ,
    \top_I.branch[28].block[15].um_I.ow[20] ,
    \top_I.branch[28].block[15].um_I.ow[19] ,
    \top_I.branch[28].block[15].um_I.ow[18] ,
    \top_I.branch[28].block[15].um_I.ow[17] ,
    \top_I.branch[28].block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[15].um_I.ow[15] ,
    \top_I.branch[28].block[15].um_I.ow[14] ,
    \top_I.branch[28].block[15].um_I.ow[13] ,
    \top_I.branch[28].block[15].um_I.ow[12] ,
    \top_I.branch[28].block[15].um_I.ow[11] ,
    \top_I.branch[28].block[15].um_I.ow[10] ,
    \top_I.branch[28].block[15].um_I.ow[9] ,
    \top_I.branch[28].block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[15].um_I.ow[7] ,
    \top_I.branch[28].block[15].um_I.ow[6] ,
    \top_I.branch[28].block[15].um_I.ow[5] ,
    \top_I.branch[28].block[15].um_I.ow[4] ,
    \top_I.branch[28].block[15].um_I.ow[3] ,
    \top_I.branch[28].block[15].um_I.ow[2] ,
    \top_I.branch[28].block[15].um_I.ow[1] ,
    \top_I.branch[28].block[15].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[1].um_I.block_28_1.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[1].um_I.block_28_1.vpwr ),
    .ctrl(\top_I.branch[28].block[1].um_I.pg_vdd ));
 tt_um_soundgen \top_I.branch[28].block[1].um_I.block_28_1.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[1].um_I.block_28_1.vpwr ),
    .clk(\top_I.branch[28].block[1].um_I.clk ),
    .ena(\top_I.branch[28].block[1].um_I.ena ),
    .rst_n(\top_I.branch[28].block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[1].um_I.iw[9] ,
    \top_I.branch[28].block[1].um_I.iw[8] ,
    \top_I.branch[28].block[1].um_I.iw[7] ,
    \top_I.branch[28].block[1].um_I.iw[6] ,
    \top_I.branch[28].block[1].um_I.iw[5] ,
    \top_I.branch[28].block[1].um_I.iw[4] ,
    \top_I.branch[28].block[1].um_I.iw[3] ,
    \top_I.branch[28].block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[1].um_I.iw[17] ,
    \top_I.branch[28].block[1].um_I.iw[16] ,
    \top_I.branch[28].block[1].um_I.iw[15] ,
    \top_I.branch[28].block[1].um_I.iw[14] ,
    \top_I.branch[28].block[1].um_I.iw[13] ,
    \top_I.branch[28].block[1].um_I.iw[12] ,
    \top_I.branch[28].block[1].um_I.iw[11] ,
    \top_I.branch[28].block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[1].um_I.ow[23] ,
    \top_I.branch[28].block[1].um_I.ow[22] ,
    \top_I.branch[28].block[1].um_I.ow[21] ,
    \top_I.branch[28].block[1].um_I.ow[20] ,
    \top_I.branch[28].block[1].um_I.ow[19] ,
    \top_I.branch[28].block[1].um_I.ow[18] ,
    \top_I.branch[28].block[1].um_I.ow[17] ,
    \top_I.branch[28].block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[1].um_I.ow[15] ,
    \top_I.branch[28].block[1].um_I.ow[14] ,
    \top_I.branch[28].block[1].um_I.ow[13] ,
    \top_I.branch[28].block[1].um_I.ow[12] ,
    \top_I.branch[28].block[1].um_I.ow[11] ,
    \top_I.branch[28].block[1].um_I.ow[10] ,
    \top_I.branch[28].block[1].um_I.ow[9] ,
    \top_I.branch[28].block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[1].um_I.ow[7] ,
    \top_I.branch[28].block[1].um_I.ow[6] ,
    \top_I.branch[28].block[1].um_I.ow[5] ,
    \top_I.branch[28].block[1].um_I.ow[4] ,
    \top_I.branch[28].block[1].um_I.ow[3] ,
    \top_I.branch[28].block[1].um_I.ow[2] ,
    \top_I.branch[28].block[1].um_I.ow[1] ,
    \top_I.branch[28].block[1].um_I.ow[0] }));
 tt_pg_vdd_2 \top_I.branch[28].block[2].um_I.block_28_2.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[2].um_I.block_28_2.vpwr ),
    .ctrl(\top_I.branch[28].block[2].um_I.pg_vdd ));
 tt_um_analog_loopback \top_I.branch[28].block[2].um_I.block_28_2.tt_um_I  (.clk(\top_I.branch[28].block[2].um_I.clk ),
    .ena(\top_I.branch[28].block[2].um_I.ena ),
    .rst_n(\top_I.branch[28].block[2].um_I.iw[1] ),
    .VPWR(\top_I.branch[28].block[2].um_I.block_28_2.vpwr ),
    .VGND(vssd1),
    .ua({_NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16}),
    .ui_in({\top_I.branch[28].block[2].um_I.iw[9] ,
    \top_I.branch[28].block[2].um_I.iw[8] ,
    \top_I.branch[28].block[2].um_I.iw[7] ,
    \top_I.branch[28].block[2].um_I.iw[6] ,
    \top_I.branch[28].block[2].um_I.iw[5] ,
    \top_I.branch[28].block[2].um_I.iw[4] ,
    \top_I.branch[28].block[2].um_I.iw[3] ,
    \top_I.branch[28].block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[2].um_I.iw[17] ,
    \top_I.branch[28].block[2].um_I.iw[16] ,
    \top_I.branch[28].block[2].um_I.iw[15] ,
    \top_I.branch[28].block[2].um_I.iw[14] ,
    \top_I.branch[28].block[2].um_I.iw[13] ,
    \top_I.branch[28].block[2].um_I.iw[12] ,
    \top_I.branch[28].block[2].um_I.iw[11] ,
    \top_I.branch[28].block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[2].um_I.ow[23] ,
    \top_I.branch[28].block[2].um_I.ow[22] ,
    \top_I.branch[28].block[2].um_I.ow[21] ,
    \top_I.branch[28].block[2].um_I.ow[20] ,
    \top_I.branch[28].block[2].um_I.ow[19] ,
    \top_I.branch[28].block[2].um_I.ow[18] ,
    \top_I.branch[28].block[2].um_I.ow[17] ,
    \top_I.branch[28].block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[2].um_I.ow[15] ,
    \top_I.branch[28].block[2].um_I.ow[14] ,
    \top_I.branch[28].block[2].um_I.ow[13] ,
    \top_I.branch[28].block[2].um_I.ow[12] ,
    \top_I.branch[28].block[2].um_I.ow[11] ,
    \top_I.branch[28].block[2].um_I.ow[10] ,
    \top_I.branch[28].block[2].um_I.ow[9] ,
    \top_I.branch[28].block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[2].um_I.ow[7] ,
    \top_I.branch[28].block[2].um_I.ow[6] ,
    \top_I.branch[28].block[2].um_I.ow[5] ,
    \top_I.branch[28].block[2].um_I.ow[4] ,
    \top_I.branch[28].block[2].um_I.ow[3] ,
    \top_I.branch[28].block[2].um_I.ow[2] ,
    \top_I.branch[28].block[2].um_I.ow[1] ,
    \top_I.branch[28].block[2].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[3].um_I.block_28_3.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[3].um_I.block_28_3.vpwr ),
    .ctrl(\top_I.branch[28].block[3].um_I.pg_vdd ));
 tt_um_urish_simon \top_I.branch[28].block[3].um_I.block_28_3.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[3].um_I.block_28_3.vpwr ),
    .clk(\top_I.branch[28].block[3].um_I.clk ),
    .ena(\top_I.branch[28].block[3].um_I.ena ),
    .rst_n(\top_I.branch[28].block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[3].um_I.iw[9] ,
    \top_I.branch[28].block[3].um_I.iw[8] ,
    \top_I.branch[28].block[3].um_I.iw[7] ,
    \top_I.branch[28].block[3].um_I.iw[6] ,
    \top_I.branch[28].block[3].um_I.iw[5] ,
    \top_I.branch[28].block[3].um_I.iw[4] ,
    \top_I.branch[28].block[3].um_I.iw[3] ,
    \top_I.branch[28].block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[3].um_I.iw[17] ,
    \top_I.branch[28].block[3].um_I.iw[16] ,
    \top_I.branch[28].block[3].um_I.iw[15] ,
    \top_I.branch[28].block[3].um_I.iw[14] ,
    \top_I.branch[28].block[3].um_I.iw[13] ,
    \top_I.branch[28].block[3].um_I.iw[12] ,
    \top_I.branch[28].block[3].um_I.iw[11] ,
    \top_I.branch[28].block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[3].um_I.ow[23] ,
    \top_I.branch[28].block[3].um_I.ow[22] ,
    \top_I.branch[28].block[3].um_I.ow[21] ,
    \top_I.branch[28].block[3].um_I.ow[20] ,
    \top_I.branch[28].block[3].um_I.ow[19] ,
    \top_I.branch[28].block[3].um_I.ow[18] ,
    \top_I.branch[28].block[3].um_I.ow[17] ,
    \top_I.branch[28].block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[3].um_I.ow[15] ,
    \top_I.branch[28].block[3].um_I.ow[14] ,
    \top_I.branch[28].block[3].um_I.ow[13] ,
    \top_I.branch[28].block[3].um_I.ow[12] ,
    \top_I.branch[28].block[3].um_I.ow[11] ,
    \top_I.branch[28].block[3].um_I.ow[10] ,
    \top_I.branch[28].block[3].um_I.ow[9] ,
    \top_I.branch[28].block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[3].um_I.ow[7] ,
    \top_I.branch[28].block[3].um_I.ow[6] ,
    \top_I.branch[28].block[3].um_I.ow[5] ,
    \top_I.branch[28].block[3].um_I.ow[4] ,
    \top_I.branch[28].block[3].um_I.ow[3] ,
    \top_I.branch[28].block[3].um_I.ow[2] ,
    \top_I.branch[28].block[3].um_I.ow[1] ,
    \top_I.branch[28].block[3].um_I.ow[0] }));
 tt_pg_vdd_2 \top_I.branch[28].block[4].um_I.block_28_4.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[4].um_I.block_28_4.vpwr ),
    .ctrl(\top_I.branch[28].block[4].um_I.pg_vdd ));
 tt_um_histefan_top \top_I.branch[28].block[4].um_I.block_28_4.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[4].um_I.block_28_4.vpwr ),
    .clk(\top_I.branch[28].block[4].um_I.clk ),
    .ena(\top_I.branch[28].block[4].um_I.ena ),
    .rst_n(\top_I.branch[28].block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[4].um_I.iw[9] ,
    \top_I.branch[28].block[4].um_I.iw[8] ,
    \top_I.branch[28].block[4].um_I.iw[7] ,
    \top_I.branch[28].block[4].um_I.iw[6] ,
    \top_I.branch[28].block[4].um_I.iw[5] ,
    \top_I.branch[28].block[4].um_I.iw[4] ,
    \top_I.branch[28].block[4].um_I.iw[3] ,
    \top_I.branch[28].block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[4].um_I.iw[17] ,
    \top_I.branch[28].block[4].um_I.iw[16] ,
    \top_I.branch[28].block[4].um_I.iw[15] ,
    \top_I.branch[28].block[4].um_I.iw[14] ,
    \top_I.branch[28].block[4].um_I.iw[13] ,
    \top_I.branch[28].block[4].um_I.iw[12] ,
    \top_I.branch[28].block[4].um_I.iw[11] ,
    \top_I.branch[28].block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[4].um_I.ow[23] ,
    \top_I.branch[28].block[4].um_I.ow[22] ,
    \top_I.branch[28].block[4].um_I.ow[21] ,
    \top_I.branch[28].block[4].um_I.ow[20] ,
    \top_I.branch[28].block[4].um_I.ow[19] ,
    \top_I.branch[28].block[4].um_I.ow[18] ,
    \top_I.branch[28].block[4].um_I.ow[17] ,
    \top_I.branch[28].block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[4].um_I.ow[15] ,
    \top_I.branch[28].block[4].um_I.ow[14] ,
    \top_I.branch[28].block[4].um_I.ow[13] ,
    \top_I.branch[28].block[4].um_I.ow[12] ,
    \top_I.branch[28].block[4].um_I.ow[11] ,
    \top_I.branch[28].block[4].um_I.ow[10] ,
    \top_I.branch[28].block[4].um_I.ow[9] ,
    \top_I.branch[28].block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[4].um_I.ow[7] ,
    \top_I.branch[28].block[4].um_I.ow[6] ,
    \top_I.branch[28].block[4].um_I.ow[5] ,
    \top_I.branch[28].block[4].um_I.ow[4] ,
    \top_I.branch[28].block[4].um_I.ow[3] ,
    \top_I.branch[28].block[4].um_I.ow[2] ,
    \top_I.branch[28].block[4].um_I.ow[1] ,
    \top_I.branch[28].block[4].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[5].um_I.block_28_5.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[5].um_I.block_28_5.vpwr ),
    .ctrl(\top_I.branch[28].block[5].um_I.pg_vdd ));
 tt_um_faramire_gate_guesser \top_I.branch[28].block[5].um_I.block_28_5.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[5].um_I.block_28_5.vpwr ),
    .clk(\top_I.branch[28].block[5].um_I.clk ),
    .ena(\top_I.branch[28].block[5].um_I.ena ),
    .rst_n(\top_I.branch[28].block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[5].um_I.iw[9] ,
    \top_I.branch[28].block[5].um_I.iw[8] ,
    \top_I.branch[28].block[5].um_I.iw[7] ,
    \top_I.branch[28].block[5].um_I.iw[6] ,
    \top_I.branch[28].block[5].um_I.iw[5] ,
    \top_I.branch[28].block[5].um_I.iw[4] ,
    \top_I.branch[28].block[5].um_I.iw[3] ,
    \top_I.branch[28].block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[5].um_I.iw[17] ,
    \top_I.branch[28].block[5].um_I.iw[16] ,
    \top_I.branch[28].block[5].um_I.iw[15] ,
    \top_I.branch[28].block[5].um_I.iw[14] ,
    \top_I.branch[28].block[5].um_I.iw[13] ,
    \top_I.branch[28].block[5].um_I.iw[12] ,
    \top_I.branch[28].block[5].um_I.iw[11] ,
    \top_I.branch[28].block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[5].um_I.ow[23] ,
    \top_I.branch[28].block[5].um_I.ow[22] ,
    \top_I.branch[28].block[5].um_I.ow[21] ,
    \top_I.branch[28].block[5].um_I.ow[20] ,
    \top_I.branch[28].block[5].um_I.ow[19] ,
    \top_I.branch[28].block[5].um_I.ow[18] ,
    \top_I.branch[28].block[5].um_I.ow[17] ,
    \top_I.branch[28].block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[5].um_I.ow[15] ,
    \top_I.branch[28].block[5].um_I.ow[14] ,
    \top_I.branch[28].block[5].um_I.ow[13] ,
    \top_I.branch[28].block[5].um_I.ow[12] ,
    \top_I.branch[28].block[5].um_I.ow[11] ,
    \top_I.branch[28].block[5].um_I.ow[10] ,
    \top_I.branch[28].block[5].um_I.ow[9] ,
    \top_I.branch[28].block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[5].um_I.ow[7] ,
    \top_I.branch[28].block[5].um_I.ow[6] ,
    \top_I.branch[28].block[5].um_I.ow[5] ,
    \top_I.branch[28].block[5].um_I.ow[4] ,
    \top_I.branch[28].block[5].um_I.ow[3] ,
    \top_I.branch[28].block[5].um_I.ow[2] ,
    \top_I.branch[28].block[5].um_I.ow[1] ,
    \top_I.branch[28].block[5].um_I.ow[0] }));
 tt_pg_vdd_2 \top_I.branch[28].block[6].um_I.block_28_6.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[6].um_I.block_28_6.vpwr ),
    .ctrl(\top_I.branch[28].block[6].um_I.pg_vdd ));
 tt_um_TT06_SAR_wulffern \top_I.branch[28].block[6].um_I.block_28_6.tt_um_I  (.clk(\top_I.branch[28].block[6].um_I.clk ),
    .ena(\top_I.branch[28].block[6].um_I.ena ),
    .rst_n(\top_I.branch[28].block[6].um_I.iw[1] ),
    .VPWR(\top_I.branch[28].block[6].um_I.block_28_6.vpwr ),
    .VGND(vssd1),
    .ua({_NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24}),
    .ui_in({\top_I.branch[28].block[6].um_I.iw[9] ,
    \top_I.branch[28].block[6].um_I.iw[8] ,
    \top_I.branch[28].block[6].um_I.iw[7] ,
    \top_I.branch[28].block[6].um_I.iw[6] ,
    \top_I.branch[28].block[6].um_I.iw[5] ,
    \top_I.branch[28].block[6].um_I.iw[4] ,
    \top_I.branch[28].block[6].um_I.iw[3] ,
    \top_I.branch[28].block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[6].um_I.iw[17] ,
    \top_I.branch[28].block[6].um_I.iw[16] ,
    \top_I.branch[28].block[6].um_I.iw[15] ,
    \top_I.branch[28].block[6].um_I.iw[14] ,
    \top_I.branch[28].block[6].um_I.iw[13] ,
    \top_I.branch[28].block[6].um_I.iw[12] ,
    \top_I.branch[28].block[6].um_I.iw[11] ,
    \top_I.branch[28].block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[6].um_I.ow[23] ,
    \top_I.branch[28].block[6].um_I.ow[22] ,
    \top_I.branch[28].block[6].um_I.ow[21] ,
    \top_I.branch[28].block[6].um_I.ow[20] ,
    \top_I.branch[28].block[6].um_I.ow[19] ,
    \top_I.branch[28].block[6].um_I.ow[18] ,
    \top_I.branch[28].block[6].um_I.ow[17] ,
    \top_I.branch[28].block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[6].um_I.ow[15] ,
    \top_I.branch[28].block[6].um_I.ow[14] ,
    \top_I.branch[28].block[6].um_I.ow[13] ,
    \top_I.branch[28].block[6].um_I.ow[12] ,
    \top_I.branch[28].block[6].um_I.ow[11] ,
    \top_I.branch[28].block[6].um_I.ow[10] ,
    \top_I.branch[28].block[6].um_I.ow[9] ,
    \top_I.branch[28].block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[6].um_I.ow[7] ,
    \top_I.branch[28].block[6].um_I.ow[6] ,
    \top_I.branch[28].block[6].um_I.ow[5] ,
    \top_I.branch[28].block[6].um_I.ow[4] ,
    \top_I.branch[28].block[6].um_I.ow[3] ,
    \top_I.branch[28].block[6].um_I.ow[2] ,
    \top_I.branch[28].block[6].um_I.ow[1] ,
    \top_I.branch[28].block[6].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[7].um_I.block_28_7.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[7].um_I.block_28_7.vpwr ),
    .ctrl(\top_I.branch[28].block[7].um_I.pg_vdd ));
 tt_um_andychip1_sn74169 \top_I.branch[28].block[7].um_I.block_28_7.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[7].um_I.block_28_7.vpwr ),
    .clk(\top_I.branch[28].block[7].um_I.clk ),
    .ena(\top_I.branch[28].block[7].um_I.ena ),
    .rst_n(\top_I.branch[28].block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[7].um_I.iw[9] ,
    \top_I.branch[28].block[7].um_I.iw[8] ,
    \top_I.branch[28].block[7].um_I.iw[7] ,
    \top_I.branch[28].block[7].um_I.iw[6] ,
    \top_I.branch[28].block[7].um_I.iw[5] ,
    \top_I.branch[28].block[7].um_I.iw[4] ,
    \top_I.branch[28].block[7].um_I.iw[3] ,
    \top_I.branch[28].block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[7].um_I.iw[17] ,
    \top_I.branch[28].block[7].um_I.iw[16] ,
    \top_I.branch[28].block[7].um_I.iw[15] ,
    \top_I.branch[28].block[7].um_I.iw[14] ,
    \top_I.branch[28].block[7].um_I.iw[13] ,
    \top_I.branch[28].block[7].um_I.iw[12] ,
    \top_I.branch[28].block[7].um_I.iw[11] ,
    \top_I.branch[28].block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[7].um_I.ow[23] ,
    \top_I.branch[28].block[7].um_I.ow[22] ,
    \top_I.branch[28].block[7].um_I.ow[21] ,
    \top_I.branch[28].block[7].um_I.ow[20] ,
    \top_I.branch[28].block[7].um_I.ow[19] ,
    \top_I.branch[28].block[7].um_I.ow[18] ,
    \top_I.branch[28].block[7].um_I.ow[17] ,
    \top_I.branch[28].block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[7].um_I.ow[15] ,
    \top_I.branch[28].block[7].um_I.ow[14] ,
    \top_I.branch[28].block[7].um_I.ow[13] ,
    \top_I.branch[28].block[7].um_I.ow[12] ,
    \top_I.branch[28].block[7].um_I.ow[11] ,
    \top_I.branch[28].block[7].um_I.ow[10] ,
    \top_I.branch[28].block[7].um_I.ow[9] ,
    \top_I.branch[28].block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[7].um_I.ow[7] ,
    \top_I.branch[28].block[7].um_I.ow[6] ,
    \top_I.branch[28].block[7].um_I.ow[5] ,
    \top_I.branch[28].block[7].um_I.ow[4] ,
    \top_I.branch[28].block[7].um_I.ow[3] ,
    \top_I.branch[28].block[7].um_I.ow[2] ,
    \top_I.branch[28].block[7].um_I.ow[1] ,
    \top_I.branch[28].block[7].um_I.ow[0] }));
 tt_pg_vdd_2 \top_I.branch[28].block[8].um_I.block_28_8.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[8].um_I.block_28_8.vpwr ),
    .ctrl(\top_I.branch[28].block[8].um_I.pg_vdd ));
 tt_um_thorkn_audiochip_v2 \top_I.branch[28].block[8].um_I.block_28_8.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[8].um_I.block_28_8.vpwr ),
    .clk(\top_I.branch[28].block[8].um_I.clk ),
    .ena(\top_I.branch[28].block[8].um_I.ena ),
    .rst_n(\top_I.branch[28].block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[8].um_I.iw[9] ,
    \top_I.branch[28].block[8].um_I.iw[8] ,
    \top_I.branch[28].block[8].um_I.iw[7] ,
    \top_I.branch[28].block[8].um_I.iw[6] ,
    \top_I.branch[28].block[8].um_I.iw[5] ,
    \top_I.branch[28].block[8].um_I.iw[4] ,
    \top_I.branch[28].block[8].um_I.iw[3] ,
    \top_I.branch[28].block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[8].um_I.iw[17] ,
    \top_I.branch[28].block[8].um_I.iw[16] ,
    \top_I.branch[28].block[8].um_I.iw[15] ,
    \top_I.branch[28].block[8].um_I.iw[14] ,
    \top_I.branch[28].block[8].um_I.iw[13] ,
    \top_I.branch[28].block[8].um_I.iw[12] ,
    \top_I.branch[28].block[8].um_I.iw[11] ,
    \top_I.branch[28].block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[8].um_I.ow[23] ,
    \top_I.branch[28].block[8].um_I.ow[22] ,
    \top_I.branch[28].block[8].um_I.ow[21] ,
    \top_I.branch[28].block[8].um_I.ow[20] ,
    \top_I.branch[28].block[8].um_I.ow[19] ,
    \top_I.branch[28].block[8].um_I.ow[18] ,
    \top_I.branch[28].block[8].um_I.ow[17] ,
    \top_I.branch[28].block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[8].um_I.ow[15] ,
    \top_I.branch[28].block[8].um_I.ow[14] ,
    \top_I.branch[28].block[8].um_I.ow[13] ,
    \top_I.branch[28].block[8].um_I.ow[12] ,
    \top_I.branch[28].block[8].um_I.ow[11] ,
    \top_I.branch[28].block[8].um_I.ow[10] ,
    \top_I.branch[28].block[8].um_I.ow[9] ,
    \top_I.branch[28].block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[8].um_I.ow[7] ,
    \top_I.branch[28].block[8].um_I.ow[6] ,
    \top_I.branch[28].block[8].um_I.ow[5] ,
    \top_I.branch[28].block[8].um_I.ow[4] ,
    \top_I.branch[28].block[8].um_I.ow[3] ,
    \top_I.branch[28].block[8].um_I.ow[2] ,
    \top_I.branch[28].block[8].um_I.ow[1] ,
    \top_I.branch[28].block[8].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[28].block[9].um_I.block_28_9.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[28].block[9].um_I.block_28_9.vpwr ),
    .ctrl(\top_I.branch[28].block[9].um_I.pg_vdd ));
 tt_um_tomkeddie_a \top_I.branch[28].block[9].um_I.block_28_9.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[28].block[9].um_I.block_28_9.vpwr ),
    .clk(\top_I.branch[28].block[9].um_I.clk ),
    .ena(\top_I.branch[28].block[9].um_I.ena ),
    .rst_n(\top_I.branch[28].block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[28].block[9].um_I.iw[9] ,
    \top_I.branch[28].block[9].um_I.iw[8] ,
    \top_I.branch[28].block[9].um_I.iw[7] ,
    \top_I.branch[28].block[9].um_I.iw[6] ,
    \top_I.branch[28].block[9].um_I.iw[5] ,
    \top_I.branch[28].block[9].um_I.iw[4] ,
    \top_I.branch[28].block[9].um_I.iw[3] ,
    \top_I.branch[28].block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[28].block[9].um_I.iw[17] ,
    \top_I.branch[28].block[9].um_I.iw[16] ,
    \top_I.branch[28].block[9].um_I.iw[15] ,
    \top_I.branch[28].block[9].um_I.iw[14] ,
    \top_I.branch[28].block[9].um_I.iw[13] ,
    \top_I.branch[28].block[9].um_I.iw[12] ,
    \top_I.branch[28].block[9].um_I.iw[11] ,
    \top_I.branch[28].block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[28].block[9].um_I.ow[23] ,
    \top_I.branch[28].block[9].um_I.ow[22] ,
    \top_I.branch[28].block[9].um_I.ow[21] ,
    \top_I.branch[28].block[9].um_I.ow[20] ,
    \top_I.branch[28].block[9].um_I.ow[19] ,
    \top_I.branch[28].block[9].um_I.ow[18] ,
    \top_I.branch[28].block[9].um_I.ow[17] ,
    \top_I.branch[28].block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[28].block[9].um_I.ow[15] ,
    \top_I.branch[28].block[9].um_I.ow[14] ,
    \top_I.branch[28].block[9].um_I.ow[13] ,
    \top_I.branch[28].block[9].um_I.ow[12] ,
    \top_I.branch[28].block[9].um_I.ow[11] ,
    \top_I.branch[28].block[9].um_I.ow[10] ,
    \top_I.branch[28].block[9].um_I.ow[9] ,
    \top_I.branch[28].block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[28].block[9].um_I.ow[7] ,
    \top_I.branch[28].block[9].um_I.ow[6] ,
    \top_I.branch[28].block[9].um_I.ow[5] ,
    \top_I.branch[28].block[9].um_I.ow[4] ,
    \top_I.branch[28].block[9].um_I.ow[3] ,
    \top_I.branch[28].block[9].um_I.ow[2] ,
    \top_I.branch[28].block[9].um_I.ow[1] ,
    \top_I.branch[28].block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[28].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[28].l_addr[1] ),
    .k_zero(\top_I.branch[28].l_addr[0] ),
    .addr({\top_I.branch[28].l_addr[1] ,
    \top_I.branch[28].l_addr[1] ,
    \top_I.branch[28].l_addr[1] ,
    \top_I.branch[28].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[28].block[15].um_I.ena ,
    \top_I.branch[28].block[14].um_I.ena ,
    \top_I.branch[28].block[13].um_I.ena ,
    \top_I.branch[28].block[12].um_I.ena ,
    \top_I.branch[28].block[11].um_I.ena ,
    \top_I.branch[28].block[10].um_I.ena ,
    \top_I.branch[28].block[9].um_I.ena ,
    \top_I.branch[28].block[8].um_I.ena ,
    \top_I.branch[28].block[7].um_I.ena ,
    \top_I.branch[28].block[6].um_I.ena ,
    \top_I.branch[28].block[5].um_I.ena ,
    \top_I.branch[28].block[4].um_I.ena ,
    \top_I.branch[28].block[3].um_I.ena ,
    \top_I.branch[28].block[2].um_I.ena ,
    \top_I.branch[28].block[1].um_I.ena ,
    \top_I.branch[28].block[0].um_I.ena }),
    .um_iw({\top_I.branch[28].block[15].um_I.iw[17] ,
    \top_I.branch[28].block[15].um_I.iw[16] ,
    \top_I.branch[28].block[15].um_I.iw[15] ,
    \top_I.branch[28].block[15].um_I.iw[14] ,
    \top_I.branch[28].block[15].um_I.iw[13] ,
    \top_I.branch[28].block[15].um_I.iw[12] ,
    \top_I.branch[28].block[15].um_I.iw[11] ,
    \top_I.branch[28].block[15].um_I.iw[10] ,
    \top_I.branch[28].block[15].um_I.iw[9] ,
    \top_I.branch[28].block[15].um_I.iw[8] ,
    \top_I.branch[28].block[15].um_I.iw[7] ,
    \top_I.branch[28].block[15].um_I.iw[6] ,
    \top_I.branch[28].block[15].um_I.iw[5] ,
    \top_I.branch[28].block[15].um_I.iw[4] ,
    \top_I.branch[28].block[15].um_I.iw[3] ,
    \top_I.branch[28].block[15].um_I.iw[2] ,
    \top_I.branch[28].block[15].um_I.iw[1] ,
    \top_I.branch[28].block[15].um_I.clk ,
    \top_I.branch[28].block[14].um_I.iw[17] ,
    \top_I.branch[28].block[14].um_I.iw[16] ,
    \top_I.branch[28].block[14].um_I.iw[15] ,
    \top_I.branch[28].block[14].um_I.iw[14] ,
    \top_I.branch[28].block[14].um_I.iw[13] ,
    \top_I.branch[28].block[14].um_I.iw[12] ,
    \top_I.branch[28].block[14].um_I.iw[11] ,
    \top_I.branch[28].block[14].um_I.iw[10] ,
    \top_I.branch[28].block[14].um_I.iw[9] ,
    \top_I.branch[28].block[14].um_I.iw[8] ,
    \top_I.branch[28].block[14].um_I.iw[7] ,
    \top_I.branch[28].block[14].um_I.iw[6] ,
    \top_I.branch[28].block[14].um_I.iw[5] ,
    \top_I.branch[28].block[14].um_I.iw[4] ,
    \top_I.branch[28].block[14].um_I.iw[3] ,
    \top_I.branch[28].block[14].um_I.iw[2] ,
    \top_I.branch[28].block[14].um_I.iw[1] ,
    \top_I.branch[28].block[14].um_I.clk ,
    \top_I.branch[28].block[13].um_I.iw[17] ,
    \top_I.branch[28].block[13].um_I.iw[16] ,
    \top_I.branch[28].block[13].um_I.iw[15] ,
    \top_I.branch[28].block[13].um_I.iw[14] ,
    \top_I.branch[28].block[13].um_I.iw[13] ,
    \top_I.branch[28].block[13].um_I.iw[12] ,
    \top_I.branch[28].block[13].um_I.iw[11] ,
    \top_I.branch[28].block[13].um_I.iw[10] ,
    \top_I.branch[28].block[13].um_I.iw[9] ,
    \top_I.branch[28].block[13].um_I.iw[8] ,
    \top_I.branch[28].block[13].um_I.iw[7] ,
    \top_I.branch[28].block[13].um_I.iw[6] ,
    \top_I.branch[28].block[13].um_I.iw[5] ,
    \top_I.branch[28].block[13].um_I.iw[4] ,
    \top_I.branch[28].block[13].um_I.iw[3] ,
    \top_I.branch[28].block[13].um_I.iw[2] ,
    \top_I.branch[28].block[13].um_I.iw[1] ,
    \top_I.branch[28].block[13].um_I.clk ,
    \top_I.branch[28].block[12].um_I.iw[17] ,
    \top_I.branch[28].block[12].um_I.iw[16] ,
    \top_I.branch[28].block[12].um_I.iw[15] ,
    \top_I.branch[28].block[12].um_I.iw[14] ,
    \top_I.branch[28].block[12].um_I.iw[13] ,
    \top_I.branch[28].block[12].um_I.iw[12] ,
    \top_I.branch[28].block[12].um_I.iw[11] ,
    \top_I.branch[28].block[12].um_I.iw[10] ,
    \top_I.branch[28].block[12].um_I.iw[9] ,
    \top_I.branch[28].block[12].um_I.iw[8] ,
    \top_I.branch[28].block[12].um_I.iw[7] ,
    \top_I.branch[28].block[12].um_I.iw[6] ,
    \top_I.branch[28].block[12].um_I.iw[5] ,
    \top_I.branch[28].block[12].um_I.iw[4] ,
    \top_I.branch[28].block[12].um_I.iw[3] ,
    \top_I.branch[28].block[12].um_I.iw[2] ,
    \top_I.branch[28].block[12].um_I.iw[1] ,
    \top_I.branch[28].block[12].um_I.clk ,
    \top_I.branch[28].block[11].um_I.iw[17] ,
    \top_I.branch[28].block[11].um_I.iw[16] ,
    \top_I.branch[28].block[11].um_I.iw[15] ,
    \top_I.branch[28].block[11].um_I.iw[14] ,
    \top_I.branch[28].block[11].um_I.iw[13] ,
    \top_I.branch[28].block[11].um_I.iw[12] ,
    \top_I.branch[28].block[11].um_I.iw[11] ,
    \top_I.branch[28].block[11].um_I.iw[10] ,
    \top_I.branch[28].block[11].um_I.iw[9] ,
    \top_I.branch[28].block[11].um_I.iw[8] ,
    \top_I.branch[28].block[11].um_I.iw[7] ,
    \top_I.branch[28].block[11].um_I.iw[6] ,
    \top_I.branch[28].block[11].um_I.iw[5] ,
    \top_I.branch[28].block[11].um_I.iw[4] ,
    \top_I.branch[28].block[11].um_I.iw[3] ,
    \top_I.branch[28].block[11].um_I.iw[2] ,
    \top_I.branch[28].block[11].um_I.iw[1] ,
    \top_I.branch[28].block[11].um_I.clk ,
    \top_I.branch[28].block[10].um_I.iw[17] ,
    \top_I.branch[28].block[10].um_I.iw[16] ,
    \top_I.branch[28].block[10].um_I.iw[15] ,
    \top_I.branch[28].block[10].um_I.iw[14] ,
    \top_I.branch[28].block[10].um_I.iw[13] ,
    \top_I.branch[28].block[10].um_I.iw[12] ,
    \top_I.branch[28].block[10].um_I.iw[11] ,
    \top_I.branch[28].block[10].um_I.iw[10] ,
    \top_I.branch[28].block[10].um_I.iw[9] ,
    \top_I.branch[28].block[10].um_I.iw[8] ,
    \top_I.branch[28].block[10].um_I.iw[7] ,
    \top_I.branch[28].block[10].um_I.iw[6] ,
    \top_I.branch[28].block[10].um_I.iw[5] ,
    \top_I.branch[28].block[10].um_I.iw[4] ,
    \top_I.branch[28].block[10].um_I.iw[3] ,
    \top_I.branch[28].block[10].um_I.iw[2] ,
    \top_I.branch[28].block[10].um_I.iw[1] ,
    \top_I.branch[28].block[10].um_I.clk ,
    \top_I.branch[28].block[9].um_I.iw[17] ,
    \top_I.branch[28].block[9].um_I.iw[16] ,
    \top_I.branch[28].block[9].um_I.iw[15] ,
    \top_I.branch[28].block[9].um_I.iw[14] ,
    \top_I.branch[28].block[9].um_I.iw[13] ,
    \top_I.branch[28].block[9].um_I.iw[12] ,
    \top_I.branch[28].block[9].um_I.iw[11] ,
    \top_I.branch[28].block[9].um_I.iw[10] ,
    \top_I.branch[28].block[9].um_I.iw[9] ,
    \top_I.branch[28].block[9].um_I.iw[8] ,
    \top_I.branch[28].block[9].um_I.iw[7] ,
    \top_I.branch[28].block[9].um_I.iw[6] ,
    \top_I.branch[28].block[9].um_I.iw[5] ,
    \top_I.branch[28].block[9].um_I.iw[4] ,
    \top_I.branch[28].block[9].um_I.iw[3] ,
    \top_I.branch[28].block[9].um_I.iw[2] ,
    \top_I.branch[28].block[9].um_I.iw[1] ,
    \top_I.branch[28].block[9].um_I.clk ,
    \top_I.branch[28].block[8].um_I.iw[17] ,
    \top_I.branch[28].block[8].um_I.iw[16] ,
    \top_I.branch[28].block[8].um_I.iw[15] ,
    \top_I.branch[28].block[8].um_I.iw[14] ,
    \top_I.branch[28].block[8].um_I.iw[13] ,
    \top_I.branch[28].block[8].um_I.iw[12] ,
    \top_I.branch[28].block[8].um_I.iw[11] ,
    \top_I.branch[28].block[8].um_I.iw[10] ,
    \top_I.branch[28].block[8].um_I.iw[9] ,
    \top_I.branch[28].block[8].um_I.iw[8] ,
    \top_I.branch[28].block[8].um_I.iw[7] ,
    \top_I.branch[28].block[8].um_I.iw[6] ,
    \top_I.branch[28].block[8].um_I.iw[5] ,
    \top_I.branch[28].block[8].um_I.iw[4] ,
    \top_I.branch[28].block[8].um_I.iw[3] ,
    \top_I.branch[28].block[8].um_I.iw[2] ,
    \top_I.branch[28].block[8].um_I.iw[1] ,
    \top_I.branch[28].block[8].um_I.clk ,
    \top_I.branch[28].block[7].um_I.iw[17] ,
    \top_I.branch[28].block[7].um_I.iw[16] ,
    \top_I.branch[28].block[7].um_I.iw[15] ,
    \top_I.branch[28].block[7].um_I.iw[14] ,
    \top_I.branch[28].block[7].um_I.iw[13] ,
    \top_I.branch[28].block[7].um_I.iw[12] ,
    \top_I.branch[28].block[7].um_I.iw[11] ,
    \top_I.branch[28].block[7].um_I.iw[10] ,
    \top_I.branch[28].block[7].um_I.iw[9] ,
    \top_I.branch[28].block[7].um_I.iw[8] ,
    \top_I.branch[28].block[7].um_I.iw[7] ,
    \top_I.branch[28].block[7].um_I.iw[6] ,
    \top_I.branch[28].block[7].um_I.iw[5] ,
    \top_I.branch[28].block[7].um_I.iw[4] ,
    \top_I.branch[28].block[7].um_I.iw[3] ,
    \top_I.branch[28].block[7].um_I.iw[2] ,
    \top_I.branch[28].block[7].um_I.iw[1] ,
    \top_I.branch[28].block[7].um_I.clk ,
    \top_I.branch[28].block[6].um_I.iw[17] ,
    \top_I.branch[28].block[6].um_I.iw[16] ,
    \top_I.branch[28].block[6].um_I.iw[15] ,
    \top_I.branch[28].block[6].um_I.iw[14] ,
    \top_I.branch[28].block[6].um_I.iw[13] ,
    \top_I.branch[28].block[6].um_I.iw[12] ,
    \top_I.branch[28].block[6].um_I.iw[11] ,
    \top_I.branch[28].block[6].um_I.iw[10] ,
    \top_I.branch[28].block[6].um_I.iw[9] ,
    \top_I.branch[28].block[6].um_I.iw[8] ,
    \top_I.branch[28].block[6].um_I.iw[7] ,
    \top_I.branch[28].block[6].um_I.iw[6] ,
    \top_I.branch[28].block[6].um_I.iw[5] ,
    \top_I.branch[28].block[6].um_I.iw[4] ,
    \top_I.branch[28].block[6].um_I.iw[3] ,
    \top_I.branch[28].block[6].um_I.iw[2] ,
    \top_I.branch[28].block[6].um_I.iw[1] ,
    \top_I.branch[28].block[6].um_I.clk ,
    \top_I.branch[28].block[5].um_I.iw[17] ,
    \top_I.branch[28].block[5].um_I.iw[16] ,
    \top_I.branch[28].block[5].um_I.iw[15] ,
    \top_I.branch[28].block[5].um_I.iw[14] ,
    \top_I.branch[28].block[5].um_I.iw[13] ,
    \top_I.branch[28].block[5].um_I.iw[12] ,
    \top_I.branch[28].block[5].um_I.iw[11] ,
    \top_I.branch[28].block[5].um_I.iw[10] ,
    \top_I.branch[28].block[5].um_I.iw[9] ,
    \top_I.branch[28].block[5].um_I.iw[8] ,
    \top_I.branch[28].block[5].um_I.iw[7] ,
    \top_I.branch[28].block[5].um_I.iw[6] ,
    \top_I.branch[28].block[5].um_I.iw[5] ,
    \top_I.branch[28].block[5].um_I.iw[4] ,
    \top_I.branch[28].block[5].um_I.iw[3] ,
    \top_I.branch[28].block[5].um_I.iw[2] ,
    \top_I.branch[28].block[5].um_I.iw[1] ,
    \top_I.branch[28].block[5].um_I.clk ,
    \top_I.branch[28].block[4].um_I.iw[17] ,
    \top_I.branch[28].block[4].um_I.iw[16] ,
    \top_I.branch[28].block[4].um_I.iw[15] ,
    \top_I.branch[28].block[4].um_I.iw[14] ,
    \top_I.branch[28].block[4].um_I.iw[13] ,
    \top_I.branch[28].block[4].um_I.iw[12] ,
    \top_I.branch[28].block[4].um_I.iw[11] ,
    \top_I.branch[28].block[4].um_I.iw[10] ,
    \top_I.branch[28].block[4].um_I.iw[9] ,
    \top_I.branch[28].block[4].um_I.iw[8] ,
    \top_I.branch[28].block[4].um_I.iw[7] ,
    \top_I.branch[28].block[4].um_I.iw[6] ,
    \top_I.branch[28].block[4].um_I.iw[5] ,
    \top_I.branch[28].block[4].um_I.iw[4] ,
    \top_I.branch[28].block[4].um_I.iw[3] ,
    \top_I.branch[28].block[4].um_I.iw[2] ,
    \top_I.branch[28].block[4].um_I.iw[1] ,
    \top_I.branch[28].block[4].um_I.clk ,
    \top_I.branch[28].block[3].um_I.iw[17] ,
    \top_I.branch[28].block[3].um_I.iw[16] ,
    \top_I.branch[28].block[3].um_I.iw[15] ,
    \top_I.branch[28].block[3].um_I.iw[14] ,
    \top_I.branch[28].block[3].um_I.iw[13] ,
    \top_I.branch[28].block[3].um_I.iw[12] ,
    \top_I.branch[28].block[3].um_I.iw[11] ,
    \top_I.branch[28].block[3].um_I.iw[10] ,
    \top_I.branch[28].block[3].um_I.iw[9] ,
    \top_I.branch[28].block[3].um_I.iw[8] ,
    \top_I.branch[28].block[3].um_I.iw[7] ,
    \top_I.branch[28].block[3].um_I.iw[6] ,
    \top_I.branch[28].block[3].um_I.iw[5] ,
    \top_I.branch[28].block[3].um_I.iw[4] ,
    \top_I.branch[28].block[3].um_I.iw[3] ,
    \top_I.branch[28].block[3].um_I.iw[2] ,
    \top_I.branch[28].block[3].um_I.iw[1] ,
    \top_I.branch[28].block[3].um_I.clk ,
    \top_I.branch[28].block[2].um_I.iw[17] ,
    \top_I.branch[28].block[2].um_I.iw[16] ,
    \top_I.branch[28].block[2].um_I.iw[15] ,
    \top_I.branch[28].block[2].um_I.iw[14] ,
    \top_I.branch[28].block[2].um_I.iw[13] ,
    \top_I.branch[28].block[2].um_I.iw[12] ,
    \top_I.branch[28].block[2].um_I.iw[11] ,
    \top_I.branch[28].block[2].um_I.iw[10] ,
    \top_I.branch[28].block[2].um_I.iw[9] ,
    \top_I.branch[28].block[2].um_I.iw[8] ,
    \top_I.branch[28].block[2].um_I.iw[7] ,
    \top_I.branch[28].block[2].um_I.iw[6] ,
    \top_I.branch[28].block[2].um_I.iw[5] ,
    \top_I.branch[28].block[2].um_I.iw[4] ,
    \top_I.branch[28].block[2].um_I.iw[3] ,
    \top_I.branch[28].block[2].um_I.iw[2] ,
    \top_I.branch[28].block[2].um_I.iw[1] ,
    \top_I.branch[28].block[2].um_I.clk ,
    \top_I.branch[28].block[1].um_I.iw[17] ,
    \top_I.branch[28].block[1].um_I.iw[16] ,
    \top_I.branch[28].block[1].um_I.iw[15] ,
    \top_I.branch[28].block[1].um_I.iw[14] ,
    \top_I.branch[28].block[1].um_I.iw[13] ,
    \top_I.branch[28].block[1].um_I.iw[12] ,
    \top_I.branch[28].block[1].um_I.iw[11] ,
    \top_I.branch[28].block[1].um_I.iw[10] ,
    \top_I.branch[28].block[1].um_I.iw[9] ,
    \top_I.branch[28].block[1].um_I.iw[8] ,
    \top_I.branch[28].block[1].um_I.iw[7] ,
    \top_I.branch[28].block[1].um_I.iw[6] ,
    \top_I.branch[28].block[1].um_I.iw[5] ,
    \top_I.branch[28].block[1].um_I.iw[4] ,
    \top_I.branch[28].block[1].um_I.iw[3] ,
    \top_I.branch[28].block[1].um_I.iw[2] ,
    \top_I.branch[28].block[1].um_I.iw[1] ,
    \top_I.branch[28].block[1].um_I.clk ,
    \top_I.branch[28].block[0].um_I.iw[17] ,
    \top_I.branch[28].block[0].um_I.iw[16] ,
    \top_I.branch[28].block[0].um_I.iw[15] ,
    \top_I.branch[28].block[0].um_I.iw[14] ,
    \top_I.branch[28].block[0].um_I.iw[13] ,
    \top_I.branch[28].block[0].um_I.iw[12] ,
    \top_I.branch[28].block[0].um_I.iw[11] ,
    \top_I.branch[28].block[0].um_I.iw[10] ,
    \top_I.branch[28].block[0].um_I.iw[9] ,
    \top_I.branch[28].block[0].um_I.iw[8] ,
    \top_I.branch[28].block[0].um_I.iw[7] ,
    \top_I.branch[28].block[0].um_I.iw[6] ,
    \top_I.branch[28].block[0].um_I.iw[5] ,
    \top_I.branch[28].block[0].um_I.iw[4] ,
    \top_I.branch[28].block[0].um_I.iw[3] ,
    \top_I.branch[28].block[0].um_I.iw[2] ,
    \top_I.branch[28].block[0].um_I.iw[1] ,
    \top_I.branch[28].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[28].block[15].um_I.k_zero ,
    \top_I.branch[28].block[14].um_I.k_zero ,
    \top_I.branch[28].block[13].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[11].um_I.k_zero ,
    \top_I.branch[28].block[10].um_I.k_zero ,
    \top_I.branch[28].block[9].um_I.k_zero ,
    \top_I.branch[28].block[8].um_I.k_zero ,
    \top_I.branch[28].block[7].um_I.k_zero ,
    \top_I.branch[28].block[6].um_I.k_zero ,
    \top_I.branch[28].block[5].um_I.k_zero ,
    \top_I.branch[28].block[4].um_I.k_zero ,
    \top_I.branch[28].block[3].um_I.k_zero ,
    \top_I.branch[28].block[2].um_I.k_zero ,
    \top_I.branch[28].block[1].um_I.k_zero ,
    \top_I.branch[28].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[28].block[15].um_I.ow[23] ,
    \top_I.branch[28].block[15].um_I.ow[22] ,
    \top_I.branch[28].block[15].um_I.ow[21] ,
    \top_I.branch[28].block[15].um_I.ow[20] ,
    \top_I.branch[28].block[15].um_I.ow[19] ,
    \top_I.branch[28].block[15].um_I.ow[18] ,
    \top_I.branch[28].block[15].um_I.ow[17] ,
    \top_I.branch[28].block[15].um_I.ow[16] ,
    \top_I.branch[28].block[15].um_I.ow[15] ,
    \top_I.branch[28].block[15].um_I.ow[14] ,
    \top_I.branch[28].block[15].um_I.ow[13] ,
    \top_I.branch[28].block[15].um_I.ow[12] ,
    \top_I.branch[28].block[15].um_I.ow[11] ,
    \top_I.branch[28].block[15].um_I.ow[10] ,
    \top_I.branch[28].block[15].um_I.ow[9] ,
    \top_I.branch[28].block[15].um_I.ow[8] ,
    \top_I.branch[28].block[15].um_I.ow[7] ,
    \top_I.branch[28].block[15].um_I.ow[6] ,
    \top_I.branch[28].block[15].um_I.ow[5] ,
    \top_I.branch[28].block[15].um_I.ow[4] ,
    \top_I.branch[28].block[15].um_I.ow[3] ,
    \top_I.branch[28].block[15].um_I.ow[2] ,
    \top_I.branch[28].block[15].um_I.ow[1] ,
    \top_I.branch[28].block[15].um_I.ow[0] ,
    \top_I.branch[28].block[14].um_I.ow[23] ,
    \top_I.branch[28].block[14].um_I.ow[22] ,
    \top_I.branch[28].block[14].um_I.ow[21] ,
    \top_I.branch[28].block[14].um_I.ow[20] ,
    \top_I.branch[28].block[14].um_I.ow[19] ,
    \top_I.branch[28].block[14].um_I.ow[18] ,
    \top_I.branch[28].block[14].um_I.ow[17] ,
    \top_I.branch[28].block[14].um_I.ow[16] ,
    \top_I.branch[28].block[14].um_I.ow[15] ,
    \top_I.branch[28].block[14].um_I.ow[14] ,
    \top_I.branch[28].block[14].um_I.ow[13] ,
    \top_I.branch[28].block[14].um_I.ow[12] ,
    \top_I.branch[28].block[14].um_I.ow[11] ,
    \top_I.branch[28].block[14].um_I.ow[10] ,
    \top_I.branch[28].block[14].um_I.ow[9] ,
    \top_I.branch[28].block[14].um_I.ow[8] ,
    \top_I.branch[28].block[14].um_I.ow[7] ,
    \top_I.branch[28].block[14].um_I.ow[6] ,
    \top_I.branch[28].block[14].um_I.ow[5] ,
    \top_I.branch[28].block[14].um_I.ow[4] ,
    \top_I.branch[28].block[14].um_I.ow[3] ,
    \top_I.branch[28].block[14].um_I.ow[2] ,
    \top_I.branch[28].block[14].um_I.ow[1] ,
    \top_I.branch[28].block[14].um_I.ow[0] ,
    \top_I.branch[28].block[13].um_I.ow[23] ,
    \top_I.branch[28].block[13].um_I.ow[22] ,
    \top_I.branch[28].block[13].um_I.ow[21] ,
    \top_I.branch[28].block[13].um_I.ow[20] ,
    \top_I.branch[28].block[13].um_I.ow[19] ,
    \top_I.branch[28].block[13].um_I.ow[18] ,
    \top_I.branch[28].block[13].um_I.ow[17] ,
    \top_I.branch[28].block[13].um_I.ow[16] ,
    \top_I.branch[28].block[13].um_I.ow[15] ,
    \top_I.branch[28].block[13].um_I.ow[14] ,
    \top_I.branch[28].block[13].um_I.ow[13] ,
    \top_I.branch[28].block[13].um_I.ow[12] ,
    \top_I.branch[28].block[13].um_I.ow[11] ,
    \top_I.branch[28].block[13].um_I.ow[10] ,
    \top_I.branch[28].block[13].um_I.ow[9] ,
    \top_I.branch[28].block[13].um_I.ow[8] ,
    \top_I.branch[28].block[13].um_I.ow[7] ,
    \top_I.branch[28].block[13].um_I.ow[6] ,
    \top_I.branch[28].block[13].um_I.ow[5] ,
    \top_I.branch[28].block[13].um_I.ow[4] ,
    \top_I.branch[28].block[13].um_I.ow[3] ,
    \top_I.branch[28].block[13].um_I.ow[2] ,
    \top_I.branch[28].block[13].um_I.ow[1] ,
    \top_I.branch[28].block[13].um_I.ow[0] ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[12].um_I.k_zero ,
    \top_I.branch[28].block[11].um_I.ow[23] ,
    \top_I.branch[28].block[11].um_I.ow[22] ,
    \top_I.branch[28].block[11].um_I.ow[21] ,
    \top_I.branch[28].block[11].um_I.ow[20] ,
    \top_I.branch[28].block[11].um_I.ow[19] ,
    \top_I.branch[28].block[11].um_I.ow[18] ,
    \top_I.branch[28].block[11].um_I.ow[17] ,
    \top_I.branch[28].block[11].um_I.ow[16] ,
    \top_I.branch[28].block[11].um_I.ow[15] ,
    \top_I.branch[28].block[11].um_I.ow[14] ,
    \top_I.branch[28].block[11].um_I.ow[13] ,
    \top_I.branch[28].block[11].um_I.ow[12] ,
    \top_I.branch[28].block[11].um_I.ow[11] ,
    \top_I.branch[28].block[11].um_I.ow[10] ,
    \top_I.branch[28].block[11].um_I.ow[9] ,
    \top_I.branch[28].block[11].um_I.ow[8] ,
    \top_I.branch[28].block[11].um_I.ow[7] ,
    \top_I.branch[28].block[11].um_I.ow[6] ,
    \top_I.branch[28].block[11].um_I.ow[5] ,
    \top_I.branch[28].block[11].um_I.ow[4] ,
    \top_I.branch[28].block[11].um_I.ow[3] ,
    \top_I.branch[28].block[11].um_I.ow[2] ,
    \top_I.branch[28].block[11].um_I.ow[1] ,
    \top_I.branch[28].block[11].um_I.ow[0] ,
    \top_I.branch[28].block[10].um_I.ow[23] ,
    \top_I.branch[28].block[10].um_I.ow[22] ,
    \top_I.branch[28].block[10].um_I.ow[21] ,
    \top_I.branch[28].block[10].um_I.ow[20] ,
    \top_I.branch[28].block[10].um_I.ow[19] ,
    \top_I.branch[28].block[10].um_I.ow[18] ,
    \top_I.branch[28].block[10].um_I.ow[17] ,
    \top_I.branch[28].block[10].um_I.ow[16] ,
    \top_I.branch[28].block[10].um_I.ow[15] ,
    \top_I.branch[28].block[10].um_I.ow[14] ,
    \top_I.branch[28].block[10].um_I.ow[13] ,
    \top_I.branch[28].block[10].um_I.ow[12] ,
    \top_I.branch[28].block[10].um_I.ow[11] ,
    \top_I.branch[28].block[10].um_I.ow[10] ,
    \top_I.branch[28].block[10].um_I.ow[9] ,
    \top_I.branch[28].block[10].um_I.ow[8] ,
    \top_I.branch[28].block[10].um_I.ow[7] ,
    \top_I.branch[28].block[10].um_I.ow[6] ,
    \top_I.branch[28].block[10].um_I.ow[5] ,
    \top_I.branch[28].block[10].um_I.ow[4] ,
    \top_I.branch[28].block[10].um_I.ow[3] ,
    \top_I.branch[28].block[10].um_I.ow[2] ,
    \top_I.branch[28].block[10].um_I.ow[1] ,
    \top_I.branch[28].block[10].um_I.ow[0] ,
    \top_I.branch[28].block[9].um_I.ow[23] ,
    \top_I.branch[28].block[9].um_I.ow[22] ,
    \top_I.branch[28].block[9].um_I.ow[21] ,
    \top_I.branch[28].block[9].um_I.ow[20] ,
    \top_I.branch[28].block[9].um_I.ow[19] ,
    \top_I.branch[28].block[9].um_I.ow[18] ,
    \top_I.branch[28].block[9].um_I.ow[17] ,
    \top_I.branch[28].block[9].um_I.ow[16] ,
    \top_I.branch[28].block[9].um_I.ow[15] ,
    \top_I.branch[28].block[9].um_I.ow[14] ,
    \top_I.branch[28].block[9].um_I.ow[13] ,
    \top_I.branch[28].block[9].um_I.ow[12] ,
    \top_I.branch[28].block[9].um_I.ow[11] ,
    \top_I.branch[28].block[9].um_I.ow[10] ,
    \top_I.branch[28].block[9].um_I.ow[9] ,
    \top_I.branch[28].block[9].um_I.ow[8] ,
    \top_I.branch[28].block[9].um_I.ow[7] ,
    \top_I.branch[28].block[9].um_I.ow[6] ,
    \top_I.branch[28].block[9].um_I.ow[5] ,
    \top_I.branch[28].block[9].um_I.ow[4] ,
    \top_I.branch[28].block[9].um_I.ow[3] ,
    \top_I.branch[28].block[9].um_I.ow[2] ,
    \top_I.branch[28].block[9].um_I.ow[1] ,
    \top_I.branch[28].block[9].um_I.ow[0] ,
    \top_I.branch[28].block[8].um_I.ow[23] ,
    \top_I.branch[28].block[8].um_I.ow[22] ,
    \top_I.branch[28].block[8].um_I.ow[21] ,
    \top_I.branch[28].block[8].um_I.ow[20] ,
    \top_I.branch[28].block[8].um_I.ow[19] ,
    \top_I.branch[28].block[8].um_I.ow[18] ,
    \top_I.branch[28].block[8].um_I.ow[17] ,
    \top_I.branch[28].block[8].um_I.ow[16] ,
    \top_I.branch[28].block[8].um_I.ow[15] ,
    \top_I.branch[28].block[8].um_I.ow[14] ,
    \top_I.branch[28].block[8].um_I.ow[13] ,
    \top_I.branch[28].block[8].um_I.ow[12] ,
    \top_I.branch[28].block[8].um_I.ow[11] ,
    \top_I.branch[28].block[8].um_I.ow[10] ,
    \top_I.branch[28].block[8].um_I.ow[9] ,
    \top_I.branch[28].block[8].um_I.ow[8] ,
    \top_I.branch[28].block[8].um_I.ow[7] ,
    \top_I.branch[28].block[8].um_I.ow[6] ,
    \top_I.branch[28].block[8].um_I.ow[5] ,
    \top_I.branch[28].block[8].um_I.ow[4] ,
    \top_I.branch[28].block[8].um_I.ow[3] ,
    \top_I.branch[28].block[8].um_I.ow[2] ,
    \top_I.branch[28].block[8].um_I.ow[1] ,
    \top_I.branch[28].block[8].um_I.ow[0] ,
    \top_I.branch[28].block[7].um_I.ow[23] ,
    \top_I.branch[28].block[7].um_I.ow[22] ,
    \top_I.branch[28].block[7].um_I.ow[21] ,
    \top_I.branch[28].block[7].um_I.ow[20] ,
    \top_I.branch[28].block[7].um_I.ow[19] ,
    \top_I.branch[28].block[7].um_I.ow[18] ,
    \top_I.branch[28].block[7].um_I.ow[17] ,
    \top_I.branch[28].block[7].um_I.ow[16] ,
    \top_I.branch[28].block[7].um_I.ow[15] ,
    \top_I.branch[28].block[7].um_I.ow[14] ,
    \top_I.branch[28].block[7].um_I.ow[13] ,
    \top_I.branch[28].block[7].um_I.ow[12] ,
    \top_I.branch[28].block[7].um_I.ow[11] ,
    \top_I.branch[28].block[7].um_I.ow[10] ,
    \top_I.branch[28].block[7].um_I.ow[9] ,
    \top_I.branch[28].block[7].um_I.ow[8] ,
    \top_I.branch[28].block[7].um_I.ow[7] ,
    \top_I.branch[28].block[7].um_I.ow[6] ,
    \top_I.branch[28].block[7].um_I.ow[5] ,
    \top_I.branch[28].block[7].um_I.ow[4] ,
    \top_I.branch[28].block[7].um_I.ow[3] ,
    \top_I.branch[28].block[7].um_I.ow[2] ,
    \top_I.branch[28].block[7].um_I.ow[1] ,
    \top_I.branch[28].block[7].um_I.ow[0] ,
    \top_I.branch[28].block[6].um_I.ow[23] ,
    \top_I.branch[28].block[6].um_I.ow[22] ,
    \top_I.branch[28].block[6].um_I.ow[21] ,
    \top_I.branch[28].block[6].um_I.ow[20] ,
    \top_I.branch[28].block[6].um_I.ow[19] ,
    \top_I.branch[28].block[6].um_I.ow[18] ,
    \top_I.branch[28].block[6].um_I.ow[17] ,
    \top_I.branch[28].block[6].um_I.ow[16] ,
    \top_I.branch[28].block[6].um_I.ow[15] ,
    \top_I.branch[28].block[6].um_I.ow[14] ,
    \top_I.branch[28].block[6].um_I.ow[13] ,
    \top_I.branch[28].block[6].um_I.ow[12] ,
    \top_I.branch[28].block[6].um_I.ow[11] ,
    \top_I.branch[28].block[6].um_I.ow[10] ,
    \top_I.branch[28].block[6].um_I.ow[9] ,
    \top_I.branch[28].block[6].um_I.ow[8] ,
    \top_I.branch[28].block[6].um_I.ow[7] ,
    \top_I.branch[28].block[6].um_I.ow[6] ,
    \top_I.branch[28].block[6].um_I.ow[5] ,
    \top_I.branch[28].block[6].um_I.ow[4] ,
    \top_I.branch[28].block[6].um_I.ow[3] ,
    \top_I.branch[28].block[6].um_I.ow[2] ,
    \top_I.branch[28].block[6].um_I.ow[1] ,
    \top_I.branch[28].block[6].um_I.ow[0] ,
    \top_I.branch[28].block[5].um_I.ow[23] ,
    \top_I.branch[28].block[5].um_I.ow[22] ,
    \top_I.branch[28].block[5].um_I.ow[21] ,
    \top_I.branch[28].block[5].um_I.ow[20] ,
    \top_I.branch[28].block[5].um_I.ow[19] ,
    \top_I.branch[28].block[5].um_I.ow[18] ,
    \top_I.branch[28].block[5].um_I.ow[17] ,
    \top_I.branch[28].block[5].um_I.ow[16] ,
    \top_I.branch[28].block[5].um_I.ow[15] ,
    \top_I.branch[28].block[5].um_I.ow[14] ,
    \top_I.branch[28].block[5].um_I.ow[13] ,
    \top_I.branch[28].block[5].um_I.ow[12] ,
    \top_I.branch[28].block[5].um_I.ow[11] ,
    \top_I.branch[28].block[5].um_I.ow[10] ,
    \top_I.branch[28].block[5].um_I.ow[9] ,
    \top_I.branch[28].block[5].um_I.ow[8] ,
    \top_I.branch[28].block[5].um_I.ow[7] ,
    \top_I.branch[28].block[5].um_I.ow[6] ,
    \top_I.branch[28].block[5].um_I.ow[5] ,
    \top_I.branch[28].block[5].um_I.ow[4] ,
    \top_I.branch[28].block[5].um_I.ow[3] ,
    \top_I.branch[28].block[5].um_I.ow[2] ,
    \top_I.branch[28].block[5].um_I.ow[1] ,
    \top_I.branch[28].block[5].um_I.ow[0] ,
    \top_I.branch[28].block[4].um_I.ow[23] ,
    \top_I.branch[28].block[4].um_I.ow[22] ,
    \top_I.branch[28].block[4].um_I.ow[21] ,
    \top_I.branch[28].block[4].um_I.ow[20] ,
    \top_I.branch[28].block[4].um_I.ow[19] ,
    \top_I.branch[28].block[4].um_I.ow[18] ,
    \top_I.branch[28].block[4].um_I.ow[17] ,
    \top_I.branch[28].block[4].um_I.ow[16] ,
    \top_I.branch[28].block[4].um_I.ow[15] ,
    \top_I.branch[28].block[4].um_I.ow[14] ,
    \top_I.branch[28].block[4].um_I.ow[13] ,
    \top_I.branch[28].block[4].um_I.ow[12] ,
    \top_I.branch[28].block[4].um_I.ow[11] ,
    \top_I.branch[28].block[4].um_I.ow[10] ,
    \top_I.branch[28].block[4].um_I.ow[9] ,
    \top_I.branch[28].block[4].um_I.ow[8] ,
    \top_I.branch[28].block[4].um_I.ow[7] ,
    \top_I.branch[28].block[4].um_I.ow[6] ,
    \top_I.branch[28].block[4].um_I.ow[5] ,
    \top_I.branch[28].block[4].um_I.ow[4] ,
    \top_I.branch[28].block[4].um_I.ow[3] ,
    \top_I.branch[28].block[4].um_I.ow[2] ,
    \top_I.branch[28].block[4].um_I.ow[1] ,
    \top_I.branch[28].block[4].um_I.ow[0] ,
    \top_I.branch[28].block[3].um_I.ow[23] ,
    \top_I.branch[28].block[3].um_I.ow[22] ,
    \top_I.branch[28].block[3].um_I.ow[21] ,
    \top_I.branch[28].block[3].um_I.ow[20] ,
    \top_I.branch[28].block[3].um_I.ow[19] ,
    \top_I.branch[28].block[3].um_I.ow[18] ,
    \top_I.branch[28].block[3].um_I.ow[17] ,
    \top_I.branch[28].block[3].um_I.ow[16] ,
    \top_I.branch[28].block[3].um_I.ow[15] ,
    \top_I.branch[28].block[3].um_I.ow[14] ,
    \top_I.branch[28].block[3].um_I.ow[13] ,
    \top_I.branch[28].block[3].um_I.ow[12] ,
    \top_I.branch[28].block[3].um_I.ow[11] ,
    \top_I.branch[28].block[3].um_I.ow[10] ,
    \top_I.branch[28].block[3].um_I.ow[9] ,
    \top_I.branch[28].block[3].um_I.ow[8] ,
    \top_I.branch[28].block[3].um_I.ow[7] ,
    \top_I.branch[28].block[3].um_I.ow[6] ,
    \top_I.branch[28].block[3].um_I.ow[5] ,
    \top_I.branch[28].block[3].um_I.ow[4] ,
    \top_I.branch[28].block[3].um_I.ow[3] ,
    \top_I.branch[28].block[3].um_I.ow[2] ,
    \top_I.branch[28].block[3].um_I.ow[1] ,
    \top_I.branch[28].block[3].um_I.ow[0] ,
    \top_I.branch[28].block[2].um_I.ow[23] ,
    \top_I.branch[28].block[2].um_I.ow[22] ,
    \top_I.branch[28].block[2].um_I.ow[21] ,
    \top_I.branch[28].block[2].um_I.ow[20] ,
    \top_I.branch[28].block[2].um_I.ow[19] ,
    \top_I.branch[28].block[2].um_I.ow[18] ,
    \top_I.branch[28].block[2].um_I.ow[17] ,
    \top_I.branch[28].block[2].um_I.ow[16] ,
    \top_I.branch[28].block[2].um_I.ow[15] ,
    \top_I.branch[28].block[2].um_I.ow[14] ,
    \top_I.branch[28].block[2].um_I.ow[13] ,
    \top_I.branch[28].block[2].um_I.ow[12] ,
    \top_I.branch[28].block[2].um_I.ow[11] ,
    \top_I.branch[28].block[2].um_I.ow[10] ,
    \top_I.branch[28].block[2].um_I.ow[9] ,
    \top_I.branch[28].block[2].um_I.ow[8] ,
    \top_I.branch[28].block[2].um_I.ow[7] ,
    \top_I.branch[28].block[2].um_I.ow[6] ,
    \top_I.branch[28].block[2].um_I.ow[5] ,
    \top_I.branch[28].block[2].um_I.ow[4] ,
    \top_I.branch[28].block[2].um_I.ow[3] ,
    \top_I.branch[28].block[2].um_I.ow[2] ,
    \top_I.branch[28].block[2].um_I.ow[1] ,
    \top_I.branch[28].block[2].um_I.ow[0] ,
    \top_I.branch[28].block[1].um_I.ow[23] ,
    \top_I.branch[28].block[1].um_I.ow[22] ,
    \top_I.branch[28].block[1].um_I.ow[21] ,
    \top_I.branch[28].block[1].um_I.ow[20] ,
    \top_I.branch[28].block[1].um_I.ow[19] ,
    \top_I.branch[28].block[1].um_I.ow[18] ,
    \top_I.branch[28].block[1].um_I.ow[17] ,
    \top_I.branch[28].block[1].um_I.ow[16] ,
    \top_I.branch[28].block[1].um_I.ow[15] ,
    \top_I.branch[28].block[1].um_I.ow[14] ,
    \top_I.branch[28].block[1].um_I.ow[13] ,
    \top_I.branch[28].block[1].um_I.ow[12] ,
    \top_I.branch[28].block[1].um_I.ow[11] ,
    \top_I.branch[28].block[1].um_I.ow[10] ,
    \top_I.branch[28].block[1].um_I.ow[9] ,
    \top_I.branch[28].block[1].um_I.ow[8] ,
    \top_I.branch[28].block[1].um_I.ow[7] ,
    \top_I.branch[28].block[1].um_I.ow[6] ,
    \top_I.branch[28].block[1].um_I.ow[5] ,
    \top_I.branch[28].block[1].um_I.ow[4] ,
    \top_I.branch[28].block[1].um_I.ow[3] ,
    \top_I.branch[28].block[1].um_I.ow[2] ,
    \top_I.branch[28].block[1].um_I.ow[1] ,
    \top_I.branch[28].block[1].um_I.ow[0] ,
    \top_I.branch[28].block[0].um_I.ow[23] ,
    \top_I.branch[28].block[0].um_I.ow[22] ,
    \top_I.branch[28].block[0].um_I.ow[21] ,
    \top_I.branch[28].block[0].um_I.ow[20] ,
    \top_I.branch[28].block[0].um_I.ow[19] ,
    \top_I.branch[28].block[0].um_I.ow[18] ,
    \top_I.branch[28].block[0].um_I.ow[17] ,
    \top_I.branch[28].block[0].um_I.ow[16] ,
    \top_I.branch[28].block[0].um_I.ow[15] ,
    \top_I.branch[28].block[0].um_I.ow[14] ,
    \top_I.branch[28].block[0].um_I.ow[13] ,
    \top_I.branch[28].block[0].um_I.ow[12] ,
    \top_I.branch[28].block[0].um_I.ow[11] ,
    \top_I.branch[28].block[0].um_I.ow[10] ,
    \top_I.branch[28].block[0].um_I.ow[9] ,
    \top_I.branch[28].block[0].um_I.ow[8] ,
    \top_I.branch[28].block[0].um_I.ow[7] ,
    \top_I.branch[28].block[0].um_I.ow[6] ,
    \top_I.branch[28].block[0].um_I.ow[5] ,
    \top_I.branch[28].block[0].um_I.ow[4] ,
    \top_I.branch[28].block[0].um_I.ow[3] ,
    \top_I.branch[28].block[0].um_I.ow[2] ,
    \top_I.branch[28].block[0].um_I.ow[1] ,
    \top_I.branch[28].block[0].um_I.ow[0] }),
    .um_pg_vdd({\top_I.branch[28].block[15].um_I.pg_vdd ,
    \top_I.branch[28].block[14].um_I.pg_vdd ,
    \top_I.branch[28].block[13].um_I.pg_vdd ,
    \top_I.branch[28].block[12].um_I.pg_vdd ,
    \top_I.branch[28].block[11].um_I.pg_vdd ,
    \top_I.branch[28].block[10].um_I.pg_vdd ,
    \top_I.branch[28].block[9].um_I.pg_vdd ,
    \top_I.branch[28].block[8].um_I.pg_vdd ,
    \top_I.branch[28].block[7].um_I.pg_vdd ,
    \top_I.branch[28].block[6].um_I.pg_vdd ,
    \top_I.branch[28].block[5].um_I.pg_vdd ,
    \top_I.branch[28].block[4].um_I.pg_vdd ,
    \top_I.branch[28].block[3].um_I.pg_vdd ,
    \top_I.branch[28].block[2].um_I.pg_vdd ,
    \top_I.branch[28].block[1].um_I.pg_vdd ,
    \top_I.branch[28].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[29].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[29].l_addr[1] ),
    .k_zero(\top_I.branch[29].l_addr[0] ),
    .addr({\top_I.branch[29].l_addr[1] ,
    \top_I.branch[29].l_addr[1] ,
    \top_I.branch[29].l_addr[1] ,
    \top_I.branch[29].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[29].block[15].um_I.ena ,
    \top_I.branch[29].block[14].um_I.ena ,
    \top_I.branch[29].block[13].um_I.ena ,
    \top_I.branch[29].block[12].um_I.ena ,
    \top_I.branch[29].block[11].um_I.ena ,
    \top_I.branch[29].block[10].um_I.ena ,
    \top_I.branch[29].block[9].um_I.ena ,
    \top_I.branch[29].block[8].um_I.ena ,
    \top_I.branch[29].block[7].um_I.ena ,
    \top_I.branch[29].block[6].um_I.ena ,
    \top_I.branch[29].block[5].um_I.ena ,
    \top_I.branch[29].block[4].um_I.ena ,
    \top_I.branch[29].block[3].um_I.ena ,
    \top_I.branch[29].block[2].um_I.ena ,
    \top_I.branch[29].block[1].um_I.ena ,
    \top_I.branch[29].block[0].um_I.ena }),
    .um_iw({\top_I.branch[29].block[15].um_I.iw[17] ,
    \top_I.branch[29].block[15].um_I.iw[16] ,
    \top_I.branch[29].block[15].um_I.iw[15] ,
    \top_I.branch[29].block[15].um_I.iw[14] ,
    \top_I.branch[29].block[15].um_I.iw[13] ,
    \top_I.branch[29].block[15].um_I.iw[12] ,
    \top_I.branch[29].block[15].um_I.iw[11] ,
    \top_I.branch[29].block[15].um_I.iw[10] ,
    \top_I.branch[29].block[15].um_I.iw[9] ,
    \top_I.branch[29].block[15].um_I.iw[8] ,
    \top_I.branch[29].block[15].um_I.iw[7] ,
    \top_I.branch[29].block[15].um_I.iw[6] ,
    \top_I.branch[29].block[15].um_I.iw[5] ,
    \top_I.branch[29].block[15].um_I.iw[4] ,
    \top_I.branch[29].block[15].um_I.iw[3] ,
    \top_I.branch[29].block[15].um_I.iw[2] ,
    \top_I.branch[29].block[15].um_I.iw[1] ,
    \top_I.branch[29].block[15].um_I.clk ,
    \top_I.branch[29].block[14].um_I.iw[17] ,
    \top_I.branch[29].block[14].um_I.iw[16] ,
    \top_I.branch[29].block[14].um_I.iw[15] ,
    \top_I.branch[29].block[14].um_I.iw[14] ,
    \top_I.branch[29].block[14].um_I.iw[13] ,
    \top_I.branch[29].block[14].um_I.iw[12] ,
    \top_I.branch[29].block[14].um_I.iw[11] ,
    \top_I.branch[29].block[14].um_I.iw[10] ,
    \top_I.branch[29].block[14].um_I.iw[9] ,
    \top_I.branch[29].block[14].um_I.iw[8] ,
    \top_I.branch[29].block[14].um_I.iw[7] ,
    \top_I.branch[29].block[14].um_I.iw[6] ,
    \top_I.branch[29].block[14].um_I.iw[5] ,
    \top_I.branch[29].block[14].um_I.iw[4] ,
    \top_I.branch[29].block[14].um_I.iw[3] ,
    \top_I.branch[29].block[14].um_I.iw[2] ,
    \top_I.branch[29].block[14].um_I.iw[1] ,
    \top_I.branch[29].block[14].um_I.clk ,
    \top_I.branch[29].block[13].um_I.iw[17] ,
    \top_I.branch[29].block[13].um_I.iw[16] ,
    \top_I.branch[29].block[13].um_I.iw[15] ,
    \top_I.branch[29].block[13].um_I.iw[14] ,
    \top_I.branch[29].block[13].um_I.iw[13] ,
    \top_I.branch[29].block[13].um_I.iw[12] ,
    \top_I.branch[29].block[13].um_I.iw[11] ,
    \top_I.branch[29].block[13].um_I.iw[10] ,
    \top_I.branch[29].block[13].um_I.iw[9] ,
    \top_I.branch[29].block[13].um_I.iw[8] ,
    \top_I.branch[29].block[13].um_I.iw[7] ,
    \top_I.branch[29].block[13].um_I.iw[6] ,
    \top_I.branch[29].block[13].um_I.iw[5] ,
    \top_I.branch[29].block[13].um_I.iw[4] ,
    \top_I.branch[29].block[13].um_I.iw[3] ,
    \top_I.branch[29].block[13].um_I.iw[2] ,
    \top_I.branch[29].block[13].um_I.iw[1] ,
    \top_I.branch[29].block[13].um_I.clk ,
    \top_I.branch[29].block[12].um_I.iw[17] ,
    \top_I.branch[29].block[12].um_I.iw[16] ,
    \top_I.branch[29].block[12].um_I.iw[15] ,
    \top_I.branch[29].block[12].um_I.iw[14] ,
    \top_I.branch[29].block[12].um_I.iw[13] ,
    \top_I.branch[29].block[12].um_I.iw[12] ,
    \top_I.branch[29].block[12].um_I.iw[11] ,
    \top_I.branch[29].block[12].um_I.iw[10] ,
    \top_I.branch[29].block[12].um_I.iw[9] ,
    \top_I.branch[29].block[12].um_I.iw[8] ,
    \top_I.branch[29].block[12].um_I.iw[7] ,
    \top_I.branch[29].block[12].um_I.iw[6] ,
    \top_I.branch[29].block[12].um_I.iw[5] ,
    \top_I.branch[29].block[12].um_I.iw[4] ,
    \top_I.branch[29].block[12].um_I.iw[3] ,
    \top_I.branch[29].block[12].um_I.iw[2] ,
    \top_I.branch[29].block[12].um_I.iw[1] ,
    \top_I.branch[29].block[12].um_I.clk ,
    \top_I.branch[29].block[11].um_I.iw[17] ,
    \top_I.branch[29].block[11].um_I.iw[16] ,
    \top_I.branch[29].block[11].um_I.iw[15] ,
    \top_I.branch[29].block[11].um_I.iw[14] ,
    \top_I.branch[29].block[11].um_I.iw[13] ,
    \top_I.branch[29].block[11].um_I.iw[12] ,
    \top_I.branch[29].block[11].um_I.iw[11] ,
    \top_I.branch[29].block[11].um_I.iw[10] ,
    \top_I.branch[29].block[11].um_I.iw[9] ,
    \top_I.branch[29].block[11].um_I.iw[8] ,
    \top_I.branch[29].block[11].um_I.iw[7] ,
    \top_I.branch[29].block[11].um_I.iw[6] ,
    \top_I.branch[29].block[11].um_I.iw[5] ,
    \top_I.branch[29].block[11].um_I.iw[4] ,
    \top_I.branch[29].block[11].um_I.iw[3] ,
    \top_I.branch[29].block[11].um_I.iw[2] ,
    \top_I.branch[29].block[11].um_I.iw[1] ,
    \top_I.branch[29].block[11].um_I.clk ,
    \top_I.branch[29].block[10].um_I.iw[17] ,
    \top_I.branch[29].block[10].um_I.iw[16] ,
    \top_I.branch[29].block[10].um_I.iw[15] ,
    \top_I.branch[29].block[10].um_I.iw[14] ,
    \top_I.branch[29].block[10].um_I.iw[13] ,
    \top_I.branch[29].block[10].um_I.iw[12] ,
    \top_I.branch[29].block[10].um_I.iw[11] ,
    \top_I.branch[29].block[10].um_I.iw[10] ,
    \top_I.branch[29].block[10].um_I.iw[9] ,
    \top_I.branch[29].block[10].um_I.iw[8] ,
    \top_I.branch[29].block[10].um_I.iw[7] ,
    \top_I.branch[29].block[10].um_I.iw[6] ,
    \top_I.branch[29].block[10].um_I.iw[5] ,
    \top_I.branch[29].block[10].um_I.iw[4] ,
    \top_I.branch[29].block[10].um_I.iw[3] ,
    \top_I.branch[29].block[10].um_I.iw[2] ,
    \top_I.branch[29].block[10].um_I.iw[1] ,
    \top_I.branch[29].block[10].um_I.clk ,
    \top_I.branch[29].block[9].um_I.iw[17] ,
    \top_I.branch[29].block[9].um_I.iw[16] ,
    \top_I.branch[29].block[9].um_I.iw[15] ,
    \top_I.branch[29].block[9].um_I.iw[14] ,
    \top_I.branch[29].block[9].um_I.iw[13] ,
    \top_I.branch[29].block[9].um_I.iw[12] ,
    \top_I.branch[29].block[9].um_I.iw[11] ,
    \top_I.branch[29].block[9].um_I.iw[10] ,
    \top_I.branch[29].block[9].um_I.iw[9] ,
    \top_I.branch[29].block[9].um_I.iw[8] ,
    \top_I.branch[29].block[9].um_I.iw[7] ,
    \top_I.branch[29].block[9].um_I.iw[6] ,
    \top_I.branch[29].block[9].um_I.iw[5] ,
    \top_I.branch[29].block[9].um_I.iw[4] ,
    \top_I.branch[29].block[9].um_I.iw[3] ,
    \top_I.branch[29].block[9].um_I.iw[2] ,
    \top_I.branch[29].block[9].um_I.iw[1] ,
    \top_I.branch[29].block[9].um_I.clk ,
    \top_I.branch[29].block[8].um_I.iw[17] ,
    \top_I.branch[29].block[8].um_I.iw[16] ,
    \top_I.branch[29].block[8].um_I.iw[15] ,
    \top_I.branch[29].block[8].um_I.iw[14] ,
    \top_I.branch[29].block[8].um_I.iw[13] ,
    \top_I.branch[29].block[8].um_I.iw[12] ,
    \top_I.branch[29].block[8].um_I.iw[11] ,
    \top_I.branch[29].block[8].um_I.iw[10] ,
    \top_I.branch[29].block[8].um_I.iw[9] ,
    \top_I.branch[29].block[8].um_I.iw[8] ,
    \top_I.branch[29].block[8].um_I.iw[7] ,
    \top_I.branch[29].block[8].um_I.iw[6] ,
    \top_I.branch[29].block[8].um_I.iw[5] ,
    \top_I.branch[29].block[8].um_I.iw[4] ,
    \top_I.branch[29].block[8].um_I.iw[3] ,
    \top_I.branch[29].block[8].um_I.iw[2] ,
    \top_I.branch[29].block[8].um_I.iw[1] ,
    \top_I.branch[29].block[8].um_I.clk ,
    \top_I.branch[29].block[7].um_I.iw[17] ,
    \top_I.branch[29].block[7].um_I.iw[16] ,
    \top_I.branch[29].block[7].um_I.iw[15] ,
    \top_I.branch[29].block[7].um_I.iw[14] ,
    \top_I.branch[29].block[7].um_I.iw[13] ,
    \top_I.branch[29].block[7].um_I.iw[12] ,
    \top_I.branch[29].block[7].um_I.iw[11] ,
    \top_I.branch[29].block[7].um_I.iw[10] ,
    \top_I.branch[29].block[7].um_I.iw[9] ,
    \top_I.branch[29].block[7].um_I.iw[8] ,
    \top_I.branch[29].block[7].um_I.iw[7] ,
    \top_I.branch[29].block[7].um_I.iw[6] ,
    \top_I.branch[29].block[7].um_I.iw[5] ,
    \top_I.branch[29].block[7].um_I.iw[4] ,
    \top_I.branch[29].block[7].um_I.iw[3] ,
    \top_I.branch[29].block[7].um_I.iw[2] ,
    \top_I.branch[29].block[7].um_I.iw[1] ,
    \top_I.branch[29].block[7].um_I.clk ,
    \top_I.branch[29].block[6].um_I.iw[17] ,
    \top_I.branch[29].block[6].um_I.iw[16] ,
    \top_I.branch[29].block[6].um_I.iw[15] ,
    \top_I.branch[29].block[6].um_I.iw[14] ,
    \top_I.branch[29].block[6].um_I.iw[13] ,
    \top_I.branch[29].block[6].um_I.iw[12] ,
    \top_I.branch[29].block[6].um_I.iw[11] ,
    \top_I.branch[29].block[6].um_I.iw[10] ,
    \top_I.branch[29].block[6].um_I.iw[9] ,
    \top_I.branch[29].block[6].um_I.iw[8] ,
    \top_I.branch[29].block[6].um_I.iw[7] ,
    \top_I.branch[29].block[6].um_I.iw[6] ,
    \top_I.branch[29].block[6].um_I.iw[5] ,
    \top_I.branch[29].block[6].um_I.iw[4] ,
    \top_I.branch[29].block[6].um_I.iw[3] ,
    \top_I.branch[29].block[6].um_I.iw[2] ,
    \top_I.branch[29].block[6].um_I.iw[1] ,
    \top_I.branch[29].block[6].um_I.clk ,
    \top_I.branch[29].block[5].um_I.iw[17] ,
    \top_I.branch[29].block[5].um_I.iw[16] ,
    \top_I.branch[29].block[5].um_I.iw[15] ,
    \top_I.branch[29].block[5].um_I.iw[14] ,
    \top_I.branch[29].block[5].um_I.iw[13] ,
    \top_I.branch[29].block[5].um_I.iw[12] ,
    \top_I.branch[29].block[5].um_I.iw[11] ,
    \top_I.branch[29].block[5].um_I.iw[10] ,
    \top_I.branch[29].block[5].um_I.iw[9] ,
    \top_I.branch[29].block[5].um_I.iw[8] ,
    \top_I.branch[29].block[5].um_I.iw[7] ,
    \top_I.branch[29].block[5].um_I.iw[6] ,
    \top_I.branch[29].block[5].um_I.iw[5] ,
    \top_I.branch[29].block[5].um_I.iw[4] ,
    \top_I.branch[29].block[5].um_I.iw[3] ,
    \top_I.branch[29].block[5].um_I.iw[2] ,
    \top_I.branch[29].block[5].um_I.iw[1] ,
    \top_I.branch[29].block[5].um_I.clk ,
    \top_I.branch[29].block[4].um_I.iw[17] ,
    \top_I.branch[29].block[4].um_I.iw[16] ,
    \top_I.branch[29].block[4].um_I.iw[15] ,
    \top_I.branch[29].block[4].um_I.iw[14] ,
    \top_I.branch[29].block[4].um_I.iw[13] ,
    \top_I.branch[29].block[4].um_I.iw[12] ,
    \top_I.branch[29].block[4].um_I.iw[11] ,
    \top_I.branch[29].block[4].um_I.iw[10] ,
    \top_I.branch[29].block[4].um_I.iw[9] ,
    \top_I.branch[29].block[4].um_I.iw[8] ,
    \top_I.branch[29].block[4].um_I.iw[7] ,
    \top_I.branch[29].block[4].um_I.iw[6] ,
    \top_I.branch[29].block[4].um_I.iw[5] ,
    \top_I.branch[29].block[4].um_I.iw[4] ,
    \top_I.branch[29].block[4].um_I.iw[3] ,
    \top_I.branch[29].block[4].um_I.iw[2] ,
    \top_I.branch[29].block[4].um_I.iw[1] ,
    \top_I.branch[29].block[4].um_I.clk ,
    \top_I.branch[29].block[3].um_I.iw[17] ,
    \top_I.branch[29].block[3].um_I.iw[16] ,
    \top_I.branch[29].block[3].um_I.iw[15] ,
    \top_I.branch[29].block[3].um_I.iw[14] ,
    \top_I.branch[29].block[3].um_I.iw[13] ,
    \top_I.branch[29].block[3].um_I.iw[12] ,
    \top_I.branch[29].block[3].um_I.iw[11] ,
    \top_I.branch[29].block[3].um_I.iw[10] ,
    \top_I.branch[29].block[3].um_I.iw[9] ,
    \top_I.branch[29].block[3].um_I.iw[8] ,
    \top_I.branch[29].block[3].um_I.iw[7] ,
    \top_I.branch[29].block[3].um_I.iw[6] ,
    \top_I.branch[29].block[3].um_I.iw[5] ,
    \top_I.branch[29].block[3].um_I.iw[4] ,
    \top_I.branch[29].block[3].um_I.iw[3] ,
    \top_I.branch[29].block[3].um_I.iw[2] ,
    \top_I.branch[29].block[3].um_I.iw[1] ,
    \top_I.branch[29].block[3].um_I.clk ,
    \top_I.branch[29].block[2].um_I.iw[17] ,
    \top_I.branch[29].block[2].um_I.iw[16] ,
    \top_I.branch[29].block[2].um_I.iw[15] ,
    \top_I.branch[29].block[2].um_I.iw[14] ,
    \top_I.branch[29].block[2].um_I.iw[13] ,
    \top_I.branch[29].block[2].um_I.iw[12] ,
    \top_I.branch[29].block[2].um_I.iw[11] ,
    \top_I.branch[29].block[2].um_I.iw[10] ,
    \top_I.branch[29].block[2].um_I.iw[9] ,
    \top_I.branch[29].block[2].um_I.iw[8] ,
    \top_I.branch[29].block[2].um_I.iw[7] ,
    \top_I.branch[29].block[2].um_I.iw[6] ,
    \top_I.branch[29].block[2].um_I.iw[5] ,
    \top_I.branch[29].block[2].um_I.iw[4] ,
    \top_I.branch[29].block[2].um_I.iw[3] ,
    \top_I.branch[29].block[2].um_I.iw[2] ,
    \top_I.branch[29].block[2].um_I.iw[1] ,
    \top_I.branch[29].block[2].um_I.clk ,
    \top_I.branch[29].block[1].um_I.iw[17] ,
    \top_I.branch[29].block[1].um_I.iw[16] ,
    \top_I.branch[29].block[1].um_I.iw[15] ,
    \top_I.branch[29].block[1].um_I.iw[14] ,
    \top_I.branch[29].block[1].um_I.iw[13] ,
    \top_I.branch[29].block[1].um_I.iw[12] ,
    \top_I.branch[29].block[1].um_I.iw[11] ,
    \top_I.branch[29].block[1].um_I.iw[10] ,
    \top_I.branch[29].block[1].um_I.iw[9] ,
    \top_I.branch[29].block[1].um_I.iw[8] ,
    \top_I.branch[29].block[1].um_I.iw[7] ,
    \top_I.branch[29].block[1].um_I.iw[6] ,
    \top_I.branch[29].block[1].um_I.iw[5] ,
    \top_I.branch[29].block[1].um_I.iw[4] ,
    \top_I.branch[29].block[1].um_I.iw[3] ,
    \top_I.branch[29].block[1].um_I.iw[2] ,
    \top_I.branch[29].block[1].um_I.iw[1] ,
    \top_I.branch[29].block[1].um_I.clk ,
    \top_I.branch[29].block[0].um_I.iw[17] ,
    \top_I.branch[29].block[0].um_I.iw[16] ,
    \top_I.branch[29].block[0].um_I.iw[15] ,
    \top_I.branch[29].block[0].um_I.iw[14] ,
    \top_I.branch[29].block[0].um_I.iw[13] ,
    \top_I.branch[29].block[0].um_I.iw[12] ,
    \top_I.branch[29].block[0].um_I.iw[11] ,
    \top_I.branch[29].block[0].um_I.iw[10] ,
    \top_I.branch[29].block[0].um_I.iw[9] ,
    \top_I.branch[29].block[0].um_I.iw[8] ,
    \top_I.branch[29].block[0].um_I.iw[7] ,
    \top_I.branch[29].block[0].um_I.iw[6] ,
    \top_I.branch[29].block[0].um_I.iw[5] ,
    \top_I.branch[29].block[0].um_I.iw[4] ,
    \top_I.branch[29].block[0].um_I.iw[3] ,
    \top_I.branch[29].block[0].um_I.iw[2] ,
    \top_I.branch[29].block[0].um_I.iw[1] ,
    \top_I.branch[29].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[15].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[14].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[13].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[12].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[11].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[10].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[9].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[8].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[7].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[6].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[5].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[4].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[3].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[2].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[1].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero ,
    \top_I.branch[29].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[29].block[15].um_I.pg_vdd ,
    \top_I.branch[29].block[14].um_I.pg_vdd ,
    \top_I.branch[29].block[13].um_I.pg_vdd ,
    \top_I.branch[29].block[12].um_I.pg_vdd ,
    \top_I.branch[29].block[11].um_I.pg_vdd ,
    \top_I.branch[29].block[10].um_I.pg_vdd ,
    \top_I.branch[29].block[9].um_I.pg_vdd ,
    \top_I.branch[29].block[8].um_I.pg_vdd ,
    \top_I.branch[29].block[7].um_I.pg_vdd ,
    \top_I.branch[29].block[6].um_I.pg_vdd ,
    \top_I.branch[29].block[5].um_I.pg_vdd ,
    \top_I.branch[29].block[4].um_I.pg_vdd ,
    \top_I.branch[29].block[3].um_I.pg_vdd ,
    \top_I.branch[29].block[2].um_I.pg_vdd ,
    \top_I.branch[29].block[1].um_I.pg_vdd ,
    \top_I.branch[29].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[2].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[2].l_addr[0] ),
    .k_zero(\top_I.branch[2].l_addr[1] ),
    .addr({\top_I.branch[2].l_addr[1] ,
    \top_I.branch[2].l_addr[1] ,
    \top_I.branch[2].l_addr[1] ,
    \top_I.branch[2].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[2].block[15].um_I.ena ,
    \top_I.branch[2].block[14].um_I.ena ,
    \top_I.branch[2].block[13].um_I.ena ,
    \top_I.branch[2].block[12].um_I.ena ,
    \top_I.branch[2].block[11].um_I.ena ,
    \top_I.branch[2].block[10].um_I.ena ,
    \top_I.branch[2].block[9].um_I.ena ,
    \top_I.branch[2].block[8].um_I.ena ,
    \top_I.branch[2].block[7].um_I.ena ,
    \top_I.branch[2].block[6].um_I.ena ,
    \top_I.branch[2].block[5].um_I.ena ,
    \top_I.branch[2].block[4].um_I.ena ,
    \top_I.branch[2].block[3].um_I.ena ,
    \top_I.branch[2].block[2].um_I.ena ,
    \top_I.branch[2].block[1].um_I.ena ,
    \top_I.branch[2].block[0].um_I.ena }),
    .um_iw({\top_I.branch[2].block[15].um_I.iw[17] ,
    \top_I.branch[2].block[15].um_I.iw[16] ,
    \top_I.branch[2].block[15].um_I.iw[15] ,
    \top_I.branch[2].block[15].um_I.iw[14] ,
    \top_I.branch[2].block[15].um_I.iw[13] ,
    \top_I.branch[2].block[15].um_I.iw[12] ,
    \top_I.branch[2].block[15].um_I.iw[11] ,
    \top_I.branch[2].block[15].um_I.iw[10] ,
    \top_I.branch[2].block[15].um_I.iw[9] ,
    \top_I.branch[2].block[15].um_I.iw[8] ,
    \top_I.branch[2].block[15].um_I.iw[7] ,
    \top_I.branch[2].block[15].um_I.iw[6] ,
    \top_I.branch[2].block[15].um_I.iw[5] ,
    \top_I.branch[2].block[15].um_I.iw[4] ,
    \top_I.branch[2].block[15].um_I.iw[3] ,
    \top_I.branch[2].block[15].um_I.iw[2] ,
    \top_I.branch[2].block[15].um_I.iw[1] ,
    \top_I.branch[2].block[15].um_I.clk ,
    \top_I.branch[2].block[14].um_I.iw[17] ,
    \top_I.branch[2].block[14].um_I.iw[16] ,
    \top_I.branch[2].block[14].um_I.iw[15] ,
    \top_I.branch[2].block[14].um_I.iw[14] ,
    \top_I.branch[2].block[14].um_I.iw[13] ,
    \top_I.branch[2].block[14].um_I.iw[12] ,
    \top_I.branch[2].block[14].um_I.iw[11] ,
    \top_I.branch[2].block[14].um_I.iw[10] ,
    \top_I.branch[2].block[14].um_I.iw[9] ,
    \top_I.branch[2].block[14].um_I.iw[8] ,
    \top_I.branch[2].block[14].um_I.iw[7] ,
    \top_I.branch[2].block[14].um_I.iw[6] ,
    \top_I.branch[2].block[14].um_I.iw[5] ,
    \top_I.branch[2].block[14].um_I.iw[4] ,
    \top_I.branch[2].block[14].um_I.iw[3] ,
    \top_I.branch[2].block[14].um_I.iw[2] ,
    \top_I.branch[2].block[14].um_I.iw[1] ,
    \top_I.branch[2].block[14].um_I.clk ,
    \top_I.branch[2].block[13].um_I.iw[17] ,
    \top_I.branch[2].block[13].um_I.iw[16] ,
    \top_I.branch[2].block[13].um_I.iw[15] ,
    \top_I.branch[2].block[13].um_I.iw[14] ,
    \top_I.branch[2].block[13].um_I.iw[13] ,
    \top_I.branch[2].block[13].um_I.iw[12] ,
    \top_I.branch[2].block[13].um_I.iw[11] ,
    \top_I.branch[2].block[13].um_I.iw[10] ,
    \top_I.branch[2].block[13].um_I.iw[9] ,
    \top_I.branch[2].block[13].um_I.iw[8] ,
    \top_I.branch[2].block[13].um_I.iw[7] ,
    \top_I.branch[2].block[13].um_I.iw[6] ,
    \top_I.branch[2].block[13].um_I.iw[5] ,
    \top_I.branch[2].block[13].um_I.iw[4] ,
    \top_I.branch[2].block[13].um_I.iw[3] ,
    \top_I.branch[2].block[13].um_I.iw[2] ,
    \top_I.branch[2].block[13].um_I.iw[1] ,
    \top_I.branch[2].block[13].um_I.clk ,
    \top_I.branch[2].block[12].um_I.iw[17] ,
    \top_I.branch[2].block[12].um_I.iw[16] ,
    \top_I.branch[2].block[12].um_I.iw[15] ,
    \top_I.branch[2].block[12].um_I.iw[14] ,
    \top_I.branch[2].block[12].um_I.iw[13] ,
    \top_I.branch[2].block[12].um_I.iw[12] ,
    \top_I.branch[2].block[12].um_I.iw[11] ,
    \top_I.branch[2].block[12].um_I.iw[10] ,
    \top_I.branch[2].block[12].um_I.iw[9] ,
    \top_I.branch[2].block[12].um_I.iw[8] ,
    \top_I.branch[2].block[12].um_I.iw[7] ,
    \top_I.branch[2].block[12].um_I.iw[6] ,
    \top_I.branch[2].block[12].um_I.iw[5] ,
    \top_I.branch[2].block[12].um_I.iw[4] ,
    \top_I.branch[2].block[12].um_I.iw[3] ,
    \top_I.branch[2].block[12].um_I.iw[2] ,
    \top_I.branch[2].block[12].um_I.iw[1] ,
    \top_I.branch[2].block[12].um_I.clk ,
    \top_I.branch[2].block[11].um_I.iw[17] ,
    \top_I.branch[2].block[11].um_I.iw[16] ,
    \top_I.branch[2].block[11].um_I.iw[15] ,
    \top_I.branch[2].block[11].um_I.iw[14] ,
    \top_I.branch[2].block[11].um_I.iw[13] ,
    \top_I.branch[2].block[11].um_I.iw[12] ,
    \top_I.branch[2].block[11].um_I.iw[11] ,
    \top_I.branch[2].block[11].um_I.iw[10] ,
    \top_I.branch[2].block[11].um_I.iw[9] ,
    \top_I.branch[2].block[11].um_I.iw[8] ,
    \top_I.branch[2].block[11].um_I.iw[7] ,
    \top_I.branch[2].block[11].um_I.iw[6] ,
    \top_I.branch[2].block[11].um_I.iw[5] ,
    \top_I.branch[2].block[11].um_I.iw[4] ,
    \top_I.branch[2].block[11].um_I.iw[3] ,
    \top_I.branch[2].block[11].um_I.iw[2] ,
    \top_I.branch[2].block[11].um_I.iw[1] ,
    \top_I.branch[2].block[11].um_I.clk ,
    \top_I.branch[2].block[10].um_I.iw[17] ,
    \top_I.branch[2].block[10].um_I.iw[16] ,
    \top_I.branch[2].block[10].um_I.iw[15] ,
    \top_I.branch[2].block[10].um_I.iw[14] ,
    \top_I.branch[2].block[10].um_I.iw[13] ,
    \top_I.branch[2].block[10].um_I.iw[12] ,
    \top_I.branch[2].block[10].um_I.iw[11] ,
    \top_I.branch[2].block[10].um_I.iw[10] ,
    \top_I.branch[2].block[10].um_I.iw[9] ,
    \top_I.branch[2].block[10].um_I.iw[8] ,
    \top_I.branch[2].block[10].um_I.iw[7] ,
    \top_I.branch[2].block[10].um_I.iw[6] ,
    \top_I.branch[2].block[10].um_I.iw[5] ,
    \top_I.branch[2].block[10].um_I.iw[4] ,
    \top_I.branch[2].block[10].um_I.iw[3] ,
    \top_I.branch[2].block[10].um_I.iw[2] ,
    \top_I.branch[2].block[10].um_I.iw[1] ,
    \top_I.branch[2].block[10].um_I.clk ,
    \top_I.branch[2].block[9].um_I.iw[17] ,
    \top_I.branch[2].block[9].um_I.iw[16] ,
    \top_I.branch[2].block[9].um_I.iw[15] ,
    \top_I.branch[2].block[9].um_I.iw[14] ,
    \top_I.branch[2].block[9].um_I.iw[13] ,
    \top_I.branch[2].block[9].um_I.iw[12] ,
    \top_I.branch[2].block[9].um_I.iw[11] ,
    \top_I.branch[2].block[9].um_I.iw[10] ,
    \top_I.branch[2].block[9].um_I.iw[9] ,
    \top_I.branch[2].block[9].um_I.iw[8] ,
    \top_I.branch[2].block[9].um_I.iw[7] ,
    \top_I.branch[2].block[9].um_I.iw[6] ,
    \top_I.branch[2].block[9].um_I.iw[5] ,
    \top_I.branch[2].block[9].um_I.iw[4] ,
    \top_I.branch[2].block[9].um_I.iw[3] ,
    \top_I.branch[2].block[9].um_I.iw[2] ,
    \top_I.branch[2].block[9].um_I.iw[1] ,
    \top_I.branch[2].block[9].um_I.clk ,
    \top_I.branch[2].block[8].um_I.iw[17] ,
    \top_I.branch[2].block[8].um_I.iw[16] ,
    \top_I.branch[2].block[8].um_I.iw[15] ,
    \top_I.branch[2].block[8].um_I.iw[14] ,
    \top_I.branch[2].block[8].um_I.iw[13] ,
    \top_I.branch[2].block[8].um_I.iw[12] ,
    \top_I.branch[2].block[8].um_I.iw[11] ,
    \top_I.branch[2].block[8].um_I.iw[10] ,
    \top_I.branch[2].block[8].um_I.iw[9] ,
    \top_I.branch[2].block[8].um_I.iw[8] ,
    \top_I.branch[2].block[8].um_I.iw[7] ,
    \top_I.branch[2].block[8].um_I.iw[6] ,
    \top_I.branch[2].block[8].um_I.iw[5] ,
    \top_I.branch[2].block[8].um_I.iw[4] ,
    \top_I.branch[2].block[8].um_I.iw[3] ,
    \top_I.branch[2].block[8].um_I.iw[2] ,
    \top_I.branch[2].block[8].um_I.iw[1] ,
    \top_I.branch[2].block[8].um_I.clk ,
    \top_I.branch[2].block[7].um_I.iw[17] ,
    \top_I.branch[2].block[7].um_I.iw[16] ,
    \top_I.branch[2].block[7].um_I.iw[15] ,
    \top_I.branch[2].block[7].um_I.iw[14] ,
    \top_I.branch[2].block[7].um_I.iw[13] ,
    \top_I.branch[2].block[7].um_I.iw[12] ,
    \top_I.branch[2].block[7].um_I.iw[11] ,
    \top_I.branch[2].block[7].um_I.iw[10] ,
    \top_I.branch[2].block[7].um_I.iw[9] ,
    \top_I.branch[2].block[7].um_I.iw[8] ,
    \top_I.branch[2].block[7].um_I.iw[7] ,
    \top_I.branch[2].block[7].um_I.iw[6] ,
    \top_I.branch[2].block[7].um_I.iw[5] ,
    \top_I.branch[2].block[7].um_I.iw[4] ,
    \top_I.branch[2].block[7].um_I.iw[3] ,
    \top_I.branch[2].block[7].um_I.iw[2] ,
    \top_I.branch[2].block[7].um_I.iw[1] ,
    \top_I.branch[2].block[7].um_I.clk ,
    \top_I.branch[2].block[6].um_I.iw[17] ,
    \top_I.branch[2].block[6].um_I.iw[16] ,
    \top_I.branch[2].block[6].um_I.iw[15] ,
    \top_I.branch[2].block[6].um_I.iw[14] ,
    \top_I.branch[2].block[6].um_I.iw[13] ,
    \top_I.branch[2].block[6].um_I.iw[12] ,
    \top_I.branch[2].block[6].um_I.iw[11] ,
    \top_I.branch[2].block[6].um_I.iw[10] ,
    \top_I.branch[2].block[6].um_I.iw[9] ,
    \top_I.branch[2].block[6].um_I.iw[8] ,
    \top_I.branch[2].block[6].um_I.iw[7] ,
    \top_I.branch[2].block[6].um_I.iw[6] ,
    \top_I.branch[2].block[6].um_I.iw[5] ,
    \top_I.branch[2].block[6].um_I.iw[4] ,
    \top_I.branch[2].block[6].um_I.iw[3] ,
    \top_I.branch[2].block[6].um_I.iw[2] ,
    \top_I.branch[2].block[6].um_I.iw[1] ,
    \top_I.branch[2].block[6].um_I.clk ,
    \top_I.branch[2].block[5].um_I.iw[17] ,
    \top_I.branch[2].block[5].um_I.iw[16] ,
    \top_I.branch[2].block[5].um_I.iw[15] ,
    \top_I.branch[2].block[5].um_I.iw[14] ,
    \top_I.branch[2].block[5].um_I.iw[13] ,
    \top_I.branch[2].block[5].um_I.iw[12] ,
    \top_I.branch[2].block[5].um_I.iw[11] ,
    \top_I.branch[2].block[5].um_I.iw[10] ,
    \top_I.branch[2].block[5].um_I.iw[9] ,
    \top_I.branch[2].block[5].um_I.iw[8] ,
    \top_I.branch[2].block[5].um_I.iw[7] ,
    \top_I.branch[2].block[5].um_I.iw[6] ,
    \top_I.branch[2].block[5].um_I.iw[5] ,
    \top_I.branch[2].block[5].um_I.iw[4] ,
    \top_I.branch[2].block[5].um_I.iw[3] ,
    \top_I.branch[2].block[5].um_I.iw[2] ,
    \top_I.branch[2].block[5].um_I.iw[1] ,
    \top_I.branch[2].block[5].um_I.clk ,
    \top_I.branch[2].block[4].um_I.iw[17] ,
    \top_I.branch[2].block[4].um_I.iw[16] ,
    \top_I.branch[2].block[4].um_I.iw[15] ,
    \top_I.branch[2].block[4].um_I.iw[14] ,
    \top_I.branch[2].block[4].um_I.iw[13] ,
    \top_I.branch[2].block[4].um_I.iw[12] ,
    \top_I.branch[2].block[4].um_I.iw[11] ,
    \top_I.branch[2].block[4].um_I.iw[10] ,
    \top_I.branch[2].block[4].um_I.iw[9] ,
    \top_I.branch[2].block[4].um_I.iw[8] ,
    \top_I.branch[2].block[4].um_I.iw[7] ,
    \top_I.branch[2].block[4].um_I.iw[6] ,
    \top_I.branch[2].block[4].um_I.iw[5] ,
    \top_I.branch[2].block[4].um_I.iw[4] ,
    \top_I.branch[2].block[4].um_I.iw[3] ,
    \top_I.branch[2].block[4].um_I.iw[2] ,
    \top_I.branch[2].block[4].um_I.iw[1] ,
    \top_I.branch[2].block[4].um_I.clk ,
    \top_I.branch[2].block[3].um_I.iw[17] ,
    \top_I.branch[2].block[3].um_I.iw[16] ,
    \top_I.branch[2].block[3].um_I.iw[15] ,
    \top_I.branch[2].block[3].um_I.iw[14] ,
    \top_I.branch[2].block[3].um_I.iw[13] ,
    \top_I.branch[2].block[3].um_I.iw[12] ,
    \top_I.branch[2].block[3].um_I.iw[11] ,
    \top_I.branch[2].block[3].um_I.iw[10] ,
    \top_I.branch[2].block[3].um_I.iw[9] ,
    \top_I.branch[2].block[3].um_I.iw[8] ,
    \top_I.branch[2].block[3].um_I.iw[7] ,
    \top_I.branch[2].block[3].um_I.iw[6] ,
    \top_I.branch[2].block[3].um_I.iw[5] ,
    \top_I.branch[2].block[3].um_I.iw[4] ,
    \top_I.branch[2].block[3].um_I.iw[3] ,
    \top_I.branch[2].block[3].um_I.iw[2] ,
    \top_I.branch[2].block[3].um_I.iw[1] ,
    \top_I.branch[2].block[3].um_I.clk ,
    \top_I.branch[2].block[2].um_I.iw[17] ,
    \top_I.branch[2].block[2].um_I.iw[16] ,
    \top_I.branch[2].block[2].um_I.iw[15] ,
    \top_I.branch[2].block[2].um_I.iw[14] ,
    \top_I.branch[2].block[2].um_I.iw[13] ,
    \top_I.branch[2].block[2].um_I.iw[12] ,
    \top_I.branch[2].block[2].um_I.iw[11] ,
    \top_I.branch[2].block[2].um_I.iw[10] ,
    \top_I.branch[2].block[2].um_I.iw[9] ,
    \top_I.branch[2].block[2].um_I.iw[8] ,
    \top_I.branch[2].block[2].um_I.iw[7] ,
    \top_I.branch[2].block[2].um_I.iw[6] ,
    \top_I.branch[2].block[2].um_I.iw[5] ,
    \top_I.branch[2].block[2].um_I.iw[4] ,
    \top_I.branch[2].block[2].um_I.iw[3] ,
    \top_I.branch[2].block[2].um_I.iw[2] ,
    \top_I.branch[2].block[2].um_I.iw[1] ,
    \top_I.branch[2].block[2].um_I.clk ,
    \top_I.branch[2].block[1].um_I.iw[17] ,
    \top_I.branch[2].block[1].um_I.iw[16] ,
    \top_I.branch[2].block[1].um_I.iw[15] ,
    \top_I.branch[2].block[1].um_I.iw[14] ,
    \top_I.branch[2].block[1].um_I.iw[13] ,
    \top_I.branch[2].block[1].um_I.iw[12] ,
    \top_I.branch[2].block[1].um_I.iw[11] ,
    \top_I.branch[2].block[1].um_I.iw[10] ,
    \top_I.branch[2].block[1].um_I.iw[9] ,
    \top_I.branch[2].block[1].um_I.iw[8] ,
    \top_I.branch[2].block[1].um_I.iw[7] ,
    \top_I.branch[2].block[1].um_I.iw[6] ,
    \top_I.branch[2].block[1].um_I.iw[5] ,
    \top_I.branch[2].block[1].um_I.iw[4] ,
    \top_I.branch[2].block[1].um_I.iw[3] ,
    \top_I.branch[2].block[1].um_I.iw[2] ,
    \top_I.branch[2].block[1].um_I.iw[1] ,
    \top_I.branch[2].block[1].um_I.clk ,
    \top_I.branch[2].block[0].um_I.iw[17] ,
    \top_I.branch[2].block[0].um_I.iw[16] ,
    \top_I.branch[2].block[0].um_I.iw[15] ,
    \top_I.branch[2].block[0].um_I.iw[14] ,
    \top_I.branch[2].block[0].um_I.iw[13] ,
    \top_I.branch[2].block[0].um_I.iw[12] ,
    \top_I.branch[2].block[0].um_I.iw[11] ,
    \top_I.branch[2].block[0].um_I.iw[10] ,
    \top_I.branch[2].block[0].um_I.iw[9] ,
    \top_I.branch[2].block[0].um_I.iw[8] ,
    \top_I.branch[2].block[0].um_I.iw[7] ,
    \top_I.branch[2].block[0].um_I.iw[6] ,
    \top_I.branch[2].block[0].um_I.iw[5] ,
    \top_I.branch[2].block[0].um_I.iw[4] ,
    \top_I.branch[2].block[0].um_I.iw[3] ,
    \top_I.branch[2].block[0].um_I.iw[2] ,
    \top_I.branch[2].block[0].um_I.iw[1] ,
    \top_I.branch[2].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[15].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[14].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[13].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[12].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[11].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[10].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[9].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[8].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[7].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[6].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[5].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[4].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[3].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[2].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[1].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero ,
    \top_I.branch[2].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[2].block[15].um_I.pg_vdd ,
    \top_I.branch[2].block[14].um_I.pg_vdd ,
    \top_I.branch[2].block[13].um_I.pg_vdd ,
    \top_I.branch[2].block[12].um_I.pg_vdd ,
    \top_I.branch[2].block[11].um_I.pg_vdd ,
    \top_I.branch[2].block[10].um_I.pg_vdd ,
    \top_I.branch[2].block[9].um_I.pg_vdd ,
    \top_I.branch[2].block[8].um_I.pg_vdd ,
    \top_I.branch[2].block[7].um_I.pg_vdd ,
    \top_I.branch[2].block[6].um_I.pg_vdd ,
    \top_I.branch[2].block[5].um_I.pg_vdd ,
    \top_I.branch[2].block[4].um_I.pg_vdd ,
    \top_I.branch[2].block[3].um_I.pg_vdd ,
    \top_I.branch[2].block[2].um_I.pg_vdd ,
    \top_I.branch[2].block[1].um_I.pg_vdd ,
    \top_I.branch[2].block[0].um_I.pg_vdd }));
 tt_pg_vdd_1 \top_I.branch[30].block[0].um_I.block_30_0.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[0].um_I.block_30_0.vpwr ),
    .ctrl(\top_I.branch[30].block[0].um_I.pg_vdd ));
 tt_um_mattvenn_rgb_mixer \top_I.branch[30].block[0].um_I.block_30_0.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[0].um_I.block_30_0.vpwr ),
    .clk(\top_I.branch[30].block[0].um_I.clk ),
    .ena(\top_I.branch[30].block[0].um_I.ena ),
    .rst_n(\top_I.branch[30].block[0].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[0].um_I.iw[9] ,
    \top_I.branch[30].block[0].um_I.iw[8] ,
    \top_I.branch[30].block[0].um_I.iw[7] ,
    \top_I.branch[30].block[0].um_I.iw[6] ,
    \top_I.branch[30].block[0].um_I.iw[5] ,
    \top_I.branch[30].block[0].um_I.iw[4] ,
    \top_I.branch[30].block[0].um_I.iw[3] ,
    \top_I.branch[30].block[0].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[0].um_I.iw[17] ,
    \top_I.branch[30].block[0].um_I.iw[16] ,
    \top_I.branch[30].block[0].um_I.iw[15] ,
    \top_I.branch[30].block[0].um_I.iw[14] ,
    \top_I.branch[30].block[0].um_I.iw[13] ,
    \top_I.branch[30].block[0].um_I.iw[12] ,
    \top_I.branch[30].block[0].um_I.iw[11] ,
    \top_I.branch[30].block[0].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[0].um_I.ow[23] ,
    \top_I.branch[30].block[0].um_I.ow[22] ,
    \top_I.branch[30].block[0].um_I.ow[21] ,
    \top_I.branch[30].block[0].um_I.ow[20] ,
    \top_I.branch[30].block[0].um_I.ow[19] ,
    \top_I.branch[30].block[0].um_I.ow[18] ,
    \top_I.branch[30].block[0].um_I.ow[17] ,
    \top_I.branch[30].block[0].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[0].um_I.ow[15] ,
    \top_I.branch[30].block[0].um_I.ow[14] ,
    \top_I.branch[30].block[0].um_I.ow[13] ,
    \top_I.branch[30].block[0].um_I.ow[12] ,
    \top_I.branch[30].block[0].um_I.ow[11] ,
    \top_I.branch[30].block[0].um_I.ow[10] ,
    \top_I.branch[30].block[0].um_I.ow[9] ,
    \top_I.branch[30].block[0].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[0].um_I.ow[7] ,
    \top_I.branch[30].block[0].um_I.ow[6] ,
    \top_I.branch[30].block[0].um_I.ow[5] ,
    \top_I.branch[30].block[0].um_I.ow[4] ,
    \top_I.branch[30].block[0].um_I.ow[3] ,
    \top_I.branch[30].block[0].um_I.ow[2] ,
    \top_I.branch[30].block[0].um_I.ow[1] ,
    \top_I.branch[30].block[0].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[11].um_I.block_30_11.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[11].um_I.block_30_11.vpwr ),
    .ctrl(\top_I.branch[30].block[11].um_I.pg_vdd ));
 tt_um_ps2_morse_encoder_top \top_I.branch[30].block[11].um_I.block_30_11.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[11].um_I.block_30_11.vpwr ),
    .clk(\top_I.branch[30].block[11].um_I.clk ),
    .ena(\top_I.branch[30].block[11].um_I.ena ),
    .rst_n(\top_I.branch[30].block[11].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[11].um_I.iw[9] ,
    \top_I.branch[30].block[11].um_I.iw[8] ,
    \top_I.branch[30].block[11].um_I.iw[7] ,
    \top_I.branch[30].block[11].um_I.iw[6] ,
    \top_I.branch[30].block[11].um_I.iw[5] ,
    \top_I.branch[30].block[11].um_I.iw[4] ,
    \top_I.branch[30].block[11].um_I.iw[3] ,
    \top_I.branch[30].block[11].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[11].um_I.iw[17] ,
    \top_I.branch[30].block[11].um_I.iw[16] ,
    \top_I.branch[30].block[11].um_I.iw[15] ,
    \top_I.branch[30].block[11].um_I.iw[14] ,
    \top_I.branch[30].block[11].um_I.iw[13] ,
    \top_I.branch[30].block[11].um_I.iw[12] ,
    \top_I.branch[30].block[11].um_I.iw[11] ,
    \top_I.branch[30].block[11].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[11].um_I.ow[23] ,
    \top_I.branch[30].block[11].um_I.ow[22] ,
    \top_I.branch[30].block[11].um_I.ow[21] ,
    \top_I.branch[30].block[11].um_I.ow[20] ,
    \top_I.branch[30].block[11].um_I.ow[19] ,
    \top_I.branch[30].block[11].um_I.ow[18] ,
    \top_I.branch[30].block[11].um_I.ow[17] ,
    \top_I.branch[30].block[11].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[11].um_I.ow[15] ,
    \top_I.branch[30].block[11].um_I.ow[14] ,
    \top_I.branch[30].block[11].um_I.ow[13] ,
    \top_I.branch[30].block[11].um_I.ow[12] ,
    \top_I.branch[30].block[11].um_I.ow[11] ,
    \top_I.branch[30].block[11].um_I.ow[10] ,
    \top_I.branch[30].block[11].um_I.ow[9] ,
    \top_I.branch[30].block[11].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[11].um_I.ow[7] ,
    \top_I.branch[30].block[11].um_I.ow[6] ,
    \top_I.branch[30].block[11].um_I.ow[5] ,
    \top_I.branch[30].block[11].um_I.ow[4] ,
    \top_I.branch[30].block[11].um_I.ow[3] ,
    \top_I.branch[30].block[11].um_I.ow[2] ,
    \top_I.branch[30].block[11].um_I.ow[1] ,
    \top_I.branch[30].block[11].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[13].um_I.block_30_13.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[13].um_I.block_30_13.vpwr ),
    .ctrl(\top_I.branch[30].block[13].um_I.pg_vdd ));
 tt_um_calculator_muehlbb \top_I.branch[30].block[13].um_I.block_30_13.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[13].um_I.block_30_13.vpwr ),
    .clk(\top_I.branch[30].block[13].um_I.clk ),
    .ena(\top_I.branch[30].block[13].um_I.ena ),
    .rst_n(\top_I.branch[30].block[13].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[13].um_I.iw[9] ,
    \top_I.branch[30].block[13].um_I.iw[8] ,
    \top_I.branch[30].block[13].um_I.iw[7] ,
    \top_I.branch[30].block[13].um_I.iw[6] ,
    \top_I.branch[30].block[13].um_I.iw[5] ,
    \top_I.branch[30].block[13].um_I.iw[4] ,
    \top_I.branch[30].block[13].um_I.iw[3] ,
    \top_I.branch[30].block[13].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[13].um_I.iw[17] ,
    \top_I.branch[30].block[13].um_I.iw[16] ,
    \top_I.branch[30].block[13].um_I.iw[15] ,
    \top_I.branch[30].block[13].um_I.iw[14] ,
    \top_I.branch[30].block[13].um_I.iw[13] ,
    \top_I.branch[30].block[13].um_I.iw[12] ,
    \top_I.branch[30].block[13].um_I.iw[11] ,
    \top_I.branch[30].block[13].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[13].um_I.ow[23] ,
    \top_I.branch[30].block[13].um_I.ow[22] ,
    \top_I.branch[30].block[13].um_I.ow[21] ,
    \top_I.branch[30].block[13].um_I.ow[20] ,
    \top_I.branch[30].block[13].um_I.ow[19] ,
    \top_I.branch[30].block[13].um_I.ow[18] ,
    \top_I.branch[30].block[13].um_I.ow[17] ,
    \top_I.branch[30].block[13].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[13].um_I.ow[15] ,
    \top_I.branch[30].block[13].um_I.ow[14] ,
    \top_I.branch[30].block[13].um_I.ow[13] ,
    \top_I.branch[30].block[13].um_I.ow[12] ,
    \top_I.branch[30].block[13].um_I.ow[11] ,
    \top_I.branch[30].block[13].um_I.ow[10] ,
    \top_I.branch[30].block[13].um_I.ow[9] ,
    \top_I.branch[30].block[13].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[13].um_I.ow[7] ,
    \top_I.branch[30].block[13].um_I.ow[6] ,
    \top_I.branch[30].block[13].um_I.ow[5] ,
    \top_I.branch[30].block[13].um_I.ow[4] ,
    \top_I.branch[30].block[13].um_I.ow[3] ,
    \top_I.branch[30].block[13].um_I.ow[2] ,
    \top_I.branch[30].block[13].um_I.ow[1] ,
    \top_I.branch[30].block[13].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[15].um_I.block_30_15.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[15].um_I.block_30_15.vpwr ),
    .ctrl(\top_I.branch[30].block[15].um_I.pg_vdd ));
 tt_um_hpretl_tt06_tempsens \top_I.branch[30].block[15].um_I.block_30_15.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[15].um_I.block_30_15.vpwr ),
    .clk(\top_I.branch[30].block[15].um_I.clk ),
    .ena(\top_I.branch[30].block[15].um_I.ena ),
    .rst_n(\top_I.branch[30].block[15].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[15].um_I.iw[9] ,
    \top_I.branch[30].block[15].um_I.iw[8] ,
    \top_I.branch[30].block[15].um_I.iw[7] ,
    \top_I.branch[30].block[15].um_I.iw[6] ,
    \top_I.branch[30].block[15].um_I.iw[5] ,
    \top_I.branch[30].block[15].um_I.iw[4] ,
    \top_I.branch[30].block[15].um_I.iw[3] ,
    \top_I.branch[30].block[15].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[15].um_I.iw[17] ,
    \top_I.branch[30].block[15].um_I.iw[16] ,
    \top_I.branch[30].block[15].um_I.iw[15] ,
    \top_I.branch[30].block[15].um_I.iw[14] ,
    \top_I.branch[30].block[15].um_I.iw[13] ,
    \top_I.branch[30].block[15].um_I.iw[12] ,
    \top_I.branch[30].block[15].um_I.iw[11] ,
    \top_I.branch[30].block[15].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[15].um_I.ow[23] ,
    \top_I.branch[30].block[15].um_I.ow[22] ,
    \top_I.branch[30].block[15].um_I.ow[21] ,
    \top_I.branch[30].block[15].um_I.ow[20] ,
    \top_I.branch[30].block[15].um_I.ow[19] ,
    \top_I.branch[30].block[15].um_I.ow[18] ,
    \top_I.branch[30].block[15].um_I.ow[17] ,
    \top_I.branch[30].block[15].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[15].um_I.ow[15] ,
    \top_I.branch[30].block[15].um_I.ow[14] ,
    \top_I.branch[30].block[15].um_I.ow[13] ,
    \top_I.branch[30].block[15].um_I.ow[12] ,
    \top_I.branch[30].block[15].um_I.ow[11] ,
    \top_I.branch[30].block[15].um_I.ow[10] ,
    \top_I.branch[30].block[15].um_I.ow[9] ,
    \top_I.branch[30].block[15].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[15].um_I.ow[7] ,
    \top_I.branch[30].block[15].um_I.ow[6] ,
    \top_I.branch[30].block[15].um_I.ow[5] ,
    \top_I.branch[30].block[15].um_I.ow[4] ,
    \top_I.branch[30].block[15].um_I.ow[3] ,
    \top_I.branch[30].block[15].um_I.ow[2] ,
    \top_I.branch[30].block[15].um_I.ow[1] ,
    \top_I.branch[30].block[15].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[1].um_I.block_30_1.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[1].um_I.block_30_1.vpwr ),
    .ctrl(\top_I.branch[30].block[1].um_I.pg_vdd ));
 tt_um_ledcontroller_Gatsch \top_I.branch[30].block[1].um_I.block_30_1.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[1].um_I.block_30_1.vpwr ),
    .clk(\top_I.branch[30].block[1].um_I.clk ),
    .ena(\top_I.branch[30].block[1].um_I.ena ),
    .rst_n(\top_I.branch[30].block[1].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[1].um_I.iw[9] ,
    \top_I.branch[30].block[1].um_I.iw[8] ,
    \top_I.branch[30].block[1].um_I.iw[7] ,
    \top_I.branch[30].block[1].um_I.iw[6] ,
    \top_I.branch[30].block[1].um_I.iw[5] ,
    \top_I.branch[30].block[1].um_I.iw[4] ,
    \top_I.branch[30].block[1].um_I.iw[3] ,
    \top_I.branch[30].block[1].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[1].um_I.iw[17] ,
    \top_I.branch[30].block[1].um_I.iw[16] ,
    \top_I.branch[30].block[1].um_I.iw[15] ,
    \top_I.branch[30].block[1].um_I.iw[14] ,
    \top_I.branch[30].block[1].um_I.iw[13] ,
    \top_I.branch[30].block[1].um_I.iw[12] ,
    \top_I.branch[30].block[1].um_I.iw[11] ,
    \top_I.branch[30].block[1].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[1].um_I.ow[23] ,
    \top_I.branch[30].block[1].um_I.ow[22] ,
    \top_I.branch[30].block[1].um_I.ow[21] ,
    \top_I.branch[30].block[1].um_I.ow[20] ,
    \top_I.branch[30].block[1].um_I.ow[19] ,
    \top_I.branch[30].block[1].um_I.ow[18] ,
    \top_I.branch[30].block[1].um_I.ow[17] ,
    \top_I.branch[30].block[1].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[1].um_I.ow[15] ,
    \top_I.branch[30].block[1].um_I.ow[14] ,
    \top_I.branch[30].block[1].um_I.ow[13] ,
    \top_I.branch[30].block[1].um_I.ow[12] ,
    \top_I.branch[30].block[1].um_I.ow[11] ,
    \top_I.branch[30].block[1].um_I.ow[10] ,
    \top_I.branch[30].block[1].um_I.ow[9] ,
    \top_I.branch[30].block[1].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[1].um_I.ow[7] ,
    \top_I.branch[30].block[1].um_I.ow[6] ,
    \top_I.branch[30].block[1].um_I.ow[5] ,
    \top_I.branch[30].block[1].um_I.ow[4] ,
    \top_I.branch[30].block[1].um_I.ow[3] ,
    \top_I.branch[30].block[1].um_I.ow[2] ,
    \top_I.branch[30].block[1].um_I.ow[1] ,
    \top_I.branch[30].block[1].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[2].um_I.block_30_2.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[2].um_I.block_30_2.vpwr ),
    .ctrl(\top_I.branch[30].block[2].um_I.pg_vdd ));
 tt_um_entwurf_integrierter_schaltungen_hadner \top_I.branch[30].block[2].um_I.block_30_2.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[2].um_I.block_30_2.vpwr ),
    .clk(\top_I.branch[30].block[2].um_I.clk ),
    .ena(\top_I.branch[30].block[2].um_I.ena ),
    .rst_n(\top_I.branch[30].block[2].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[2].um_I.iw[9] ,
    \top_I.branch[30].block[2].um_I.iw[8] ,
    \top_I.branch[30].block[2].um_I.iw[7] ,
    \top_I.branch[30].block[2].um_I.iw[6] ,
    \top_I.branch[30].block[2].um_I.iw[5] ,
    \top_I.branch[30].block[2].um_I.iw[4] ,
    \top_I.branch[30].block[2].um_I.iw[3] ,
    \top_I.branch[30].block[2].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[2].um_I.iw[17] ,
    \top_I.branch[30].block[2].um_I.iw[16] ,
    \top_I.branch[30].block[2].um_I.iw[15] ,
    \top_I.branch[30].block[2].um_I.iw[14] ,
    \top_I.branch[30].block[2].um_I.iw[13] ,
    \top_I.branch[30].block[2].um_I.iw[12] ,
    \top_I.branch[30].block[2].um_I.iw[11] ,
    \top_I.branch[30].block[2].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[2].um_I.ow[23] ,
    \top_I.branch[30].block[2].um_I.ow[22] ,
    \top_I.branch[30].block[2].um_I.ow[21] ,
    \top_I.branch[30].block[2].um_I.ow[20] ,
    \top_I.branch[30].block[2].um_I.ow[19] ,
    \top_I.branch[30].block[2].um_I.ow[18] ,
    \top_I.branch[30].block[2].um_I.ow[17] ,
    \top_I.branch[30].block[2].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[2].um_I.ow[15] ,
    \top_I.branch[30].block[2].um_I.ow[14] ,
    \top_I.branch[30].block[2].um_I.ow[13] ,
    \top_I.branch[30].block[2].um_I.ow[12] ,
    \top_I.branch[30].block[2].um_I.ow[11] ,
    \top_I.branch[30].block[2].um_I.ow[10] ,
    \top_I.branch[30].block[2].um_I.ow[9] ,
    \top_I.branch[30].block[2].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[2].um_I.ow[7] ,
    \top_I.branch[30].block[2].um_I.ow[6] ,
    \top_I.branch[30].block[2].um_I.ow[5] ,
    \top_I.branch[30].block[2].um_I.ow[4] ,
    \top_I.branch[30].block[2].um_I.ow[3] ,
    \top_I.branch[30].block[2].um_I.ow[2] ,
    \top_I.branch[30].block[2].um_I.ow[1] ,
    \top_I.branch[30].block[2].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[3].um_I.block_30_3.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[3].um_I.block_30_3.vpwr ),
    .ctrl(\top_I.branch[30].block[3].um_I.pg_vdd ));
 tt_um_digitaler_filter_rathmayr \top_I.branch[30].block[3].um_I.block_30_3.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[3].um_I.block_30_3.vpwr ),
    .clk(\top_I.branch[30].block[3].um_I.clk ),
    .ena(\top_I.branch[30].block[3].um_I.ena ),
    .rst_n(\top_I.branch[30].block[3].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[3].um_I.iw[9] ,
    \top_I.branch[30].block[3].um_I.iw[8] ,
    \top_I.branch[30].block[3].um_I.iw[7] ,
    \top_I.branch[30].block[3].um_I.iw[6] ,
    \top_I.branch[30].block[3].um_I.iw[5] ,
    \top_I.branch[30].block[3].um_I.iw[4] ,
    \top_I.branch[30].block[3].um_I.iw[3] ,
    \top_I.branch[30].block[3].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[3].um_I.iw[17] ,
    \top_I.branch[30].block[3].um_I.iw[16] ,
    \top_I.branch[30].block[3].um_I.iw[15] ,
    \top_I.branch[30].block[3].um_I.iw[14] ,
    \top_I.branch[30].block[3].um_I.iw[13] ,
    \top_I.branch[30].block[3].um_I.iw[12] ,
    \top_I.branch[30].block[3].um_I.iw[11] ,
    \top_I.branch[30].block[3].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[3].um_I.ow[23] ,
    \top_I.branch[30].block[3].um_I.ow[22] ,
    \top_I.branch[30].block[3].um_I.ow[21] ,
    \top_I.branch[30].block[3].um_I.ow[20] ,
    \top_I.branch[30].block[3].um_I.ow[19] ,
    \top_I.branch[30].block[3].um_I.ow[18] ,
    \top_I.branch[30].block[3].um_I.ow[17] ,
    \top_I.branch[30].block[3].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[3].um_I.ow[15] ,
    \top_I.branch[30].block[3].um_I.ow[14] ,
    \top_I.branch[30].block[3].um_I.ow[13] ,
    \top_I.branch[30].block[3].um_I.ow[12] ,
    \top_I.branch[30].block[3].um_I.ow[11] ,
    \top_I.branch[30].block[3].um_I.ow[10] ,
    \top_I.branch[30].block[3].um_I.ow[9] ,
    \top_I.branch[30].block[3].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[3].um_I.ow[7] ,
    \top_I.branch[30].block[3].um_I.ow[6] ,
    \top_I.branch[30].block[3].um_I.ow[5] ,
    \top_I.branch[30].block[3].um_I.ow[4] ,
    \top_I.branch[30].block[3].um_I.ow[3] ,
    \top_I.branch[30].block[3].um_I.ow[2] ,
    \top_I.branch[30].block[3].um_I.ow[1] ,
    \top_I.branch[30].block[3].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[4].um_I.block_30_4.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[4].um_I.block_30_4.vpwr ),
    .ctrl(\top_I.branch[30].block[4].um_I.pg_vdd ));
 tt_um_seven_segment_fun1 \top_I.branch[30].block[4].um_I.block_30_4.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[4].um_I.block_30_4.vpwr ),
    .clk(\top_I.branch[30].block[4].um_I.clk ),
    .ena(\top_I.branch[30].block[4].um_I.ena ),
    .rst_n(\top_I.branch[30].block[4].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[4].um_I.iw[9] ,
    \top_I.branch[30].block[4].um_I.iw[8] ,
    \top_I.branch[30].block[4].um_I.iw[7] ,
    \top_I.branch[30].block[4].um_I.iw[6] ,
    \top_I.branch[30].block[4].um_I.iw[5] ,
    \top_I.branch[30].block[4].um_I.iw[4] ,
    \top_I.branch[30].block[4].um_I.iw[3] ,
    \top_I.branch[30].block[4].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[4].um_I.iw[17] ,
    \top_I.branch[30].block[4].um_I.iw[16] ,
    \top_I.branch[30].block[4].um_I.iw[15] ,
    \top_I.branch[30].block[4].um_I.iw[14] ,
    \top_I.branch[30].block[4].um_I.iw[13] ,
    \top_I.branch[30].block[4].um_I.iw[12] ,
    \top_I.branch[30].block[4].um_I.iw[11] ,
    \top_I.branch[30].block[4].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[4].um_I.ow[23] ,
    \top_I.branch[30].block[4].um_I.ow[22] ,
    \top_I.branch[30].block[4].um_I.ow[21] ,
    \top_I.branch[30].block[4].um_I.ow[20] ,
    \top_I.branch[30].block[4].um_I.ow[19] ,
    \top_I.branch[30].block[4].um_I.ow[18] ,
    \top_I.branch[30].block[4].um_I.ow[17] ,
    \top_I.branch[30].block[4].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[4].um_I.ow[15] ,
    \top_I.branch[30].block[4].um_I.ow[14] ,
    \top_I.branch[30].block[4].um_I.ow[13] ,
    \top_I.branch[30].block[4].um_I.ow[12] ,
    \top_I.branch[30].block[4].um_I.ow[11] ,
    \top_I.branch[30].block[4].um_I.ow[10] ,
    \top_I.branch[30].block[4].um_I.ow[9] ,
    \top_I.branch[30].block[4].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[4].um_I.ow[7] ,
    \top_I.branch[30].block[4].um_I.ow[6] ,
    \top_I.branch[30].block[4].um_I.ow[5] ,
    \top_I.branch[30].block[4].um_I.ow[4] ,
    \top_I.branch[30].block[4].um_I.ow[3] ,
    \top_I.branch[30].block[4].um_I.ow[2] ,
    \top_I.branch[30].block[4].um_I.ow[1] ,
    \top_I.branch[30].block[4].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[5].um_I.block_30_5.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[5].um_I.block_30_5.vpwr ),
    .ctrl(\top_I.branch[30].block[5].um_I.pg_vdd ));
 tt_um_mayrmichael_wave_generator \top_I.branch[30].block[5].um_I.block_30_5.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[5].um_I.block_30_5.vpwr ),
    .clk(\top_I.branch[30].block[5].um_I.clk ),
    .ena(\top_I.branch[30].block[5].um_I.ena ),
    .rst_n(\top_I.branch[30].block[5].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[5].um_I.iw[9] ,
    \top_I.branch[30].block[5].um_I.iw[8] ,
    \top_I.branch[30].block[5].um_I.iw[7] ,
    \top_I.branch[30].block[5].um_I.iw[6] ,
    \top_I.branch[30].block[5].um_I.iw[5] ,
    \top_I.branch[30].block[5].um_I.iw[4] ,
    \top_I.branch[30].block[5].um_I.iw[3] ,
    \top_I.branch[30].block[5].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[5].um_I.iw[17] ,
    \top_I.branch[30].block[5].um_I.iw[16] ,
    \top_I.branch[30].block[5].um_I.iw[15] ,
    \top_I.branch[30].block[5].um_I.iw[14] ,
    \top_I.branch[30].block[5].um_I.iw[13] ,
    \top_I.branch[30].block[5].um_I.iw[12] ,
    \top_I.branch[30].block[5].um_I.iw[11] ,
    \top_I.branch[30].block[5].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[5].um_I.ow[23] ,
    \top_I.branch[30].block[5].um_I.ow[22] ,
    \top_I.branch[30].block[5].um_I.ow[21] ,
    \top_I.branch[30].block[5].um_I.ow[20] ,
    \top_I.branch[30].block[5].um_I.ow[19] ,
    \top_I.branch[30].block[5].um_I.ow[18] ,
    \top_I.branch[30].block[5].um_I.ow[17] ,
    \top_I.branch[30].block[5].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[5].um_I.ow[15] ,
    \top_I.branch[30].block[5].um_I.ow[14] ,
    \top_I.branch[30].block[5].um_I.ow[13] ,
    \top_I.branch[30].block[5].um_I.ow[12] ,
    \top_I.branch[30].block[5].um_I.ow[11] ,
    \top_I.branch[30].block[5].um_I.ow[10] ,
    \top_I.branch[30].block[5].um_I.ow[9] ,
    \top_I.branch[30].block[5].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[5].um_I.ow[7] ,
    \top_I.branch[30].block[5].um_I.ow[6] ,
    \top_I.branch[30].block[5].um_I.ow[5] ,
    \top_I.branch[30].block[5].um_I.ow[4] ,
    \top_I.branch[30].block[5].um_I.ow[3] ,
    \top_I.branch[30].block[5].um_I.ow[2] ,
    \top_I.branch[30].block[5].um_I.ow[1] ,
    \top_I.branch[30].block[5].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[6].um_I.block_30_6.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[6].um_I.block_30_6.vpwr ),
    .ctrl(\top_I.branch[30].block[6].um_I.pg_vdd ));
 tt_um_moving_average_master \top_I.branch[30].block[6].um_I.block_30_6.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[6].um_I.block_30_6.vpwr ),
    .clk(\top_I.branch[30].block[6].um_I.clk ),
    .ena(\top_I.branch[30].block[6].um_I.ena ),
    .rst_n(\top_I.branch[30].block[6].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[6].um_I.iw[9] ,
    \top_I.branch[30].block[6].um_I.iw[8] ,
    \top_I.branch[30].block[6].um_I.iw[7] ,
    \top_I.branch[30].block[6].um_I.iw[6] ,
    \top_I.branch[30].block[6].um_I.iw[5] ,
    \top_I.branch[30].block[6].um_I.iw[4] ,
    \top_I.branch[30].block[6].um_I.iw[3] ,
    \top_I.branch[30].block[6].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[6].um_I.iw[17] ,
    \top_I.branch[30].block[6].um_I.iw[16] ,
    \top_I.branch[30].block[6].um_I.iw[15] ,
    \top_I.branch[30].block[6].um_I.iw[14] ,
    \top_I.branch[30].block[6].um_I.iw[13] ,
    \top_I.branch[30].block[6].um_I.iw[12] ,
    \top_I.branch[30].block[6].um_I.iw[11] ,
    \top_I.branch[30].block[6].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[6].um_I.ow[23] ,
    \top_I.branch[30].block[6].um_I.ow[22] ,
    \top_I.branch[30].block[6].um_I.ow[21] ,
    \top_I.branch[30].block[6].um_I.ow[20] ,
    \top_I.branch[30].block[6].um_I.ow[19] ,
    \top_I.branch[30].block[6].um_I.ow[18] ,
    \top_I.branch[30].block[6].um_I.ow[17] ,
    \top_I.branch[30].block[6].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[6].um_I.ow[15] ,
    \top_I.branch[30].block[6].um_I.ow[14] ,
    \top_I.branch[30].block[6].um_I.ow[13] ,
    \top_I.branch[30].block[6].um_I.ow[12] ,
    \top_I.branch[30].block[6].um_I.ow[11] ,
    \top_I.branch[30].block[6].um_I.ow[10] ,
    \top_I.branch[30].block[6].um_I.ow[9] ,
    \top_I.branch[30].block[6].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[6].um_I.ow[7] ,
    \top_I.branch[30].block[6].um_I.ow[6] ,
    \top_I.branch[30].block[6].um_I.ow[5] ,
    \top_I.branch[30].block[6].um_I.ow[4] ,
    \top_I.branch[30].block[6].um_I.ow[3] ,
    \top_I.branch[30].block[6].um_I.ow[2] ,
    \top_I.branch[30].block[6].um_I.ow[1] ,
    \top_I.branch[30].block[6].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[7].um_I.block_30_7.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[7].um_I.block_30_7.vpwr ),
    .ctrl(\top_I.branch[30].block[7].um_I.pg_vdd ));
 tt_um_advanced_counter \top_I.branch[30].block[7].um_I.block_30_7.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[7].um_I.block_30_7.vpwr ),
    .clk(\top_I.branch[30].block[7].um_I.clk ),
    .ena(\top_I.branch[30].block[7].um_I.ena ),
    .rst_n(\top_I.branch[30].block[7].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[7].um_I.iw[9] ,
    \top_I.branch[30].block[7].um_I.iw[8] ,
    \top_I.branch[30].block[7].um_I.iw[7] ,
    \top_I.branch[30].block[7].um_I.iw[6] ,
    \top_I.branch[30].block[7].um_I.iw[5] ,
    \top_I.branch[30].block[7].um_I.iw[4] ,
    \top_I.branch[30].block[7].um_I.iw[3] ,
    \top_I.branch[30].block[7].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[7].um_I.iw[17] ,
    \top_I.branch[30].block[7].um_I.iw[16] ,
    \top_I.branch[30].block[7].um_I.iw[15] ,
    \top_I.branch[30].block[7].um_I.iw[14] ,
    \top_I.branch[30].block[7].um_I.iw[13] ,
    \top_I.branch[30].block[7].um_I.iw[12] ,
    \top_I.branch[30].block[7].um_I.iw[11] ,
    \top_I.branch[30].block[7].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[7].um_I.ow[23] ,
    \top_I.branch[30].block[7].um_I.ow[22] ,
    \top_I.branch[30].block[7].um_I.ow[21] ,
    \top_I.branch[30].block[7].um_I.ow[20] ,
    \top_I.branch[30].block[7].um_I.ow[19] ,
    \top_I.branch[30].block[7].um_I.ow[18] ,
    \top_I.branch[30].block[7].um_I.ow[17] ,
    \top_I.branch[30].block[7].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[7].um_I.ow[15] ,
    \top_I.branch[30].block[7].um_I.ow[14] ,
    \top_I.branch[30].block[7].um_I.ow[13] ,
    \top_I.branch[30].block[7].um_I.ow[12] ,
    \top_I.branch[30].block[7].um_I.ow[11] ,
    \top_I.branch[30].block[7].um_I.ow[10] ,
    \top_I.branch[30].block[7].um_I.ow[9] ,
    \top_I.branch[30].block[7].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[7].um_I.ow[7] ,
    \top_I.branch[30].block[7].um_I.ow[6] ,
    \top_I.branch[30].block[7].um_I.ow[5] ,
    \top_I.branch[30].block[7].um_I.ow[4] ,
    \top_I.branch[30].block[7].um_I.ow[3] ,
    \top_I.branch[30].block[7].um_I.ow[2] ,
    \top_I.branch[30].block[7].um_I.ow[1] ,
    \top_I.branch[30].block[7].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[8].um_I.block_30_8.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[8].um_I.block_30_8.vpwr ),
    .ctrl(\top_I.branch[30].block[8].um_I.pg_vdd ));
 tt_um_rgbled_decoder \top_I.branch[30].block[8].um_I.block_30_8.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[8].um_I.block_30_8.vpwr ),
    .clk(\top_I.branch[30].block[8].um_I.clk ),
    .ena(\top_I.branch[30].block[8].um_I.ena ),
    .rst_n(\top_I.branch[30].block[8].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[8].um_I.iw[9] ,
    \top_I.branch[30].block[8].um_I.iw[8] ,
    \top_I.branch[30].block[8].um_I.iw[7] ,
    \top_I.branch[30].block[8].um_I.iw[6] ,
    \top_I.branch[30].block[8].um_I.iw[5] ,
    \top_I.branch[30].block[8].um_I.iw[4] ,
    \top_I.branch[30].block[8].um_I.iw[3] ,
    \top_I.branch[30].block[8].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[8].um_I.iw[17] ,
    \top_I.branch[30].block[8].um_I.iw[16] ,
    \top_I.branch[30].block[8].um_I.iw[15] ,
    \top_I.branch[30].block[8].um_I.iw[14] ,
    \top_I.branch[30].block[8].um_I.iw[13] ,
    \top_I.branch[30].block[8].um_I.iw[12] ,
    \top_I.branch[30].block[8].um_I.iw[11] ,
    \top_I.branch[30].block[8].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[8].um_I.ow[23] ,
    \top_I.branch[30].block[8].um_I.ow[22] ,
    \top_I.branch[30].block[8].um_I.ow[21] ,
    \top_I.branch[30].block[8].um_I.ow[20] ,
    \top_I.branch[30].block[8].um_I.ow[19] ,
    \top_I.branch[30].block[8].um_I.ow[18] ,
    \top_I.branch[30].block[8].um_I.ow[17] ,
    \top_I.branch[30].block[8].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[8].um_I.ow[15] ,
    \top_I.branch[30].block[8].um_I.ow[14] ,
    \top_I.branch[30].block[8].um_I.ow[13] ,
    \top_I.branch[30].block[8].um_I.ow[12] ,
    \top_I.branch[30].block[8].um_I.ow[11] ,
    \top_I.branch[30].block[8].um_I.ow[10] ,
    \top_I.branch[30].block[8].um_I.ow[9] ,
    \top_I.branch[30].block[8].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[8].um_I.ow[7] ,
    \top_I.branch[30].block[8].um_I.ow[6] ,
    \top_I.branch[30].block[8].um_I.ow[5] ,
    \top_I.branch[30].block[8].um_I.ow[4] ,
    \top_I.branch[30].block[8].um_I.ow[3] ,
    \top_I.branch[30].block[8].um_I.ow[2] ,
    \top_I.branch[30].block[8].um_I.ow[1] ,
    \top_I.branch[30].block[8].um_I.ow[0] }));
 tt_pg_vdd_1 \top_I.branch[30].block[9].um_I.block_30_9.tt_pg_vdd_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .GPWR(\top_I.branch[30].block[9].um_I.block_30_9.vpwr ),
    .ctrl(\top_I.branch[30].block[9].um_I.pg_vdd ));
 tt_um_FanCTRL_DomnikBrandstetter \top_I.branch[30].block[9].um_I.block_30_9.tt_um_I  (.VGND(vssd1),
    .VPWR(\top_I.branch[30].block[9].um_I.block_30_9.vpwr ),
    .clk(\top_I.branch[30].block[9].um_I.clk ),
    .ena(\top_I.branch[30].block[9].um_I.ena ),
    .rst_n(\top_I.branch[30].block[9].um_I.iw[1] ),
    .ui_in({\top_I.branch[30].block[9].um_I.iw[9] ,
    \top_I.branch[30].block[9].um_I.iw[8] ,
    \top_I.branch[30].block[9].um_I.iw[7] ,
    \top_I.branch[30].block[9].um_I.iw[6] ,
    \top_I.branch[30].block[9].um_I.iw[5] ,
    \top_I.branch[30].block[9].um_I.iw[4] ,
    \top_I.branch[30].block[9].um_I.iw[3] ,
    \top_I.branch[30].block[9].um_I.iw[2] }),
    .uio_in({\top_I.branch[30].block[9].um_I.iw[17] ,
    \top_I.branch[30].block[9].um_I.iw[16] ,
    \top_I.branch[30].block[9].um_I.iw[15] ,
    \top_I.branch[30].block[9].um_I.iw[14] ,
    \top_I.branch[30].block[9].um_I.iw[13] ,
    \top_I.branch[30].block[9].um_I.iw[12] ,
    \top_I.branch[30].block[9].um_I.iw[11] ,
    \top_I.branch[30].block[9].um_I.iw[10] }),
    .uio_oe({\top_I.branch[30].block[9].um_I.ow[23] ,
    \top_I.branch[30].block[9].um_I.ow[22] ,
    \top_I.branch[30].block[9].um_I.ow[21] ,
    \top_I.branch[30].block[9].um_I.ow[20] ,
    \top_I.branch[30].block[9].um_I.ow[19] ,
    \top_I.branch[30].block[9].um_I.ow[18] ,
    \top_I.branch[30].block[9].um_I.ow[17] ,
    \top_I.branch[30].block[9].um_I.ow[16] }),
    .uio_out({\top_I.branch[30].block[9].um_I.ow[15] ,
    \top_I.branch[30].block[9].um_I.ow[14] ,
    \top_I.branch[30].block[9].um_I.ow[13] ,
    \top_I.branch[30].block[9].um_I.ow[12] ,
    \top_I.branch[30].block[9].um_I.ow[11] ,
    \top_I.branch[30].block[9].um_I.ow[10] ,
    \top_I.branch[30].block[9].um_I.ow[9] ,
    \top_I.branch[30].block[9].um_I.ow[8] }),
    .uo_out({\top_I.branch[30].block[9].um_I.ow[7] ,
    \top_I.branch[30].block[9].um_I.ow[6] ,
    \top_I.branch[30].block[9].um_I.ow[5] ,
    \top_I.branch[30].block[9].um_I.ow[4] ,
    \top_I.branch[30].block[9].um_I.ow[3] ,
    \top_I.branch[30].block[9].um_I.ow[2] ,
    \top_I.branch[30].block[9].um_I.ow[1] ,
    \top_I.branch[30].block[9].um_I.ow[0] }));
 tt_mux \top_I.branch[30].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[30].l_addr[0] ),
    .k_zero(\top_I.branch[30].l_k_zero ),
    .addr({\top_I.branch[30].l_addr[0] ,
    \top_I.branch[30].l_addr[0] ,
    \top_I.branch[30].l_addr[0] ,
    \top_I.branch[30].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[30].block[15].um_I.ena ,
    \top_I.branch[30].block[14].um_I.ena ,
    \top_I.branch[30].block[13].um_I.ena ,
    \top_I.branch[30].block[12].um_I.ena ,
    \top_I.branch[30].block[11].um_I.ena ,
    \top_I.branch[30].block[10].um_I.ena ,
    \top_I.branch[30].block[9].um_I.ena ,
    \top_I.branch[30].block[8].um_I.ena ,
    \top_I.branch[30].block[7].um_I.ena ,
    \top_I.branch[30].block[6].um_I.ena ,
    \top_I.branch[30].block[5].um_I.ena ,
    \top_I.branch[30].block[4].um_I.ena ,
    \top_I.branch[30].block[3].um_I.ena ,
    \top_I.branch[30].block[2].um_I.ena ,
    \top_I.branch[30].block[1].um_I.ena ,
    \top_I.branch[30].block[0].um_I.ena }),
    .um_iw({\top_I.branch[30].block[15].um_I.iw[17] ,
    \top_I.branch[30].block[15].um_I.iw[16] ,
    \top_I.branch[30].block[15].um_I.iw[15] ,
    \top_I.branch[30].block[15].um_I.iw[14] ,
    \top_I.branch[30].block[15].um_I.iw[13] ,
    \top_I.branch[30].block[15].um_I.iw[12] ,
    \top_I.branch[30].block[15].um_I.iw[11] ,
    \top_I.branch[30].block[15].um_I.iw[10] ,
    \top_I.branch[30].block[15].um_I.iw[9] ,
    \top_I.branch[30].block[15].um_I.iw[8] ,
    \top_I.branch[30].block[15].um_I.iw[7] ,
    \top_I.branch[30].block[15].um_I.iw[6] ,
    \top_I.branch[30].block[15].um_I.iw[5] ,
    \top_I.branch[30].block[15].um_I.iw[4] ,
    \top_I.branch[30].block[15].um_I.iw[3] ,
    \top_I.branch[30].block[15].um_I.iw[2] ,
    \top_I.branch[30].block[15].um_I.iw[1] ,
    \top_I.branch[30].block[15].um_I.clk ,
    \top_I.branch[30].block[14].um_I.iw[17] ,
    \top_I.branch[30].block[14].um_I.iw[16] ,
    \top_I.branch[30].block[14].um_I.iw[15] ,
    \top_I.branch[30].block[14].um_I.iw[14] ,
    \top_I.branch[30].block[14].um_I.iw[13] ,
    \top_I.branch[30].block[14].um_I.iw[12] ,
    \top_I.branch[30].block[14].um_I.iw[11] ,
    \top_I.branch[30].block[14].um_I.iw[10] ,
    \top_I.branch[30].block[14].um_I.iw[9] ,
    \top_I.branch[30].block[14].um_I.iw[8] ,
    \top_I.branch[30].block[14].um_I.iw[7] ,
    \top_I.branch[30].block[14].um_I.iw[6] ,
    \top_I.branch[30].block[14].um_I.iw[5] ,
    \top_I.branch[30].block[14].um_I.iw[4] ,
    \top_I.branch[30].block[14].um_I.iw[3] ,
    \top_I.branch[30].block[14].um_I.iw[2] ,
    \top_I.branch[30].block[14].um_I.iw[1] ,
    \top_I.branch[30].block[14].um_I.clk ,
    \top_I.branch[30].block[13].um_I.iw[17] ,
    \top_I.branch[30].block[13].um_I.iw[16] ,
    \top_I.branch[30].block[13].um_I.iw[15] ,
    \top_I.branch[30].block[13].um_I.iw[14] ,
    \top_I.branch[30].block[13].um_I.iw[13] ,
    \top_I.branch[30].block[13].um_I.iw[12] ,
    \top_I.branch[30].block[13].um_I.iw[11] ,
    \top_I.branch[30].block[13].um_I.iw[10] ,
    \top_I.branch[30].block[13].um_I.iw[9] ,
    \top_I.branch[30].block[13].um_I.iw[8] ,
    \top_I.branch[30].block[13].um_I.iw[7] ,
    \top_I.branch[30].block[13].um_I.iw[6] ,
    \top_I.branch[30].block[13].um_I.iw[5] ,
    \top_I.branch[30].block[13].um_I.iw[4] ,
    \top_I.branch[30].block[13].um_I.iw[3] ,
    \top_I.branch[30].block[13].um_I.iw[2] ,
    \top_I.branch[30].block[13].um_I.iw[1] ,
    \top_I.branch[30].block[13].um_I.clk ,
    \top_I.branch[30].block[12].um_I.iw[17] ,
    \top_I.branch[30].block[12].um_I.iw[16] ,
    \top_I.branch[30].block[12].um_I.iw[15] ,
    \top_I.branch[30].block[12].um_I.iw[14] ,
    \top_I.branch[30].block[12].um_I.iw[13] ,
    \top_I.branch[30].block[12].um_I.iw[12] ,
    \top_I.branch[30].block[12].um_I.iw[11] ,
    \top_I.branch[30].block[12].um_I.iw[10] ,
    \top_I.branch[30].block[12].um_I.iw[9] ,
    \top_I.branch[30].block[12].um_I.iw[8] ,
    \top_I.branch[30].block[12].um_I.iw[7] ,
    \top_I.branch[30].block[12].um_I.iw[6] ,
    \top_I.branch[30].block[12].um_I.iw[5] ,
    \top_I.branch[30].block[12].um_I.iw[4] ,
    \top_I.branch[30].block[12].um_I.iw[3] ,
    \top_I.branch[30].block[12].um_I.iw[2] ,
    \top_I.branch[30].block[12].um_I.iw[1] ,
    \top_I.branch[30].block[12].um_I.clk ,
    \top_I.branch[30].block[11].um_I.iw[17] ,
    \top_I.branch[30].block[11].um_I.iw[16] ,
    \top_I.branch[30].block[11].um_I.iw[15] ,
    \top_I.branch[30].block[11].um_I.iw[14] ,
    \top_I.branch[30].block[11].um_I.iw[13] ,
    \top_I.branch[30].block[11].um_I.iw[12] ,
    \top_I.branch[30].block[11].um_I.iw[11] ,
    \top_I.branch[30].block[11].um_I.iw[10] ,
    \top_I.branch[30].block[11].um_I.iw[9] ,
    \top_I.branch[30].block[11].um_I.iw[8] ,
    \top_I.branch[30].block[11].um_I.iw[7] ,
    \top_I.branch[30].block[11].um_I.iw[6] ,
    \top_I.branch[30].block[11].um_I.iw[5] ,
    \top_I.branch[30].block[11].um_I.iw[4] ,
    \top_I.branch[30].block[11].um_I.iw[3] ,
    \top_I.branch[30].block[11].um_I.iw[2] ,
    \top_I.branch[30].block[11].um_I.iw[1] ,
    \top_I.branch[30].block[11].um_I.clk ,
    \top_I.branch[30].block[10].um_I.iw[17] ,
    \top_I.branch[30].block[10].um_I.iw[16] ,
    \top_I.branch[30].block[10].um_I.iw[15] ,
    \top_I.branch[30].block[10].um_I.iw[14] ,
    \top_I.branch[30].block[10].um_I.iw[13] ,
    \top_I.branch[30].block[10].um_I.iw[12] ,
    \top_I.branch[30].block[10].um_I.iw[11] ,
    \top_I.branch[30].block[10].um_I.iw[10] ,
    \top_I.branch[30].block[10].um_I.iw[9] ,
    \top_I.branch[30].block[10].um_I.iw[8] ,
    \top_I.branch[30].block[10].um_I.iw[7] ,
    \top_I.branch[30].block[10].um_I.iw[6] ,
    \top_I.branch[30].block[10].um_I.iw[5] ,
    \top_I.branch[30].block[10].um_I.iw[4] ,
    \top_I.branch[30].block[10].um_I.iw[3] ,
    \top_I.branch[30].block[10].um_I.iw[2] ,
    \top_I.branch[30].block[10].um_I.iw[1] ,
    \top_I.branch[30].block[10].um_I.clk ,
    \top_I.branch[30].block[9].um_I.iw[17] ,
    \top_I.branch[30].block[9].um_I.iw[16] ,
    \top_I.branch[30].block[9].um_I.iw[15] ,
    \top_I.branch[30].block[9].um_I.iw[14] ,
    \top_I.branch[30].block[9].um_I.iw[13] ,
    \top_I.branch[30].block[9].um_I.iw[12] ,
    \top_I.branch[30].block[9].um_I.iw[11] ,
    \top_I.branch[30].block[9].um_I.iw[10] ,
    \top_I.branch[30].block[9].um_I.iw[9] ,
    \top_I.branch[30].block[9].um_I.iw[8] ,
    \top_I.branch[30].block[9].um_I.iw[7] ,
    \top_I.branch[30].block[9].um_I.iw[6] ,
    \top_I.branch[30].block[9].um_I.iw[5] ,
    \top_I.branch[30].block[9].um_I.iw[4] ,
    \top_I.branch[30].block[9].um_I.iw[3] ,
    \top_I.branch[30].block[9].um_I.iw[2] ,
    \top_I.branch[30].block[9].um_I.iw[1] ,
    \top_I.branch[30].block[9].um_I.clk ,
    \top_I.branch[30].block[8].um_I.iw[17] ,
    \top_I.branch[30].block[8].um_I.iw[16] ,
    \top_I.branch[30].block[8].um_I.iw[15] ,
    \top_I.branch[30].block[8].um_I.iw[14] ,
    \top_I.branch[30].block[8].um_I.iw[13] ,
    \top_I.branch[30].block[8].um_I.iw[12] ,
    \top_I.branch[30].block[8].um_I.iw[11] ,
    \top_I.branch[30].block[8].um_I.iw[10] ,
    \top_I.branch[30].block[8].um_I.iw[9] ,
    \top_I.branch[30].block[8].um_I.iw[8] ,
    \top_I.branch[30].block[8].um_I.iw[7] ,
    \top_I.branch[30].block[8].um_I.iw[6] ,
    \top_I.branch[30].block[8].um_I.iw[5] ,
    \top_I.branch[30].block[8].um_I.iw[4] ,
    \top_I.branch[30].block[8].um_I.iw[3] ,
    \top_I.branch[30].block[8].um_I.iw[2] ,
    \top_I.branch[30].block[8].um_I.iw[1] ,
    \top_I.branch[30].block[8].um_I.clk ,
    \top_I.branch[30].block[7].um_I.iw[17] ,
    \top_I.branch[30].block[7].um_I.iw[16] ,
    \top_I.branch[30].block[7].um_I.iw[15] ,
    \top_I.branch[30].block[7].um_I.iw[14] ,
    \top_I.branch[30].block[7].um_I.iw[13] ,
    \top_I.branch[30].block[7].um_I.iw[12] ,
    \top_I.branch[30].block[7].um_I.iw[11] ,
    \top_I.branch[30].block[7].um_I.iw[10] ,
    \top_I.branch[30].block[7].um_I.iw[9] ,
    \top_I.branch[30].block[7].um_I.iw[8] ,
    \top_I.branch[30].block[7].um_I.iw[7] ,
    \top_I.branch[30].block[7].um_I.iw[6] ,
    \top_I.branch[30].block[7].um_I.iw[5] ,
    \top_I.branch[30].block[7].um_I.iw[4] ,
    \top_I.branch[30].block[7].um_I.iw[3] ,
    \top_I.branch[30].block[7].um_I.iw[2] ,
    \top_I.branch[30].block[7].um_I.iw[1] ,
    \top_I.branch[30].block[7].um_I.clk ,
    \top_I.branch[30].block[6].um_I.iw[17] ,
    \top_I.branch[30].block[6].um_I.iw[16] ,
    \top_I.branch[30].block[6].um_I.iw[15] ,
    \top_I.branch[30].block[6].um_I.iw[14] ,
    \top_I.branch[30].block[6].um_I.iw[13] ,
    \top_I.branch[30].block[6].um_I.iw[12] ,
    \top_I.branch[30].block[6].um_I.iw[11] ,
    \top_I.branch[30].block[6].um_I.iw[10] ,
    \top_I.branch[30].block[6].um_I.iw[9] ,
    \top_I.branch[30].block[6].um_I.iw[8] ,
    \top_I.branch[30].block[6].um_I.iw[7] ,
    \top_I.branch[30].block[6].um_I.iw[6] ,
    \top_I.branch[30].block[6].um_I.iw[5] ,
    \top_I.branch[30].block[6].um_I.iw[4] ,
    \top_I.branch[30].block[6].um_I.iw[3] ,
    \top_I.branch[30].block[6].um_I.iw[2] ,
    \top_I.branch[30].block[6].um_I.iw[1] ,
    \top_I.branch[30].block[6].um_I.clk ,
    \top_I.branch[30].block[5].um_I.iw[17] ,
    \top_I.branch[30].block[5].um_I.iw[16] ,
    \top_I.branch[30].block[5].um_I.iw[15] ,
    \top_I.branch[30].block[5].um_I.iw[14] ,
    \top_I.branch[30].block[5].um_I.iw[13] ,
    \top_I.branch[30].block[5].um_I.iw[12] ,
    \top_I.branch[30].block[5].um_I.iw[11] ,
    \top_I.branch[30].block[5].um_I.iw[10] ,
    \top_I.branch[30].block[5].um_I.iw[9] ,
    \top_I.branch[30].block[5].um_I.iw[8] ,
    \top_I.branch[30].block[5].um_I.iw[7] ,
    \top_I.branch[30].block[5].um_I.iw[6] ,
    \top_I.branch[30].block[5].um_I.iw[5] ,
    \top_I.branch[30].block[5].um_I.iw[4] ,
    \top_I.branch[30].block[5].um_I.iw[3] ,
    \top_I.branch[30].block[5].um_I.iw[2] ,
    \top_I.branch[30].block[5].um_I.iw[1] ,
    \top_I.branch[30].block[5].um_I.clk ,
    \top_I.branch[30].block[4].um_I.iw[17] ,
    \top_I.branch[30].block[4].um_I.iw[16] ,
    \top_I.branch[30].block[4].um_I.iw[15] ,
    \top_I.branch[30].block[4].um_I.iw[14] ,
    \top_I.branch[30].block[4].um_I.iw[13] ,
    \top_I.branch[30].block[4].um_I.iw[12] ,
    \top_I.branch[30].block[4].um_I.iw[11] ,
    \top_I.branch[30].block[4].um_I.iw[10] ,
    \top_I.branch[30].block[4].um_I.iw[9] ,
    \top_I.branch[30].block[4].um_I.iw[8] ,
    \top_I.branch[30].block[4].um_I.iw[7] ,
    \top_I.branch[30].block[4].um_I.iw[6] ,
    \top_I.branch[30].block[4].um_I.iw[5] ,
    \top_I.branch[30].block[4].um_I.iw[4] ,
    \top_I.branch[30].block[4].um_I.iw[3] ,
    \top_I.branch[30].block[4].um_I.iw[2] ,
    \top_I.branch[30].block[4].um_I.iw[1] ,
    \top_I.branch[30].block[4].um_I.clk ,
    \top_I.branch[30].block[3].um_I.iw[17] ,
    \top_I.branch[30].block[3].um_I.iw[16] ,
    \top_I.branch[30].block[3].um_I.iw[15] ,
    \top_I.branch[30].block[3].um_I.iw[14] ,
    \top_I.branch[30].block[3].um_I.iw[13] ,
    \top_I.branch[30].block[3].um_I.iw[12] ,
    \top_I.branch[30].block[3].um_I.iw[11] ,
    \top_I.branch[30].block[3].um_I.iw[10] ,
    \top_I.branch[30].block[3].um_I.iw[9] ,
    \top_I.branch[30].block[3].um_I.iw[8] ,
    \top_I.branch[30].block[3].um_I.iw[7] ,
    \top_I.branch[30].block[3].um_I.iw[6] ,
    \top_I.branch[30].block[3].um_I.iw[5] ,
    \top_I.branch[30].block[3].um_I.iw[4] ,
    \top_I.branch[30].block[3].um_I.iw[3] ,
    \top_I.branch[30].block[3].um_I.iw[2] ,
    \top_I.branch[30].block[3].um_I.iw[1] ,
    \top_I.branch[30].block[3].um_I.clk ,
    \top_I.branch[30].block[2].um_I.iw[17] ,
    \top_I.branch[30].block[2].um_I.iw[16] ,
    \top_I.branch[30].block[2].um_I.iw[15] ,
    \top_I.branch[30].block[2].um_I.iw[14] ,
    \top_I.branch[30].block[2].um_I.iw[13] ,
    \top_I.branch[30].block[2].um_I.iw[12] ,
    \top_I.branch[30].block[2].um_I.iw[11] ,
    \top_I.branch[30].block[2].um_I.iw[10] ,
    \top_I.branch[30].block[2].um_I.iw[9] ,
    \top_I.branch[30].block[2].um_I.iw[8] ,
    \top_I.branch[30].block[2].um_I.iw[7] ,
    \top_I.branch[30].block[2].um_I.iw[6] ,
    \top_I.branch[30].block[2].um_I.iw[5] ,
    \top_I.branch[30].block[2].um_I.iw[4] ,
    \top_I.branch[30].block[2].um_I.iw[3] ,
    \top_I.branch[30].block[2].um_I.iw[2] ,
    \top_I.branch[30].block[2].um_I.iw[1] ,
    \top_I.branch[30].block[2].um_I.clk ,
    \top_I.branch[30].block[1].um_I.iw[17] ,
    \top_I.branch[30].block[1].um_I.iw[16] ,
    \top_I.branch[30].block[1].um_I.iw[15] ,
    \top_I.branch[30].block[1].um_I.iw[14] ,
    \top_I.branch[30].block[1].um_I.iw[13] ,
    \top_I.branch[30].block[1].um_I.iw[12] ,
    \top_I.branch[30].block[1].um_I.iw[11] ,
    \top_I.branch[30].block[1].um_I.iw[10] ,
    \top_I.branch[30].block[1].um_I.iw[9] ,
    \top_I.branch[30].block[1].um_I.iw[8] ,
    \top_I.branch[30].block[1].um_I.iw[7] ,
    \top_I.branch[30].block[1].um_I.iw[6] ,
    \top_I.branch[30].block[1].um_I.iw[5] ,
    \top_I.branch[30].block[1].um_I.iw[4] ,
    \top_I.branch[30].block[1].um_I.iw[3] ,
    \top_I.branch[30].block[1].um_I.iw[2] ,
    \top_I.branch[30].block[1].um_I.iw[1] ,
    \top_I.branch[30].block[1].um_I.clk ,
    \top_I.branch[30].block[0].um_I.iw[17] ,
    \top_I.branch[30].block[0].um_I.iw[16] ,
    \top_I.branch[30].block[0].um_I.iw[15] ,
    \top_I.branch[30].block[0].um_I.iw[14] ,
    \top_I.branch[30].block[0].um_I.iw[13] ,
    \top_I.branch[30].block[0].um_I.iw[12] ,
    \top_I.branch[30].block[0].um_I.iw[11] ,
    \top_I.branch[30].block[0].um_I.iw[10] ,
    \top_I.branch[30].block[0].um_I.iw[9] ,
    \top_I.branch[30].block[0].um_I.iw[8] ,
    \top_I.branch[30].block[0].um_I.iw[7] ,
    \top_I.branch[30].block[0].um_I.iw[6] ,
    \top_I.branch[30].block[0].um_I.iw[5] ,
    \top_I.branch[30].block[0].um_I.iw[4] ,
    \top_I.branch[30].block[0].um_I.iw[3] ,
    \top_I.branch[30].block[0].um_I.iw[2] ,
    \top_I.branch[30].block[0].um_I.iw[1] ,
    \top_I.branch[30].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[30].block[15].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[13].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[11].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[9].um_I.k_zero ,
    \top_I.branch[30].block[8].um_I.k_zero ,
    \top_I.branch[30].block[7].um_I.k_zero ,
    \top_I.branch[30].block[6].um_I.k_zero ,
    \top_I.branch[30].block[5].um_I.k_zero ,
    \top_I.branch[30].block[4].um_I.k_zero ,
    \top_I.branch[30].block[3].um_I.k_zero ,
    \top_I.branch[30].block[2].um_I.k_zero ,
    \top_I.branch[30].block[1].um_I.k_zero ,
    \top_I.branch[30].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[30].block[15].um_I.ow[23] ,
    \top_I.branch[30].block[15].um_I.ow[22] ,
    \top_I.branch[30].block[15].um_I.ow[21] ,
    \top_I.branch[30].block[15].um_I.ow[20] ,
    \top_I.branch[30].block[15].um_I.ow[19] ,
    \top_I.branch[30].block[15].um_I.ow[18] ,
    \top_I.branch[30].block[15].um_I.ow[17] ,
    \top_I.branch[30].block[15].um_I.ow[16] ,
    \top_I.branch[30].block[15].um_I.ow[15] ,
    \top_I.branch[30].block[15].um_I.ow[14] ,
    \top_I.branch[30].block[15].um_I.ow[13] ,
    \top_I.branch[30].block[15].um_I.ow[12] ,
    \top_I.branch[30].block[15].um_I.ow[11] ,
    \top_I.branch[30].block[15].um_I.ow[10] ,
    \top_I.branch[30].block[15].um_I.ow[9] ,
    \top_I.branch[30].block[15].um_I.ow[8] ,
    \top_I.branch[30].block[15].um_I.ow[7] ,
    \top_I.branch[30].block[15].um_I.ow[6] ,
    \top_I.branch[30].block[15].um_I.ow[5] ,
    \top_I.branch[30].block[15].um_I.ow[4] ,
    \top_I.branch[30].block[15].um_I.ow[3] ,
    \top_I.branch[30].block[15].um_I.ow[2] ,
    \top_I.branch[30].block[15].um_I.ow[1] ,
    \top_I.branch[30].block[15].um_I.ow[0] ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[14].um_I.k_zero ,
    \top_I.branch[30].block[13].um_I.ow[23] ,
    \top_I.branch[30].block[13].um_I.ow[22] ,
    \top_I.branch[30].block[13].um_I.ow[21] ,
    \top_I.branch[30].block[13].um_I.ow[20] ,
    \top_I.branch[30].block[13].um_I.ow[19] ,
    \top_I.branch[30].block[13].um_I.ow[18] ,
    \top_I.branch[30].block[13].um_I.ow[17] ,
    \top_I.branch[30].block[13].um_I.ow[16] ,
    \top_I.branch[30].block[13].um_I.ow[15] ,
    \top_I.branch[30].block[13].um_I.ow[14] ,
    \top_I.branch[30].block[13].um_I.ow[13] ,
    \top_I.branch[30].block[13].um_I.ow[12] ,
    \top_I.branch[30].block[13].um_I.ow[11] ,
    \top_I.branch[30].block[13].um_I.ow[10] ,
    \top_I.branch[30].block[13].um_I.ow[9] ,
    \top_I.branch[30].block[13].um_I.ow[8] ,
    \top_I.branch[30].block[13].um_I.ow[7] ,
    \top_I.branch[30].block[13].um_I.ow[6] ,
    \top_I.branch[30].block[13].um_I.ow[5] ,
    \top_I.branch[30].block[13].um_I.ow[4] ,
    \top_I.branch[30].block[13].um_I.ow[3] ,
    \top_I.branch[30].block[13].um_I.ow[2] ,
    \top_I.branch[30].block[13].um_I.ow[1] ,
    \top_I.branch[30].block[13].um_I.ow[0] ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[12].um_I.k_zero ,
    \top_I.branch[30].block[11].um_I.ow[23] ,
    \top_I.branch[30].block[11].um_I.ow[22] ,
    \top_I.branch[30].block[11].um_I.ow[21] ,
    \top_I.branch[30].block[11].um_I.ow[20] ,
    \top_I.branch[30].block[11].um_I.ow[19] ,
    \top_I.branch[30].block[11].um_I.ow[18] ,
    \top_I.branch[30].block[11].um_I.ow[17] ,
    \top_I.branch[30].block[11].um_I.ow[16] ,
    \top_I.branch[30].block[11].um_I.ow[15] ,
    \top_I.branch[30].block[11].um_I.ow[14] ,
    \top_I.branch[30].block[11].um_I.ow[13] ,
    \top_I.branch[30].block[11].um_I.ow[12] ,
    \top_I.branch[30].block[11].um_I.ow[11] ,
    \top_I.branch[30].block[11].um_I.ow[10] ,
    \top_I.branch[30].block[11].um_I.ow[9] ,
    \top_I.branch[30].block[11].um_I.ow[8] ,
    \top_I.branch[30].block[11].um_I.ow[7] ,
    \top_I.branch[30].block[11].um_I.ow[6] ,
    \top_I.branch[30].block[11].um_I.ow[5] ,
    \top_I.branch[30].block[11].um_I.ow[4] ,
    \top_I.branch[30].block[11].um_I.ow[3] ,
    \top_I.branch[30].block[11].um_I.ow[2] ,
    \top_I.branch[30].block[11].um_I.ow[1] ,
    \top_I.branch[30].block[11].um_I.ow[0] ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[10].um_I.k_zero ,
    \top_I.branch[30].block[9].um_I.ow[23] ,
    \top_I.branch[30].block[9].um_I.ow[22] ,
    \top_I.branch[30].block[9].um_I.ow[21] ,
    \top_I.branch[30].block[9].um_I.ow[20] ,
    \top_I.branch[30].block[9].um_I.ow[19] ,
    \top_I.branch[30].block[9].um_I.ow[18] ,
    \top_I.branch[30].block[9].um_I.ow[17] ,
    \top_I.branch[30].block[9].um_I.ow[16] ,
    \top_I.branch[30].block[9].um_I.ow[15] ,
    \top_I.branch[30].block[9].um_I.ow[14] ,
    \top_I.branch[30].block[9].um_I.ow[13] ,
    \top_I.branch[30].block[9].um_I.ow[12] ,
    \top_I.branch[30].block[9].um_I.ow[11] ,
    \top_I.branch[30].block[9].um_I.ow[10] ,
    \top_I.branch[30].block[9].um_I.ow[9] ,
    \top_I.branch[30].block[9].um_I.ow[8] ,
    \top_I.branch[30].block[9].um_I.ow[7] ,
    \top_I.branch[30].block[9].um_I.ow[6] ,
    \top_I.branch[30].block[9].um_I.ow[5] ,
    \top_I.branch[30].block[9].um_I.ow[4] ,
    \top_I.branch[30].block[9].um_I.ow[3] ,
    \top_I.branch[30].block[9].um_I.ow[2] ,
    \top_I.branch[30].block[9].um_I.ow[1] ,
    \top_I.branch[30].block[9].um_I.ow[0] ,
    \top_I.branch[30].block[8].um_I.ow[23] ,
    \top_I.branch[30].block[8].um_I.ow[22] ,
    \top_I.branch[30].block[8].um_I.ow[21] ,
    \top_I.branch[30].block[8].um_I.ow[20] ,
    \top_I.branch[30].block[8].um_I.ow[19] ,
    \top_I.branch[30].block[8].um_I.ow[18] ,
    \top_I.branch[30].block[8].um_I.ow[17] ,
    \top_I.branch[30].block[8].um_I.ow[16] ,
    \top_I.branch[30].block[8].um_I.ow[15] ,
    \top_I.branch[30].block[8].um_I.ow[14] ,
    \top_I.branch[30].block[8].um_I.ow[13] ,
    \top_I.branch[30].block[8].um_I.ow[12] ,
    \top_I.branch[30].block[8].um_I.ow[11] ,
    \top_I.branch[30].block[8].um_I.ow[10] ,
    \top_I.branch[30].block[8].um_I.ow[9] ,
    \top_I.branch[30].block[8].um_I.ow[8] ,
    \top_I.branch[30].block[8].um_I.ow[7] ,
    \top_I.branch[30].block[8].um_I.ow[6] ,
    \top_I.branch[30].block[8].um_I.ow[5] ,
    \top_I.branch[30].block[8].um_I.ow[4] ,
    \top_I.branch[30].block[8].um_I.ow[3] ,
    \top_I.branch[30].block[8].um_I.ow[2] ,
    \top_I.branch[30].block[8].um_I.ow[1] ,
    \top_I.branch[30].block[8].um_I.ow[0] ,
    \top_I.branch[30].block[7].um_I.ow[23] ,
    \top_I.branch[30].block[7].um_I.ow[22] ,
    \top_I.branch[30].block[7].um_I.ow[21] ,
    \top_I.branch[30].block[7].um_I.ow[20] ,
    \top_I.branch[30].block[7].um_I.ow[19] ,
    \top_I.branch[30].block[7].um_I.ow[18] ,
    \top_I.branch[30].block[7].um_I.ow[17] ,
    \top_I.branch[30].block[7].um_I.ow[16] ,
    \top_I.branch[30].block[7].um_I.ow[15] ,
    \top_I.branch[30].block[7].um_I.ow[14] ,
    \top_I.branch[30].block[7].um_I.ow[13] ,
    \top_I.branch[30].block[7].um_I.ow[12] ,
    \top_I.branch[30].block[7].um_I.ow[11] ,
    \top_I.branch[30].block[7].um_I.ow[10] ,
    \top_I.branch[30].block[7].um_I.ow[9] ,
    \top_I.branch[30].block[7].um_I.ow[8] ,
    \top_I.branch[30].block[7].um_I.ow[7] ,
    \top_I.branch[30].block[7].um_I.ow[6] ,
    \top_I.branch[30].block[7].um_I.ow[5] ,
    \top_I.branch[30].block[7].um_I.ow[4] ,
    \top_I.branch[30].block[7].um_I.ow[3] ,
    \top_I.branch[30].block[7].um_I.ow[2] ,
    \top_I.branch[30].block[7].um_I.ow[1] ,
    \top_I.branch[30].block[7].um_I.ow[0] ,
    \top_I.branch[30].block[6].um_I.ow[23] ,
    \top_I.branch[30].block[6].um_I.ow[22] ,
    \top_I.branch[30].block[6].um_I.ow[21] ,
    \top_I.branch[30].block[6].um_I.ow[20] ,
    \top_I.branch[30].block[6].um_I.ow[19] ,
    \top_I.branch[30].block[6].um_I.ow[18] ,
    \top_I.branch[30].block[6].um_I.ow[17] ,
    \top_I.branch[30].block[6].um_I.ow[16] ,
    \top_I.branch[30].block[6].um_I.ow[15] ,
    \top_I.branch[30].block[6].um_I.ow[14] ,
    \top_I.branch[30].block[6].um_I.ow[13] ,
    \top_I.branch[30].block[6].um_I.ow[12] ,
    \top_I.branch[30].block[6].um_I.ow[11] ,
    \top_I.branch[30].block[6].um_I.ow[10] ,
    \top_I.branch[30].block[6].um_I.ow[9] ,
    \top_I.branch[30].block[6].um_I.ow[8] ,
    \top_I.branch[30].block[6].um_I.ow[7] ,
    \top_I.branch[30].block[6].um_I.ow[6] ,
    \top_I.branch[30].block[6].um_I.ow[5] ,
    \top_I.branch[30].block[6].um_I.ow[4] ,
    \top_I.branch[30].block[6].um_I.ow[3] ,
    \top_I.branch[30].block[6].um_I.ow[2] ,
    \top_I.branch[30].block[6].um_I.ow[1] ,
    \top_I.branch[30].block[6].um_I.ow[0] ,
    \top_I.branch[30].block[5].um_I.ow[23] ,
    \top_I.branch[30].block[5].um_I.ow[22] ,
    \top_I.branch[30].block[5].um_I.ow[21] ,
    \top_I.branch[30].block[5].um_I.ow[20] ,
    \top_I.branch[30].block[5].um_I.ow[19] ,
    \top_I.branch[30].block[5].um_I.ow[18] ,
    \top_I.branch[30].block[5].um_I.ow[17] ,
    \top_I.branch[30].block[5].um_I.ow[16] ,
    \top_I.branch[30].block[5].um_I.ow[15] ,
    \top_I.branch[30].block[5].um_I.ow[14] ,
    \top_I.branch[30].block[5].um_I.ow[13] ,
    \top_I.branch[30].block[5].um_I.ow[12] ,
    \top_I.branch[30].block[5].um_I.ow[11] ,
    \top_I.branch[30].block[5].um_I.ow[10] ,
    \top_I.branch[30].block[5].um_I.ow[9] ,
    \top_I.branch[30].block[5].um_I.ow[8] ,
    \top_I.branch[30].block[5].um_I.ow[7] ,
    \top_I.branch[30].block[5].um_I.ow[6] ,
    \top_I.branch[30].block[5].um_I.ow[5] ,
    \top_I.branch[30].block[5].um_I.ow[4] ,
    \top_I.branch[30].block[5].um_I.ow[3] ,
    \top_I.branch[30].block[5].um_I.ow[2] ,
    \top_I.branch[30].block[5].um_I.ow[1] ,
    \top_I.branch[30].block[5].um_I.ow[0] ,
    \top_I.branch[30].block[4].um_I.ow[23] ,
    \top_I.branch[30].block[4].um_I.ow[22] ,
    \top_I.branch[30].block[4].um_I.ow[21] ,
    \top_I.branch[30].block[4].um_I.ow[20] ,
    \top_I.branch[30].block[4].um_I.ow[19] ,
    \top_I.branch[30].block[4].um_I.ow[18] ,
    \top_I.branch[30].block[4].um_I.ow[17] ,
    \top_I.branch[30].block[4].um_I.ow[16] ,
    \top_I.branch[30].block[4].um_I.ow[15] ,
    \top_I.branch[30].block[4].um_I.ow[14] ,
    \top_I.branch[30].block[4].um_I.ow[13] ,
    \top_I.branch[30].block[4].um_I.ow[12] ,
    \top_I.branch[30].block[4].um_I.ow[11] ,
    \top_I.branch[30].block[4].um_I.ow[10] ,
    \top_I.branch[30].block[4].um_I.ow[9] ,
    \top_I.branch[30].block[4].um_I.ow[8] ,
    \top_I.branch[30].block[4].um_I.ow[7] ,
    \top_I.branch[30].block[4].um_I.ow[6] ,
    \top_I.branch[30].block[4].um_I.ow[5] ,
    \top_I.branch[30].block[4].um_I.ow[4] ,
    \top_I.branch[30].block[4].um_I.ow[3] ,
    \top_I.branch[30].block[4].um_I.ow[2] ,
    \top_I.branch[30].block[4].um_I.ow[1] ,
    \top_I.branch[30].block[4].um_I.ow[0] ,
    \top_I.branch[30].block[3].um_I.ow[23] ,
    \top_I.branch[30].block[3].um_I.ow[22] ,
    \top_I.branch[30].block[3].um_I.ow[21] ,
    \top_I.branch[30].block[3].um_I.ow[20] ,
    \top_I.branch[30].block[3].um_I.ow[19] ,
    \top_I.branch[30].block[3].um_I.ow[18] ,
    \top_I.branch[30].block[3].um_I.ow[17] ,
    \top_I.branch[30].block[3].um_I.ow[16] ,
    \top_I.branch[30].block[3].um_I.ow[15] ,
    \top_I.branch[30].block[3].um_I.ow[14] ,
    \top_I.branch[30].block[3].um_I.ow[13] ,
    \top_I.branch[30].block[3].um_I.ow[12] ,
    \top_I.branch[30].block[3].um_I.ow[11] ,
    \top_I.branch[30].block[3].um_I.ow[10] ,
    \top_I.branch[30].block[3].um_I.ow[9] ,
    \top_I.branch[30].block[3].um_I.ow[8] ,
    \top_I.branch[30].block[3].um_I.ow[7] ,
    \top_I.branch[30].block[3].um_I.ow[6] ,
    \top_I.branch[30].block[3].um_I.ow[5] ,
    \top_I.branch[30].block[3].um_I.ow[4] ,
    \top_I.branch[30].block[3].um_I.ow[3] ,
    \top_I.branch[30].block[3].um_I.ow[2] ,
    \top_I.branch[30].block[3].um_I.ow[1] ,
    \top_I.branch[30].block[3].um_I.ow[0] ,
    \top_I.branch[30].block[2].um_I.ow[23] ,
    \top_I.branch[30].block[2].um_I.ow[22] ,
    \top_I.branch[30].block[2].um_I.ow[21] ,
    \top_I.branch[30].block[2].um_I.ow[20] ,
    \top_I.branch[30].block[2].um_I.ow[19] ,
    \top_I.branch[30].block[2].um_I.ow[18] ,
    \top_I.branch[30].block[2].um_I.ow[17] ,
    \top_I.branch[30].block[2].um_I.ow[16] ,
    \top_I.branch[30].block[2].um_I.ow[15] ,
    \top_I.branch[30].block[2].um_I.ow[14] ,
    \top_I.branch[30].block[2].um_I.ow[13] ,
    \top_I.branch[30].block[2].um_I.ow[12] ,
    \top_I.branch[30].block[2].um_I.ow[11] ,
    \top_I.branch[30].block[2].um_I.ow[10] ,
    \top_I.branch[30].block[2].um_I.ow[9] ,
    \top_I.branch[30].block[2].um_I.ow[8] ,
    \top_I.branch[30].block[2].um_I.ow[7] ,
    \top_I.branch[30].block[2].um_I.ow[6] ,
    \top_I.branch[30].block[2].um_I.ow[5] ,
    \top_I.branch[30].block[2].um_I.ow[4] ,
    \top_I.branch[30].block[2].um_I.ow[3] ,
    \top_I.branch[30].block[2].um_I.ow[2] ,
    \top_I.branch[30].block[2].um_I.ow[1] ,
    \top_I.branch[30].block[2].um_I.ow[0] ,
    \top_I.branch[30].block[1].um_I.ow[23] ,
    \top_I.branch[30].block[1].um_I.ow[22] ,
    \top_I.branch[30].block[1].um_I.ow[21] ,
    \top_I.branch[30].block[1].um_I.ow[20] ,
    \top_I.branch[30].block[1].um_I.ow[19] ,
    \top_I.branch[30].block[1].um_I.ow[18] ,
    \top_I.branch[30].block[1].um_I.ow[17] ,
    \top_I.branch[30].block[1].um_I.ow[16] ,
    \top_I.branch[30].block[1].um_I.ow[15] ,
    \top_I.branch[30].block[1].um_I.ow[14] ,
    \top_I.branch[30].block[1].um_I.ow[13] ,
    \top_I.branch[30].block[1].um_I.ow[12] ,
    \top_I.branch[30].block[1].um_I.ow[11] ,
    \top_I.branch[30].block[1].um_I.ow[10] ,
    \top_I.branch[30].block[1].um_I.ow[9] ,
    \top_I.branch[30].block[1].um_I.ow[8] ,
    \top_I.branch[30].block[1].um_I.ow[7] ,
    \top_I.branch[30].block[1].um_I.ow[6] ,
    \top_I.branch[30].block[1].um_I.ow[5] ,
    \top_I.branch[30].block[1].um_I.ow[4] ,
    \top_I.branch[30].block[1].um_I.ow[3] ,
    \top_I.branch[30].block[1].um_I.ow[2] ,
    \top_I.branch[30].block[1].um_I.ow[1] ,
    \top_I.branch[30].block[1].um_I.ow[0] ,
    \top_I.branch[30].block[0].um_I.ow[23] ,
    \top_I.branch[30].block[0].um_I.ow[22] ,
    \top_I.branch[30].block[0].um_I.ow[21] ,
    \top_I.branch[30].block[0].um_I.ow[20] ,
    \top_I.branch[30].block[0].um_I.ow[19] ,
    \top_I.branch[30].block[0].um_I.ow[18] ,
    \top_I.branch[30].block[0].um_I.ow[17] ,
    \top_I.branch[30].block[0].um_I.ow[16] ,
    \top_I.branch[30].block[0].um_I.ow[15] ,
    \top_I.branch[30].block[0].um_I.ow[14] ,
    \top_I.branch[30].block[0].um_I.ow[13] ,
    \top_I.branch[30].block[0].um_I.ow[12] ,
    \top_I.branch[30].block[0].um_I.ow[11] ,
    \top_I.branch[30].block[0].um_I.ow[10] ,
    \top_I.branch[30].block[0].um_I.ow[9] ,
    \top_I.branch[30].block[0].um_I.ow[8] ,
    \top_I.branch[30].block[0].um_I.ow[7] ,
    \top_I.branch[30].block[0].um_I.ow[6] ,
    \top_I.branch[30].block[0].um_I.ow[5] ,
    \top_I.branch[30].block[0].um_I.ow[4] ,
    \top_I.branch[30].block[0].um_I.ow[3] ,
    \top_I.branch[30].block[0].um_I.ow[2] ,
    \top_I.branch[30].block[0].um_I.ow[1] ,
    \top_I.branch[30].block[0].um_I.ow[0] }),
    .um_pg_vdd({\top_I.branch[30].block[15].um_I.pg_vdd ,
    \top_I.branch[30].block[14].um_I.pg_vdd ,
    \top_I.branch[30].block[13].um_I.pg_vdd ,
    \top_I.branch[30].block[12].um_I.pg_vdd ,
    \top_I.branch[30].block[11].um_I.pg_vdd ,
    \top_I.branch[30].block[10].um_I.pg_vdd ,
    \top_I.branch[30].block[9].um_I.pg_vdd ,
    \top_I.branch[30].block[8].um_I.pg_vdd ,
    \top_I.branch[30].block[7].um_I.pg_vdd ,
    \top_I.branch[30].block[6].um_I.pg_vdd ,
    \top_I.branch[30].block[5].um_I.pg_vdd ,
    \top_I.branch[30].block[4].um_I.pg_vdd ,
    \top_I.branch[30].block[3].um_I.pg_vdd ,
    \top_I.branch[30].block[2].um_I.pg_vdd ,
    \top_I.branch[30].block[1].um_I.pg_vdd ,
    \top_I.branch[30].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[31].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[31].l_addr[0] ),
    .k_zero(\top_I.branch[31].l_k_zero ),
    .addr({\top_I.branch[31].l_addr[0] ,
    \top_I.branch[31].l_addr[0] ,
    \top_I.branch[31].l_addr[0] ,
    \top_I.branch[31].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[31].block[15].um_I.ena ,
    \top_I.branch[31].block[14].um_I.ena ,
    \top_I.branch[31].block[13].um_I.ena ,
    \top_I.branch[31].block[12].um_I.ena ,
    \top_I.branch[31].block[11].um_I.ena ,
    \top_I.branch[31].block[10].um_I.ena ,
    \top_I.branch[31].block[9].um_I.ena ,
    \top_I.branch[31].block[8].um_I.ena ,
    \top_I.branch[31].block[7].um_I.ena ,
    \top_I.branch[31].block[6].um_I.ena ,
    \top_I.branch[31].block[5].um_I.ena ,
    \top_I.branch[31].block[4].um_I.ena ,
    \top_I.branch[31].block[3].um_I.ena ,
    \top_I.branch[31].block[2].um_I.ena ,
    \top_I.branch[31].block[1].um_I.ena ,
    \top_I.branch[31].block[0].um_I.ena }),
    .um_iw({\top_I.branch[31].block[15].um_I.iw[17] ,
    \top_I.branch[31].block[15].um_I.iw[16] ,
    \top_I.branch[31].block[15].um_I.iw[15] ,
    \top_I.branch[31].block[15].um_I.iw[14] ,
    \top_I.branch[31].block[15].um_I.iw[13] ,
    \top_I.branch[31].block[15].um_I.iw[12] ,
    \top_I.branch[31].block[15].um_I.iw[11] ,
    \top_I.branch[31].block[15].um_I.iw[10] ,
    \top_I.branch[31].block[15].um_I.iw[9] ,
    \top_I.branch[31].block[15].um_I.iw[8] ,
    \top_I.branch[31].block[15].um_I.iw[7] ,
    \top_I.branch[31].block[15].um_I.iw[6] ,
    \top_I.branch[31].block[15].um_I.iw[5] ,
    \top_I.branch[31].block[15].um_I.iw[4] ,
    \top_I.branch[31].block[15].um_I.iw[3] ,
    \top_I.branch[31].block[15].um_I.iw[2] ,
    \top_I.branch[31].block[15].um_I.iw[1] ,
    \top_I.branch[31].block[15].um_I.clk ,
    \top_I.branch[31].block[14].um_I.iw[17] ,
    \top_I.branch[31].block[14].um_I.iw[16] ,
    \top_I.branch[31].block[14].um_I.iw[15] ,
    \top_I.branch[31].block[14].um_I.iw[14] ,
    \top_I.branch[31].block[14].um_I.iw[13] ,
    \top_I.branch[31].block[14].um_I.iw[12] ,
    \top_I.branch[31].block[14].um_I.iw[11] ,
    \top_I.branch[31].block[14].um_I.iw[10] ,
    \top_I.branch[31].block[14].um_I.iw[9] ,
    \top_I.branch[31].block[14].um_I.iw[8] ,
    \top_I.branch[31].block[14].um_I.iw[7] ,
    \top_I.branch[31].block[14].um_I.iw[6] ,
    \top_I.branch[31].block[14].um_I.iw[5] ,
    \top_I.branch[31].block[14].um_I.iw[4] ,
    \top_I.branch[31].block[14].um_I.iw[3] ,
    \top_I.branch[31].block[14].um_I.iw[2] ,
    \top_I.branch[31].block[14].um_I.iw[1] ,
    \top_I.branch[31].block[14].um_I.clk ,
    \top_I.branch[31].block[13].um_I.iw[17] ,
    \top_I.branch[31].block[13].um_I.iw[16] ,
    \top_I.branch[31].block[13].um_I.iw[15] ,
    \top_I.branch[31].block[13].um_I.iw[14] ,
    \top_I.branch[31].block[13].um_I.iw[13] ,
    \top_I.branch[31].block[13].um_I.iw[12] ,
    \top_I.branch[31].block[13].um_I.iw[11] ,
    \top_I.branch[31].block[13].um_I.iw[10] ,
    \top_I.branch[31].block[13].um_I.iw[9] ,
    \top_I.branch[31].block[13].um_I.iw[8] ,
    \top_I.branch[31].block[13].um_I.iw[7] ,
    \top_I.branch[31].block[13].um_I.iw[6] ,
    \top_I.branch[31].block[13].um_I.iw[5] ,
    \top_I.branch[31].block[13].um_I.iw[4] ,
    \top_I.branch[31].block[13].um_I.iw[3] ,
    \top_I.branch[31].block[13].um_I.iw[2] ,
    \top_I.branch[31].block[13].um_I.iw[1] ,
    \top_I.branch[31].block[13].um_I.clk ,
    \top_I.branch[31].block[12].um_I.iw[17] ,
    \top_I.branch[31].block[12].um_I.iw[16] ,
    \top_I.branch[31].block[12].um_I.iw[15] ,
    \top_I.branch[31].block[12].um_I.iw[14] ,
    \top_I.branch[31].block[12].um_I.iw[13] ,
    \top_I.branch[31].block[12].um_I.iw[12] ,
    \top_I.branch[31].block[12].um_I.iw[11] ,
    \top_I.branch[31].block[12].um_I.iw[10] ,
    \top_I.branch[31].block[12].um_I.iw[9] ,
    \top_I.branch[31].block[12].um_I.iw[8] ,
    \top_I.branch[31].block[12].um_I.iw[7] ,
    \top_I.branch[31].block[12].um_I.iw[6] ,
    \top_I.branch[31].block[12].um_I.iw[5] ,
    \top_I.branch[31].block[12].um_I.iw[4] ,
    \top_I.branch[31].block[12].um_I.iw[3] ,
    \top_I.branch[31].block[12].um_I.iw[2] ,
    \top_I.branch[31].block[12].um_I.iw[1] ,
    \top_I.branch[31].block[12].um_I.clk ,
    \top_I.branch[31].block[11].um_I.iw[17] ,
    \top_I.branch[31].block[11].um_I.iw[16] ,
    \top_I.branch[31].block[11].um_I.iw[15] ,
    \top_I.branch[31].block[11].um_I.iw[14] ,
    \top_I.branch[31].block[11].um_I.iw[13] ,
    \top_I.branch[31].block[11].um_I.iw[12] ,
    \top_I.branch[31].block[11].um_I.iw[11] ,
    \top_I.branch[31].block[11].um_I.iw[10] ,
    \top_I.branch[31].block[11].um_I.iw[9] ,
    \top_I.branch[31].block[11].um_I.iw[8] ,
    \top_I.branch[31].block[11].um_I.iw[7] ,
    \top_I.branch[31].block[11].um_I.iw[6] ,
    \top_I.branch[31].block[11].um_I.iw[5] ,
    \top_I.branch[31].block[11].um_I.iw[4] ,
    \top_I.branch[31].block[11].um_I.iw[3] ,
    \top_I.branch[31].block[11].um_I.iw[2] ,
    \top_I.branch[31].block[11].um_I.iw[1] ,
    \top_I.branch[31].block[11].um_I.clk ,
    \top_I.branch[31].block[10].um_I.iw[17] ,
    \top_I.branch[31].block[10].um_I.iw[16] ,
    \top_I.branch[31].block[10].um_I.iw[15] ,
    \top_I.branch[31].block[10].um_I.iw[14] ,
    \top_I.branch[31].block[10].um_I.iw[13] ,
    \top_I.branch[31].block[10].um_I.iw[12] ,
    \top_I.branch[31].block[10].um_I.iw[11] ,
    \top_I.branch[31].block[10].um_I.iw[10] ,
    \top_I.branch[31].block[10].um_I.iw[9] ,
    \top_I.branch[31].block[10].um_I.iw[8] ,
    \top_I.branch[31].block[10].um_I.iw[7] ,
    \top_I.branch[31].block[10].um_I.iw[6] ,
    \top_I.branch[31].block[10].um_I.iw[5] ,
    \top_I.branch[31].block[10].um_I.iw[4] ,
    \top_I.branch[31].block[10].um_I.iw[3] ,
    \top_I.branch[31].block[10].um_I.iw[2] ,
    \top_I.branch[31].block[10].um_I.iw[1] ,
    \top_I.branch[31].block[10].um_I.clk ,
    \top_I.branch[31].block[9].um_I.iw[17] ,
    \top_I.branch[31].block[9].um_I.iw[16] ,
    \top_I.branch[31].block[9].um_I.iw[15] ,
    \top_I.branch[31].block[9].um_I.iw[14] ,
    \top_I.branch[31].block[9].um_I.iw[13] ,
    \top_I.branch[31].block[9].um_I.iw[12] ,
    \top_I.branch[31].block[9].um_I.iw[11] ,
    \top_I.branch[31].block[9].um_I.iw[10] ,
    \top_I.branch[31].block[9].um_I.iw[9] ,
    \top_I.branch[31].block[9].um_I.iw[8] ,
    \top_I.branch[31].block[9].um_I.iw[7] ,
    \top_I.branch[31].block[9].um_I.iw[6] ,
    \top_I.branch[31].block[9].um_I.iw[5] ,
    \top_I.branch[31].block[9].um_I.iw[4] ,
    \top_I.branch[31].block[9].um_I.iw[3] ,
    \top_I.branch[31].block[9].um_I.iw[2] ,
    \top_I.branch[31].block[9].um_I.iw[1] ,
    \top_I.branch[31].block[9].um_I.clk ,
    \top_I.branch[31].block[8].um_I.iw[17] ,
    \top_I.branch[31].block[8].um_I.iw[16] ,
    \top_I.branch[31].block[8].um_I.iw[15] ,
    \top_I.branch[31].block[8].um_I.iw[14] ,
    \top_I.branch[31].block[8].um_I.iw[13] ,
    \top_I.branch[31].block[8].um_I.iw[12] ,
    \top_I.branch[31].block[8].um_I.iw[11] ,
    \top_I.branch[31].block[8].um_I.iw[10] ,
    \top_I.branch[31].block[8].um_I.iw[9] ,
    \top_I.branch[31].block[8].um_I.iw[8] ,
    \top_I.branch[31].block[8].um_I.iw[7] ,
    \top_I.branch[31].block[8].um_I.iw[6] ,
    \top_I.branch[31].block[8].um_I.iw[5] ,
    \top_I.branch[31].block[8].um_I.iw[4] ,
    \top_I.branch[31].block[8].um_I.iw[3] ,
    \top_I.branch[31].block[8].um_I.iw[2] ,
    \top_I.branch[31].block[8].um_I.iw[1] ,
    \top_I.branch[31].block[8].um_I.clk ,
    \top_I.branch[31].block[7].um_I.iw[17] ,
    \top_I.branch[31].block[7].um_I.iw[16] ,
    \top_I.branch[31].block[7].um_I.iw[15] ,
    \top_I.branch[31].block[7].um_I.iw[14] ,
    \top_I.branch[31].block[7].um_I.iw[13] ,
    \top_I.branch[31].block[7].um_I.iw[12] ,
    \top_I.branch[31].block[7].um_I.iw[11] ,
    \top_I.branch[31].block[7].um_I.iw[10] ,
    \top_I.branch[31].block[7].um_I.iw[9] ,
    \top_I.branch[31].block[7].um_I.iw[8] ,
    \top_I.branch[31].block[7].um_I.iw[7] ,
    \top_I.branch[31].block[7].um_I.iw[6] ,
    \top_I.branch[31].block[7].um_I.iw[5] ,
    \top_I.branch[31].block[7].um_I.iw[4] ,
    \top_I.branch[31].block[7].um_I.iw[3] ,
    \top_I.branch[31].block[7].um_I.iw[2] ,
    \top_I.branch[31].block[7].um_I.iw[1] ,
    \top_I.branch[31].block[7].um_I.clk ,
    \top_I.branch[31].block[6].um_I.iw[17] ,
    \top_I.branch[31].block[6].um_I.iw[16] ,
    \top_I.branch[31].block[6].um_I.iw[15] ,
    \top_I.branch[31].block[6].um_I.iw[14] ,
    \top_I.branch[31].block[6].um_I.iw[13] ,
    \top_I.branch[31].block[6].um_I.iw[12] ,
    \top_I.branch[31].block[6].um_I.iw[11] ,
    \top_I.branch[31].block[6].um_I.iw[10] ,
    \top_I.branch[31].block[6].um_I.iw[9] ,
    \top_I.branch[31].block[6].um_I.iw[8] ,
    \top_I.branch[31].block[6].um_I.iw[7] ,
    \top_I.branch[31].block[6].um_I.iw[6] ,
    \top_I.branch[31].block[6].um_I.iw[5] ,
    \top_I.branch[31].block[6].um_I.iw[4] ,
    \top_I.branch[31].block[6].um_I.iw[3] ,
    \top_I.branch[31].block[6].um_I.iw[2] ,
    \top_I.branch[31].block[6].um_I.iw[1] ,
    \top_I.branch[31].block[6].um_I.clk ,
    \top_I.branch[31].block[5].um_I.iw[17] ,
    \top_I.branch[31].block[5].um_I.iw[16] ,
    \top_I.branch[31].block[5].um_I.iw[15] ,
    \top_I.branch[31].block[5].um_I.iw[14] ,
    \top_I.branch[31].block[5].um_I.iw[13] ,
    \top_I.branch[31].block[5].um_I.iw[12] ,
    \top_I.branch[31].block[5].um_I.iw[11] ,
    \top_I.branch[31].block[5].um_I.iw[10] ,
    \top_I.branch[31].block[5].um_I.iw[9] ,
    \top_I.branch[31].block[5].um_I.iw[8] ,
    \top_I.branch[31].block[5].um_I.iw[7] ,
    \top_I.branch[31].block[5].um_I.iw[6] ,
    \top_I.branch[31].block[5].um_I.iw[5] ,
    \top_I.branch[31].block[5].um_I.iw[4] ,
    \top_I.branch[31].block[5].um_I.iw[3] ,
    \top_I.branch[31].block[5].um_I.iw[2] ,
    \top_I.branch[31].block[5].um_I.iw[1] ,
    \top_I.branch[31].block[5].um_I.clk ,
    \top_I.branch[31].block[4].um_I.iw[17] ,
    \top_I.branch[31].block[4].um_I.iw[16] ,
    \top_I.branch[31].block[4].um_I.iw[15] ,
    \top_I.branch[31].block[4].um_I.iw[14] ,
    \top_I.branch[31].block[4].um_I.iw[13] ,
    \top_I.branch[31].block[4].um_I.iw[12] ,
    \top_I.branch[31].block[4].um_I.iw[11] ,
    \top_I.branch[31].block[4].um_I.iw[10] ,
    \top_I.branch[31].block[4].um_I.iw[9] ,
    \top_I.branch[31].block[4].um_I.iw[8] ,
    \top_I.branch[31].block[4].um_I.iw[7] ,
    \top_I.branch[31].block[4].um_I.iw[6] ,
    \top_I.branch[31].block[4].um_I.iw[5] ,
    \top_I.branch[31].block[4].um_I.iw[4] ,
    \top_I.branch[31].block[4].um_I.iw[3] ,
    \top_I.branch[31].block[4].um_I.iw[2] ,
    \top_I.branch[31].block[4].um_I.iw[1] ,
    \top_I.branch[31].block[4].um_I.clk ,
    \top_I.branch[31].block[3].um_I.iw[17] ,
    \top_I.branch[31].block[3].um_I.iw[16] ,
    \top_I.branch[31].block[3].um_I.iw[15] ,
    \top_I.branch[31].block[3].um_I.iw[14] ,
    \top_I.branch[31].block[3].um_I.iw[13] ,
    \top_I.branch[31].block[3].um_I.iw[12] ,
    \top_I.branch[31].block[3].um_I.iw[11] ,
    \top_I.branch[31].block[3].um_I.iw[10] ,
    \top_I.branch[31].block[3].um_I.iw[9] ,
    \top_I.branch[31].block[3].um_I.iw[8] ,
    \top_I.branch[31].block[3].um_I.iw[7] ,
    \top_I.branch[31].block[3].um_I.iw[6] ,
    \top_I.branch[31].block[3].um_I.iw[5] ,
    \top_I.branch[31].block[3].um_I.iw[4] ,
    \top_I.branch[31].block[3].um_I.iw[3] ,
    \top_I.branch[31].block[3].um_I.iw[2] ,
    \top_I.branch[31].block[3].um_I.iw[1] ,
    \top_I.branch[31].block[3].um_I.clk ,
    \top_I.branch[31].block[2].um_I.iw[17] ,
    \top_I.branch[31].block[2].um_I.iw[16] ,
    \top_I.branch[31].block[2].um_I.iw[15] ,
    \top_I.branch[31].block[2].um_I.iw[14] ,
    \top_I.branch[31].block[2].um_I.iw[13] ,
    \top_I.branch[31].block[2].um_I.iw[12] ,
    \top_I.branch[31].block[2].um_I.iw[11] ,
    \top_I.branch[31].block[2].um_I.iw[10] ,
    \top_I.branch[31].block[2].um_I.iw[9] ,
    \top_I.branch[31].block[2].um_I.iw[8] ,
    \top_I.branch[31].block[2].um_I.iw[7] ,
    \top_I.branch[31].block[2].um_I.iw[6] ,
    \top_I.branch[31].block[2].um_I.iw[5] ,
    \top_I.branch[31].block[2].um_I.iw[4] ,
    \top_I.branch[31].block[2].um_I.iw[3] ,
    \top_I.branch[31].block[2].um_I.iw[2] ,
    \top_I.branch[31].block[2].um_I.iw[1] ,
    \top_I.branch[31].block[2].um_I.clk ,
    \top_I.branch[31].block[1].um_I.iw[17] ,
    \top_I.branch[31].block[1].um_I.iw[16] ,
    \top_I.branch[31].block[1].um_I.iw[15] ,
    \top_I.branch[31].block[1].um_I.iw[14] ,
    \top_I.branch[31].block[1].um_I.iw[13] ,
    \top_I.branch[31].block[1].um_I.iw[12] ,
    \top_I.branch[31].block[1].um_I.iw[11] ,
    \top_I.branch[31].block[1].um_I.iw[10] ,
    \top_I.branch[31].block[1].um_I.iw[9] ,
    \top_I.branch[31].block[1].um_I.iw[8] ,
    \top_I.branch[31].block[1].um_I.iw[7] ,
    \top_I.branch[31].block[1].um_I.iw[6] ,
    \top_I.branch[31].block[1].um_I.iw[5] ,
    \top_I.branch[31].block[1].um_I.iw[4] ,
    \top_I.branch[31].block[1].um_I.iw[3] ,
    \top_I.branch[31].block[1].um_I.iw[2] ,
    \top_I.branch[31].block[1].um_I.iw[1] ,
    \top_I.branch[31].block[1].um_I.clk ,
    \top_I.branch[31].block[0].um_I.iw[17] ,
    \top_I.branch[31].block[0].um_I.iw[16] ,
    \top_I.branch[31].block[0].um_I.iw[15] ,
    \top_I.branch[31].block[0].um_I.iw[14] ,
    \top_I.branch[31].block[0].um_I.iw[13] ,
    \top_I.branch[31].block[0].um_I.iw[12] ,
    \top_I.branch[31].block[0].um_I.iw[11] ,
    \top_I.branch[31].block[0].um_I.iw[10] ,
    \top_I.branch[31].block[0].um_I.iw[9] ,
    \top_I.branch[31].block[0].um_I.iw[8] ,
    \top_I.branch[31].block[0].um_I.iw[7] ,
    \top_I.branch[31].block[0].um_I.iw[6] ,
    \top_I.branch[31].block[0].um_I.iw[5] ,
    \top_I.branch[31].block[0].um_I.iw[4] ,
    \top_I.branch[31].block[0].um_I.iw[3] ,
    \top_I.branch[31].block[0].um_I.iw[2] ,
    \top_I.branch[31].block[0].um_I.iw[1] ,
    \top_I.branch[31].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[15].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[14].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[13].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[12].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[11].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[10].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[9].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[8].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[7].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[6].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[5].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[4].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[3].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[2].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[1].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero ,
    \top_I.branch[31].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[31].block[15].um_I.pg_vdd ,
    \top_I.branch[31].block[14].um_I.pg_vdd ,
    \top_I.branch[31].block[13].um_I.pg_vdd ,
    \top_I.branch[31].block[12].um_I.pg_vdd ,
    \top_I.branch[31].block[11].um_I.pg_vdd ,
    \top_I.branch[31].block[10].um_I.pg_vdd ,
    \top_I.branch[31].block[9].um_I.pg_vdd ,
    \top_I.branch[31].block[8].um_I.pg_vdd ,
    \top_I.branch[31].block[7].um_I.pg_vdd ,
    \top_I.branch[31].block[6].um_I.pg_vdd ,
    \top_I.branch[31].block[5].um_I.pg_vdd ,
    \top_I.branch[31].block[4].um_I.pg_vdd ,
    \top_I.branch[31].block[3].um_I.pg_vdd ,
    \top_I.branch[31].block[2].um_I.pg_vdd ,
    \top_I.branch[31].block[1].um_I.pg_vdd ,
    \top_I.branch[31].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[3].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[3].l_addr[0] ),
    .k_zero(\top_I.branch[3].l_addr[1] ),
    .addr({\top_I.branch[3].l_addr[1] ,
    \top_I.branch[3].l_addr[1] ,
    \top_I.branch[3].l_addr[1] ,
    \top_I.branch[3].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[3].block[15].um_I.ena ,
    \top_I.branch[3].block[14].um_I.ena ,
    \top_I.branch[3].block[13].um_I.ena ,
    \top_I.branch[3].block[12].um_I.ena ,
    \top_I.branch[3].block[11].um_I.ena ,
    \top_I.branch[3].block[10].um_I.ena ,
    \top_I.branch[3].block[9].um_I.ena ,
    \top_I.branch[3].block[8].um_I.ena ,
    \top_I.branch[3].block[7].um_I.ena ,
    \top_I.branch[3].block[6].um_I.ena ,
    \top_I.branch[3].block[5].um_I.ena ,
    \top_I.branch[3].block[4].um_I.ena ,
    \top_I.branch[3].block[3].um_I.ena ,
    \top_I.branch[3].block[2].um_I.ena ,
    \top_I.branch[3].block[1].um_I.ena ,
    \top_I.branch[3].block[0].um_I.ena }),
    .um_iw({\top_I.branch[3].block[15].um_I.iw[17] ,
    \top_I.branch[3].block[15].um_I.iw[16] ,
    \top_I.branch[3].block[15].um_I.iw[15] ,
    \top_I.branch[3].block[15].um_I.iw[14] ,
    \top_I.branch[3].block[15].um_I.iw[13] ,
    \top_I.branch[3].block[15].um_I.iw[12] ,
    \top_I.branch[3].block[15].um_I.iw[11] ,
    \top_I.branch[3].block[15].um_I.iw[10] ,
    \top_I.branch[3].block[15].um_I.iw[9] ,
    \top_I.branch[3].block[15].um_I.iw[8] ,
    \top_I.branch[3].block[15].um_I.iw[7] ,
    \top_I.branch[3].block[15].um_I.iw[6] ,
    \top_I.branch[3].block[15].um_I.iw[5] ,
    \top_I.branch[3].block[15].um_I.iw[4] ,
    \top_I.branch[3].block[15].um_I.iw[3] ,
    \top_I.branch[3].block[15].um_I.iw[2] ,
    \top_I.branch[3].block[15].um_I.iw[1] ,
    \top_I.branch[3].block[15].um_I.clk ,
    \top_I.branch[3].block[14].um_I.iw[17] ,
    \top_I.branch[3].block[14].um_I.iw[16] ,
    \top_I.branch[3].block[14].um_I.iw[15] ,
    \top_I.branch[3].block[14].um_I.iw[14] ,
    \top_I.branch[3].block[14].um_I.iw[13] ,
    \top_I.branch[3].block[14].um_I.iw[12] ,
    \top_I.branch[3].block[14].um_I.iw[11] ,
    \top_I.branch[3].block[14].um_I.iw[10] ,
    \top_I.branch[3].block[14].um_I.iw[9] ,
    \top_I.branch[3].block[14].um_I.iw[8] ,
    \top_I.branch[3].block[14].um_I.iw[7] ,
    \top_I.branch[3].block[14].um_I.iw[6] ,
    \top_I.branch[3].block[14].um_I.iw[5] ,
    \top_I.branch[3].block[14].um_I.iw[4] ,
    \top_I.branch[3].block[14].um_I.iw[3] ,
    \top_I.branch[3].block[14].um_I.iw[2] ,
    \top_I.branch[3].block[14].um_I.iw[1] ,
    \top_I.branch[3].block[14].um_I.clk ,
    \top_I.branch[3].block[13].um_I.iw[17] ,
    \top_I.branch[3].block[13].um_I.iw[16] ,
    \top_I.branch[3].block[13].um_I.iw[15] ,
    \top_I.branch[3].block[13].um_I.iw[14] ,
    \top_I.branch[3].block[13].um_I.iw[13] ,
    \top_I.branch[3].block[13].um_I.iw[12] ,
    \top_I.branch[3].block[13].um_I.iw[11] ,
    \top_I.branch[3].block[13].um_I.iw[10] ,
    \top_I.branch[3].block[13].um_I.iw[9] ,
    \top_I.branch[3].block[13].um_I.iw[8] ,
    \top_I.branch[3].block[13].um_I.iw[7] ,
    \top_I.branch[3].block[13].um_I.iw[6] ,
    \top_I.branch[3].block[13].um_I.iw[5] ,
    \top_I.branch[3].block[13].um_I.iw[4] ,
    \top_I.branch[3].block[13].um_I.iw[3] ,
    \top_I.branch[3].block[13].um_I.iw[2] ,
    \top_I.branch[3].block[13].um_I.iw[1] ,
    \top_I.branch[3].block[13].um_I.clk ,
    \top_I.branch[3].block[12].um_I.iw[17] ,
    \top_I.branch[3].block[12].um_I.iw[16] ,
    \top_I.branch[3].block[12].um_I.iw[15] ,
    \top_I.branch[3].block[12].um_I.iw[14] ,
    \top_I.branch[3].block[12].um_I.iw[13] ,
    \top_I.branch[3].block[12].um_I.iw[12] ,
    \top_I.branch[3].block[12].um_I.iw[11] ,
    \top_I.branch[3].block[12].um_I.iw[10] ,
    \top_I.branch[3].block[12].um_I.iw[9] ,
    \top_I.branch[3].block[12].um_I.iw[8] ,
    \top_I.branch[3].block[12].um_I.iw[7] ,
    \top_I.branch[3].block[12].um_I.iw[6] ,
    \top_I.branch[3].block[12].um_I.iw[5] ,
    \top_I.branch[3].block[12].um_I.iw[4] ,
    \top_I.branch[3].block[12].um_I.iw[3] ,
    \top_I.branch[3].block[12].um_I.iw[2] ,
    \top_I.branch[3].block[12].um_I.iw[1] ,
    \top_I.branch[3].block[12].um_I.clk ,
    \top_I.branch[3].block[11].um_I.iw[17] ,
    \top_I.branch[3].block[11].um_I.iw[16] ,
    \top_I.branch[3].block[11].um_I.iw[15] ,
    \top_I.branch[3].block[11].um_I.iw[14] ,
    \top_I.branch[3].block[11].um_I.iw[13] ,
    \top_I.branch[3].block[11].um_I.iw[12] ,
    \top_I.branch[3].block[11].um_I.iw[11] ,
    \top_I.branch[3].block[11].um_I.iw[10] ,
    \top_I.branch[3].block[11].um_I.iw[9] ,
    \top_I.branch[3].block[11].um_I.iw[8] ,
    \top_I.branch[3].block[11].um_I.iw[7] ,
    \top_I.branch[3].block[11].um_I.iw[6] ,
    \top_I.branch[3].block[11].um_I.iw[5] ,
    \top_I.branch[3].block[11].um_I.iw[4] ,
    \top_I.branch[3].block[11].um_I.iw[3] ,
    \top_I.branch[3].block[11].um_I.iw[2] ,
    \top_I.branch[3].block[11].um_I.iw[1] ,
    \top_I.branch[3].block[11].um_I.clk ,
    \top_I.branch[3].block[10].um_I.iw[17] ,
    \top_I.branch[3].block[10].um_I.iw[16] ,
    \top_I.branch[3].block[10].um_I.iw[15] ,
    \top_I.branch[3].block[10].um_I.iw[14] ,
    \top_I.branch[3].block[10].um_I.iw[13] ,
    \top_I.branch[3].block[10].um_I.iw[12] ,
    \top_I.branch[3].block[10].um_I.iw[11] ,
    \top_I.branch[3].block[10].um_I.iw[10] ,
    \top_I.branch[3].block[10].um_I.iw[9] ,
    \top_I.branch[3].block[10].um_I.iw[8] ,
    \top_I.branch[3].block[10].um_I.iw[7] ,
    \top_I.branch[3].block[10].um_I.iw[6] ,
    \top_I.branch[3].block[10].um_I.iw[5] ,
    \top_I.branch[3].block[10].um_I.iw[4] ,
    \top_I.branch[3].block[10].um_I.iw[3] ,
    \top_I.branch[3].block[10].um_I.iw[2] ,
    \top_I.branch[3].block[10].um_I.iw[1] ,
    \top_I.branch[3].block[10].um_I.clk ,
    \top_I.branch[3].block[9].um_I.iw[17] ,
    \top_I.branch[3].block[9].um_I.iw[16] ,
    \top_I.branch[3].block[9].um_I.iw[15] ,
    \top_I.branch[3].block[9].um_I.iw[14] ,
    \top_I.branch[3].block[9].um_I.iw[13] ,
    \top_I.branch[3].block[9].um_I.iw[12] ,
    \top_I.branch[3].block[9].um_I.iw[11] ,
    \top_I.branch[3].block[9].um_I.iw[10] ,
    \top_I.branch[3].block[9].um_I.iw[9] ,
    \top_I.branch[3].block[9].um_I.iw[8] ,
    \top_I.branch[3].block[9].um_I.iw[7] ,
    \top_I.branch[3].block[9].um_I.iw[6] ,
    \top_I.branch[3].block[9].um_I.iw[5] ,
    \top_I.branch[3].block[9].um_I.iw[4] ,
    \top_I.branch[3].block[9].um_I.iw[3] ,
    \top_I.branch[3].block[9].um_I.iw[2] ,
    \top_I.branch[3].block[9].um_I.iw[1] ,
    \top_I.branch[3].block[9].um_I.clk ,
    \top_I.branch[3].block[8].um_I.iw[17] ,
    \top_I.branch[3].block[8].um_I.iw[16] ,
    \top_I.branch[3].block[8].um_I.iw[15] ,
    \top_I.branch[3].block[8].um_I.iw[14] ,
    \top_I.branch[3].block[8].um_I.iw[13] ,
    \top_I.branch[3].block[8].um_I.iw[12] ,
    \top_I.branch[3].block[8].um_I.iw[11] ,
    \top_I.branch[3].block[8].um_I.iw[10] ,
    \top_I.branch[3].block[8].um_I.iw[9] ,
    \top_I.branch[3].block[8].um_I.iw[8] ,
    \top_I.branch[3].block[8].um_I.iw[7] ,
    \top_I.branch[3].block[8].um_I.iw[6] ,
    \top_I.branch[3].block[8].um_I.iw[5] ,
    \top_I.branch[3].block[8].um_I.iw[4] ,
    \top_I.branch[3].block[8].um_I.iw[3] ,
    \top_I.branch[3].block[8].um_I.iw[2] ,
    \top_I.branch[3].block[8].um_I.iw[1] ,
    \top_I.branch[3].block[8].um_I.clk ,
    \top_I.branch[3].block[7].um_I.iw[17] ,
    \top_I.branch[3].block[7].um_I.iw[16] ,
    \top_I.branch[3].block[7].um_I.iw[15] ,
    \top_I.branch[3].block[7].um_I.iw[14] ,
    \top_I.branch[3].block[7].um_I.iw[13] ,
    \top_I.branch[3].block[7].um_I.iw[12] ,
    \top_I.branch[3].block[7].um_I.iw[11] ,
    \top_I.branch[3].block[7].um_I.iw[10] ,
    \top_I.branch[3].block[7].um_I.iw[9] ,
    \top_I.branch[3].block[7].um_I.iw[8] ,
    \top_I.branch[3].block[7].um_I.iw[7] ,
    \top_I.branch[3].block[7].um_I.iw[6] ,
    \top_I.branch[3].block[7].um_I.iw[5] ,
    \top_I.branch[3].block[7].um_I.iw[4] ,
    \top_I.branch[3].block[7].um_I.iw[3] ,
    \top_I.branch[3].block[7].um_I.iw[2] ,
    \top_I.branch[3].block[7].um_I.iw[1] ,
    \top_I.branch[3].block[7].um_I.clk ,
    \top_I.branch[3].block[6].um_I.iw[17] ,
    \top_I.branch[3].block[6].um_I.iw[16] ,
    \top_I.branch[3].block[6].um_I.iw[15] ,
    \top_I.branch[3].block[6].um_I.iw[14] ,
    \top_I.branch[3].block[6].um_I.iw[13] ,
    \top_I.branch[3].block[6].um_I.iw[12] ,
    \top_I.branch[3].block[6].um_I.iw[11] ,
    \top_I.branch[3].block[6].um_I.iw[10] ,
    \top_I.branch[3].block[6].um_I.iw[9] ,
    \top_I.branch[3].block[6].um_I.iw[8] ,
    \top_I.branch[3].block[6].um_I.iw[7] ,
    \top_I.branch[3].block[6].um_I.iw[6] ,
    \top_I.branch[3].block[6].um_I.iw[5] ,
    \top_I.branch[3].block[6].um_I.iw[4] ,
    \top_I.branch[3].block[6].um_I.iw[3] ,
    \top_I.branch[3].block[6].um_I.iw[2] ,
    \top_I.branch[3].block[6].um_I.iw[1] ,
    \top_I.branch[3].block[6].um_I.clk ,
    \top_I.branch[3].block[5].um_I.iw[17] ,
    \top_I.branch[3].block[5].um_I.iw[16] ,
    \top_I.branch[3].block[5].um_I.iw[15] ,
    \top_I.branch[3].block[5].um_I.iw[14] ,
    \top_I.branch[3].block[5].um_I.iw[13] ,
    \top_I.branch[3].block[5].um_I.iw[12] ,
    \top_I.branch[3].block[5].um_I.iw[11] ,
    \top_I.branch[3].block[5].um_I.iw[10] ,
    \top_I.branch[3].block[5].um_I.iw[9] ,
    \top_I.branch[3].block[5].um_I.iw[8] ,
    \top_I.branch[3].block[5].um_I.iw[7] ,
    \top_I.branch[3].block[5].um_I.iw[6] ,
    \top_I.branch[3].block[5].um_I.iw[5] ,
    \top_I.branch[3].block[5].um_I.iw[4] ,
    \top_I.branch[3].block[5].um_I.iw[3] ,
    \top_I.branch[3].block[5].um_I.iw[2] ,
    \top_I.branch[3].block[5].um_I.iw[1] ,
    \top_I.branch[3].block[5].um_I.clk ,
    \top_I.branch[3].block[4].um_I.iw[17] ,
    \top_I.branch[3].block[4].um_I.iw[16] ,
    \top_I.branch[3].block[4].um_I.iw[15] ,
    \top_I.branch[3].block[4].um_I.iw[14] ,
    \top_I.branch[3].block[4].um_I.iw[13] ,
    \top_I.branch[3].block[4].um_I.iw[12] ,
    \top_I.branch[3].block[4].um_I.iw[11] ,
    \top_I.branch[3].block[4].um_I.iw[10] ,
    \top_I.branch[3].block[4].um_I.iw[9] ,
    \top_I.branch[3].block[4].um_I.iw[8] ,
    \top_I.branch[3].block[4].um_I.iw[7] ,
    \top_I.branch[3].block[4].um_I.iw[6] ,
    \top_I.branch[3].block[4].um_I.iw[5] ,
    \top_I.branch[3].block[4].um_I.iw[4] ,
    \top_I.branch[3].block[4].um_I.iw[3] ,
    \top_I.branch[3].block[4].um_I.iw[2] ,
    \top_I.branch[3].block[4].um_I.iw[1] ,
    \top_I.branch[3].block[4].um_I.clk ,
    \top_I.branch[3].block[3].um_I.iw[17] ,
    \top_I.branch[3].block[3].um_I.iw[16] ,
    \top_I.branch[3].block[3].um_I.iw[15] ,
    \top_I.branch[3].block[3].um_I.iw[14] ,
    \top_I.branch[3].block[3].um_I.iw[13] ,
    \top_I.branch[3].block[3].um_I.iw[12] ,
    \top_I.branch[3].block[3].um_I.iw[11] ,
    \top_I.branch[3].block[3].um_I.iw[10] ,
    \top_I.branch[3].block[3].um_I.iw[9] ,
    \top_I.branch[3].block[3].um_I.iw[8] ,
    \top_I.branch[3].block[3].um_I.iw[7] ,
    \top_I.branch[3].block[3].um_I.iw[6] ,
    \top_I.branch[3].block[3].um_I.iw[5] ,
    \top_I.branch[3].block[3].um_I.iw[4] ,
    \top_I.branch[3].block[3].um_I.iw[3] ,
    \top_I.branch[3].block[3].um_I.iw[2] ,
    \top_I.branch[3].block[3].um_I.iw[1] ,
    \top_I.branch[3].block[3].um_I.clk ,
    \top_I.branch[3].block[2].um_I.iw[17] ,
    \top_I.branch[3].block[2].um_I.iw[16] ,
    \top_I.branch[3].block[2].um_I.iw[15] ,
    \top_I.branch[3].block[2].um_I.iw[14] ,
    \top_I.branch[3].block[2].um_I.iw[13] ,
    \top_I.branch[3].block[2].um_I.iw[12] ,
    \top_I.branch[3].block[2].um_I.iw[11] ,
    \top_I.branch[3].block[2].um_I.iw[10] ,
    \top_I.branch[3].block[2].um_I.iw[9] ,
    \top_I.branch[3].block[2].um_I.iw[8] ,
    \top_I.branch[3].block[2].um_I.iw[7] ,
    \top_I.branch[3].block[2].um_I.iw[6] ,
    \top_I.branch[3].block[2].um_I.iw[5] ,
    \top_I.branch[3].block[2].um_I.iw[4] ,
    \top_I.branch[3].block[2].um_I.iw[3] ,
    \top_I.branch[3].block[2].um_I.iw[2] ,
    \top_I.branch[3].block[2].um_I.iw[1] ,
    \top_I.branch[3].block[2].um_I.clk ,
    \top_I.branch[3].block[1].um_I.iw[17] ,
    \top_I.branch[3].block[1].um_I.iw[16] ,
    \top_I.branch[3].block[1].um_I.iw[15] ,
    \top_I.branch[3].block[1].um_I.iw[14] ,
    \top_I.branch[3].block[1].um_I.iw[13] ,
    \top_I.branch[3].block[1].um_I.iw[12] ,
    \top_I.branch[3].block[1].um_I.iw[11] ,
    \top_I.branch[3].block[1].um_I.iw[10] ,
    \top_I.branch[3].block[1].um_I.iw[9] ,
    \top_I.branch[3].block[1].um_I.iw[8] ,
    \top_I.branch[3].block[1].um_I.iw[7] ,
    \top_I.branch[3].block[1].um_I.iw[6] ,
    \top_I.branch[3].block[1].um_I.iw[5] ,
    \top_I.branch[3].block[1].um_I.iw[4] ,
    \top_I.branch[3].block[1].um_I.iw[3] ,
    \top_I.branch[3].block[1].um_I.iw[2] ,
    \top_I.branch[3].block[1].um_I.iw[1] ,
    \top_I.branch[3].block[1].um_I.clk ,
    \top_I.branch[3].block[0].um_I.iw[17] ,
    \top_I.branch[3].block[0].um_I.iw[16] ,
    \top_I.branch[3].block[0].um_I.iw[15] ,
    \top_I.branch[3].block[0].um_I.iw[14] ,
    \top_I.branch[3].block[0].um_I.iw[13] ,
    \top_I.branch[3].block[0].um_I.iw[12] ,
    \top_I.branch[3].block[0].um_I.iw[11] ,
    \top_I.branch[3].block[0].um_I.iw[10] ,
    \top_I.branch[3].block[0].um_I.iw[9] ,
    \top_I.branch[3].block[0].um_I.iw[8] ,
    \top_I.branch[3].block[0].um_I.iw[7] ,
    \top_I.branch[3].block[0].um_I.iw[6] ,
    \top_I.branch[3].block[0].um_I.iw[5] ,
    \top_I.branch[3].block[0].um_I.iw[4] ,
    \top_I.branch[3].block[0].um_I.iw[3] ,
    \top_I.branch[3].block[0].um_I.iw[2] ,
    \top_I.branch[3].block[0].um_I.iw[1] ,
    \top_I.branch[3].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[15].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[14].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[13].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[12].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[11].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[10].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[9].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[8].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[7].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[6].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[5].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[4].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[3].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[2].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[1].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero ,
    \top_I.branch[3].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[3].block[15].um_I.pg_vdd ,
    \top_I.branch[3].block[14].um_I.pg_vdd ,
    \top_I.branch[3].block[13].um_I.pg_vdd ,
    \top_I.branch[3].block[12].um_I.pg_vdd ,
    \top_I.branch[3].block[11].um_I.pg_vdd ,
    \top_I.branch[3].block[10].um_I.pg_vdd ,
    \top_I.branch[3].block[9].um_I.pg_vdd ,
    \top_I.branch[3].block[8].um_I.pg_vdd ,
    \top_I.branch[3].block[7].um_I.pg_vdd ,
    \top_I.branch[3].block[6].um_I.pg_vdd ,
    \top_I.branch[3].block[5].um_I.pg_vdd ,
    \top_I.branch[3].block[4].um_I.pg_vdd ,
    \top_I.branch[3].block[3].um_I.pg_vdd ,
    \top_I.branch[3].block[2].um_I.pg_vdd ,
    \top_I.branch[3].block[1].um_I.pg_vdd ,
    \top_I.branch[3].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[4].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[4].l_addr[1] ),
    .k_zero(\top_I.branch[4].l_addr[0] ),
    .addr({\top_I.branch[4].l_addr[0] ,
    \top_I.branch[4].l_addr[0] ,
    \top_I.branch[4].l_addr[1] ,
    \top_I.branch[4].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[4].block[15].um_I.ena ,
    \top_I.branch[4].block[14].um_I.ena ,
    \top_I.branch[4].block[13].um_I.ena ,
    \top_I.branch[4].block[12].um_I.ena ,
    \top_I.branch[4].block[11].um_I.ena ,
    \top_I.branch[4].block[10].um_I.ena ,
    \top_I.branch[4].block[9].um_I.ena ,
    \top_I.branch[4].block[8].um_I.ena ,
    \top_I.branch[4].block[7].um_I.ena ,
    \top_I.branch[4].block[6].um_I.ena ,
    \top_I.branch[4].block[5].um_I.ena ,
    \top_I.branch[4].block[4].um_I.ena ,
    \top_I.branch[4].block[3].um_I.ena ,
    \top_I.branch[4].block[2].um_I.ena ,
    \top_I.branch[4].block[1].um_I.ena ,
    \top_I.branch[4].block[0].um_I.ena }),
    .um_iw({\top_I.branch[4].block[15].um_I.iw[17] ,
    \top_I.branch[4].block[15].um_I.iw[16] ,
    \top_I.branch[4].block[15].um_I.iw[15] ,
    \top_I.branch[4].block[15].um_I.iw[14] ,
    \top_I.branch[4].block[15].um_I.iw[13] ,
    \top_I.branch[4].block[15].um_I.iw[12] ,
    \top_I.branch[4].block[15].um_I.iw[11] ,
    \top_I.branch[4].block[15].um_I.iw[10] ,
    \top_I.branch[4].block[15].um_I.iw[9] ,
    \top_I.branch[4].block[15].um_I.iw[8] ,
    \top_I.branch[4].block[15].um_I.iw[7] ,
    \top_I.branch[4].block[15].um_I.iw[6] ,
    \top_I.branch[4].block[15].um_I.iw[5] ,
    \top_I.branch[4].block[15].um_I.iw[4] ,
    \top_I.branch[4].block[15].um_I.iw[3] ,
    \top_I.branch[4].block[15].um_I.iw[2] ,
    \top_I.branch[4].block[15].um_I.iw[1] ,
    \top_I.branch[4].block[15].um_I.clk ,
    \top_I.branch[4].block[14].um_I.iw[17] ,
    \top_I.branch[4].block[14].um_I.iw[16] ,
    \top_I.branch[4].block[14].um_I.iw[15] ,
    \top_I.branch[4].block[14].um_I.iw[14] ,
    \top_I.branch[4].block[14].um_I.iw[13] ,
    \top_I.branch[4].block[14].um_I.iw[12] ,
    \top_I.branch[4].block[14].um_I.iw[11] ,
    \top_I.branch[4].block[14].um_I.iw[10] ,
    \top_I.branch[4].block[14].um_I.iw[9] ,
    \top_I.branch[4].block[14].um_I.iw[8] ,
    \top_I.branch[4].block[14].um_I.iw[7] ,
    \top_I.branch[4].block[14].um_I.iw[6] ,
    \top_I.branch[4].block[14].um_I.iw[5] ,
    \top_I.branch[4].block[14].um_I.iw[4] ,
    \top_I.branch[4].block[14].um_I.iw[3] ,
    \top_I.branch[4].block[14].um_I.iw[2] ,
    \top_I.branch[4].block[14].um_I.iw[1] ,
    \top_I.branch[4].block[14].um_I.clk ,
    \top_I.branch[4].block[13].um_I.iw[17] ,
    \top_I.branch[4].block[13].um_I.iw[16] ,
    \top_I.branch[4].block[13].um_I.iw[15] ,
    \top_I.branch[4].block[13].um_I.iw[14] ,
    \top_I.branch[4].block[13].um_I.iw[13] ,
    \top_I.branch[4].block[13].um_I.iw[12] ,
    \top_I.branch[4].block[13].um_I.iw[11] ,
    \top_I.branch[4].block[13].um_I.iw[10] ,
    \top_I.branch[4].block[13].um_I.iw[9] ,
    \top_I.branch[4].block[13].um_I.iw[8] ,
    \top_I.branch[4].block[13].um_I.iw[7] ,
    \top_I.branch[4].block[13].um_I.iw[6] ,
    \top_I.branch[4].block[13].um_I.iw[5] ,
    \top_I.branch[4].block[13].um_I.iw[4] ,
    \top_I.branch[4].block[13].um_I.iw[3] ,
    \top_I.branch[4].block[13].um_I.iw[2] ,
    \top_I.branch[4].block[13].um_I.iw[1] ,
    \top_I.branch[4].block[13].um_I.clk ,
    \top_I.branch[4].block[12].um_I.iw[17] ,
    \top_I.branch[4].block[12].um_I.iw[16] ,
    \top_I.branch[4].block[12].um_I.iw[15] ,
    \top_I.branch[4].block[12].um_I.iw[14] ,
    \top_I.branch[4].block[12].um_I.iw[13] ,
    \top_I.branch[4].block[12].um_I.iw[12] ,
    \top_I.branch[4].block[12].um_I.iw[11] ,
    \top_I.branch[4].block[12].um_I.iw[10] ,
    \top_I.branch[4].block[12].um_I.iw[9] ,
    \top_I.branch[4].block[12].um_I.iw[8] ,
    \top_I.branch[4].block[12].um_I.iw[7] ,
    \top_I.branch[4].block[12].um_I.iw[6] ,
    \top_I.branch[4].block[12].um_I.iw[5] ,
    \top_I.branch[4].block[12].um_I.iw[4] ,
    \top_I.branch[4].block[12].um_I.iw[3] ,
    \top_I.branch[4].block[12].um_I.iw[2] ,
    \top_I.branch[4].block[12].um_I.iw[1] ,
    \top_I.branch[4].block[12].um_I.clk ,
    \top_I.branch[4].block[11].um_I.iw[17] ,
    \top_I.branch[4].block[11].um_I.iw[16] ,
    \top_I.branch[4].block[11].um_I.iw[15] ,
    \top_I.branch[4].block[11].um_I.iw[14] ,
    \top_I.branch[4].block[11].um_I.iw[13] ,
    \top_I.branch[4].block[11].um_I.iw[12] ,
    \top_I.branch[4].block[11].um_I.iw[11] ,
    \top_I.branch[4].block[11].um_I.iw[10] ,
    \top_I.branch[4].block[11].um_I.iw[9] ,
    \top_I.branch[4].block[11].um_I.iw[8] ,
    \top_I.branch[4].block[11].um_I.iw[7] ,
    \top_I.branch[4].block[11].um_I.iw[6] ,
    \top_I.branch[4].block[11].um_I.iw[5] ,
    \top_I.branch[4].block[11].um_I.iw[4] ,
    \top_I.branch[4].block[11].um_I.iw[3] ,
    \top_I.branch[4].block[11].um_I.iw[2] ,
    \top_I.branch[4].block[11].um_I.iw[1] ,
    \top_I.branch[4].block[11].um_I.clk ,
    \top_I.branch[4].block[10].um_I.iw[17] ,
    \top_I.branch[4].block[10].um_I.iw[16] ,
    \top_I.branch[4].block[10].um_I.iw[15] ,
    \top_I.branch[4].block[10].um_I.iw[14] ,
    \top_I.branch[4].block[10].um_I.iw[13] ,
    \top_I.branch[4].block[10].um_I.iw[12] ,
    \top_I.branch[4].block[10].um_I.iw[11] ,
    \top_I.branch[4].block[10].um_I.iw[10] ,
    \top_I.branch[4].block[10].um_I.iw[9] ,
    \top_I.branch[4].block[10].um_I.iw[8] ,
    \top_I.branch[4].block[10].um_I.iw[7] ,
    \top_I.branch[4].block[10].um_I.iw[6] ,
    \top_I.branch[4].block[10].um_I.iw[5] ,
    \top_I.branch[4].block[10].um_I.iw[4] ,
    \top_I.branch[4].block[10].um_I.iw[3] ,
    \top_I.branch[4].block[10].um_I.iw[2] ,
    \top_I.branch[4].block[10].um_I.iw[1] ,
    \top_I.branch[4].block[10].um_I.clk ,
    \top_I.branch[4].block[9].um_I.iw[17] ,
    \top_I.branch[4].block[9].um_I.iw[16] ,
    \top_I.branch[4].block[9].um_I.iw[15] ,
    \top_I.branch[4].block[9].um_I.iw[14] ,
    \top_I.branch[4].block[9].um_I.iw[13] ,
    \top_I.branch[4].block[9].um_I.iw[12] ,
    \top_I.branch[4].block[9].um_I.iw[11] ,
    \top_I.branch[4].block[9].um_I.iw[10] ,
    \top_I.branch[4].block[9].um_I.iw[9] ,
    \top_I.branch[4].block[9].um_I.iw[8] ,
    \top_I.branch[4].block[9].um_I.iw[7] ,
    \top_I.branch[4].block[9].um_I.iw[6] ,
    \top_I.branch[4].block[9].um_I.iw[5] ,
    \top_I.branch[4].block[9].um_I.iw[4] ,
    \top_I.branch[4].block[9].um_I.iw[3] ,
    \top_I.branch[4].block[9].um_I.iw[2] ,
    \top_I.branch[4].block[9].um_I.iw[1] ,
    \top_I.branch[4].block[9].um_I.clk ,
    \top_I.branch[4].block[8].um_I.iw[17] ,
    \top_I.branch[4].block[8].um_I.iw[16] ,
    \top_I.branch[4].block[8].um_I.iw[15] ,
    \top_I.branch[4].block[8].um_I.iw[14] ,
    \top_I.branch[4].block[8].um_I.iw[13] ,
    \top_I.branch[4].block[8].um_I.iw[12] ,
    \top_I.branch[4].block[8].um_I.iw[11] ,
    \top_I.branch[4].block[8].um_I.iw[10] ,
    \top_I.branch[4].block[8].um_I.iw[9] ,
    \top_I.branch[4].block[8].um_I.iw[8] ,
    \top_I.branch[4].block[8].um_I.iw[7] ,
    \top_I.branch[4].block[8].um_I.iw[6] ,
    \top_I.branch[4].block[8].um_I.iw[5] ,
    \top_I.branch[4].block[8].um_I.iw[4] ,
    \top_I.branch[4].block[8].um_I.iw[3] ,
    \top_I.branch[4].block[8].um_I.iw[2] ,
    \top_I.branch[4].block[8].um_I.iw[1] ,
    \top_I.branch[4].block[8].um_I.clk ,
    \top_I.branch[4].block[7].um_I.iw[17] ,
    \top_I.branch[4].block[7].um_I.iw[16] ,
    \top_I.branch[4].block[7].um_I.iw[15] ,
    \top_I.branch[4].block[7].um_I.iw[14] ,
    \top_I.branch[4].block[7].um_I.iw[13] ,
    \top_I.branch[4].block[7].um_I.iw[12] ,
    \top_I.branch[4].block[7].um_I.iw[11] ,
    \top_I.branch[4].block[7].um_I.iw[10] ,
    \top_I.branch[4].block[7].um_I.iw[9] ,
    \top_I.branch[4].block[7].um_I.iw[8] ,
    \top_I.branch[4].block[7].um_I.iw[7] ,
    \top_I.branch[4].block[7].um_I.iw[6] ,
    \top_I.branch[4].block[7].um_I.iw[5] ,
    \top_I.branch[4].block[7].um_I.iw[4] ,
    \top_I.branch[4].block[7].um_I.iw[3] ,
    \top_I.branch[4].block[7].um_I.iw[2] ,
    \top_I.branch[4].block[7].um_I.iw[1] ,
    \top_I.branch[4].block[7].um_I.clk ,
    \top_I.branch[4].block[6].um_I.iw[17] ,
    \top_I.branch[4].block[6].um_I.iw[16] ,
    \top_I.branch[4].block[6].um_I.iw[15] ,
    \top_I.branch[4].block[6].um_I.iw[14] ,
    \top_I.branch[4].block[6].um_I.iw[13] ,
    \top_I.branch[4].block[6].um_I.iw[12] ,
    \top_I.branch[4].block[6].um_I.iw[11] ,
    \top_I.branch[4].block[6].um_I.iw[10] ,
    \top_I.branch[4].block[6].um_I.iw[9] ,
    \top_I.branch[4].block[6].um_I.iw[8] ,
    \top_I.branch[4].block[6].um_I.iw[7] ,
    \top_I.branch[4].block[6].um_I.iw[6] ,
    \top_I.branch[4].block[6].um_I.iw[5] ,
    \top_I.branch[4].block[6].um_I.iw[4] ,
    \top_I.branch[4].block[6].um_I.iw[3] ,
    \top_I.branch[4].block[6].um_I.iw[2] ,
    \top_I.branch[4].block[6].um_I.iw[1] ,
    \top_I.branch[4].block[6].um_I.clk ,
    \top_I.branch[4].block[5].um_I.iw[17] ,
    \top_I.branch[4].block[5].um_I.iw[16] ,
    \top_I.branch[4].block[5].um_I.iw[15] ,
    \top_I.branch[4].block[5].um_I.iw[14] ,
    \top_I.branch[4].block[5].um_I.iw[13] ,
    \top_I.branch[4].block[5].um_I.iw[12] ,
    \top_I.branch[4].block[5].um_I.iw[11] ,
    \top_I.branch[4].block[5].um_I.iw[10] ,
    \top_I.branch[4].block[5].um_I.iw[9] ,
    \top_I.branch[4].block[5].um_I.iw[8] ,
    \top_I.branch[4].block[5].um_I.iw[7] ,
    \top_I.branch[4].block[5].um_I.iw[6] ,
    \top_I.branch[4].block[5].um_I.iw[5] ,
    \top_I.branch[4].block[5].um_I.iw[4] ,
    \top_I.branch[4].block[5].um_I.iw[3] ,
    \top_I.branch[4].block[5].um_I.iw[2] ,
    \top_I.branch[4].block[5].um_I.iw[1] ,
    \top_I.branch[4].block[5].um_I.clk ,
    \top_I.branch[4].block[4].um_I.iw[17] ,
    \top_I.branch[4].block[4].um_I.iw[16] ,
    \top_I.branch[4].block[4].um_I.iw[15] ,
    \top_I.branch[4].block[4].um_I.iw[14] ,
    \top_I.branch[4].block[4].um_I.iw[13] ,
    \top_I.branch[4].block[4].um_I.iw[12] ,
    \top_I.branch[4].block[4].um_I.iw[11] ,
    \top_I.branch[4].block[4].um_I.iw[10] ,
    \top_I.branch[4].block[4].um_I.iw[9] ,
    \top_I.branch[4].block[4].um_I.iw[8] ,
    \top_I.branch[4].block[4].um_I.iw[7] ,
    \top_I.branch[4].block[4].um_I.iw[6] ,
    \top_I.branch[4].block[4].um_I.iw[5] ,
    \top_I.branch[4].block[4].um_I.iw[4] ,
    \top_I.branch[4].block[4].um_I.iw[3] ,
    \top_I.branch[4].block[4].um_I.iw[2] ,
    \top_I.branch[4].block[4].um_I.iw[1] ,
    \top_I.branch[4].block[4].um_I.clk ,
    \top_I.branch[4].block[3].um_I.iw[17] ,
    \top_I.branch[4].block[3].um_I.iw[16] ,
    \top_I.branch[4].block[3].um_I.iw[15] ,
    \top_I.branch[4].block[3].um_I.iw[14] ,
    \top_I.branch[4].block[3].um_I.iw[13] ,
    \top_I.branch[4].block[3].um_I.iw[12] ,
    \top_I.branch[4].block[3].um_I.iw[11] ,
    \top_I.branch[4].block[3].um_I.iw[10] ,
    \top_I.branch[4].block[3].um_I.iw[9] ,
    \top_I.branch[4].block[3].um_I.iw[8] ,
    \top_I.branch[4].block[3].um_I.iw[7] ,
    \top_I.branch[4].block[3].um_I.iw[6] ,
    \top_I.branch[4].block[3].um_I.iw[5] ,
    \top_I.branch[4].block[3].um_I.iw[4] ,
    \top_I.branch[4].block[3].um_I.iw[3] ,
    \top_I.branch[4].block[3].um_I.iw[2] ,
    \top_I.branch[4].block[3].um_I.iw[1] ,
    \top_I.branch[4].block[3].um_I.clk ,
    \top_I.branch[4].block[2].um_I.iw[17] ,
    \top_I.branch[4].block[2].um_I.iw[16] ,
    \top_I.branch[4].block[2].um_I.iw[15] ,
    \top_I.branch[4].block[2].um_I.iw[14] ,
    \top_I.branch[4].block[2].um_I.iw[13] ,
    \top_I.branch[4].block[2].um_I.iw[12] ,
    \top_I.branch[4].block[2].um_I.iw[11] ,
    \top_I.branch[4].block[2].um_I.iw[10] ,
    \top_I.branch[4].block[2].um_I.iw[9] ,
    \top_I.branch[4].block[2].um_I.iw[8] ,
    \top_I.branch[4].block[2].um_I.iw[7] ,
    \top_I.branch[4].block[2].um_I.iw[6] ,
    \top_I.branch[4].block[2].um_I.iw[5] ,
    \top_I.branch[4].block[2].um_I.iw[4] ,
    \top_I.branch[4].block[2].um_I.iw[3] ,
    \top_I.branch[4].block[2].um_I.iw[2] ,
    \top_I.branch[4].block[2].um_I.iw[1] ,
    \top_I.branch[4].block[2].um_I.clk ,
    \top_I.branch[4].block[1].um_I.iw[17] ,
    \top_I.branch[4].block[1].um_I.iw[16] ,
    \top_I.branch[4].block[1].um_I.iw[15] ,
    \top_I.branch[4].block[1].um_I.iw[14] ,
    \top_I.branch[4].block[1].um_I.iw[13] ,
    \top_I.branch[4].block[1].um_I.iw[12] ,
    \top_I.branch[4].block[1].um_I.iw[11] ,
    \top_I.branch[4].block[1].um_I.iw[10] ,
    \top_I.branch[4].block[1].um_I.iw[9] ,
    \top_I.branch[4].block[1].um_I.iw[8] ,
    \top_I.branch[4].block[1].um_I.iw[7] ,
    \top_I.branch[4].block[1].um_I.iw[6] ,
    \top_I.branch[4].block[1].um_I.iw[5] ,
    \top_I.branch[4].block[1].um_I.iw[4] ,
    \top_I.branch[4].block[1].um_I.iw[3] ,
    \top_I.branch[4].block[1].um_I.iw[2] ,
    \top_I.branch[4].block[1].um_I.iw[1] ,
    \top_I.branch[4].block[1].um_I.clk ,
    \top_I.branch[4].block[0].um_I.iw[17] ,
    \top_I.branch[4].block[0].um_I.iw[16] ,
    \top_I.branch[4].block[0].um_I.iw[15] ,
    \top_I.branch[4].block[0].um_I.iw[14] ,
    \top_I.branch[4].block[0].um_I.iw[13] ,
    \top_I.branch[4].block[0].um_I.iw[12] ,
    \top_I.branch[4].block[0].um_I.iw[11] ,
    \top_I.branch[4].block[0].um_I.iw[10] ,
    \top_I.branch[4].block[0].um_I.iw[9] ,
    \top_I.branch[4].block[0].um_I.iw[8] ,
    \top_I.branch[4].block[0].um_I.iw[7] ,
    \top_I.branch[4].block[0].um_I.iw[6] ,
    \top_I.branch[4].block[0].um_I.iw[5] ,
    \top_I.branch[4].block[0].um_I.iw[4] ,
    \top_I.branch[4].block[0].um_I.iw[3] ,
    \top_I.branch[4].block[0].um_I.iw[2] ,
    \top_I.branch[4].block[0].um_I.iw[1] ,
    \top_I.branch[4].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[15].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[14].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[13].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[12].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[11].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[10].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[9].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[8].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[7].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[6].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[5].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[4].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[3].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[2].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[1].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero ,
    \top_I.branch[4].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[4].block[15].um_I.pg_vdd ,
    \top_I.branch[4].block[14].um_I.pg_vdd ,
    \top_I.branch[4].block[13].um_I.pg_vdd ,
    \top_I.branch[4].block[12].um_I.pg_vdd ,
    \top_I.branch[4].block[11].um_I.pg_vdd ,
    \top_I.branch[4].block[10].um_I.pg_vdd ,
    \top_I.branch[4].block[9].um_I.pg_vdd ,
    \top_I.branch[4].block[8].um_I.pg_vdd ,
    \top_I.branch[4].block[7].um_I.pg_vdd ,
    \top_I.branch[4].block[6].um_I.pg_vdd ,
    \top_I.branch[4].block[5].um_I.pg_vdd ,
    \top_I.branch[4].block[4].um_I.pg_vdd ,
    \top_I.branch[4].block[3].um_I.pg_vdd ,
    \top_I.branch[4].block[2].um_I.pg_vdd ,
    \top_I.branch[4].block[1].um_I.pg_vdd ,
    \top_I.branch[4].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[5].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[5].l_addr[1] ),
    .k_zero(\top_I.branch[5].l_addr[0] ),
    .addr({\top_I.branch[5].l_addr[0] ,
    \top_I.branch[5].l_addr[0] ,
    \top_I.branch[5].l_addr[1] ,
    \top_I.branch[5].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[5].block[15].um_I.ena ,
    \top_I.branch[5].block[14].um_I.ena ,
    \top_I.branch[5].block[13].um_I.ena ,
    \top_I.branch[5].block[12].um_I.ena ,
    \top_I.branch[5].block[11].um_I.ena ,
    \top_I.branch[5].block[10].um_I.ena ,
    \top_I.branch[5].block[9].um_I.ena ,
    \top_I.branch[5].block[8].um_I.ena ,
    \top_I.branch[5].block[7].um_I.ena ,
    \top_I.branch[5].block[6].um_I.ena ,
    \top_I.branch[5].block[5].um_I.ena ,
    \top_I.branch[5].block[4].um_I.ena ,
    \top_I.branch[5].block[3].um_I.ena ,
    \top_I.branch[5].block[2].um_I.ena ,
    \top_I.branch[5].block[1].um_I.ena ,
    \top_I.branch[5].block[0].um_I.ena }),
    .um_iw({\top_I.branch[5].block[15].um_I.iw[17] ,
    \top_I.branch[5].block[15].um_I.iw[16] ,
    \top_I.branch[5].block[15].um_I.iw[15] ,
    \top_I.branch[5].block[15].um_I.iw[14] ,
    \top_I.branch[5].block[15].um_I.iw[13] ,
    \top_I.branch[5].block[15].um_I.iw[12] ,
    \top_I.branch[5].block[15].um_I.iw[11] ,
    \top_I.branch[5].block[15].um_I.iw[10] ,
    \top_I.branch[5].block[15].um_I.iw[9] ,
    \top_I.branch[5].block[15].um_I.iw[8] ,
    \top_I.branch[5].block[15].um_I.iw[7] ,
    \top_I.branch[5].block[15].um_I.iw[6] ,
    \top_I.branch[5].block[15].um_I.iw[5] ,
    \top_I.branch[5].block[15].um_I.iw[4] ,
    \top_I.branch[5].block[15].um_I.iw[3] ,
    \top_I.branch[5].block[15].um_I.iw[2] ,
    \top_I.branch[5].block[15].um_I.iw[1] ,
    \top_I.branch[5].block[15].um_I.clk ,
    \top_I.branch[5].block[14].um_I.iw[17] ,
    \top_I.branch[5].block[14].um_I.iw[16] ,
    \top_I.branch[5].block[14].um_I.iw[15] ,
    \top_I.branch[5].block[14].um_I.iw[14] ,
    \top_I.branch[5].block[14].um_I.iw[13] ,
    \top_I.branch[5].block[14].um_I.iw[12] ,
    \top_I.branch[5].block[14].um_I.iw[11] ,
    \top_I.branch[5].block[14].um_I.iw[10] ,
    \top_I.branch[5].block[14].um_I.iw[9] ,
    \top_I.branch[5].block[14].um_I.iw[8] ,
    \top_I.branch[5].block[14].um_I.iw[7] ,
    \top_I.branch[5].block[14].um_I.iw[6] ,
    \top_I.branch[5].block[14].um_I.iw[5] ,
    \top_I.branch[5].block[14].um_I.iw[4] ,
    \top_I.branch[5].block[14].um_I.iw[3] ,
    \top_I.branch[5].block[14].um_I.iw[2] ,
    \top_I.branch[5].block[14].um_I.iw[1] ,
    \top_I.branch[5].block[14].um_I.clk ,
    \top_I.branch[5].block[13].um_I.iw[17] ,
    \top_I.branch[5].block[13].um_I.iw[16] ,
    \top_I.branch[5].block[13].um_I.iw[15] ,
    \top_I.branch[5].block[13].um_I.iw[14] ,
    \top_I.branch[5].block[13].um_I.iw[13] ,
    \top_I.branch[5].block[13].um_I.iw[12] ,
    \top_I.branch[5].block[13].um_I.iw[11] ,
    \top_I.branch[5].block[13].um_I.iw[10] ,
    \top_I.branch[5].block[13].um_I.iw[9] ,
    \top_I.branch[5].block[13].um_I.iw[8] ,
    \top_I.branch[5].block[13].um_I.iw[7] ,
    \top_I.branch[5].block[13].um_I.iw[6] ,
    \top_I.branch[5].block[13].um_I.iw[5] ,
    \top_I.branch[5].block[13].um_I.iw[4] ,
    \top_I.branch[5].block[13].um_I.iw[3] ,
    \top_I.branch[5].block[13].um_I.iw[2] ,
    \top_I.branch[5].block[13].um_I.iw[1] ,
    \top_I.branch[5].block[13].um_I.clk ,
    \top_I.branch[5].block[12].um_I.iw[17] ,
    \top_I.branch[5].block[12].um_I.iw[16] ,
    \top_I.branch[5].block[12].um_I.iw[15] ,
    \top_I.branch[5].block[12].um_I.iw[14] ,
    \top_I.branch[5].block[12].um_I.iw[13] ,
    \top_I.branch[5].block[12].um_I.iw[12] ,
    \top_I.branch[5].block[12].um_I.iw[11] ,
    \top_I.branch[5].block[12].um_I.iw[10] ,
    \top_I.branch[5].block[12].um_I.iw[9] ,
    \top_I.branch[5].block[12].um_I.iw[8] ,
    \top_I.branch[5].block[12].um_I.iw[7] ,
    \top_I.branch[5].block[12].um_I.iw[6] ,
    \top_I.branch[5].block[12].um_I.iw[5] ,
    \top_I.branch[5].block[12].um_I.iw[4] ,
    \top_I.branch[5].block[12].um_I.iw[3] ,
    \top_I.branch[5].block[12].um_I.iw[2] ,
    \top_I.branch[5].block[12].um_I.iw[1] ,
    \top_I.branch[5].block[12].um_I.clk ,
    \top_I.branch[5].block[11].um_I.iw[17] ,
    \top_I.branch[5].block[11].um_I.iw[16] ,
    \top_I.branch[5].block[11].um_I.iw[15] ,
    \top_I.branch[5].block[11].um_I.iw[14] ,
    \top_I.branch[5].block[11].um_I.iw[13] ,
    \top_I.branch[5].block[11].um_I.iw[12] ,
    \top_I.branch[5].block[11].um_I.iw[11] ,
    \top_I.branch[5].block[11].um_I.iw[10] ,
    \top_I.branch[5].block[11].um_I.iw[9] ,
    \top_I.branch[5].block[11].um_I.iw[8] ,
    \top_I.branch[5].block[11].um_I.iw[7] ,
    \top_I.branch[5].block[11].um_I.iw[6] ,
    \top_I.branch[5].block[11].um_I.iw[5] ,
    \top_I.branch[5].block[11].um_I.iw[4] ,
    \top_I.branch[5].block[11].um_I.iw[3] ,
    \top_I.branch[5].block[11].um_I.iw[2] ,
    \top_I.branch[5].block[11].um_I.iw[1] ,
    \top_I.branch[5].block[11].um_I.clk ,
    \top_I.branch[5].block[10].um_I.iw[17] ,
    \top_I.branch[5].block[10].um_I.iw[16] ,
    \top_I.branch[5].block[10].um_I.iw[15] ,
    \top_I.branch[5].block[10].um_I.iw[14] ,
    \top_I.branch[5].block[10].um_I.iw[13] ,
    \top_I.branch[5].block[10].um_I.iw[12] ,
    \top_I.branch[5].block[10].um_I.iw[11] ,
    \top_I.branch[5].block[10].um_I.iw[10] ,
    \top_I.branch[5].block[10].um_I.iw[9] ,
    \top_I.branch[5].block[10].um_I.iw[8] ,
    \top_I.branch[5].block[10].um_I.iw[7] ,
    \top_I.branch[5].block[10].um_I.iw[6] ,
    \top_I.branch[5].block[10].um_I.iw[5] ,
    \top_I.branch[5].block[10].um_I.iw[4] ,
    \top_I.branch[5].block[10].um_I.iw[3] ,
    \top_I.branch[5].block[10].um_I.iw[2] ,
    \top_I.branch[5].block[10].um_I.iw[1] ,
    \top_I.branch[5].block[10].um_I.clk ,
    \top_I.branch[5].block[9].um_I.iw[17] ,
    \top_I.branch[5].block[9].um_I.iw[16] ,
    \top_I.branch[5].block[9].um_I.iw[15] ,
    \top_I.branch[5].block[9].um_I.iw[14] ,
    \top_I.branch[5].block[9].um_I.iw[13] ,
    \top_I.branch[5].block[9].um_I.iw[12] ,
    \top_I.branch[5].block[9].um_I.iw[11] ,
    \top_I.branch[5].block[9].um_I.iw[10] ,
    \top_I.branch[5].block[9].um_I.iw[9] ,
    \top_I.branch[5].block[9].um_I.iw[8] ,
    \top_I.branch[5].block[9].um_I.iw[7] ,
    \top_I.branch[5].block[9].um_I.iw[6] ,
    \top_I.branch[5].block[9].um_I.iw[5] ,
    \top_I.branch[5].block[9].um_I.iw[4] ,
    \top_I.branch[5].block[9].um_I.iw[3] ,
    \top_I.branch[5].block[9].um_I.iw[2] ,
    \top_I.branch[5].block[9].um_I.iw[1] ,
    \top_I.branch[5].block[9].um_I.clk ,
    \top_I.branch[5].block[8].um_I.iw[17] ,
    \top_I.branch[5].block[8].um_I.iw[16] ,
    \top_I.branch[5].block[8].um_I.iw[15] ,
    \top_I.branch[5].block[8].um_I.iw[14] ,
    \top_I.branch[5].block[8].um_I.iw[13] ,
    \top_I.branch[5].block[8].um_I.iw[12] ,
    \top_I.branch[5].block[8].um_I.iw[11] ,
    \top_I.branch[5].block[8].um_I.iw[10] ,
    \top_I.branch[5].block[8].um_I.iw[9] ,
    \top_I.branch[5].block[8].um_I.iw[8] ,
    \top_I.branch[5].block[8].um_I.iw[7] ,
    \top_I.branch[5].block[8].um_I.iw[6] ,
    \top_I.branch[5].block[8].um_I.iw[5] ,
    \top_I.branch[5].block[8].um_I.iw[4] ,
    \top_I.branch[5].block[8].um_I.iw[3] ,
    \top_I.branch[5].block[8].um_I.iw[2] ,
    \top_I.branch[5].block[8].um_I.iw[1] ,
    \top_I.branch[5].block[8].um_I.clk ,
    \top_I.branch[5].block[7].um_I.iw[17] ,
    \top_I.branch[5].block[7].um_I.iw[16] ,
    \top_I.branch[5].block[7].um_I.iw[15] ,
    \top_I.branch[5].block[7].um_I.iw[14] ,
    \top_I.branch[5].block[7].um_I.iw[13] ,
    \top_I.branch[5].block[7].um_I.iw[12] ,
    \top_I.branch[5].block[7].um_I.iw[11] ,
    \top_I.branch[5].block[7].um_I.iw[10] ,
    \top_I.branch[5].block[7].um_I.iw[9] ,
    \top_I.branch[5].block[7].um_I.iw[8] ,
    \top_I.branch[5].block[7].um_I.iw[7] ,
    \top_I.branch[5].block[7].um_I.iw[6] ,
    \top_I.branch[5].block[7].um_I.iw[5] ,
    \top_I.branch[5].block[7].um_I.iw[4] ,
    \top_I.branch[5].block[7].um_I.iw[3] ,
    \top_I.branch[5].block[7].um_I.iw[2] ,
    \top_I.branch[5].block[7].um_I.iw[1] ,
    \top_I.branch[5].block[7].um_I.clk ,
    \top_I.branch[5].block[6].um_I.iw[17] ,
    \top_I.branch[5].block[6].um_I.iw[16] ,
    \top_I.branch[5].block[6].um_I.iw[15] ,
    \top_I.branch[5].block[6].um_I.iw[14] ,
    \top_I.branch[5].block[6].um_I.iw[13] ,
    \top_I.branch[5].block[6].um_I.iw[12] ,
    \top_I.branch[5].block[6].um_I.iw[11] ,
    \top_I.branch[5].block[6].um_I.iw[10] ,
    \top_I.branch[5].block[6].um_I.iw[9] ,
    \top_I.branch[5].block[6].um_I.iw[8] ,
    \top_I.branch[5].block[6].um_I.iw[7] ,
    \top_I.branch[5].block[6].um_I.iw[6] ,
    \top_I.branch[5].block[6].um_I.iw[5] ,
    \top_I.branch[5].block[6].um_I.iw[4] ,
    \top_I.branch[5].block[6].um_I.iw[3] ,
    \top_I.branch[5].block[6].um_I.iw[2] ,
    \top_I.branch[5].block[6].um_I.iw[1] ,
    \top_I.branch[5].block[6].um_I.clk ,
    \top_I.branch[5].block[5].um_I.iw[17] ,
    \top_I.branch[5].block[5].um_I.iw[16] ,
    \top_I.branch[5].block[5].um_I.iw[15] ,
    \top_I.branch[5].block[5].um_I.iw[14] ,
    \top_I.branch[5].block[5].um_I.iw[13] ,
    \top_I.branch[5].block[5].um_I.iw[12] ,
    \top_I.branch[5].block[5].um_I.iw[11] ,
    \top_I.branch[5].block[5].um_I.iw[10] ,
    \top_I.branch[5].block[5].um_I.iw[9] ,
    \top_I.branch[5].block[5].um_I.iw[8] ,
    \top_I.branch[5].block[5].um_I.iw[7] ,
    \top_I.branch[5].block[5].um_I.iw[6] ,
    \top_I.branch[5].block[5].um_I.iw[5] ,
    \top_I.branch[5].block[5].um_I.iw[4] ,
    \top_I.branch[5].block[5].um_I.iw[3] ,
    \top_I.branch[5].block[5].um_I.iw[2] ,
    \top_I.branch[5].block[5].um_I.iw[1] ,
    \top_I.branch[5].block[5].um_I.clk ,
    \top_I.branch[5].block[4].um_I.iw[17] ,
    \top_I.branch[5].block[4].um_I.iw[16] ,
    \top_I.branch[5].block[4].um_I.iw[15] ,
    \top_I.branch[5].block[4].um_I.iw[14] ,
    \top_I.branch[5].block[4].um_I.iw[13] ,
    \top_I.branch[5].block[4].um_I.iw[12] ,
    \top_I.branch[5].block[4].um_I.iw[11] ,
    \top_I.branch[5].block[4].um_I.iw[10] ,
    \top_I.branch[5].block[4].um_I.iw[9] ,
    \top_I.branch[5].block[4].um_I.iw[8] ,
    \top_I.branch[5].block[4].um_I.iw[7] ,
    \top_I.branch[5].block[4].um_I.iw[6] ,
    \top_I.branch[5].block[4].um_I.iw[5] ,
    \top_I.branch[5].block[4].um_I.iw[4] ,
    \top_I.branch[5].block[4].um_I.iw[3] ,
    \top_I.branch[5].block[4].um_I.iw[2] ,
    \top_I.branch[5].block[4].um_I.iw[1] ,
    \top_I.branch[5].block[4].um_I.clk ,
    \top_I.branch[5].block[3].um_I.iw[17] ,
    \top_I.branch[5].block[3].um_I.iw[16] ,
    \top_I.branch[5].block[3].um_I.iw[15] ,
    \top_I.branch[5].block[3].um_I.iw[14] ,
    \top_I.branch[5].block[3].um_I.iw[13] ,
    \top_I.branch[5].block[3].um_I.iw[12] ,
    \top_I.branch[5].block[3].um_I.iw[11] ,
    \top_I.branch[5].block[3].um_I.iw[10] ,
    \top_I.branch[5].block[3].um_I.iw[9] ,
    \top_I.branch[5].block[3].um_I.iw[8] ,
    \top_I.branch[5].block[3].um_I.iw[7] ,
    \top_I.branch[5].block[3].um_I.iw[6] ,
    \top_I.branch[5].block[3].um_I.iw[5] ,
    \top_I.branch[5].block[3].um_I.iw[4] ,
    \top_I.branch[5].block[3].um_I.iw[3] ,
    \top_I.branch[5].block[3].um_I.iw[2] ,
    \top_I.branch[5].block[3].um_I.iw[1] ,
    \top_I.branch[5].block[3].um_I.clk ,
    \top_I.branch[5].block[2].um_I.iw[17] ,
    \top_I.branch[5].block[2].um_I.iw[16] ,
    \top_I.branch[5].block[2].um_I.iw[15] ,
    \top_I.branch[5].block[2].um_I.iw[14] ,
    \top_I.branch[5].block[2].um_I.iw[13] ,
    \top_I.branch[5].block[2].um_I.iw[12] ,
    \top_I.branch[5].block[2].um_I.iw[11] ,
    \top_I.branch[5].block[2].um_I.iw[10] ,
    \top_I.branch[5].block[2].um_I.iw[9] ,
    \top_I.branch[5].block[2].um_I.iw[8] ,
    \top_I.branch[5].block[2].um_I.iw[7] ,
    \top_I.branch[5].block[2].um_I.iw[6] ,
    \top_I.branch[5].block[2].um_I.iw[5] ,
    \top_I.branch[5].block[2].um_I.iw[4] ,
    \top_I.branch[5].block[2].um_I.iw[3] ,
    \top_I.branch[5].block[2].um_I.iw[2] ,
    \top_I.branch[5].block[2].um_I.iw[1] ,
    \top_I.branch[5].block[2].um_I.clk ,
    \top_I.branch[5].block[1].um_I.iw[17] ,
    \top_I.branch[5].block[1].um_I.iw[16] ,
    \top_I.branch[5].block[1].um_I.iw[15] ,
    \top_I.branch[5].block[1].um_I.iw[14] ,
    \top_I.branch[5].block[1].um_I.iw[13] ,
    \top_I.branch[5].block[1].um_I.iw[12] ,
    \top_I.branch[5].block[1].um_I.iw[11] ,
    \top_I.branch[5].block[1].um_I.iw[10] ,
    \top_I.branch[5].block[1].um_I.iw[9] ,
    \top_I.branch[5].block[1].um_I.iw[8] ,
    \top_I.branch[5].block[1].um_I.iw[7] ,
    \top_I.branch[5].block[1].um_I.iw[6] ,
    \top_I.branch[5].block[1].um_I.iw[5] ,
    \top_I.branch[5].block[1].um_I.iw[4] ,
    \top_I.branch[5].block[1].um_I.iw[3] ,
    \top_I.branch[5].block[1].um_I.iw[2] ,
    \top_I.branch[5].block[1].um_I.iw[1] ,
    \top_I.branch[5].block[1].um_I.clk ,
    \top_I.branch[5].block[0].um_I.iw[17] ,
    \top_I.branch[5].block[0].um_I.iw[16] ,
    \top_I.branch[5].block[0].um_I.iw[15] ,
    \top_I.branch[5].block[0].um_I.iw[14] ,
    \top_I.branch[5].block[0].um_I.iw[13] ,
    \top_I.branch[5].block[0].um_I.iw[12] ,
    \top_I.branch[5].block[0].um_I.iw[11] ,
    \top_I.branch[5].block[0].um_I.iw[10] ,
    \top_I.branch[5].block[0].um_I.iw[9] ,
    \top_I.branch[5].block[0].um_I.iw[8] ,
    \top_I.branch[5].block[0].um_I.iw[7] ,
    \top_I.branch[5].block[0].um_I.iw[6] ,
    \top_I.branch[5].block[0].um_I.iw[5] ,
    \top_I.branch[5].block[0].um_I.iw[4] ,
    \top_I.branch[5].block[0].um_I.iw[3] ,
    \top_I.branch[5].block[0].um_I.iw[2] ,
    \top_I.branch[5].block[0].um_I.iw[1] ,
    \top_I.branch[5].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[15].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[14].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[13].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[12].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[11].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[10].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[9].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[8].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[7].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[6].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[5].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[4].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[3].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[2].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[1].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero ,
    \top_I.branch[5].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[5].block[15].um_I.pg_vdd ,
    \top_I.branch[5].block[14].um_I.pg_vdd ,
    \top_I.branch[5].block[13].um_I.pg_vdd ,
    \top_I.branch[5].block[12].um_I.pg_vdd ,
    \top_I.branch[5].block[11].um_I.pg_vdd ,
    \top_I.branch[5].block[10].um_I.pg_vdd ,
    \top_I.branch[5].block[9].um_I.pg_vdd ,
    \top_I.branch[5].block[8].um_I.pg_vdd ,
    \top_I.branch[5].block[7].um_I.pg_vdd ,
    \top_I.branch[5].block[6].um_I.pg_vdd ,
    \top_I.branch[5].block[5].um_I.pg_vdd ,
    \top_I.branch[5].block[4].um_I.pg_vdd ,
    \top_I.branch[5].block[3].um_I.pg_vdd ,
    \top_I.branch[5].block[2].um_I.pg_vdd ,
    \top_I.branch[5].block[1].um_I.pg_vdd ,
    \top_I.branch[5].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[6].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[6].l_addr[0] ),
    .k_zero(\top_I.branch[6].l_addr[2] ),
    .addr({\top_I.branch[6].l_addr[2] ,
    \top_I.branch[6].l_addr[2] ,
    \top_I.branch[6].l_addr[0] ,
    \top_I.branch[6].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[6].block[15].um_I.ena ,
    \top_I.branch[6].block[14].um_I.ena ,
    \top_I.branch[6].block[13].um_I.ena ,
    \top_I.branch[6].block[12].um_I.ena ,
    \top_I.branch[6].block[11].um_I.ena ,
    \top_I.branch[6].block[10].um_I.ena ,
    \top_I.branch[6].block[9].um_I.ena ,
    \top_I.branch[6].block[8].um_I.ena ,
    \top_I.branch[6].block[7].um_I.ena ,
    \top_I.branch[6].block[6].um_I.ena ,
    \top_I.branch[6].block[5].um_I.ena ,
    \top_I.branch[6].block[4].um_I.ena ,
    \top_I.branch[6].block[3].um_I.ena ,
    \top_I.branch[6].block[2].um_I.ena ,
    \top_I.branch[6].block[1].um_I.ena ,
    \top_I.branch[6].block[0].um_I.ena }),
    .um_iw({\top_I.branch[6].block[15].um_I.iw[17] ,
    \top_I.branch[6].block[15].um_I.iw[16] ,
    \top_I.branch[6].block[15].um_I.iw[15] ,
    \top_I.branch[6].block[15].um_I.iw[14] ,
    \top_I.branch[6].block[15].um_I.iw[13] ,
    \top_I.branch[6].block[15].um_I.iw[12] ,
    \top_I.branch[6].block[15].um_I.iw[11] ,
    \top_I.branch[6].block[15].um_I.iw[10] ,
    \top_I.branch[6].block[15].um_I.iw[9] ,
    \top_I.branch[6].block[15].um_I.iw[8] ,
    \top_I.branch[6].block[15].um_I.iw[7] ,
    \top_I.branch[6].block[15].um_I.iw[6] ,
    \top_I.branch[6].block[15].um_I.iw[5] ,
    \top_I.branch[6].block[15].um_I.iw[4] ,
    \top_I.branch[6].block[15].um_I.iw[3] ,
    \top_I.branch[6].block[15].um_I.iw[2] ,
    \top_I.branch[6].block[15].um_I.iw[1] ,
    \top_I.branch[6].block[15].um_I.clk ,
    \top_I.branch[6].block[14].um_I.iw[17] ,
    \top_I.branch[6].block[14].um_I.iw[16] ,
    \top_I.branch[6].block[14].um_I.iw[15] ,
    \top_I.branch[6].block[14].um_I.iw[14] ,
    \top_I.branch[6].block[14].um_I.iw[13] ,
    \top_I.branch[6].block[14].um_I.iw[12] ,
    \top_I.branch[6].block[14].um_I.iw[11] ,
    \top_I.branch[6].block[14].um_I.iw[10] ,
    \top_I.branch[6].block[14].um_I.iw[9] ,
    \top_I.branch[6].block[14].um_I.iw[8] ,
    \top_I.branch[6].block[14].um_I.iw[7] ,
    \top_I.branch[6].block[14].um_I.iw[6] ,
    \top_I.branch[6].block[14].um_I.iw[5] ,
    \top_I.branch[6].block[14].um_I.iw[4] ,
    \top_I.branch[6].block[14].um_I.iw[3] ,
    \top_I.branch[6].block[14].um_I.iw[2] ,
    \top_I.branch[6].block[14].um_I.iw[1] ,
    \top_I.branch[6].block[14].um_I.clk ,
    \top_I.branch[6].block[13].um_I.iw[17] ,
    \top_I.branch[6].block[13].um_I.iw[16] ,
    \top_I.branch[6].block[13].um_I.iw[15] ,
    \top_I.branch[6].block[13].um_I.iw[14] ,
    \top_I.branch[6].block[13].um_I.iw[13] ,
    \top_I.branch[6].block[13].um_I.iw[12] ,
    \top_I.branch[6].block[13].um_I.iw[11] ,
    \top_I.branch[6].block[13].um_I.iw[10] ,
    \top_I.branch[6].block[13].um_I.iw[9] ,
    \top_I.branch[6].block[13].um_I.iw[8] ,
    \top_I.branch[6].block[13].um_I.iw[7] ,
    \top_I.branch[6].block[13].um_I.iw[6] ,
    \top_I.branch[6].block[13].um_I.iw[5] ,
    \top_I.branch[6].block[13].um_I.iw[4] ,
    \top_I.branch[6].block[13].um_I.iw[3] ,
    \top_I.branch[6].block[13].um_I.iw[2] ,
    \top_I.branch[6].block[13].um_I.iw[1] ,
    \top_I.branch[6].block[13].um_I.clk ,
    \top_I.branch[6].block[12].um_I.iw[17] ,
    \top_I.branch[6].block[12].um_I.iw[16] ,
    \top_I.branch[6].block[12].um_I.iw[15] ,
    \top_I.branch[6].block[12].um_I.iw[14] ,
    \top_I.branch[6].block[12].um_I.iw[13] ,
    \top_I.branch[6].block[12].um_I.iw[12] ,
    \top_I.branch[6].block[12].um_I.iw[11] ,
    \top_I.branch[6].block[12].um_I.iw[10] ,
    \top_I.branch[6].block[12].um_I.iw[9] ,
    \top_I.branch[6].block[12].um_I.iw[8] ,
    \top_I.branch[6].block[12].um_I.iw[7] ,
    \top_I.branch[6].block[12].um_I.iw[6] ,
    \top_I.branch[6].block[12].um_I.iw[5] ,
    \top_I.branch[6].block[12].um_I.iw[4] ,
    \top_I.branch[6].block[12].um_I.iw[3] ,
    \top_I.branch[6].block[12].um_I.iw[2] ,
    \top_I.branch[6].block[12].um_I.iw[1] ,
    \top_I.branch[6].block[12].um_I.clk ,
    \top_I.branch[6].block[11].um_I.iw[17] ,
    \top_I.branch[6].block[11].um_I.iw[16] ,
    \top_I.branch[6].block[11].um_I.iw[15] ,
    \top_I.branch[6].block[11].um_I.iw[14] ,
    \top_I.branch[6].block[11].um_I.iw[13] ,
    \top_I.branch[6].block[11].um_I.iw[12] ,
    \top_I.branch[6].block[11].um_I.iw[11] ,
    \top_I.branch[6].block[11].um_I.iw[10] ,
    \top_I.branch[6].block[11].um_I.iw[9] ,
    \top_I.branch[6].block[11].um_I.iw[8] ,
    \top_I.branch[6].block[11].um_I.iw[7] ,
    \top_I.branch[6].block[11].um_I.iw[6] ,
    \top_I.branch[6].block[11].um_I.iw[5] ,
    \top_I.branch[6].block[11].um_I.iw[4] ,
    \top_I.branch[6].block[11].um_I.iw[3] ,
    \top_I.branch[6].block[11].um_I.iw[2] ,
    \top_I.branch[6].block[11].um_I.iw[1] ,
    \top_I.branch[6].block[11].um_I.clk ,
    \top_I.branch[6].block[10].um_I.iw[17] ,
    \top_I.branch[6].block[10].um_I.iw[16] ,
    \top_I.branch[6].block[10].um_I.iw[15] ,
    \top_I.branch[6].block[10].um_I.iw[14] ,
    \top_I.branch[6].block[10].um_I.iw[13] ,
    \top_I.branch[6].block[10].um_I.iw[12] ,
    \top_I.branch[6].block[10].um_I.iw[11] ,
    \top_I.branch[6].block[10].um_I.iw[10] ,
    \top_I.branch[6].block[10].um_I.iw[9] ,
    \top_I.branch[6].block[10].um_I.iw[8] ,
    \top_I.branch[6].block[10].um_I.iw[7] ,
    \top_I.branch[6].block[10].um_I.iw[6] ,
    \top_I.branch[6].block[10].um_I.iw[5] ,
    \top_I.branch[6].block[10].um_I.iw[4] ,
    \top_I.branch[6].block[10].um_I.iw[3] ,
    \top_I.branch[6].block[10].um_I.iw[2] ,
    \top_I.branch[6].block[10].um_I.iw[1] ,
    \top_I.branch[6].block[10].um_I.clk ,
    \top_I.branch[6].block[9].um_I.iw[17] ,
    \top_I.branch[6].block[9].um_I.iw[16] ,
    \top_I.branch[6].block[9].um_I.iw[15] ,
    \top_I.branch[6].block[9].um_I.iw[14] ,
    \top_I.branch[6].block[9].um_I.iw[13] ,
    \top_I.branch[6].block[9].um_I.iw[12] ,
    \top_I.branch[6].block[9].um_I.iw[11] ,
    \top_I.branch[6].block[9].um_I.iw[10] ,
    \top_I.branch[6].block[9].um_I.iw[9] ,
    \top_I.branch[6].block[9].um_I.iw[8] ,
    \top_I.branch[6].block[9].um_I.iw[7] ,
    \top_I.branch[6].block[9].um_I.iw[6] ,
    \top_I.branch[6].block[9].um_I.iw[5] ,
    \top_I.branch[6].block[9].um_I.iw[4] ,
    \top_I.branch[6].block[9].um_I.iw[3] ,
    \top_I.branch[6].block[9].um_I.iw[2] ,
    \top_I.branch[6].block[9].um_I.iw[1] ,
    \top_I.branch[6].block[9].um_I.clk ,
    \top_I.branch[6].block[8].um_I.iw[17] ,
    \top_I.branch[6].block[8].um_I.iw[16] ,
    \top_I.branch[6].block[8].um_I.iw[15] ,
    \top_I.branch[6].block[8].um_I.iw[14] ,
    \top_I.branch[6].block[8].um_I.iw[13] ,
    \top_I.branch[6].block[8].um_I.iw[12] ,
    \top_I.branch[6].block[8].um_I.iw[11] ,
    \top_I.branch[6].block[8].um_I.iw[10] ,
    \top_I.branch[6].block[8].um_I.iw[9] ,
    \top_I.branch[6].block[8].um_I.iw[8] ,
    \top_I.branch[6].block[8].um_I.iw[7] ,
    \top_I.branch[6].block[8].um_I.iw[6] ,
    \top_I.branch[6].block[8].um_I.iw[5] ,
    \top_I.branch[6].block[8].um_I.iw[4] ,
    \top_I.branch[6].block[8].um_I.iw[3] ,
    \top_I.branch[6].block[8].um_I.iw[2] ,
    \top_I.branch[6].block[8].um_I.iw[1] ,
    \top_I.branch[6].block[8].um_I.clk ,
    \top_I.branch[6].block[7].um_I.iw[17] ,
    \top_I.branch[6].block[7].um_I.iw[16] ,
    \top_I.branch[6].block[7].um_I.iw[15] ,
    \top_I.branch[6].block[7].um_I.iw[14] ,
    \top_I.branch[6].block[7].um_I.iw[13] ,
    \top_I.branch[6].block[7].um_I.iw[12] ,
    \top_I.branch[6].block[7].um_I.iw[11] ,
    \top_I.branch[6].block[7].um_I.iw[10] ,
    \top_I.branch[6].block[7].um_I.iw[9] ,
    \top_I.branch[6].block[7].um_I.iw[8] ,
    \top_I.branch[6].block[7].um_I.iw[7] ,
    \top_I.branch[6].block[7].um_I.iw[6] ,
    \top_I.branch[6].block[7].um_I.iw[5] ,
    \top_I.branch[6].block[7].um_I.iw[4] ,
    \top_I.branch[6].block[7].um_I.iw[3] ,
    \top_I.branch[6].block[7].um_I.iw[2] ,
    \top_I.branch[6].block[7].um_I.iw[1] ,
    \top_I.branch[6].block[7].um_I.clk ,
    \top_I.branch[6].block[6].um_I.iw[17] ,
    \top_I.branch[6].block[6].um_I.iw[16] ,
    \top_I.branch[6].block[6].um_I.iw[15] ,
    \top_I.branch[6].block[6].um_I.iw[14] ,
    \top_I.branch[6].block[6].um_I.iw[13] ,
    \top_I.branch[6].block[6].um_I.iw[12] ,
    \top_I.branch[6].block[6].um_I.iw[11] ,
    \top_I.branch[6].block[6].um_I.iw[10] ,
    \top_I.branch[6].block[6].um_I.iw[9] ,
    \top_I.branch[6].block[6].um_I.iw[8] ,
    \top_I.branch[6].block[6].um_I.iw[7] ,
    \top_I.branch[6].block[6].um_I.iw[6] ,
    \top_I.branch[6].block[6].um_I.iw[5] ,
    \top_I.branch[6].block[6].um_I.iw[4] ,
    \top_I.branch[6].block[6].um_I.iw[3] ,
    \top_I.branch[6].block[6].um_I.iw[2] ,
    \top_I.branch[6].block[6].um_I.iw[1] ,
    \top_I.branch[6].block[6].um_I.clk ,
    \top_I.branch[6].block[5].um_I.iw[17] ,
    \top_I.branch[6].block[5].um_I.iw[16] ,
    \top_I.branch[6].block[5].um_I.iw[15] ,
    \top_I.branch[6].block[5].um_I.iw[14] ,
    \top_I.branch[6].block[5].um_I.iw[13] ,
    \top_I.branch[6].block[5].um_I.iw[12] ,
    \top_I.branch[6].block[5].um_I.iw[11] ,
    \top_I.branch[6].block[5].um_I.iw[10] ,
    \top_I.branch[6].block[5].um_I.iw[9] ,
    \top_I.branch[6].block[5].um_I.iw[8] ,
    \top_I.branch[6].block[5].um_I.iw[7] ,
    \top_I.branch[6].block[5].um_I.iw[6] ,
    \top_I.branch[6].block[5].um_I.iw[5] ,
    \top_I.branch[6].block[5].um_I.iw[4] ,
    \top_I.branch[6].block[5].um_I.iw[3] ,
    \top_I.branch[6].block[5].um_I.iw[2] ,
    \top_I.branch[6].block[5].um_I.iw[1] ,
    \top_I.branch[6].block[5].um_I.clk ,
    \top_I.branch[6].block[4].um_I.iw[17] ,
    \top_I.branch[6].block[4].um_I.iw[16] ,
    \top_I.branch[6].block[4].um_I.iw[15] ,
    \top_I.branch[6].block[4].um_I.iw[14] ,
    \top_I.branch[6].block[4].um_I.iw[13] ,
    \top_I.branch[6].block[4].um_I.iw[12] ,
    \top_I.branch[6].block[4].um_I.iw[11] ,
    \top_I.branch[6].block[4].um_I.iw[10] ,
    \top_I.branch[6].block[4].um_I.iw[9] ,
    \top_I.branch[6].block[4].um_I.iw[8] ,
    \top_I.branch[6].block[4].um_I.iw[7] ,
    \top_I.branch[6].block[4].um_I.iw[6] ,
    \top_I.branch[6].block[4].um_I.iw[5] ,
    \top_I.branch[6].block[4].um_I.iw[4] ,
    \top_I.branch[6].block[4].um_I.iw[3] ,
    \top_I.branch[6].block[4].um_I.iw[2] ,
    \top_I.branch[6].block[4].um_I.iw[1] ,
    \top_I.branch[6].block[4].um_I.clk ,
    \top_I.branch[6].block[3].um_I.iw[17] ,
    \top_I.branch[6].block[3].um_I.iw[16] ,
    \top_I.branch[6].block[3].um_I.iw[15] ,
    \top_I.branch[6].block[3].um_I.iw[14] ,
    \top_I.branch[6].block[3].um_I.iw[13] ,
    \top_I.branch[6].block[3].um_I.iw[12] ,
    \top_I.branch[6].block[3].um_I.iw[11] ,
    \top_I.branch[6].block[3].um_I.iw[10] ,
    \top_I.branch[6].block[3].um_I.iw[9] ,
    \top_I.branch[6].block[3].um_I.iw[8] ,
    \top_I.branch[6].block[3].um_I.iw[7] ,
    \top_I.branch[6].block[3].um_I.iw[6] ,
    \top_I.branch[6].block[3].um_I.iw[5] ,
    \top_I.branch[6].block[3].um_I.iw[4] ,
    \top_I.branch[6].block[3].um_I.iw[3] ,
    \top_I.branch[6].block[3].um_I.iw[2] ,
    \top_I.branch[6].block[3].um_I.iw[1] ,
    \top_I.branch[6].block[3].um_I.clk ,
    \top_I.branch[6].block[2].um_I.iw[17] ,
    \top_I.branch[6].block[2].um_I.iw[16] ,
    \top_I.branch[6].block[2].um_I.iw[15] ,
    \top_I.branch[6].block[2].um_I.iw[14] ,
    \top_I.branch[6].block[2].um_I.iw[13] ,
    \top_I.branch[6].block[2].um_I.iw[12] ,
    \top_I.branch[6].block[2].um_I.iw[11] ,
    \top_I.branch[6].block[2].um_I.iw[10] ,
    \top_I.branch[6].block[2].um_I.iw[9] ,
    \top_I.branch[6].block[2].um_I.iw[8] ,
    \top_I.branch[6].block[2].um_I.iw[7] ,
    \top_I.branch[6].block[2].um_I.iw[6] ,
    \top_I.branch[6].block[2].um_I.iw[5] ,
    \top_I.branch[6].block[2].um_I.iw[4] ,
    \top_I.branch[6].block[2].um_I.iw[3] ,
    \top_I.branch[6].block[2].um_I.iw[2] ,
    \top_I.branch[6].block[2].um_I.iw[1] ,
    \top_I.branch[6].block[2].um_I.clk ,
    \top_I.branch[6].block[1].um_I.iw[17] ,
    \top_I.branch[6].block[1].um_I.iw[16] ,
    \top_I.branch[6].block[1].um_I.iw[15] ,
    \top_I.branch[6].block[1].um_I.iw[14] ,
    \top_I.branch[6].block[1].um_I.iw[13] ,
    \top_I.branch[6].block[1].um_I.iw[12] ,
    \top_I.branch[6].block[1].um_I.iw[11] ,
    \top_I.branch[6].block[1].um_I.iw[10] ,
    \top_I.branch[6].block[1].um_I.iw[9] ,
    \top_I.branch[6].block[1].um_I.iw[8] ,
    \top_I.branch[6].block[1].um_I.iw[7] ,
    \top_I.branch[6].block[1].um_I.iw[6] ,
    \top_I.branch[6].block[1].um_I.iw[5] ,
    \top_I.branch[6].block[1].um_I.iw[4] ,
    \top_I.branch[6].block[1].um_I.iw[3] ,
    \top_I.branch[6].block[1].um_I.iw[2] ,
    \top_I.branch[6].block[1].um_I.iw[1] ,
    \top_I.branch[6].block[1].um_I.clk ,
    \top_I.branch[6].block[0].um_I.iw[17] ,
    \top_I.branch[6].block[0].um_I.iw[16] ,
    \top_I.branch[6].block[0].um_I.iw[15] ,
    \top_I.branch[6].block[0].um_I.iw[14] ,
    \top_I.branch[6].block[0].um_I.iw[13] ,
    \top_I.branch[6].block[0].um_I.iw[12] ,
    \top_I.branch[6].block[0].um_I.iw[11] ,
    \top_I.branch[6].block[0].um_I.iw[10] ,
    \top_I.branch[6].block[0].um_I.iw[9] ,
    \top_I.branch[6].block[0].um_I.iw[8] ,
    \top_I.branch[6].block[0].um_I.iw[7] ,
    \top_I.branch[6].block[0].um_I.iw[6] ,
    \top_I.branch[6].block[0].um_I.iw[5] ,
    \top_I.branch[6].block[0].um_I.iw[4] ,
    \top_I.branch[6].block[0].um_I.iw[3] ,
    \top_I.branch[6].block[0].um_I.iw[2] ,
    \top_I.branch[6].block[0].um_I.iw[1] ,
    \top_I.branch[6].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[15].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[14].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[13].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[12].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[11].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[10].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[9].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[8].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[7].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[6].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[5].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[4].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[3].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[2].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[1].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero ,
    \top_I.branch[6].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[6].block[15].um_I.pg_vdd ,
    \top_I.branch[6].block[14].um_I.pg_vdd ,
    \top_I.branch[6].block[13].um_I.pg_vdd ,
    \top_I.branch[6].block[12].um_I.pg_vdd ,
    \top_I.branch[6].block[11].um_I.pg_vdd ,
    \top_I.branch[6].block[10].um_I.pg_vdd ,
    \top_I.branch[6].block[9].um_I.pg_vdd ,
    \top_I.branch[6].block[8].um_I.pg_vdd ,
    \top_I.branch[6].block[7].um_I.pg_vdd ,
    \top_I.branch[6].block[6].um_I.pg_vdd ,
    \top_I.branch[6].block[5].um_I.pg_vdd ,
    \top_I.branch[6].block[4].um_I.pg_vdd ,
    \top_I.branch[6].block[3].um_I.pg_vdd ,
    \top_I.branch[6].block[2].um_I.pg_vdd ,
    \top_I.branch[6].block[1].um_I.pg_vdd ,
    \top_I.branch[6].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[7].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[7].l_addr[0] ),
    .k_zero(\top_I.branch[7].l_addr[2] ),
    .addr({\top_I.branch[7].l_addr[2] ,
    \top_I.branch[7].l_addr[2] ,
    \top_I.branch[7].l_addr[0] ,
    \top_I.branch[7].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[7].block[15].um_I.ena ,
    \top_I.branch[7].block[14].um_I.ena ,
    \top_I.branch[7].block[13].um_I.ena ,
    \top_I.branch[7].block[12].um_I.ena ,
    \top_I.branch[7].block[11].um_I.ena ,
    \top_I.branch[7].block[10].um_I.ena ,
    \top_I.branch[7].block[9].um_I.ena ,
    \top_I.branch[7].block[8].um_I.ena ,
    \top_I.branch[7].block[7].um_I.ena ,
    \top_I.branch[7].block[6].um_I.ena ,
    \top_I.branch[7].block[5].um_I.ena ,
    \top_I.branch[7].block[4].um_I.ena ,
    \top_I.branch[7].block[3].um_I.ena ,
    \top_I.branch[7].block[2].um_I.ena ,
    \top_I.branch[7].block[1].um_I.ena ,
    \top_I.branch[7].block[0].um_I.ena }),
    .um_iw({\top_I.branch[7].block[15].um_I.iw[17] ,
    \top_I.branch[7].block[15].um_I.iw[16] ,
    \top_I.branch[7].block[15].um_I.iw[15] ,
    \top_I.branch[7].block[15].um_I.iw[14] ,
    \top_I.branch[7].block[15].um_I.iw[13] ,
    \top_I.branch[7].block[15].um_I.iw[12] ,
    \top_I.branch[7].block[15].um_I.iw[11] ,
    \top_I.branch[7].block[15].um_I.iw[10] ,
    \top_I.branch[7].block[15].um_I.iw[9] ,
    \top_I.branch[7].block[15].um_I.iw[8] ,
    \top_I.branch[7].block[15].um_I.iw[7] ,
    \top_I.branch[7].block[15].um_I.iw[6] ,
    \top_I.branch[7].block[15].um_I.iw[5] ,
    \top_I.branch[7].block[15].um_I.iw[4] ,
    \top_I.branch[7].block[15].um_I.iw[3] ,
    \top_I.branch[7].block[15].um_I.iw[2] ,
    \top_I.branch[7].block[15].um_I.iw[1] ,
    \top_I.branch[7].block[15].um_I.clk ,
    \top_I.branch[7].block[14].um_I.iw[17] ,
    \top_I.branch[7].block[14].um_I.iw[16] ,
    \top_I.branch[7].block[14].um_I.iw[15] ,
    \top_I.branch[7].block[14].um_I.iw[14] ,
    \top_I.branch[7].block[14].um_I.iw[13] ,
    \top_I.branch[7].block[14].um_I.iw[12] ,
    \top_I.branch[7].block[14].um_I.iw[11] ,
    \top_I.branch[7].block[14].um_I.iw[10] ,
    \top_I.branch[7].block[14].um_I.iw[9] ,
    \top_I.branch[7].block[14].um_I.iw[8] ,
    \top_I.branch[7].block[14].um_I.iw[7] ,
    \top_I.branch[7].block[14].um_I.iw[6] ,
    \top_I.branch[7].block[14].um_I.iw[5] ,
    \top_I.branch[7].block[14].um_I.iw[4] ,
    \top_I.branch[7].block[14].um_I.iw[3] ,
    \top_I.branch[7].block[14].um_I.iw[2] ,
    \top_I.branch[7].block[14].um_I.iw[1] ,
    \top_I.branch[7].block[14].um_I.clk ,
    \top_I.branch[7].block[13].um_I.iw[17] ,
    \top_I.branch[7].block[13].um_I.iw[16] ,
    \top_I.branch[7].block[13].um_I.iw[15] ,
    \top_I.branch[7].block[13].um_I.iw[14] ,
    \top_I.branch[7].block[13].um_I.iw[13] ,
    \top_I.branch[7].block[13].um_I.iw[12] ,
    \top_I.branch[7].block[13].um_I.iw[11] ,
    \top_I.branch[7].block[13].um_I.iw[10] ,
    \top_I.branch[7].block[13].um_I.iw[9] ,
    \top_I.branch[7].block[13].um_I.iw[8] ,
    \top_I.branch[7].block[13].um_I.iw[7] ,
    \top_I.branch[7].block[13].um_I.iw[6] ,
    \top_I.branch[7].block[13].um_I.iw[5] ,
    \top_I.branch[7].block[13].um_I.iw[4] ,
    \top_I.branch[7].block[13].um_I.iw[3] ,
    \top_I.branch[7].block[13].um_I.iw[2] ,
    \top_I.branch[7].block[13].um_I.iw[1] ,
    \top_I.branch[7].block[13].um_I.clk ,
    \top_I.branch[7].block[12].um_I.iw[17] ,
    \top_I.branch[7].block[12].um_I.iw[16] ,
    \top_I.branch[7].block[12].um_I.iw[15] ,
    \top_I.branch[7].block[12].um_I.iw[14] ,
    \top_I.branch[7].block[12].um_I.iw[13] ,
    \top_I.branch[7].block[12].um_I.iw[12] ,
    \top_I.branch[7].block[12].um_I.iw[11] ,
    \top_I.branch[7].block[12].um_I.iw[10] ,
    \top_I.branch[7].block[12].um_I.iw[9] ,
    \top_I.branch[7].block[12].um_I.iw[8] ,
    \top_I.branch[7].block[12].um_I.iw[7] ,
    \top_I.branch[7].block[12].um_I.iw[6] ,
    \top_I.branch[7].block[12].um_I.iw[5] ,
    \top_I.branch[7].block[12].um_I.iw[4] ,
    \top_I.branch[7].block[12].um_I.iw[3] ,
    \top_I.branch[7].block[12].um_I.iw[2] ,
    \top_I.branch[7].block[12].um_I.iw[1] ,
    \top_I.branch[7].block[12].um_I.clk ,
    \top_I.branch[7].block[11].um_I.iw[17] ,
    \top_I.branch[7].block[11].um_I.iw[16] ,
    \top_I.branch[7].block[11].um_I.iw[15] ,
    \top_I.branch[7].block[11].um_I.iw[14] ,
    \top_I.branch[7].block[11].um_I.iw[13] ,
    \top_I.branch[7].block[11].um_I.iw[12] ,
    \top_I.branch[7].block[11].um_I.iw[11] ,
    \top_I.branch[7].block[11].um_I.iw[10] ,
    \top_I.branch[7].block[11].um_I.iw[9] ,
    \top_I.branch[7].block[11].um_I.iw[8] ,
    \top_I.branch[7].block[11].um_I.iw[7] ,
    \top_I.branch[7].block[11].um_I.iw[6] ,
    \top_I.branch[7].block[11].um_I.iw[5] ,
    \top_I.branch[7].block[11].um_I.iw[4] ,
    \top_I.branch[7].block[11].um_I.iw[3] ,
    \top_I.branch[7].block[11].um_I.iw[2] ,
    \top_I.branch[7].block[11].um_I.iw[1] ,
    \top_I.branch[7].block[11].um_I.clk ,
    \top_I.branch[7].block[10].um_I.iw[17] ,
    \top_I.branch[7].block[10].um_I.iw[16] ,
    \top_I.branch[7].block[10].um_I.iw[15] ,
    \top_I.branch[7].block[10].um_I.iw[14] ,
    \top_I.branch[7].block[10].um_I.iw[13] ,
    \top_I.branch[7].block[10].um_I.iw[12] ,
    \top_I.branch[7].block[10].um_I.iw[11] ,
    \top_I.branch[7].block[10].um_I.iw[10] ,
    \top_I.branch[7].block[10].um_I.iw[9] ,
    \top_I.branch[7].block[10].um_I.iw[8] ,
    \top_I.branch[7].block[10].um_I.iw[7] ,
    \top_I.branch[7].block[10].um_I.iw[6] ,
    \top_I.branch[7].block[10].um_I.iw[5] ,
    \top_I.branch[7].block[10].um_I.iw[4] ,
    \top_I.branch[7].block[10].um_I.iw[3] ,
    \top_I.branch[7].block[10].um_I.iw[2] ,
    \top_I.branch[7].block[10].um_I.iw[1] ,
    \top_I.branch[7].block[10].um_I.clk ,
    \top_I.branch[7].block[9].um_I.iw[17] ,
    \top_I.branch[7].block[9].um_I.iw[16] ,
    \top_I.branch[7].block[9].um_I.iw[15] ,
    \top_I.branch[7].block[9].um_I.iw[14] ,
    \top_I.branch[7].block[9].um_I.iw[13] ,
    \top_I.branch[7].block[9].um_I.iw[12] ,
    \top_I.branch[7].block[9].um_I.iw[11] ,
    \top_I.branch[7].block[9].um_I.iw[10] ,
    \top_I.branch[7].block[9].um_I.iw[9] ,
    \top_I.branch[7].block[9].um_I.iw[8] ,
    \top_I.branch[7].block[9].um_I.iw[7] ,
    \top_I.branch[7].block[9].um_I.iw[6] ,
    \top_I.branch[7].block[9].um_I.iw[5] ,
    \top_I.branch[7].block[9].um_I.iw[4] ,
    \top_I.branch[7].block[9].um_I.iw[3] ,
    \top_I.branch[7].block[9].um_I.iw[2] ,
    \top_I.branch[7].block[9].um_I.iw[1] ,
    \top_I.branch[7].block[9].um_I.clk ,
    \top_I.branch[7].block[8].um_I.iw[17] ,
    \top_I.branch[7].block[8].um_I.iw[16] ,
    \top_I.branch[7].block[8].um_I.iw[15] ,
    \top_I.branch[7].block[8].um_I.iw[14] ,
    \top_I.branch[7].block[8].um_I.iw[13] ,
    \top_I.branch[7].block[8].um_I.iw[12] ,
    \top_I.branch[7].block[8].um_I.iw[11] ,
    \top_I.branch[7].block[8].um_I.iw[10] ,
    \top_I.branch[7].block[8].um_I.iw[9] ,
    \top_I.branch[7].block[8].um_I.iw[8] ,
    \top_I.branch[7].block[8].um_I.iw[7] ,
    \top_I.branch[7].block[8].um_I.iw[6] ,
    \top_I.branch[7].block[8].um_I.iw[5] ,
    \top_I.branch[7].block[8].um_I.iw[4] ,
    \top_I.branch[7].block[8].um_I.iw[3] ,
    \top_I.branch[7].block[8].um_I.iw[2] ,
    \top_I.branch[7].block[8].um_I.iw[1] ,
    \top_I.branch[7].block[8].um_I.clk ,
    \top_I.branch[7].block[7].um_I.iw[17] ,
    \top_I.branch[7].block[7].um_I.iw[16] ,
    \top_I.branch[7].block[7].um_I.iw[15] ,
    \top_I.branch[7].block[7].um_I.iw[14] ,
    \top_I.branch[7].block[7].um_I.iw[13] ,
    \top_I.branch[7].block[7].um_I.iw[12] ,
    \top_I.branch[7].block[7].um_I.iw[11] ,
    \top_I.branch[7].block[7].um_I.iw[10] ,
    \top_I.branch[7].block[7].um_I.iw[9] ,
    \top_I.branch[7].block[7].um_I.iw[8] ,
    \top_I.branch[7].block[7].um_I.iw[7] ,
    \top_I.branch[7].block[7].um_I.iw[6] ,
    \top_I.branch[7].block[7].um_I.iw[5] ,
    \top_I.branch[7].block[7].um_I.iw[4] ,
    \top_I.branch[7].block[7].um_I.iw[3] ,
    \top_I.branch[7].block[7].um_I.iw[2] ,
    \top_I.branch[7].block[7].um_I.iw[1] ,
    \top_I.branch[7].block[7].um_I.clk ,
    \top_I.branch[7].block[6].um_I.iw[17] ,
    \top_I.branch[7].block[6].um_I.iw[16] ,
    \top_I.branch[7].block[6].um_I.iw[15] ,
    \top_I.branch[7].block[6].um_I.iw[14] ,
    \top_I.branch[7].block[6].um_I.iw[13] ,
    \top_I.branch[7].block[6].um_I.iw[12] ,
    \top_I.branch[7].block[6].um_I.iw[11] ,
    \top_I.branch[7].block[6].um_I.iw[10] ,
    \top_I.branch[7].block[6].um_I.iw[9] ,
    \top_I.branch[7].block[6].um_I.iw[8] ,
    \top_I.branch[7].block[6].um_I.iw[7] ,
    \top_I.branch[7].block[6].um_I.iw[6] ,
    \top_I.branch[7].block[6].um_I.iw[5] ,
    \top_I.branch[7].block[6].um_I.iw[4] ,
    \top_I.branch[7].block[6].um_I.iw[3] ,
    \top_I.branch[7].block[6].um_I.iw[2] ,
    \top_I.branch[7].block[6].um_I.iw[1] ,
    \top_I.branch[7].block[6].um_I.clk ,
    \top_I.branch[7].block[5].um_I.iw[17] ,
    \top_I.branch[7].block[5].um_I.iw[16] ,
    \top_I.branch[7].block[5].um_I.iw[15] ,
    \top_I.branch[7].block[5].um_I.iw[14] ,
    \top_I.branch[7].block[5].um_I.iw[13] ,
    \top_I.branch[7].block[5].um_I.iw[12] ,
    \top_I.branch[7].block[5].um_I.iw[11] ,
    \top_I.branch[7].block[5].um_I.iw[10] ,
    \top_I.branch[7].block[5].um_I.iw[9] ,
    \top_I.branch[7].block[5].um_I.iw[8] ,
    \top_I.branch[7].block[5].um_I.iw[7] ,
    \top_I.branch[7].block[5].um_I.iw[6] ,
    \top_I.branch[7].block[5].um_I.iw[5] ,
    \top_I.branch[7].block[5].um_I.iw[4] ,
    \top_I.branch[7].block[5].um_I.iw[3] ,
    \top_I.branch[7].block[5].um_I.iw[2] ,
    \top_I.branch[7].block[5].um_I.iw[1] ,
    \top_I.branch[7].block[5].um_I.clk ,
    \top_I.branch[7].block[4].um_I.iw[17] ,
    \top_I.branch[7].block[4].um_I.iw[16] ,
    \top_I.branch[7].block[4].um_I.iw[15] ,
    \top_I.branch[7].block[4].um_I.iw[14] ,
    \top_I.branch[7].block[4].um_I.iw[13] ,
    \top_I.branch[7].block[4].um_I.iw[12] ,
    \top_I.branch[7].block[4].um_I.iw[11] ,
    \top_I.branch[7].block[4].um_I.iw[10] ,
    \top_I.branch[7].block[4].um_I.iw[9] ,
    \top_I.branch[7].block[4].um_I.iw[8] ,
    \top_I.branch[7].block[4].um_I.iw[7] ,
    \top_I.branch[7].block[4].um_I.iw[6] ,
    \top_I.branch[7].block[4].um_I.iw[5] ,
    \top_I.branch[7].block[4].um_I.iw[4] ,
    \top_I.branch[7].block[4].um_I.iw[3] ,
    \top_I.branch[7].block[4].um_I.iw[2] ,
    \top_I.branch[7].block[4].um_I.iw[1] ,
    \top_I.branch[7].block[4].um_I.clk ,
    \top_I.branch[7].block[3].um_I.iw[17] ,
    \top_I.branch[7].block[3].um_I.iw[16] ,
    \top_I.branch[7].block[3].um_I.iw[15] ,
    \top_I.branch[7].block[3].um_I.iw[14] ,
    \top_I.branch[7].block[3].um_I.iw[13] ,
    \top_I.branch[7].block[3].um_I.iw[12] ,
    \top_I.branch[7].block[3].um_I.iw[11] ,
    \top_I.branch[7].block[3].um_I.iw[10] ,
    \top_I.branch[7].block[3].um_I.iw[9] ,
    \top_I.branch[7].block[3].um_I.iw[8] ,
    \top_I.branch[7].block[3].um_I.iw[7] ,
    \top_I.branch[7].block[3].um_I.iw[6] ,
    \top_I.branch[7].block[3].um_I.iw[5] ,
    \top_I.branch[7].block[3].um_I.iw[4] ,
    \top_I.branch[7].block[3].um_I.iw[3] ,
    \top_I.branch[7].block[3].um_I.iw[2] ,
    \top_I.branch[7].block[3].um_I.iw[1] ,
    \top_I.branch[7].block[3].um_I.clk ,
    \top_I.branch[7].block[2].um_I.iw[17] ,
    \top_I.branch[7].block[2].um_I.iw[16] ,
    \top_I.branch[7].block[2].um_I.iw[15] ,
    \top_I.branch[7].block[2].um_I.iw[14] ,
    \top_I.branch[7].block[2].um_I.iw[13] ,
    \top_I.branch[7].block[2].um_I.iw[12] ,
    \top_I.branch[7].block[2].um_I.iw[11] ,
    \top_I.branch[7].block[2].um_I.iw[10] ,
    \top_I.branch[7].block[2].um_I.iw[9] ,
    \top_I.branch[7].block[2].um_I.iw[8] ,
    \top_I.branch[7].block[2].um_I.iw[7] ,
    \top_I.branch[7].block[2].um_I.iw[6] ,
    \top_I.branch[7].block[2].um_I.iw[5] ,
    \top_I.branch[7].block[2].um_I.iw[4] ,
    \top_I.branch[7].block[2].um_I.iw[3] ,
    \top_I.branch[7].block[2].um_I.iw[2] ,
    \top_I.branch[7].block[2].um_I.iw[1] ,
    \top_I.branch[7].block[2].um_I.clk ,
    \top_I.branch[7].block[1].um_I.iw[17] ,
    \top_I.branch[7].block[1].um_I.iw[16] ,
    \top_I.branch[7].block[1].um_I.iw[15] ,
    \top_I.branch[7].block[1].um_I.iw[14] ,
    \top_I.branch[7].block[1].um_I.iw[13] ,
    \top_I.branch[7].block[1].um_I.iw[12] ,
    \top_I.branch[7].block[1].um_I.iw[11] ,
    \top_I.branch[7].block[1].um_I.iw[10] ,
    \top_I.branch[7].block[1].um_I.iw[9] ,
    \top_I.branch[7].block[1].um_I.iw[8] ,
    \top_I.branch[7].block[1].um_I.iw[7] ,
    \top_I.branch[7].block[1].um_I.iw[6] ,
    \top_I.branch[7].block[1].um_I.iw[5] ,
    \top_I.branch[7].block[1].um_I.iw[4] ,
    \top_I.branch[7].block[1].um_I.iw[3] ,
    \top_I.branch[7].block[1].um_I.iw[2] ,
    \top_I.branch[7].block[1].um_I.iw[1] ,
    \top_I.branch[7].block[1].um_I.clk ,
    \top_I.branch[7].block[0].um_I.iw[17] ,
    \top_I.branch[7].block[0].um_I.iw[16] ,
    \top_I.branch[7].block[0].um_I.iw[15] ,
    \top_I.branch[7].block[0].um_I.iw[14] ,
    \top_I.branch[7].block[0].um_I.iw[13] ,
    \top_I.branch[7].block[0].um_I.iw[12] ,
    \top_I.branch[7].block[0].um_I.iw[11] ,
    \top_I.branch[7].block[0].um_I.iw[10] ,
    \top_I.branch[7].block[0].um_I.iw[9] ,
    \top_I.branch[7].block[0].um_I.iw[8] ,
    \top_I.branch[7].block[0].um_I.iw[7] ,
    \top_I.branch[7].block[0].um_I.iw[6] ,
    \top_I.branch[7].block[0].um_I.iw[5] ,
    \top_I.branch[7].block[0].um_I.iw[4] ,
    \top_I.branch[7].block[0].um_I.iw[3] ,
    \top_I.branch[7].block[0].um_I.iw[2] ,
    \top_I.branch[7].block[0].um_I.iw[1] ,
    \top_I.branch[7].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[15].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[14].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[13].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[12].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[11].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[10].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[9].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[8].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[7].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[6].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[5].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[4].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[3].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[2].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[1].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero ,
    \top_I.branch[7].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[7].block[15].um_I.pg_vdd ,
    \top_I.branch[7].block[14].um_I.pg_vdd ,
    \top_I.branch[7].block[13].um_I.pg_vdd ,
    \top_I.branch[7].block[12].um_I.pg_vdd ,
    \top_I.branch[7].block[11].um_I.pg_vdd ,
    \top_I.branch[7].block[10].um_I.pg_vdd ,
    \top_I.branch[7].block[9].um_I.pg_vdd ,
    \top_I.branch[7].block[8].um_I.pg_vdd ,
    \top_I.branch[7].block[7].um_I.pg_vdd ,
    \top_I.branch[7].block[6].um_I.pg_vdd ,
    \top_I.branch[7].block[5].um_I.pg_vdd ,
    \top_I.branch[7].block[4].um_I.pg_vdd ,
    \top_I.branch[7].block[3].um_I.pg_vdd ,
    \top_I.branch[7].block[2].um_I.pg_vdd ,
    \top_I.branch[7].block[1].um_I.pg_vdd ,
    \top_I.branch[7].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[8].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[8].l_addr[2] ),
    .k_zero(\top_I.branch[8].l_addr[0] ),
    .addr({\top_I.branch[8].l_addr[0] ,
    \top_I.branch[8].l_addr[2] ,
    \top_I.branch[8].l_addr[0] ,
    \top_I.branch[8].l_addr[0] }),
    .spine_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .um_ena({\top_I.branch[8].block[15].um_I.ena ,
    \top_I.branch[8].block[14].um_I.ena ,
    \top_I.branch[8].block[13].um_I.ena ,
    \top_I.branch[8].block[12].um_I.ena ,
    \top_I.branch[8].block[11].um_I.ena ,
    \top_I.branch[8].block[10].um_I.ena ,
    \top_I.branch[8].block[9].um_I.ena ,
    \top_I.branch[8].block[8].um_I.ena ,
    \top_I.branch[8].block[7].um_I.ena ,
    \top_I.branch[8].block[6].um_I.ena ,
    \top_I.branch[8].block[5].um_I.ena ,
    \top_I.branch[8].block[4].um_I.ena ,
    \top_I.branch[8].block[3].um_I.ena ,
    \top_I.branch[8].block[2].um_I.ena ,
    \top_I.branch[8].block[1].um_I.ena ,
    \top_I.branch[8].block[0].um_I.ena }),
    .um_iw({\top_I.branch[8].block[15].um_I.iw[17] ,
    \top_I.branch[8].block[15].um_I.iw[16] ,
    \top_I.branch[8].block[15].um_I.iw[15] ,
    \top_I.branch[8].block[15].um_I.iw[14] ,
    \top_I.branch[8].block[15].um_I.iw[13] ,
    \top_I.branch[8].block[15].um_I.iw[12] ,
    \top_I.branch[8].block[15].um_I.iw[11] ,
    \top_I.branch[8].block[15].um_I.iw[10] ,
    \top_I.branch[8].block[15].um_I.iw[9] ,
    \top_I.branch[8].block[15].um_I.iw[8] ,
    \top_I.branch[8].block[15].um_I.iw[7] ,
    \top_I.branch[8].block[15].um_I.iw[6] ,
    \top_I.branch[8].block[15].um_I.iw[5] ,
    \top_I.branch[8].block[15].um_I.iw[4] ,
    \top_I.branch[8].block[15].um_I.iw[3] ,
    \top_I.branch[8].block[15].um_I.iw[2] ,
    \top_I.branch[8].block[15].um_I.iw[1] ,
    \top_I.branch[8].block[15].um_I.clk ,
    \top_I.branch[8].block[14].um_I.iw[17] ,
    \top_I.branch[8].block[14].um_I.iw[16] ,
    \top_I.branch[8].block[14].um_I.iw[15] ,
    \top_I.branch[8].block[14].um_I.iw[14] ,
    \top_I.branch[8].block[14].um_I.iw[13] ,
    \top_I.branch[8].block[14].um_I.iw[12] ,
    \top_I.branch[8].block[14].um_I.iw[11] ,
    \top_I.branch[8].block[14].um_I.iw[10] ,
    \top_I.branch[8].block[14].um_I.iw[9] ,
    \top_I.branch[8].block[14].um_I.iw[8] ,
    \top_I.branch[8].block[14].um_I.iw[7] ,
    \top_I.branch[8].block[14].um_I.iw[6] ,
    \top_I.branch[8].block[14].um_I.iw[5] ,
    \top_I.branch[8].block[14].um_I.iw[4] ,
    \top_I.branch[8].block[14].um_I.iw[3] ,
    \top_I.branch[8].block[14].um_I.iw[2] ,
    \top_I.branch[8].block[14].um_I.iw[1] ,
    \top_I.branch[8].block[14].um_I.clk ,
    \top_I.branch[8].block[13].um_I.iw[17] ,
    \top_I.branch[8].block[13].um_I.iw[16] ,
    \top_I.branch[8].block[13].um_I.iw[15] ,
    \top_I.branch[8].block[13].um_I.iw[14] ,
    \top_I.branch[8].block[13].um_I.iw[13] ,
    \top_I.branch[8].block[13].um_I.iw[12] ,
    \top_I.branch[8].block[13].um_I.iw[11] ,
    \top_I.branch[8].block[13].um_I.iw[10] ,
    \top_I.branch[8].block[13].um_I.iw[9] ,
    \top_I.branch[8].block[13].um_I.iw[8] ,
    \top_I.branch[8].block[13].um_I.iw[7] ,
    \top_I.branch[8].block[13].um_I.iw[6] ,
    \top_I.branch[8].block[13].um_I.iw[5] ,
    \top_I.branch[8].block[13].um_I.iw[4] ,
    \top_I.branch[8].block[13].um_I.iw[3] ,
    \top_I.branch[8].block[13].um_I.iw[2] ,
    \top_I.branch[8].block[13].um_I.iw[1] ,
    \top_I.branch[8].block[13].um_I.clk ,
    \top_I.branch[8].block[12].um_I.iw[17] ,
    \top_I.branch[8].block[12].um_I.iw[16] ,
    \top_I.branch[8].block[12].um_I.iw[15] ,
    \top_I.branch[8].block[12].um_I.iw[14] ,
    \top_I.branch[8].block[12].um_I.iw[13] ,
    \top_I.branch[8].block[12].um_I.iw[12] ,
    \top_I.branch[8].block[12].um_I.iw[11] ,
    \top_I.branch[8].block[12].um_I.iw[10] ,
    \top_I.branch[8].block[12].um_I.iw[9] ,
    \top_I.branch[8].block[12].um_I.iw[8] ,
    \top_I.branch[8].block[12].um_I.iw[7] ,
    \top_I.branch[8].block[12].um_I.iw[6] ,
    \top_I.branch[8].block[12].um_I.iw[5] ,
    \top_I.branch[8].block[12].um_I.iw[4] ,
    \top_I.branch[8].block[12].um_I.iw[3] ,
    \top_I.branch[8].block[12].um_I.iw[2] ,
    \top_I.branch[8].block[12].um_I.iw[1] ,
    \top_I.branch[8].block[12].um_I.clk ,
    \top_I.branch[8].block[11].um_I.iw[17] ,
    \top_I.branch[8].block[11].um_I.iw[16] ,
    \top_I.branch[8].block[11].um_I.iw[15] ,
    \top_I.branch[8].block[11].um_I.iw[14] ,
    \top_I.branch[8].block[11].um_I.iw[13] ,
    \top_I.branch[8].block[11].um_I.iw[12] ,
    \top_I.branch[8].block[11].um_I.iw[11] ,
    \top_I.branch[8].block[11].um_I.iw[10] ,
    \top_I.branch[8].block[11].um_I.iw[9] ,
    \top_I.branch[8].block[11].um_I.iw[8] ,
    \top_I.branch[8].block[11].um_I.iw[7] ,
    \top_I.branch[8].block[11].um_I.iw[6] ,
    \top_I.branch[8].block[11].um_I.iw[5] ,
    \top_I.branch[8].block[11].um_I.iw[4] ,
    \top_I.branch[8].block[11].um_I.iw[3] ,
    \top_I.branch[8].block[11].um_I.iw[2] ,
    \top_I.branch[8].block[11].um_I.iw[1] ,
    \top_I.branch[8].block[11].um_I.clk ,
    \top_I.branch[8].block[10].um_I.iw[17] ,
    \top_I.branch[8].block[10].um_I.iw[16] ,
    \top_I.branch[8].block[10].um_I.iw[15] ,
    \top_I.branch[8].block[10].um_I.iw[14] ,
    \top_I.branch[8].block[10].um_I.iw[13] ,
    \top_I.branch[8].block[10].um_I.iw[12] ,
    \top_I.branch[8].block[10].um_I.iw[11] ,
    \top_I.branch[8].block[10].um_I.iw[10] ,
    \top_I.branch[8].block[10].um_I.iw[9] ,
    \top_I.branch[8].block[10].um_I.iw[8] ,
    \top_I.branch[8].block[10].um_I.iw[7] ,
    \top_I.branch[8].block[10].um_I.iw[6] ,
    \top_I.branch[8].block[10].um_I.iw[5] ,
    \top_I.branch[8].block[10].um_I.iw[4] ,
    \top_I.branch[8].block[10].um_I.iw[3] ,
    \top_I.branch[8].block[10].um_I.iw[2] ,
    \top_I.branch[8].block[10].um_I.iw[1] ,
    \top_I.branch[8].block[10].um_I.clk ,
    \top_I.branch[8].block[9].um_I.iw[17] ,
    \top_I.branch[8].block[9].um_I.iw[16] ,
    \top_I.branch[8].block[9].um_I.iw[15] ,
    \top_I.branch[8].block[9].um_I.iw[14] ,
    \top_I.branch[8].block[9].um_I.iw[13] ,
    \top_I.branch[8].block[9].um_I.iw[12] ,
    \top_I.branch[8].block[9].um_I.iw[11] ,
    \top_I.branch[8].block[9].um_I.iw[10] ,
    \top_I.branch[8].block[9].um_I.iw[9] ,
    \top_I.branch[8].block[9].um_I.iw[8] ,
    \top_I.branch[8].block[9].um_I.iw[7] ,
    \top_I.branch[8].block[9].um_I.iw[6] ,
    \top_I.branch[8].block[9].um_I.iw[5] ,
    \top_I.branch[8].block[9].um_I.iw[4] ,
    \top_I.branch[8].block[9].um_I.iw[3] ,
    \top_I.branch[8].block[9].um_I.iw[2] ,
    \top_I.branch[8].block[9].um_I.iw[1] ,
    \top_I.branch[8].block[9].um_I.clk ,
    \top_I.branch[8].block[8].um_I.iw[17] ,
    \top_I.branch[8].block[8].um_I.iw[16] ,
    \top_I.branch[8].block[8].um_I.iw[15] ,
    \top_I.branch[8].block[8].um_I.iw[14] ,
    \top_I.branch[8].block[8].um_I.iw[13] ,
    \top_I.branch[8].block[8].um_I.iw[12] ,
    \top_I.branch[8].block[8].um_I.iw[11] ,
    \top_I.branch[8].block[8].um_I.iw[10] ,
    \top_I.branch[8].block[8].um_I.iw[9] ,
    \top_I.branch[8].block[8].um_I.iw[8] ,
    \top_I.branch[8].block[8].um_I.iw[7] ,
    \top_I.branch[8].block[8].um_I.iw[6] ,
    \top_I.branch[8].block[8].um_I.iw[5] ,
    \top_I.branch[8].block[8].um_I.iw[4] ,
    \top_I.branch[8].block[8].um_I.iw[3] ,
    \top_I.branch[8].block[8].um_I.iw[2] ,
    \top_I.branch[8].block[8].um_I.iw[1] ,
    \top_I.branch[8].block[8].um_I.clk ,
    \top_I.branch[8].block[7].um_I.iw[17] ,
    \top_I.branch[8].block[7].um_I.iw[16] ,
    \top_I.branch[8].block[7].um_I.iw[15] ,
    \top_I.branch[8].block[7].um_I.iw[14] ,
    \top_I.branch[8].block[7].um_I.iw[13] ,
    \top_I.branch[8].block[7].um_I.iw[12] ,
    \top_I.branch[8].block[7].um_I.iw[11] ,
    \top_I.branch[8].block[7].um_I.iw[10] ,
    \top_I.branch[8].block[7].um_I.iw[9] ,
    \top_I.branch[8].block[7].um_I.iw[8] ,
    \top_I.branch[8].block[7].um_I.iw[7] ,
    \top_I.branch[8].block[7].um_I.iw[6] ,
    \top_I.branch[8].block[7].um_I.iw[5] ,
    \top_I.branch[8].block[7].um_I.iw[4] ,
    \top_I.branch[8].block[7].um_I.iw[3] ,
    \top_I.branch[8].block[7].um_I.iw[2] ,
    \top_I.branch[8].block[7].um_I.iw[1] ,
    \top_I.branch[8].block[7].um_I.clk ,
    \top_I.branch[8].block[6].um_I.iw[17] ,
    \top_I.branch[8].block[6].um_I.iw[16] ,
    \top_I.branch[8].block[6].um_I.iw[15] ,
    \top_I.branch[8].block[6].um_I.iw[14] ,
    \top_I.branch[8].block[6].um_I.iw[13] ,
    \top_I.branch[8].block[6].um_I.iw[12] ,
    \top_I.branch[8].block[6].um_I.iw[11] ,
    \top_I.branch[8].block[6].um_I.iw[10] ,
    \top_I.branch[8].block[6].um_I.iw[9] ,
    \top_I.branch[8].block[6].um_I.iw[8] ,
    \top_I.branch[8].block[6].um_I.iw[7] ,
    \top_I.branch[8].block[6].um_I.iw[6] ,
    \top_I.branch[8].block[6].um_I.iw[5] ,
    \top_I.branch[8].block[6].um_I.iw[4] ,
    \top_I.branch[8].block[6].um_I.iw[3] ,
    \top_I.branch[8].block[6].um_I.iw[2] ,
    \top_I.branch[8].block[6].um_I.iw[1] ,
    \top_I.branch[8].block[6].um_I.clk ,
    \top_I.branch[8].block[5].um_I.iw[17] ,
    \top_I.branch[8].block[5].um_I.iw[16] ,
    \top_I.branch[8].block[5].um_I.iw[15] ,
    \top_I.branch[8].block[5].um_I.iw[14] ,
    \top_I.branch[8].block[5].um_I.iw[13] ,
    \top_I.branch[8].block[5].um_I.iw[12] ,
    \top_I.branch[8].block[5].um_I.iw[11] ,
    \top_I.branch[8].block[5].um_I.iw[10] ,
    \top_I.branch[8].block[5].um_I.iw[9] ,
    \top_I.branch[8].block[5].um_I.iw[8] ,
    \top_I.branch[8].block[5].um_I.iw[7] ,
    \top_I.branch[8].block[5].um_I.iw[6] ,
    \top_I.branch[8].block[5].um_I.iw[5] ,
    \top_I.branch[8].block[5].um_I.iw[4] ,
    \top_I.branch[8].block[5].um_I.iw[3] ,
    \top_I.branch[8].block[5].um_I.iw[2] ,
    \top_I.branch[8].block[5].um_I.iw[1] ,
    \top_I.branch[8].block[5].um_I.clk ,
    \top_I.branch[8].block[4].um_I.iw[17] ,
    \top_I.branch[8].block[4].um_I.iw[16] ,
    \top_I.branch[8].block[4].um_I.iw[15] ,
    \top_I.branch[8].block[4].um_I.iw[14] ,
    \top_I.branch[8].block[4].um_I.iw[13] ,
    \top_I.branch[8].block[4].um_I.iw[12] ,
    \top_I.branch[8].block[4].um_I.iw[11] ,
    \top_I.branch[8].block[4].um_I.iw[10] ,
    \top_I.branch[8].block[4].um_I.iw[9] ,
    \top_I.branch[8].block[4].um_I.iw[8] ,
    \top_I.branch[8].block[4].um_I.iw[7] ,
    \top_I.branch[8].block[4].um_I.iw[6] ,
    \top_I.branch[8].block[4].um_I.iw[5] ,
    \top_I.branch[8].block[4].um_I.iw[4] ,
    \top_I.branch[8].block[4].um_I.iw[3] ,
    \top_I.branch[8].block[4].um_I.iw[2] ,
    \top_I.branch[8].block[4].um_I.iw[1] ,
    \top_I.branch[8].block[4].um_I.clk ,
    \top_I.branch[8].block[3].um_I.iw[17] ,
    \top_I.branch[8].block[3].um_I.iw[16] ,
    \top_I.branch[8].block[3].um_I.iw[15] ,
    \top_I.branch[8].block[3].um_I.iw[14] ,
    \top_I.branch[8].block[3].um_I.iw[13] ,
    \top_I.branch[8].block[3].um_I.iw[12] ,
    \top_I.branch[8].block[3].um_I.iw[11] ,
    \top_I.branch[8].block[3].um_I.iw[10] ,
    \top_I.branch[8].block[3].um_I.iw[9] ,
    \top_I.branch[8].block[3].um_I.iw[8] ,
    \top_I.branch[8].block[3].um_I.iw[7] ,
    \top_I.branch[8].block[3].um_I.iw[6] ,
    \top_I.branch[8].block[3].um_I.iw[5] ,
    \top_I.branch[8].block[3].um_I.iw[4] ,
    \top_I.branch[8].block[3].um_I.iw[3] ,
    \top_I.branch[8].block[3].um_I.iw[2] ,
    \top_I.branch[8].block[3].um_I.iw[1] ,
    \top_I.branch[8].block[3].um_I.clk ,
    \top_I.branch[8].block[2].um_I.iw[17] ,
    \top_I.branch[8].block[2].um_I.iw[16] ,
    \top_I.branch[8].block[2].um_I.iw[15] ,
    \top_I.branch[8].block[2].um_I.iw[14] ,
    \top_I.branch[8].block[2].um_I.iw[13] ,
    \top_I.branch[8].block[2].um_I.iw[12] ,
    \top_I.branch[8].block[2].um_I.iw[11] ,
    \top_I.branch[8].block[2].um_I.iw[10] ,
    \top_I.branch[8].block[2].um_I.iw[9] ,
    \top_I.branch[8].block[2].um_I.iw[8] ,
    \top_I.branch[8].block[2].um_I.iw[7] ,
    \top_I.branch[8].block[2].um_I.iw[6] ,
    \top_I.branch[8].block[2].um_I.iw[5] ,
    \top_I.branch[8].block[2].um_I.iw[4] ,
    \top_I.branch[8].block[2].um_I.iw[3] ,
    \top_I.branch[8].block[2].um_I.iw[2] ,
    \top_I.branch[8].block[2].um_I.iw[1] ,
    \top_I.branch[8].block[2].um_I.clk ,
    \top_I.branch[8].block[1].um_I.iw[17] ,
    \top_I.branch[8].block[1].um_I.iw[16] ,
    \top_I.branch[8].block[1].um_I.iw[15] ,
    \top_I.branch[8].block[1].um_I.iw[14] ,
    \top_I.branch[8].block[1].um_I.iw[13] ,
    \top_I.branch[8].block[1].um_I.iw[12] ,
    \top_I.branch[8].block[1].um_I.iw[11] ,
    \top_I.branch[8].block[1].um_I.iw[10] ,
    \top_I.branch[8].block[1].um_I.iw[9] ,
    \top_I.branch[8].block[1].um_I.iw[8] ,
    \top_I.branch[8].block[1].um_I.iw[7] ,
    \top_I.branch[8].block[1].um_I.iw[6] ,
    \top_I.branch[8].block[1].um_I.iw[5] ,
    \top_I.branch[8].block[1].um_I.iw[4] ,
    \top_I.branch[8].block[1].um_I.iw[3] ,
    \top_I.branch[8].block[1].um_I.iw[2] ,
    \top_I.branch[8].block[1].um_I.iw[1] ,
    \top_I.branch[8].block[1].um_I.clk ,
    \top_I.branch[8].block[0].um_I.iw[17] ,
    \top_I.branch[8].block[0].um_I.iw[16] ,
    \top_I.branch[8].block[0].um_I.iw[15] ,
    \top_I.branch[8].block[0].um_I.iw[14] ,
    \top_I.branch[8].block[0].um_I.iw[13] ,
    \top_I.branch[8].block[0].um_I.iw[12] ,
    \top_I.branch[8].block[0].um_I.iw[11] ,
    \top_I.branch[8].block[0].um_I.iw[10] ,
    \top_I.branch[8].block[0].um_I.iw[9] ,
    \top_I.branch[8].block[0].um_I.iw[8] ,
    \top_I.branch[8].block[0].um_I.iw[7] ,
    \top_I.branch[8].block[0].um_I.iw[6] ,
    \top_I.branch[8].block[0].um_I.iw[5] ,
    \top_I.branch[8].block[0].um_I.iw[4] ,
    \top_I.branch[8].block[0].um_I.iw[3] ,
    \top_I.branch[8].block[0].um_I.iw[2] ,
    \top_I.branch[8].block[0].um_I.iw[1] ,
    \top_I.branch[8].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[15].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[14].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[13].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[12].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[11].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[10].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[9].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[8].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[7].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[6].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[5].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[4].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[3].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[2].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[1].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero ,
    \top_I.branch[8].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[8].block[15].um_I.pg_vdd ,
    \top_I.branch[8].block[14].um_I.pg_vdd ,
    \top_I.branch[8].block[13].um_I.pg_vdd ,
    \top_I.branch[8].block[12].um_I.pg_vdd ,
    \top_I.branch[8].block[11].um_I.pg_vdd ,
    \top_I.branch[8].block[10].um_I.pg_vdd ,
    \top_I.branch[8].block[9].um_I.pg_vdd ,
    \top_I.branch[8].block[8].um_I.pg_vdd ,
    \top_I.branch[8].block[7].um_I.pg_vdd ,
    \top_I.branch[8].block[6].um_I.pg_vdd ,
    \top_I.branch[8].block[5].um_I.pg_vdd ,
    \top_I.branch[8].block[4].um_I.pg_vdd ,
    \top_I.branch[8].block[3].um_I.pg_vdd ,
    \top_I.branch[8].block[2].um_I.pg_vdd ,
    \top_I.branch[8].block[1].um_I.pg_vdd ,
    \top_I.branch[8].block[0].um_I.pg_vdd }));
 tt_mux \top_I.branch[9].mux_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .k_one(\top_I.branch[9].l_addr[2] ),
    .k_zero(\top_I.branch[9].l_addr[0] ),
    .addr({\top_I.branch[9].l_addr[0] ,
    \top_I.branch[9].l_addr[2] ,
    \top_I.branch[9].l_addr[0] ,
    \top_I.branch[9].l_addr[0] }),
    .spine_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }),
    .um_ena({\top_I.branch[9].block[15].um_I.ena ,
    \top_I.branch[9].block[14].um_I.ena ,
    \top_I.branch[9].block[13].um_I.ena ,
    \top_I.branch[9].block[12].um_I.ena ,
    \top_I.branch[9].block[11].um_I.ena ,
    \top_I.branch[9].block[10].um_I.ena ,
    \top_I.branch[9].block[9].um_I.ena ,
    \top_I.branch[9].block[8].um_I.ena ,
    \top_I.branch[9].block[7].um_I.ena ,
    \top_I.branch[9].block[6].um_I.ena ,
    \top_I.branch[9].block[5].um_I.ena ,
    \top_I.branch[9].block[4].um_I.ena ,
    \top_I.branch[9].block[3].um_I.ena ,
    \top_I.branch[9].block[2].um_I.ena ,
    \top_I.branch[9].block[1].um_I.ena ,
    \top_I.branch[9].block[0].um_I.ena }),
    .um_iw({\top_I.branch[9].block[15].um_I.iw[17] ,
    \top_I.branch[9].block[15].um_I.iw[16] ,
    \top_I.branch[9].block[15].um_I.iw[15] ,
    \top_I.branch[9].block[15].um_I.iw[14] ,
    \top_I.branch[9].block[15].um_I.iw[13] ,
    \top_I.branch[9].block[15].um_I.iw[12] ,
    \top_I.branch[9].block[15].um_I.iw[11] ,
    \top_I.branch[9].block[15].um_I.iw[10] ,
    \top_I.branch[9].block[15].um_I.iw[9] ,
    \top_I.branch[9].block[15].um_I.iw[8] ,
    \top_I.branch[9].block[15].um_I.iw[7] ,
    \top_I.branch[9].block[15].um_I.iw[6] ,
    \top_I.branch[9].block[15].um_I.iw[5] ,
    \top_I.branch[9].block[15].um_I.iw[4] ,
    \top_I.branch[9].block[15].um_I.iw[3] ,
    \top_I.branch[9].block[15].um_I.iw[2] ,
    \top_I.branch[9].block[15].um_I.iw[1] ,
    \top_I.branch[9].block[15].um_I.clk ,
    \top_I.branch[9].block[14].um_I.iw[17] ,
    \top_I.branch[9].block[14].um_I.iw[16] ,
    \top_I.branch[9].block[14].um_I.iw[15] ,
    \top_I.branch[9].block[14].um_I.iw[14] ,
    \top_I.branch[9].block[14].um_I.iw[13] ,
    \top_I.branch[9].block[14].um_I.iw[12] ,
    \top_I.branch[9].block[14].um_I.iw[11] ,
    \top_I.branch[9].block[14].um_I.iw[10] ,
    \top_I.branch[9].block[14].um_I.iw[9] ,
    \top_I.branch[9].block[14].um_I.iw[8] ,
    \top_I.branch[9].block[14].um_I.iw[7] ,
    \top_I.branch[9].block[14].um_I.iw[6] ,
    \top_I.branch[9].block[14].um_I.iw[5] ,
    \top_I.branch[9].block[14].um_I.iw[4] ,
    \top_I.branch[9].block[14].um_I.iw[3] ,
    \top_I.branch[9].block[14].um_I.iw[2] ,
    \top_I.branch[9].block[14].um_I.iw[1] ,
    \top_I.branch[9].block[14].um_I.clk ,
    \top_I.branch[9].block[13].um_I.iw[17] ,
    \top_I.branch[9].block[13].um_I.iw[16] ,
    \top_I.branch[9].block[13].um_I.iw[15] ,
    \top_I.branch[9].block[13].um_I.iw[14] ,
    \top_I.branch[9].block[13].um_I.iw[13] ,
    \top_I.branch[9].block[13].um_I.iw[12] ,
    \top_I.branch[9].block[13].um_I.iw[11] ,
    \top_I.branch[9].block[13].um_I.iw[10] ,
    \top_I.branch[9].block[13].um_I.iw[9] ,
    \top_I.branch[9].block[13].um_I.iw[8] ,
    \top_I.branch[9].block[13].um_I.iw[7] ,
    \top_I.branch[9].block[13].um_I.iw[6] ,
    \top_I.branch[9].block[13].um_I.iw[5] ,
    \top_I.branch[9].block[13].um_I.iw[4] ,
    \top_I.branch[9].block[13].um_I.iw[3] ,
    \top_I.branch[9].block[13].um_I.iw[2] ,
    \top_I.branch[9].block[13].um_I.iw[1] ,
    \top_I.branch[9].block[13].um_I.clk ,
    \top_I.branch[9].block[12].um_I.iw[17] ,
    \top_I.branch[9].block[12].um_I.iw[16] ,
    \top_I.branch[9].block[12].um_I.iw[15] ,
    \top_I.branch[9].block[12].um_I.iw[14] ,
    \top_I.branch[9].block[12].um_I.iw[13] ,
    \top_I.branch[9].block[12].um_I.iw[12] ,
    \top_I.branch[9].block[12].um_I.iw[11] ,
    \top_I.branch[9].block[12].um_I.iw[10] ,
    \top_I.branch[9].block[12].um_I.iw[9] ,
    \top_I.branch[9].block[12].um_I.iw[8] ,
    \top_I.branch[9].block[12].um_I.iw[7] ,
    \top_I.branch[9].block[12].um_I.iw[6] ,
    \top_I.branch[9].block[12].um_I.iw[5] ,
    \top_I.branch[9].block[12].um_I.iw[4] ,
    \top_I.branch[9].block[12].um_I.iw[3] ,
    \top_I.branch[9].block[12].um_I.iw[2] ,
    \top_I.branch[9].block[12].um_I.iw[1] ,
    \top_I.branch[9].block[12].um_I.clk ,
    \top_I.branch[9].block[11].um_I.iw[17] ,
    \top_I.branch[9].block[11].um_I.iw[16] ,
    \top_I.branch[9].block[11].um_I.iw[15] ,
    \top_I.branch[9].block[11].um_I.iw[14] ,
    \top_I.branch[9].block[11].um_I.iw[13] ,
    \top_I.branch[9].block[11].um_I.iw[12] ,
    \top_I.branch[9].block[11].um_I.iw[11] ,
    \top_I.branch[9].block[11].um_I.iw[10] ,
    \top_I.branch[9].block[11].um_I.iw[9] ,
    \top_I.branch[9].block[11].um_I.iw[8] ,
    \top_I.branch[9].block[11].um_I.iw[7] ,
    \top_I.branch[9].block[11].um_I.iw[6] ,
    \top_I.branch[9].block[11].um_I.iw[5] ,
    \top_I.branch[9].block[11].um_I.iw[4] ,
    \top_I.branch[9].block[11].um_I.iw[3] ,
    \top_I.branch[9].block[11].um_I.iw[2] ,
    \top_I.branch[9].block[11].um_I.iw[1] ,
    \top_I.branch[9].block[11].um_I.clk ,
    \top_I.branch[9].block[10].um_I.iw[17] ,
    \top_I.branch[9].block[10].um_I.iw[16] ,
    \top_I.branch[9].block[10].um_I.iw[15] ,
    \top_I.branch[9].block[10].um_I.iw[14] ,
    \top_I.branch[9].block[10].um_I.iw[13] ,
    \top_I.branch[9].block[10].um_I.iw[12] ,
    \top_I.branch[9].block[10].um_I.iw[11] ,
    \top_I.branch[9].block[10].um_I.iw[10] ,
    \top_I.branch[9].block[10].um_I.iw[9] ,
    \top_I.branch[9].block[10].um_I.iw[8] ,
    \top_I.branch[9].block[10].um_I.iw[7] ,
    \top_I.branch[9].block[10].um_I.iw[6] ,
    \top_I.branch[9].block[10].um_I.iw[5] ,
    \top_I.branch[9].block[10].um_I.iw[4] ,
    \top_I.branch[9].block[10].um_I.iw[3] ,
    \top_I.branch[9].block[10].um_I.iw[2] ,
    \top_I.branch[9].block[10].um_I.iw[1] ,
    \top_I.branch[9].block[10].um_I.clk ,
    \top_I.branch[9].block[9].um_I.iw[17] ,
    \top_I.branch[9].block[9].um_I.iw[16] ,
    \top_I.branch[9].block[9].um_I.iw[15] ,
    \top_I.branch[9].block[9].um_I.iw[14] ,
    \top_I.branch[9].block[9].um_I.iw[13] ,
    \top_I.branch[9].block[9].um_I.iw[12] ,
    \top_I.branch[9].block[9].um_I.iw[11] ,
    \top_I.branch[9].block[9].um_I.iw[10] ,
    \top_I.branch[9].block[9].um_I.iw[9] ,
    \top_I.branch[9].block[9].um_I.iw[8] ,
    \top_I.branch[9].block[9].um_I.iw[7] ,
    \top_I.branch[9].block[9].um_I.iw[6] ,
    \top_I.branch[9].block[9].um_I.iw[5] ,
    \top_I.branch[9].block[9].um_I.iw[4] ,
    \top_I.branch[9].block[9].um_I.iw[3] ,
    \top_I.branch[9].block[9].um_I.iw[2] ,
    \top_I.branch[9].block[9].um_I.iw[1] ,
    \top_I.branch[9].block[9].um_I.clk ,
    \top_I.branch[9].block[8].um_I.iw[17] ,
    \top_I.branch[9].block[8].um_I.iw[16] ,
    \top_I.branch[9].block[8].um_I.iw[15] ,
    \top_I.branch[9].block[8].um_I.iw[14] ,
    \top_I.branch[9].block[8].um_I.iw[13] ,
    \top_I.branch[9].block[8].um_I.iw[12] ,
    \top_I.branch[9].block[8].um_I.iw[11] ,
    \top_I.branch[9].block[8].um_I.iw[10] ,
    \top_I.branch[9].block[8].um_I.iw[9] ,
    \top_I.branch[9].block[8].um_I.iw[8] ,
    \top_I.branch[9].block[8].um_I.iw[7] ,
    \top_I.branch[9].block[8].um_I.iw[6] ,
    \top_I.branch[9].block[8].um_I.iw[5] ,
    \top_I.branch[9].block[8].um_I.iw[4] ,
    \top_I.branch[9].block[8].um_I.iw[3] ,
    \top_I.branch[9].block[8].um_I.iw[2] ,
    \top_I.branch[9].block[8].um_I.iw[1] ,
    \top_I.branch[9].block[8].um_I.clk ,
    \top_I.branch[9].block[7].um_I.iw[17] ,
    \top_I.branch[9].block[7].um_I.iw[16] ,
    \top_I.branch[9].block[7].um_I.iw[15] ,
    \top_I.branch[9].block[7].um_I.iw[14] ,
    \top_I.branch[9].block[7].um_I.iw[13] ,
    \top_I.branch[9].block[7].um_I.iw[12] ,
    \top_I.branch[9].block[7].um_I.iw[11] ,
    \top_I.branch[9].block[7].um_I.iw[10] ,
    \top_I.branch[9].block[7].um_I.iw[9] ,
    \top_I.branch[9].block[7].um_I.iw[8] ,
    \top_I.branch[9].block[7].um_I.iw[7] ,
    \top_I.branch[9].block[7].um_I.iw[6] ,
    \top_I.branch[9].block[7].um_I.iw[5] ,
    \top_I.branch[9].block[7].um_I.iw[4] ,
    \top_I.branch[9].block[7].um_I.iw[3] ,
    \top_I.branch[9].block[7].um_I.iw[2] ,
    \top_I.branch[9].block[7].um_I.iw[1] ,
    \top_I.branch[9].block[7].um_I.clk ,
    \top_I.branch[9].block[6].um_I.iw[17] ,
    \top_I.branch[9].block[6].um_I.iw[16] ,
    \top_I.branch[9].block[6].um_I.iw[15] ,
    \top_I.branch[9].block[6].um_I.iw[14] ,
    \top_I.branch[9].block[6].um_I.iw[13] ,
    \top_I.branch[9].block[6].um_I.iw[12] ,
    \top_I.branch[9].block[6].um_I.iw[11] ,
    \top_I.branch[9].block[6].um_I.iw[10] ,
    \top_I.branch[9].block[6].um_I.iw[9] ,
    \top_I.branch[9].block[6].um_I.iw[8] ,
    \top_I.branch[9].block[6].um_I.iw[7] ,
    \top_I.branch[9].block[6].um_I.iw[6] ,
    \top_I.branch[9].block[6].um_I.iw[5] ,
    \top_I.branch[9].block[6].um_I.iw[4] ,
    \top_I.branch[9].block[6].um_I.iw[3] ,
    \top_I.branch[9].block[6].um_I.iw[2] ,
    \top_I.branch[9].block[6].um_I.iw[1] ,
    \top_I.branch[9].block[6].um_I.clk ,
    \top_I.branch[9].block[5].um_I.iw[17] ,
    \top_I.branch[9].block[5].um_I.iw[16] ,
    \top_I.branch[9].block[5].um_I.iw[15] ,
    \top_I.branch[9].block[5].um_I.iw[14] ,
    \top_I.branch[9].block[5].um_I.iw[13] ,
    \top_I.branch[9].block[5].um_I.iw[12] ,
    \top_I.branch[9].block[5].um_I.iw[11] ,
    \top_I.branch[9].block[5].um_I.iw[10] ,
    \top_I.branch[9].block[5].um_I.iw[9] ,
    \top_I.branch[9].block[5].um_I.iw[8] ,
    \top_I.branch[9].block[5].um_I.iw[7] ,
    \top_I.branch[9].block[5].um_I.iw[6] ,
    \top_I.branch[9].block[5].um_I.iw[5] ,
    \top_I.branch[9].block[5].um_I.iw[4] ,
    \top_I.branch[9].block[5].um_I.iw[3] ,
    \top_I.branch[9].block[5].um_I.iw[2] ,
    \top_I.branch[9].block[5].um_I.iw[1] ,
    \top_I.branch[9].block[5].um_I.clk ,
    \top_I.branch[9].block[4].um_I.iw[17] ,
    \top_I.branch[9].block[4].um_I.iw[16] ,
    \top_I.branch[9].block[4].um_I.iw[15] ,
    \top_I.branch[9].block[4].um_I.iw[14] ,
    \top_I.branch[9].block[4].um_I.iw[13] ,
    \top_I.branch[9].block[4].um_I.iw[12] ,
    \top_I.branch[9].block[4].um_I.iw[11] ,
    \top_I.branch[9].block[4].um_I.iw[10] ,
    \top_I.branch[9].block[4].um_I.iw[9] ,
    \top_I.branch[9].block[4].um_I.iw[8] ,
    \top_I.branch[9].block[4].um_I.iw[7] ,
    \top_I.branch[9].block[4].um_I.iw[6] ,
    \top_I.branch[9].block[4].um_I.iw[5] ,
    \top_I.branch[9].block[4].um_I.iw[4] ,
    \top_I.branch[9].block[4].um_I.iw[3] ,
    \top_I.branch[9].block[4].um_I.iw[2] ,
    \top_I.branch[9].block[4].um_I.iw[1] ,
    \top_I.branch[9].block[4].um_I.clk ,
    \top_I.branch[9].block[3].um_I.iw[17] ,
    \top_I.branch[9].block[3].um_I.iw[16] ,
    \top_I.branch[9].block[3].um_I.iw[15] ,
    \top_I.branch[9].block[3].um_I.iw[14] ,
    \top_I.branch[9].block[3].um_I.iw[13] ,
    \top_I.branch[9].block[3].um_I.iw[12] ,
    \top_I.branch[9].block[3].um_I.iw[11] ,
    \top_I.branch[9].block[3].um_I.iw[10] ,
    \top_I.branch[9].block[3].um_I.iw[9] ,
    \top_I.branch[9].block[3].um_I.iw[8] ,
    \top_I.branch[9].block[3].um_I.iw[7] ,
    \top_I.branch[9].block[3].um_I.iw[6] ,
    \top_I.branch[9].block[3].um_I.iw[5] ,
    \top_I.branch[9].block[3].um_I.iw[4] ,
    \top_I.branch[9].block[3].um_I.iw[3] ,
    \top_I.branch[9].block[3].um_I.iw[2] ,
    \top_I.branch[9].block[3].um_I.iw[1] ,
    \top_I.branch[9].block[3].um_I.clk ,
    \top_I.branch[9].block[2].um_I.iw[17] ,
    \top_I.branch[9].block[2].um_I.iw[16] ,
    \top_I.branch[9].block[2].um_I.iw[15] ,
    \top_I.branch[9].block[2].um_I.iw[14] ,
    \top_I.branch[9].block[2].um_I.iw[13] ,
    \top_I.branch[9].block[2].um_I.iw[12] ,
    \top_I.branch[9].block[2].um_I.iw[11] ,
    \top_I.branch[9].block[2].um_I.iw[10] ,
    \top_I.branch[9].block[2].um_I.iw[9] ,
    \top_I.branch[9].block[2].um_I.iw[8] ,
    \top_I.branch[9].block[2].um_I.iw[7] ,
    \top_I.branch[9].block[2].um_I.iw[6] ,
    \top_I.branch[9].block[2].um_I.iw[5] ,
    \top_I.branch[9].block[2].um_I.iw[4] ,
    \top_I.branch[9].block[2].um_I.iw[3] ,
    \top_I.branch[9].block[2].um_I.iw[2] ,
    \top_I.branch[9].block[2].um_I.iw[1] ,
    \top_I.branch[9].block[2].um_I.clk ,
    \top_I.branch[9].block[1].um_I.iw[17] ,
    \top_I.branch[9].block[1].um_I.iw[16] ,
    \top_I.branch[9].block[1].um_I.iw[15] ,
    \top_I.branch[9].block[1].um_I.iw[14] ,
    \top_I.branch[9].block[1].um_I.iw[13] ,
    \top_I.branch[9].block[1].um_I.iw[12] ,
    \top_I.branch[9].block[1].um_I.iw[11] ,
    \top_I.branch[9].block[1].um_I.iw[10] ,
    \top_I.branch[9].block[1].um_I.iw[9] ,
    \top_I.branch[9].block[1].um_I.iw[8] ,
    \top_I.branch[9].block[1].um_I.iw[7] ,
    \top_I.branch[9].block[1].um_I.iw[6] ,
    \top_I.branch[9].block[1].um_I.iw[5] ,
    \top_I.branch[9].block[1].um_I.iw[4] ,
    \top_I.branch[9].block[1].um_I.iw[3] ,
    \top_I.branch[9].block[1].um_I.iw[2] ,
    \top_I.branch[9].block[1].um_I.iw[1] ,
    \top_I.branch[9].block[1].um_I.clk ,
    \top_I.branch[9].block[0].um_I.iw[17] ,
    \top_I.branch[9].block[0].um_I.iw[16] ,
    \top_I.branch[9].block[0].um_I.iw[15] ,
    \top_I.branch[9].block[0].um_I.iw[14] ,
    \top_I.branch[9].block[0].um_I.iw[13] ,
    \top_I.branch[9].block[0].um_I.iw[12] ,
    \top_I.branch[9].block[0].um_I.iw[11] ,
    \top_I.branch[9].block[0].um_I.iw[10] ,
    \top_I.branch[9].block[0].um_I.iw[9] ,
    \top_I.branch[9].block[0].um_I.iw[8] ,
    \top_I.branch[9].block[0].um_I.iw[7] ,
    \top_I.branch[9].block[0].um_I.iw[6] ,
    \top_I.branch[9].block[0].um_I.iw[5] ,
    \top_I.branch[9].block[0].um_I.iw[4] ,
    \top_I.branch[9].block[0].um_I.iw[3] ,
    \top_I.branch[9].block[0].um_I.iw[2] ,
    \top_I.branch[9].block[0].um_I.iw[1] ,
    \top_I.branch[9].block[0].um_I.clk }),
    .um_k_zero({\top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero }),
    .um_ow({\top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[15].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[14].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[13].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[12].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[11].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[10].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[9].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[8].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[7].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[6].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[5].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[4].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[3].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[2].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[1].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero ,
    \top_I.branch[9].block[0].um_I.k_zero }),
    .um_pg_vdd({\top_I.branch[9].block[15].um_I.pg_vdd ,
    \top_I.branch[9].block[14].um_I.pg_vdd ,
    \top_I.branch[9].block[13].um_I.pg_vdd ,
    \top_I.branch[9].block[12].um_I.pg_vdd ,
    \top_I.branch[9].block[11].um_I.pg_vdd ,
    \top_I.branch[9].block[10].um_I.pg_vdd ,
    \top_I.branch[9].block[9].um_I.pg_vdd ,
    \top_I.branch[9].block[8].um_I.pg_vdd ,
    \top_I.branch[9].block[7].um_I.pg_vdd ,
    \top_I.branch[9].block[6].um_I.pg_vdd ,
    \top_I.branch[9].block[5].um_I.pg_vdd ,
    \top_I.branch[9].block[4].um_I.pg_vdd ,
    \top_I.branch[9].block[3].um_I.pg_vdd ,
    \top_I.branch[9].block[2].um_I.pg_vdd ,
    \top_I.branch[9].block[1].um_I.pg_vdd ,
    \top_I.branch[9].block[0].um_I.pg_vdd }));
 tt_ctrl \top_I.ctrl_I  (.VGND(vssd1),
    .VPWR(vccd1),
    .ctrl_ena(gpio_in[38]),
    .ctrl_sel_inc(gpio_in[39]),
    .ctrl_sel_rst_n(gpio_in[40]),
    .k_one(\gpio[0].gpio_I.gpio_dm0 ),
    .k_zero(\gpio[0].gpio_I.gpio_analog_en ),
    .pad_ui_in({gpio_in[13],
    gpio_in[6],
    gpio_in[5],
    gpio_in[4],
    gpio_in[3],
    gpio_in[2],
    gpio_in[1],
    gpio_in[0],
    gpio_in[15],
    gpio_in[14]}),
    .pad_uio_in({gpio_in[23],
    gpio_in[22],
    gpio_in[21],
    gpio_in[20],
    gpio_in[19],
    gpio_in[18],
    gpio_in[17],
    gpio_in[16]}),
    .pad_uio_oe_n({gpio_oeb[23],
    gpio_oeb[22],
    gpio_oeb[21],
    gpio_oeb[20],
    gpio_oeb[19],
    gpio_oeb[18],
    gpio_oeb[17],
    gpio_oeb[16]}),
    .pad_uio_out({gpio_out[23],
    gpio_out[22],
    gpio_out[21],
    gpio_out[20],
    gpio_out[19],
    gpio_out[18],
    gpio_out[17],
    gpio_out[16]}),
    .pad_uo_out({gpio_out[31],
    gpio_out[30],
    gpio_out[29],
    gpio_out[28],
    gpio_out[27],
    gpio_out[26],
    gpio_out[25],
    gpio_out[24]}),
    .spine_bot_iw({\top_I.branch[0].l_spine_iw[29] ,
    \top_I.branch[0].l_spine_iw[28] ,
    \top_I.branch[0].l_spine_iw[27] ,
    \top_I.branch[0].l_spine_iw[26] ,
    \top_I.branch[0].l_spine_iw[25] ,
    \top_I.branch[0].l_spine_iw[24] ,
    \top_I.branch[0].l_spine_iw[23] ,
    \top_I.branch[0].l_spine_iw[22] ,
    \top_I.branch[0].l_spine_iw[21] ,
    \top_I.branch[0].l_spine_iw[20] ,
    \top_I.branch[0].l_spine_iw[19] ,
    \top_I.branch[0].l_spine_iw[18] ,
    \top_I.branch[0].l_spine_iw[17] ,
    \top_I.branch[0].l_spine_iw[16] ,
    \top_I.branch[0].l_spine_iw[15] ,
    \top_I.branch[0].l_spine_iw[14] ,
    \top_I.branch[0].l_spine_iw[13] ,
    \top_I.branch[0].l_spine_iw[12] ,
    \top_I.branch[0].l_spine_iw[11] ,
    \top_I.branch[0].l_spine_iw[10] ,
    \top_I.branch[0].l_spine_iw[9] ,
    \top_I.branch[0].l_spine_iw[8] ,
    \top_I.branch[0].l_spine_iw[7] ,
    \top_I.branch[0].l_spine_iw[6] ,
    \top_I.branch[0].l_spine_iw[5] ,
    \top_I.branch[0].l_spine_iw[4] ,
    \top_I.branch[0].l_spine_iw[3] ,
    \top_I.branch[0].l_spine_iw[2] ,
    \top_I.branch[0].l_spine_iw[1] ,
    \top_I.branch[0].l_spine_iw[0] }),
    .spine_bot_ow({\top_I.branch[0].l_spine_ow[25] ,
    \top_I.branch[0].l_spine_ow[24] ,
    \top_I.branch[0].l_spine_ow[23] ,
    \top_I.branch[0].l_spine_ow[22] ,
    \top_I.branch[0].l_spine_ow[21] ,
    \top_I.branch[0].l_spine_ow[20] ,
    \top_I.branch[0].l_spine_ow[19] ,
    \top_I.branch[0].l_spine_ow[18] ,
    \top_I.branch[0].l_spine_ow[17] ,
    \top_I.branch[0].l_spine_ow[16] ,
    \top_I.branch[0].l_spine_ow[15] ,
    \top_I.branch[0].l_spine_ow[14] ,
    \top_I.branch[0].l_spine_ow[13] ,
    \top_I.branch[0].l_spine_ow[12] ,
    \top_I.branch[0].l_spine_ow[11] ,
    \top_I.branch[0].l_spine_ow[10] ,
    \top_I.branch[0].l_spine_ow[9] ,
    \top_I.branch[0].l_spine_ow[8] ,
    \top_I.branch[0].l_spine_ow[7] ,
    \top_I.branch[0].l_spine_ow[6] ,
    \top_I.branch[0].l_spine_ow[5] ,
    \top_I.branch[0].l_spine_ow[4] ,
    \top_I.branch[0].l_spine_ow[3] ,
    \top_I.branch[0].l_spine_ow[2] ,
    \top_I.branch[0].l_spine_ow[1] ,
    \top_I.branch[0].l_spine_ow[0] }),
    .spine_top_iw({\top_I.branch[11].l_spine_iw[29] ,
    \top_I.branch[11].l_spine_iw[28] ,
    \top_I.branch[11].l_spine_iw[27] ,
    \top_I.branch[11].l_spine_iw[26] ,
    \top_I.branch[11].l_spine_iw[25] ,
    \top_I.branch[11].l_spine_iw[24] ,
    \top_I.branch[11].l_spine_iw[23] ,
    \top_I.branch[11].l_spine_iw[22] ,
    \top_I.branch[11].l_spine_iw[21] ,
    \top_I.branch[11].l_spine_iw[20] ,
    \top_I.branch[11].l_spine_iw[19] ,
    \top_I.branch[11].l_spine_iw[18] ,
    \top_I.branch[11].l_spine_iw[17] ,
    \top_I.branch[11].l_spine_iw[16] ,
    \top_I.branch[11].l_spine_iw[15] ,
    \top_I.branch[11].l_spine_iw[14] ,
    \top_I.branch[11].l_spine_iw[13] ,
    \top_I.branch[11].l_spine_iw[12] ,
    \top_I.branch[11].l_spine_iw[11] ,
    \top_I.branch[11].l_spine_iw[10] ,
    \top_I.branch[11].l_spine_iw[9] ,
    \top_I.branch[11].l_spine_iw[8] ,
    \top_I.branch[11].l_spine_iw[7] ,
    \top_I.branch[11].l_spine_iw[6] ,
    \top_I.branch[11].l_spine_iw[5] ,
    \top_I.branch[11].l_spine_iw[4] ,
    \top_I.branch[11].l_spine_iw[3] ,
    \top_I.branch[11].l_spine_iw[2] ,
    \top_I.branch[11].l_spine_iw[1] ,
    \top_I.branch[11].l_spine_iw[0] }),
    .spine_top_ow({\top_I.branch[11].l_spine_ow[25] ,
    \top_I.branch[11].l_spine_ow[24] ,
    \top_I.branch[11].l_spine_ow[23] ,
    \top_I.branch[11].l_spine_ow[22] ,
    \top_I.branch[11].l_spine_ow[21] ,
    \top_I.branch[11].l_spine_ow[20] ,
    \top_I.branch[11].l_spine_ow[19] ,
    \top_I.branch[11].l_spine_ow[18] ,
    \top_I.branch[11].l_spine_ow[17] ,
    \top_I.branch[11].l_spine_ow[16] ,
    \top_I.branch[11].l_spine_ow[15] ,
    \top_I.branch[11].l_spine_ow[14] ,
    \top_I.branch[11].l_spine_ow[13] ,
    \top_I.branch[11].l_spine_ow[12] ,
    \top_I.branch[11].l_spine_ow[11] ,
    \top_I.branch[11].l_spine_ow[10] ,
    \top_I.branch[11].l_spine_ow[9] ,
    \top_I.branch[11].l_spine_ow[8] ,
    \top_I.branch[11].l_spine_ow[7] ,
    \top_I.branch[11].l_spine_ow[6] ,
    \top_I.branch[11].l_spine_ow[5] ,
    \top_I.branch[11].l_spine_ow[4] ,
    \top_I.branch[11].l_spine_ow[3] ,
    \top_I.branch[11].l_spine_ow[2] ,
    \top_I.branch[11].l_spine_ow[1] ,
    \top_I.branch[11].l_spine_ow[0] }));
 assign gpio_analog_en[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_en[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_pol[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_analog_sel[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm1[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm2[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_holdover[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_ib_mode_sel[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_inp_dis[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_oeb[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_out[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_slow_sel[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[0] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[10] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[11] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[12] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[13] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[14] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[15] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[16] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[17] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[18] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[19] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[1] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[20] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[21] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[22] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[23] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[24] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[25] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[26] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[27] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[28] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[29] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[2] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[30] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[31] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[32] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[33] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[34] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[35] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[36] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[37] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[38] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[39] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[3] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[40] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[41] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[42] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[43] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[4] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[5] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[6] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[7] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[8] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_vtrip_sel[9] = \gpio[0].gpio_I.gpio_analog_en ;
 assign gpio_dm0[0] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[13] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[14] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[15] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[1] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[2] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[38] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[39] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[3] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[40] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[41] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[42] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[43] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[4] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[5] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm0[6] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[16] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[17] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[18] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[19] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[20] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[21] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[22] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[23] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[24] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[25] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[26] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[27] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[28] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[29] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[30] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm1[31] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[16] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[17] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[18] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[19] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[20] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[21] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[22] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[23] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[24] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[25] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[26] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[27] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[28] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[29] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[30] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_dm2[31] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[10] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[11] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[12] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[24] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[25] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[26] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[27] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[28] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[29] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[30] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[31] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[32] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[33] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[34] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[35] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[36] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[37] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[7] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[8] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_inp_dis[9] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[0] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[10] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[11] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[12] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[13] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[14] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[15] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[1] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[2] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[32] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[33] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[34] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[35] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[36] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[37] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[38] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[39] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[3] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[40] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[41] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[42] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[43] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[4] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[5] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[6] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[7] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[8] = \gpio[0].gpio_I.gpio_dm0 ;
 assign gpio_oeb[9] = \gpio[0].gpio_I.gpio_dm0 ;
endmodule
