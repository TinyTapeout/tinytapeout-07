VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_twin_tee_opamp_osc
  CLASS BLOCK ;
  FOREIGN tt_um_twin_tee_opamp_osc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 4.060000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 403.149292 ;
    ANTENNADIFFAREA 132.837051 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 61.335 207.485 61.505 207.675 ;
        RECT 62.715 207.485 62.885 207.675 ;
        RECT 68.235 207.485 68.405 207.675 ;
        RECT 61.195 206.675 62.565 207.485 ;
        RECT 62.575 206.675 68.085 207.485 ;
        RECT 68.095 206.675 69.925 207.485 ;
        RECT 70.080 207.455 70.250 207.675 ;
        RECT 73.305 207.530 73.465 207.640 ;
        RECT 74.680 207.485 74.850 207.675 ;
        RECT 77.895 207.485 78.065 207.675 ;
        RECT 79.735 207.485 79.905 207.675 ;
        RECT 83.415 207.485 83.585 207.675 ;
        RECT 86.185 207.530 86.345 207.640 ;
        RECT 87.565 207.530 87.725 207.640 ;
        RECT 89.855 207.485 90.025 207.675 ;
        RECT 91.695 207.485 91.865 207.675 ;
        RECT 92.155 207.485 92.325 207.675 ;
        RECT 95.830 207.485 96.000 207.675 ;
        RECT 96.300 207.485 96.470 207.675 ;
        RECT 99.515 207.505 99.685 207.675 ;
        RECT 99.515 207.485 99.665 207.505 ;
        RECT 100.435 207.485 100.605 207.675 ;
        RECT 111.015 207.485 111.185 207.675 ;
        RECT 112.395 207.505 112.565 207.675 ;
        RECT 113.325 207.530 113.485 207.640 ;
        RECT 115.155 207.485 115.325 207.675 ;
        RECT 72.210 207.455 73.145 207.485 ;
        RECT 70.080 207.255 73.145 207.455 ;
        RECT 69.935 206.775 73.145 207.255 ;
        RECT 69.935 206.575 70.865 206.775 ;
        RECT 72.195 206.575 73.145 206.775 ;
        RECT 74.085 206.615 74.515 207.400 ;
        RECT 74.535 206.575 77.455 207.485 ;
        RECT 77.755 206.805 79.585 207.485 ;
        RECT 79.705 206.805 83.170 207.485 ;
        RECT 78.240 206.575 79.585 206.805 ;
        RECT 82.250 206.575 83.170 206.805 ;
        RECT 83.275 206.575 86.025 207.485 ;
        RECT 86.965 206.615 87.395 207.400 ;
        RECT 88.335 206.805 90.165 207.485 ;
        RECT 90.175 206.805 92.005 207.485 ;
        RECT 92.015 206.805 94.305 207.485 ;
        RECT 88.335 206.575 89.680 206.805 ;
        RECT 90.175 206.575 91.520 206.805 ;
        RECT 93.385 206.575 94.305 206.805 ;
        RECT 94.375 206.575 96.145 207.485 ;
        RECT 96.155 206.575 97.505 207.485 ;
        RECT 97.735 206.665 99.665 207.485 ;
        RECT 97.735 206.575 98.685 206.665 ;
        RECT 99.845 206.615 100.275 207.400 ;
        RECT 100.295 206.805 107.605 207.485 ;
        RECT 103.810 206.585 104.720 206.805 ;
        RECT 106.255 206.575 107.605 206.805 ;
        RECT 107.750 206.805 111.215 207.485 ;
        RECT 107.750 206.575 108.670 206.805 ;
        RECT 112.725 206.615 113.155 207.400 ;
        RECT 114.095 206.675 115.465 207.485 ;
      LAYER nwell ;
        RECT 61.000 203.455 115.660 206.285 ;
      LAYER pwell ;
        RECT 61.195 202.255 62.565 203.065 ;
        RECT 62.575 202.255 64.405 203.065 ;
        RECT 64.415 202.935 65.760 203.165 ;
        RECT 66.255 202.935 67.600 203.165 ;
        RECT 70.750 202.935 71.670 203.165 ;
        RECT 64.415 202.255 66.245 202.935 ;
        RECT 66.255 202.255 68.085 202.935 ;
        RECT 68.205 202.255 71.670 202.935 ;
        RECT 72.235 202.935 73.580 203.165 ;
        RECT 72.235 202.255 74.065 202.935 ;
        RECT 74.085 202.340 74.515 203.125 ;
        RECT 74.535 202.255 76.350 203.165 ;
        RECT 76.375 202.255 79.295 203.165 ;
        RECT 79.690 202.935 80.610 203.165 ;
        RECT 79.690 202.255 83.155 202.935 ;
        RECT 83.285 202.255 84.635 203.165 ;
        RECT 88.170 202.935 89.080 203.155 ;
        RECT 90.615 202.935 91.965 203.165 ;
        RECT 84.655 202.255 91.965 202.935 ;
        RECT 92.110 202.935 93.030 203.165 ;
        RECT 95.895 203.075 96.845 203.165 ;
        RECT 92.110 202.255 95.575 202.935 ;
        RECT 95.895 202.255 97.825 203.075 ;
        RECT 97.995 202.255 99.810 203.165 ;
        RECT 99.845 202.340 100.275 203.125 ;
        RECT 100.390 202.935 101.310 203.165 ;
        RECT 104.895 202.935 105.815 203.165 ;
        RECT 108.645 202.935 109.575 203.155 ;
        RECT 100.390 202.255 103.855 202.935 ;
        RECT 104.895 202.255 114.085 202.935 ;
        RECT 114.095 202.255 115.465 203.065 ;
        RECT 61.335 202.045 61.505 202.255 ;
        RECT 62.715 202.065 62.885 202.255 ;
        RECT 64.550 202.045 64.720 202.235 ;
        RECT 65.935 202.065 66.105 202.255 ;
        RECT 66.395 202.045 66.565 202.235 ;
        RECT 67.775 202.065 67.945 202.255 ;
        RECT 68.235 202.065 68.405 202.255 ;
        RECT 71.910 202.095 72.030 202.205 ;
        RECT 73.755 202.045 73.925 202.255 ;
        RECT 74.210 202.045 74.380 202.235 ;
        RECT 76.055 202.065 76.225 202.255 ;
        RECT 76.520 202.065 76.690 202.255 ;
        RECT 82.495 202.045 82.665 202.235 ;
        RECT 82.955 202.065 83.125 202.255 ;
        RECT 83.870 202.045 84.040 202.235 ;
        RECT 84.335 202.045 84.505 202.255 ;
        RECT 84.795 202.065 84.965 202.255 ;
        RECT 87.555 202.045 87.725 202.235 ;
        RECT 93.535 202.045 93.705 202.235 ;
        RECT 93.995 202.045 94.165 202.235 ;
        RECT 95.375 202.065 95.545 202.255 ;
        RECT 97.675 202.235 97.825 202.255 ;
        RECT 97.675 202.065 97.845 202.235 ;
        RECT 99.515 202.065 99.685 202.255 ;
        RECT 103.655 202.065 103.825 202.255 ;
        RECT 104.125 202.100 104.285 202.210 ;
        RECT 104.575 202.045 104.745 202.235 ;
        RECT 105.035 202.045 105.205 202.235 ;
        RECT 111.040 202.065 111.210 202.235 ;
        RECT 111.040 202.045 111.150 202.065 ;
        RECT 111.480 202.045 111.650 202.235 ;
        RECT 113.325 202.090 113.485 202.200 ;
        RECT 113.775 202.065 113.945 202.255 ;
        RECT 115.155 202.045 115.325 202.255 ;
        RECT 61.195 201.235 62.565 202.045 ;
        RECT 63.515 201.135 64.865 202.045 ;
        RECT 64.875 201.135 66.690 202.045 ;
        RECT 66.755 201.365 74.065 202.045 ;
        RECT 66.755 201.135 68.105 201.365 ;
        RECT 69.640 201.145 70.550 201.365 ;
        RECT 74.095 201.135 75.445 202.045 ;
        RECT 75.495 201.365 82.805 202.045 ;
        RECT 75.495 201.135 76.845 201.365 ;
        RECT 78.380 201.145 79.290 201.365 ;
        RECT 82.835 201.135 84.185 202.045 ;
        RECT 84.195 201.135 86.945 202.045 ;
        RECT 86.965 201.175 87.395 201.960 ;
        RECT 87.415 201.135 90.165 202.045 ;
        RECT 90.270 201.365 93.735 202.045 ;
        RECT 93.855 201.365 101.165 202.045 ;
        RECT 90.270 201.135 91.190 201.365 ;
        RECT 97.370 201.145 98.280 201.365 ;
        RECT 99.815 201.135 101.165 201.365 ;
        RECT 101.310 201.365 104.775 202.045 ;
        RECT 104.895 201.365 106.725 202.045 ;
        RECT 101.310 201.135 102.230 201.365 ;
        RECT 105.380 201.135 106.725 201.365 ;
        RECT 106.735 201.365 111.150 202.045 ;
        RECT 106.735 201.135 110.665 201.365 ;
        RECT 111.335 201.135 112.685 202.045 ;
        RECT 112.725 201.175 113.155 201.960 ;
        RECT 114.095 201.235 115.465 202.045 ;
      LAYER nwell ;
        RECT 61.000 198.015 115.660 200.845 ;
      LAYER pwell ;
        RECT 61.195 196.815 62.565 197.625 ;
        RECT 63.505 196.815 64.855 197.725 ;
        RECT 64.915 197.495 66.265 197.725 ;
        RECT 67.800 197.495 68.710 197.715 ;
        RECT 72.235 197.495 73.580 197.725 ;
        RECT 64.915 196.815 72.225 197.495 ;
        RECT 72.235 196.815 74.065 197.495 ;
        RECT 74.085 196.900 74.515 197.685 ;
        RECT 78.970 197.495 79.880 197.715 ;
        RECT 81.415 197.495 82.765 197.725 ;
        RECT 75.455 196.815 82.765 197.495 ;
        RECT 82.815 197.495 84.160 197.725 ;
        RECT 82.815 196.815 84.645 197.495 ;
        RECT 84.670 196.815 86.485 197.725 ;
        RECT 90.010 197.495 90.920 197.715 ;
        RECT 92.455 197.495 93.805 197.725 ;
        RECT 86.495 196.815 93.805 197.495 ;
        RECT 93.855 197.495 94.990 197.725 ;
        RECT 97.075 197.495 97.995 197.725 ;
        RECT 93.855 196.815 97.065 197.495 ;
        RECT 97.075 196.815 99.365 197.495 ;
        RECT 99.845 196.900 100.275 197.685 ;
        RECT 100.295 196.815 103.045 197.725 ;
        RECT 106.570 197.495 107.480 197.715 ;
        RECT 109.015 197.495 110.365 197.725 ;
        RECT 103.055 196.815 110.365 197.495 ;
        RECT 110.510 197.495 111.430 197.725 ;
        RECT 110.510 196.815 113.975 197.495 ;
        RECT 114.095 196.815 115.465 197.625 ;
        RECT 61.335 196.605 61.505 196.815 ;
        RECT 62.715 196.605 62.885 196.795 ;
        RECT 64.555 196.625 64.725 196.815 ;
        RECT 68.235 196.605 68.405 196.795 ;
        RECT 70.070 196.655 70.190 196.765 ;
        RECT 70.540 196.605 70.710 196.795 ;
        RECT 71.915 196.625 72.085 196.815 ;
        RECT 73.755 196.625 73.925 196.815 ;
        RECT 74.685 196.660 74.845 196.770 ;
        RECT 75.595 196.625 75.765 196.815 ;
        RECT 76.515 196.605 76.685 196.795 ;
        RECT 84.335 196.625 84.505 196.815 ;
        RECT 84.795 196.625 84.965 196.815 ;
        RECT 85.715 196.605 85.885 196.795 ;
        RECT 86.185 196.650 86.345 196.760 ;
        RECT 86.635 196.625 86.805 196.815 ;
        RECT 88.475 196.605 88.645 196.795 ;
        RECT 96.755 196.625 96.925 196.815 ;
        RECT 97.675 196.605 97.845 196.795 ;
        RECT 98.130 196.655 98.250 196.765 ;
        RECT 98.595 196.605 98.765 196.795 ;
        RECT 99.055 196.625 99.225 196.815 ;
        RECT 99.510 196.655 99.630 196.765 ;
        RECT 101.355 196.605 101.525 196.795 ;
        RECT 102.735 196.625 102.905 196.815 ;
        RECT 103.195 196.625 103.365 196.815 ;
        RECT 112.395 196.625 112.565 196.795 ;
        RECT 113.325 196.650 113.485 196.760 ;
        RECT 113.775 196.625 113.945 196.815 ;
        RECT 112.395 196.605 112.545 196.625 ;
        RECT 115.155 196.605 115.325 196.815 ;
        RECT 61.195 195.795 62.565 196.605 ;
        RECT 62.575 195.795 68.085 196.605 ;
        RECT 68.095 195.795 69.925 196.605 ;
        RECT 70.395 195.695 73.315 196.605 ;
        RECT 74.535 195.925 76.825 196.605 ;
        RECT 76.920 195.925 86.025 196.605 ;
        RECT 74.535 195.695 75.455 195.925 ;
        RECT 86.965 195.735 87.395 196.520 ;
        RECT 87.415 195.825 88.785 196.605 ;
        RECT 88.880 195.925 97.985 196.605 ;
        RECT 98.455 195.695 101.205 196.605 ;
        RECT 101.215 195.925 110.320 196.605 ;
        RECT 110.615 195.785 112.545 196.605 ;
        RECT 110.615 195.695 111.565 195.785 ;
        RECT 112.725 195.735 113.155 196.520 ;
        RECT 114.095 195.795 115.465 196.605 ;
      LAYER nwell ;
        RECT 61.000 192.575 115.660 195.405 ;
      LAYER pwell ;
        RECT 61.195 191.375 62.565 192.185 ;
        RECT 62.575 191.375 68.085 192.185 ;
        RECT 68.095 191.375 71.765 192.185 ;
        RECT 72.695 191.375 74.065 192.155 ;
        RECT 74.085 191.460 74.515 192.245 ;
        RECT 74.555 191.375 75.905 192.285 ;
        RECT 75.975 191.375 77.745 192.285 ;
        RECT 77.755 191.375 79.570 192.285 ;
        RECT 79.690 192.055 80.610 192.285 ;
        RECT 85.350 192.055 86.485 192.285 ;
        RECT 79.690 191.375 83.155 192.055 ;
        RECT 83.275 191.375 86.485 192.055 ;
        RECT 86.495 191.375 88.325 192.055 ;
        RECT 88.335 191.375 91.085 192.285 ;
        RECT 91.275 191.605 93.610 192.285 ;
        RECT 94.995 192.195 95.945 192.285 ;
        RECT 91.275 191.375 93.125 191.605 ;
        RECT 94.015 191.375 95.945 192.195 ;
        RECT 97.075 191.375 99.825 192.285 ;
        RECT 99.845 191.460 100.275 192.245 ;
        RECT 100.295 191.375 103.045 192.285 ;
        RECT 106.570 192.055 107.480 192.275 ;
        RECT 109.015 192.055 110.365 192.285 ;
        RECT 103.055 191.375 110.365 192.055 ;
        RECT 110.510 192.055 111.430 192.285 ;
        RECT 110.510 191.375 113.975 192.055 ;
        RECT 114.095 191.375 115.465 192.185 ;
        RECT 61.335 191.165 61.505 191.375 ;
        RECT 62.715 191.165 62.885 191.375 ;
        RECT 68.235 191.165 68.405 191.375 ;
        RECT 70.990 191.215 71.110 191.325 ;
        RECT 71.455 191.165 71.625 191.355 ;
        RECT 71.925 191.220 72.085 191.330 ;
        RECT 73.755 191.185 73.925 191.375 ;
        RECT 74.215 191.165 74.385 191.355 ;
        RECT 75.590 191.185 75.760 191.375 ;
        RECT 77.430 191.185 77.600 191.375 ;
        RECT 79.275 191.185 79.445 191.375 ;
        RECT 81.585 191.210 81.745 191.320 ;
        RECT 82.955 191.185 83.125 191.375 ;
        RECT 83.415 191.185 83.585 191.375 ;
        RECT 85.715 191.165 85.885 191.355 ;
        RECT 86.185 191.210 86.345 191.320 ;
        RECT 88.015 191.185 88.185 191.375 ;
        RECT 88.475 191.185 88.645 191.375 ;
        RECT 91.275 191.355 91.405 191.375 ;
        RECT 94.015 191.355 94.165 191.375 ;
        RECT 90.775 191.165 90.945 191.355 ;
        RECT 91.235 191.185 91.405 191.355 ;
        RECT 93.995 191.185 94.165 191.355 ;
        RECT 95.375 191.165 95.545 191.355 ;
        RECT 95.840 191.165 96.010 191.355 ;
        RECT 96.305 191.220 96.465 191.330 ;
        RECT 97.215 191.185 97.385 191.375 ;
        RECT 99.055 191.165 99.225 191.355 ;
        RECT 100.435 191.185 100.605 191.375 ;
        RECT 102.285 191.210 102.445 191.320 ;
        RECT 103.195 191.185 103.365 191.375 ;
        RECT 106.415 191.165 106.585 191.355 ;
        RECT 106.875 191.165 107.045 191.355 ;
        RECT 112.395 191.165 112.565 191.355 ;
        RECT 113.325 191.210 113.485 191.320 ;
        RECT 113.775 191.185 113.945 191.375 ;
        RECT 115.155 191.165 115.325 191.375 ;
        RECT 61.195 190.355 62.565 191.165 ;
        RECT 62.575 190.355 68.085 191.165 ;
        RECT 68.095 190.355 70.845 191.165 ;
        RECT 71.315 190.255 74.065 191.165 ;
        RECT 74.075 190.485 81.385 191.165 ;
        RECT 77.590 190.265 78.500 190.485 ;
        RECT 80.035 190.255 81.385 190.485 ;
        RECT 82.450 190.485 85.915 191.165 ;
        RECT 82.450 190.255 83.370 190.485 ;
        RECT 86.965 190.295 87.395 191.080 ;
        RECT 87.510 190.485 90.975 191.165 ;
        RECT 92.110 190.485 95.575 191.165 ;
        RECT 87.510 190.255 88.430 190.485 ;
        RECT 92.110 190.255 93.030 190.485 ;
        RECT 95.695 190.255 98.615 191.165 ;
        RECT 98.915 190.485 102.125 191.165 ;
        RECT 100.990 190.255 102.125 190.485 ;
        RECT 103.150 190.485 106.615 191.165 ;
        RECT 103.150 190.255 104.070 190.485 ;
        RECT 106.735 190.255 109.485 191.165 ;
        RECT 109.495 190.485 112.705 191.165 ;
        RECT 109.495 190.255 110.630 190.485 ;
        RECT 112.725 190.295 113.155 191.080 ;
        RECT 114.095 190.355 115.465 191.165 ;
      LAYER nwell ;
        RECT 61.000 187.135 115.660 189.965 ;
      LAYER pwell ;
        RECT 61.195 185.935 62.565 186.745 ;
        RECT 62.575 185.935 66.245 186.745 ;
        RECT 69.370 186.615 70.290 186.845 ;
        RECT 66.825 185.935 70.290 186.615 ;
        RECT 70.490 186.615 71.410 186.845 ;
        RECT 70.490 185.935 73.955 186.615 ;
        RECT 74.085 186.020 74.515 186.805 ;
        RECT 75.905 186.615 76.825 186.845 ;
        RECT 80.350 186.615 81.260 186.835 ;
        RECT 82.795 186.615 84.145 186.845 ;
        RECT 74.535 185.935 76.825 186.615 ;
        RECT 76.835 185.935 84.145 186.615 ;
        RECT 84.195 185.935 86.010 186.845 ;
        RECT 90.010 186.615 90.920 186.835 ;
        RECT 92.455 186.615 93.805 186.845 ;
        RECT 86.495 185.935 93.805 186.615 ;
        RECT 93.855 185.935 95.670 186.845 ;
        RECT 98.810 186.615 99.730 186.845 ;
        RECT 96.265 185.935 99.730 186.615 ;
        RECT 99.845 186.020 100.275 186.805 ;
        RECT 100.295 186.615 104.225 186.845 ;
        RECT 100.295 185.935 104.710 186.615 ;
        RECT 104.895 185.935 106.245 186.845 ;
        RECT 106.370 186.615 107.290 186.845 ;
        RECT 112.610 186.615 113.530 186.845 ;
        RECT 106.370 185.935 109.835 186.615 ;
        RECT 110.065 185.935 113.530 186.615 ;
        RECT 114.095 185.935 115.465 186.745 ;
        RECT 61.335 185.725 61.505 185.935 ;
        RECT 62.715 185.725 62.885 185.935 ;
        RECT 66.390 185.775 66.510 185.885 ;
        RECT 66.855 185.745 67.025 185.935 ;
        RECT 68.235 185.725 68.405 185.915 ;
        RECT 69.615 185.725 69.785 185.915 ;
        RECT 73.755 185.745 73.925 185.935 ;
        RECT 74.675 185.745 74.845 185.935 ;
        RECT 76.975 185.725 77.145 185.935 ;
        RECT 85.250 185.725 85.420 185.915 ;
        RECT 85.715 185.725 85.885 185.935 ;
        RECT 86.170 185.775 86.290 185.885 ;
        RECT 86.635 185.745 86.805 185.935 ;
        RECT 87.555 185.725 87.725 185.915 ;
        RECT 89.850 185.725 90.020 185.915 ;
        RECT 90.315 185.725 90.485 185.915 ;
        RECT 95.375 185.745 95.545 185.935 ;
        RECT 95.830 185.775 95.950 185.885 ;
        RECT 96.295 185.745 96.465 185.935 ;
        RECT 104.600 185.915 104.710 185.935 ;
        RECT 105.040 185.915 105.210 185.935 ;
        RECT 97.675 185.725 97.845 185.915 ;
        RECT 104.600 185.745 104.770 185.915 ;
        RECT 105.035 185.745 105.210 185.915 ;
        RECT 109.635 185.745 109.805 185.935 ;
        RECT 110.095 185.745 110.265 185.935 ;
        RECT 112.390 185.775 112.510 185.885 ;
        RECT 113.325 185.770 113.485 185.880 ;
        RECT 113.770 185.775 113.890 185.885 ;
        RECT 105.035 185.725 105.205 185.745 ;
        RECT 115.155 185.725 115.325 185.935 ;
        RECT 61.195 184.915 62.565 185.725 ;
        RECT 62.575 184.915 68.085 185.725 ;
        RECT 68.095 184.915 69.465 185.725 ;
        RECT 69.475 185.045 76.785 185.725 ;
        RECT 76.835 185.045 84.145 185.725 ;
        RECT 72.990 184.825 73.900 185.045 ;
        RECT 75.435 184.815 76.785 185.045 ;
        RECT 80.350 184.825 81.260 185.045 ;
        RECT 82.795 184.815 84.145 185.045 ;
        RECT 84.215 184.815 85.565 185.725 ;
        RECT 85.575 184.915 86.945 185.725 ;
        RECT 86.965 184.855 87.395 185.640 ;
        RECT 87.415 184.915 88.785 185.725 ;
        RECT 88.815 184.815 90.165 185.725 ;
        RECT 90.175 185.045 97.485 185.725 ;
        RECT 97.535 185.045 104.845 185.725 ;
        RECT 104.895 185.045 112.205 185.725 ;
        RECT 93.690 184.825 94.600 185.045 ;
        RECT 96.135 184.815 97.485 185.045 ;
        RECT 101.050 184.825 101.960 185.045 ;
        RECT 103.495 184.815 104.845 185.045 ;
        RECT 108.410 184.825 109.320 185.045 ;
        RECT 110.855 184.815 112.205 185.045 ;
        RECT 112.725 184.855 113.155 185.640 ;
        RECT 114.095 184.915 115.465 185.725 ;
      LAYER nwell ;
        RECT 61.000 181.695 115.660 184.525 ;
      LAYER pwell ;
        RECT 61.195 180.495 62.565 181.305 ;
        RECT 62.575 180.495 68.085 181.305 ;
        RECT 68.095 180.495 73.605 181.305 ;
        RECT 74.085 180.580 74.515 181.365 ;
        RECT 74.535 180.495 76.365 181.305 ;
        RECT 76.850 180.495 78.665 181.405 ;
        RECT 79.135 180.495 81.885 181.405 ;
        RECT 82.910 181.175 83.830 181.405 ;
        RECT 90.930 181.175 91.840 181.395 ;
        RECT 93.375 181.175 94.725 181.405 ;
        RECT 98.350 181.175 99.270 181.405 ;
        RECT 82.910 180.495 86.375 181.175 ;
        RECT 87.415 180.495 94.725 181.175 ;
        RECT 95.805 180.495 99.270 181.175 ;
        RECT 99.845 180.580 100.275 181.365 ;
        RECT 101.215 181.175 102.560 181.405 ;
        RECT 101.215 180.495 103.045 181.175 ;
        RECT 103.055 180.495 105.805 181.405 ;
        RECT 105.855 181.175 107.205 181.405 ;
        RECT 108.740 181.175 109.650 181.395 ;
        RECT 105.855 180.495 113.165 181.175 ;
        RECT 114.095 180.495 115.465 181.305 ;
        RECT 61.335 180.285 61.505 180.495 ;
        RECT 62.715 180.285 62.885 180.495 ;
        RECT 68.235 180.285 68.405 180.495 ;
        RECT 73.755 180.445 73.925 180.475 ;
        RECT 73.750 180.335 73.925 180.445 ;
        RECT 73.755 180.285 73.925 180.335 ;
        RECT 74.675 180.305 74.845 180.495 ;
        RECT 76.510 180.335 76.630 180.445 ;
        RECT 76.975 180.305 77.145 180.495 ;
        RECT 78.810 180.335 78.930 180.445 ;
        RECT 79.275 180.285 79.445 180.495 ;
        RECT 82.045 180.340 82.205 180.450 ;
        RECT 84.795 180.285 84.965 180.475 ;
        RECT 86.175 180.305 86.345 180.495 ;
        RECT 86.645 180.445 86.805 180.450 ;
        RECT 86.630 180.340 86.805 180.445 ;
        RECT 86.630 180.335 86.750 180.340 ;
        RECT 87.555 180.285 87.725 180.495 ;
        RECT 93.075 180.285 93.245 180.475 ;
        RECT 94.915 180.305 95.085 180.475 ;
        RECT 95.835 180.305 96.005 180.495 ;
        RECT 102.735 180.475 102.905 180.495 ;
        RECT 94.935 180.285 95.085 180.305 ;
        RECT 97.215 180.285 97.385 180.475 ;
        RECT 99.510 180.335 99.630 180.445 ;
        RECT 100.445 180.340 100.605 180.450 ;
        RECT 100.905 180.330 101.065 180.440 ;
        RECT 102.730 180.305 102.905 180.475 ;
        RECT 103.195 180.305 103.365 180.495 ;
        RECT 102.730 180.285 102.900 180.305 ;
        RECT 105.495 180.285 105.665 180.475 ;
        RECT 105.955 180.285 106.125 180.475 ;
        RECT 107.335 180.285 107.505 180.475 ;
        RECT 111.015 180.285 111.185 180.475 ;
        RECT 112.855 180.305 113.025 180.495 ;
        RECT 113.325 180.330 113.485 180.450 ;
        RECT 115.155 180.285 115.325 180.495 ;
        RECT 61.195 179.475 62.565 180.285 ;
        RECT 62.575 179.475 68.085 180.285 ;
        RECT 68.095 179.475 73.605 180.285 ;
        RECT 73.615 179.475 79.125 180.285 ;
        RECT 79.135 179.475 84.645 180.285 ;
        RECT 84.655 179.475 86.485 180.285 ;
        RECT 86.965 179.415 87.395 180.200 ;
        RECT 87.415 179.475 92.925 180.285 ;
        RECT 92.935 179.475 94.765 180.285 ;
        RECT 94.935 179.465 96.865 180.285 ;
        RECT 97.075 179.475 100.745 180.285 ;
        RECT 95.915 179.375 96.865 179.465 ;
        RECT 101.695 179.375 103.045 180.285 ;
        RECT 103.975 179.375 105.790 180.285 ;
        RECT 105.815 179.475 107.185 180.285 ;
        RECT 107.305 179.605 110.770 180.285 ;
        RECT 109.850 179.375 110.770 179.605 ;
        RECT 110.890 179.375 112.705 180.285 ;
        RECT 112.725 179.415 113.155 180.200 ;
        RECT 114.095 179.475 115.465 180.285 ;
      LAYER nwell ;
        RECT 61.000 176.255 115.660 179.085 ;
      LAYER pwell ;
        RECT 61.195 175.055 62.565 175.865 ;
        RECT 62.575 175.055 68.085 175.865 ;
        RECT 68.095 175.055 73.605 175.865 ;
        RECT 74.085 175.140 74.515 175.925 ;
        RECT 74.535 175.055 80.045 175.865 ;
        RECT 80.055 175.055 85.565 175.865 ;
        RECT 85.575 175.055 91.085 175.865 ;
        RECT 91.095 175.055 96.605 175.865 ;
        RECT 96.615 175.055 99.365 175.865 ;
        RECT 99.845 175.140 100.275 175.925 ;
        RECT 109.255 175.875 110.205 175.965 ;
        RECT 100.295 175.055 105.805 175.865 ;
        RECT 105.815 175.055 107.645 175.865 ;
        RECT 108.275 175.055 110.205 175.875 ;
        RECT 110.415 175.735 111.335 175.965 ;
        RECT 110.415 175.055 112.705 175.735 ;
        RECT 112.715 175.055 114.085 175.865 ;
        RECT 114.095 175.055 115.465 175.865 ;
        RECT 61.335 174.845 61.505 175.055 ;
        RECT 62.715 174.845 62.885 175.055 ;
        RECT 68.235 174.845 68.405 175.055 ;
        RECT 73.755 175.005 73.925 175.035 ;
        RECT 73.750 174.895 73.925 175.005 ;
        RECT 73.755 174.845 73.925 174.895 ;
        RECT 74.675 174.865 74.845 175.055 ;
        RECT 79.275 174.845 79.445 175.035 ;
        RECT 80.195 174.865 80.365 175.055 ;
        RECT 84.795 174.845 84.965 175.035 ;
        RECT 85.715 174.865 85.885 175.055 ;
        RECT 86.630 174.895 86.750 175.005 ;
        RECT 87.555 174.845 87.725 175.035 ;
        RECT 91.235 174.865 91.405 175.055 ;
        RECT 93.075 174.845 93.245 175.035 ;
        RECT 96.755 174.865 96.925 175.055 ;
        RECT 98.595 174.845 98.765 175.035 ;
        RECT 99.510 174.895 99.630 175.005 ;
        RECT 100.435 174.865 100.605 175.055 ;
        RECT 104.115 174.845 104.285 175.035 ;
        RECT 105.955 174.865 106.125 175.055 ;
        RECT 108.275 175.035 108.425 175.055 ;
        RECT 112.395 175.035 112.565 175.055 ;
        RECT 107.790 174.895 107.910 175.005 ;
        RECT 108.255 174.865 108.425 175.035 ;
        RECT 109.635 174.845 109.805 175.035 ;
        RECT 112.390 174.865 112.565 175.035 ;
        RECT 112.855 174.865 113.025 175.055 ;
        RECT 113.325 174.890 113.485 175.000 ;
        RECT 112.390 174.845 112.560 174.865 ;
        RECT 115.155 174.845 115.325 175.055 ;
        RECT 61.195 174.035 62.565 174.845 ;
        RECT 62.575 174.035 68.085 174.845 ;
        RECT 68.095 174.035 73.605 174.845 ;
        RECT 73.615 174.035 79.125 174.845 ;
        RECT 79.135 174.035 84.645 174.845 ;
        RECT 84.655 174.035 86.485 174.845 ;
        RECT 86.965 173.975 87.395 174.760 ;
        RECT 87.415 174.035 92.925 174.845 ;
        RECT 92.935 174.035 98.445 174.845 ;
        RECT 98.455 174.035 103.965 174.845 ;
        RECT 103.975 174.035 109.485 174.845 ;
        RECT 109.495 174.035 110.865 174.845 ;
        RECT 110.935 173.935 112.705 174.845 ;
        RECT 112.725 173.975 113.155 174.760 ;
        RECT 114.095 174.035 115.465 174.845 ;
      LAYER nwell ;
        RECT 61.000 170.815 115.660 173.645 ;
      LAYER pwell ;
        RECT 61.195 169.615 62.565 170.425 ;
        RECT 62.575 169.615 68.085 170.425 ;
        RECT 68.095 169.615 73.605 170.425 ;
        RECT 74.085 169.700 74.515 170.485 ;
        RECT 74.535 169.615 80.045 170.425 ;
        RECT 80.055 169.615 85.565 170.425 ;
        RECT 85.575 169.615 91.085 170.425 ;
        RECT 91.095 169.615 96.605 170.425 ;
        RECT 96.615 169.615 99.365 170.425 ;
        RECT 99.845 169.700 100.275 170.485 ;
        RECT 100.295 169.615 105.805 170.425 ;
        RECT 105.815 169.615 111.325 170.425 ;
        RECT 111.335 169.615 114.085 170.425 ;
        RECT 114.095 169.615 115.465 170.425 ;
        RECT 61.335 169.405 61.505 169.615 ;
        RECT 62.715 169.405 62.885 169.615 ;
        RECT 68.235 169.405 68.405 169.615 ;
        RECT 73.755 169.565 73.925 169.595 ;
        RECT 73.750 169.455 73.925 169.565 ;
        RECT 73.755 169.405 73.925 169.455 ;
        RECT 74.675 169.425 74.845 169.615 ;
        RECT 79.275 169.405 79.445 169.595 ;
        RECT 80.195 169.425 80.365 169.615 ;
        RECT 84.795 169.405 84.965 169.595 ;
        RECT 85.715 169.425 85.885 169.615 ;
        RECT 86.630 169.455 86.750 169.565 ;
        RECT 87.555 169.405 87.725 169.595 ;
        RECT 91.235 169.425 91.405 169.615 ;
        RECT 93.075 169.405 93.245 169.595 ;
        RECT 96.755 169.425 96.925 169.615 ;
        RECT 98.595 169.405 98.765 169.595 ;
        RECT 99.510 169.455 99.630 169.565 ;
        RECT 100.435 169.425 100.605 169.615 ;
        RECT 104.115 169.405 104.285 169.595 ;
        RECT 105.955 169.425 106.125 169.615 ;
        RECT 109.635 169.405 109.805 169.595 ;
        RECT 111.475 169.425 111.645 169.615 ;
        RECT 112.390 169.455 112.510 169.565 ;
        RECT 113.325 169.450 113.485 169.560 ;
        RECT 115.155 169.405 115.325 169.615 ;
        RECT 61.195 168.595 62.565 169.405 ;
        RECT 62.575 168.595 68.085 169.405 ;
        RECT 68.095 168.595 73.605 169.405 ;
        RECT 73.615 168.595 79.125 169.405 ;
        RECT 79.135 168.595 84.645 169.405 ;
        RECT 84.655 168.595 86.485 169.405 ;
        RECT 86.965 168.535 87.395 169.320 ;
        RECT 87.415 168.595 92.925 169.405 ;
        RECT 92.935 168.595 98.445 169.405 ;
        RECT 98.455 168.595 103.965 169.405 ;
        RECT 103.975 168.595 109.485 169.405 ;
        RECT 109.495 168.595 112.245 169.405 ;
        RECT 112.725 168.535 113.155 169.320 ;
        RECT 114.095 168.595 115.465 169.405 ;
      LAYER nwell ;
        RECT 61.000 165.375 115.660 168.205 ;
      LAYER pwell ;
        RECT 61.195 164.175 62.565 164.985 ;
        RECT 62.575 164.175 68.085 164.985 ;
        RECT 68.095 164.175 73.605 164.985 ;
        RECT 74.085 164.260 74.515 165.045 ;
        RECT 74.535 164.175 80.045 164.985 ;
        RECT 80.055 164.175 85.565 164.985 ;
        RECT 85.575 164.175 91.085 164.985 ;
        RECT 91.095 164.175 96.605 164.985 ;
        RECT 96.615 164.175 99.365 164.985 ;
        RECT 99.845 164.260 100.275 165.045 ;
        RECT 100.295 164.175 105.805 164.985 ;
        RECT 105.815 164.175 111.325 164.985 ;
        RECT 111.335 164.175 114.085 164.985 ;
        RECT 114.095 164.175 115.465 164.985 ;
        RECT 61.335 163.965 61.505 164.175 ;
        RECT 62.715 163.965 62.885 164.175 ;
        RECT 68.235 163.965 68.405 164.175 ;
        RECT 73.755 164.125 73.925 164.155 ;
        RECT 73.750 164.015 73.925 164.125 ;
        RECT 73.755 163.965 73.925 164.015 ;
        RECT 74.675 163.985 74.845 164.175 ;
        RECT 79.275 163.965 79.445 164.155 ;
        RECT 80.195 163.985 80.365 164.175 ;
        RECT 84.795 163.965 84.965 164.155 ;
        RECT 85.715 163.985 85.885 164.175 ;
        RECT 86.630 164.015 86.750 164.125 ;
        RECT 87.555 163.965 87.725 164.155 ;
        RECT 91.235 163.985 91.405 164.175 ;
        RECT 93.075 163.965 93.245 164.155 ;
        RECT 96.755 163.985 96.925 164.175 ;
        RECT 98.595 163.965 98.765 164.155 ;
        RECT 99.510 164.015 99.630 164.125 ;
        RECT 100.435 163.985 100.605 164.175 ;
        RECT 104.115 163.965 104.285 164.155 ;
        RECT 105.955 163.985 106.125 164.175 ;
        RECT 109.635 163.965 109.805 164.155 ;
        RECT 111.475 163.985 111.645 164.175 ;
        RECT 112.390 164.015 112.510 164.125 ;
        RECT 113.325 164.010 113.485 164.120 ;
        RECT 115.155 163.965 115.325 164.175 ;
        RECT 61.195 163.155 62.565 163.965 ;
        RECT 62.575 163.155 68.085 163.965 ;
        RECT 68.095 163.155 73.605 163.965 ;
        RECT 73.615 163.155 79.125 163.965 ;
        RECT 79.135 163.155 84.645 163.965 ;
        RECT 84.655 163.155 86.485 163.965 ;
        RECT 86.965 163.095 87.395 163.880 ;
        RECT 87.415 163.155 92.925 163.965 ;
        RECT 92.935 163.155 98.445 163.965 ;
        RECT 98.455 163.155 103.965 163.965 ;
        RECT 103.975 163.155 109.485 163.965 ;
        RECT 109.495 163.155 112.245 163.965 ;
        RECT 112.725 163.095 113.155 163.880 ;
        RECT 114.095 163.155 115.465 163.965 ;
      LAYER nwell ;
        RECT 61.000 159.935 115.660 162.765 ;
      LAYER pwell ;
        RECT 61.195 158.735 62.565 159.545 ;
        RECT 62.575 158.735 68.085 159.545 ;
        RECT 68.095 158.735 73.605 159.545 ;
        RECT 74.085 158.820 74.515 159.605 ;
        RECT 74.535 158.735 80.045 159.545 ;
        RECT 80.055 158.735 85.565 159.545 ;
        RECT 85.575 158.735 91.085 159.545 ;
        RECT 91.095 158.735 96.605 159.545 ;
        RECT 96.615 158.735 99.365 159.545 ;
        RECT 99.845 158.820 100.275 159.605 ;
        RECT 100.295 158.735 105.805 159.545 ;
        RECT 105.815 158.735 111.325 159.545 ;
        RECT 111.335 158.735 114.085 159.545 ;
        RECT 114.095 158.735 115.465 159.545 ;
        RECT 61.335 158.525 61.505 158.735 ;
        RECT 62.715 158.525 62.885 158.735 ;
        RECT 68.235 158.525 68.405 158.735 ;
        RECT 73.755 158.685 73.925 158.715 ;
        RECT 73.750 158.575 73.925 158.685 ;
        RECT 73.755 158.525 73.925 158.575 ;
        RECT 74.675 158.545 74.845 158.735 ;
        RECT 79.275 158.525 79.445 158.715 ;
        RECT 80.195 158.545 80.365 158.735 ;
        RECT 84.795 158.525 84.965 158.715 ;
        RECT 85.715 158.545 85.885 158.735 ;
        RECT 86.630 158.575 86.750 158.685 ;
        RECT 87.555 158.525 87.725 158.715 ;
        RECT 91.235 158.545 91.405 158.735 ;
        RECT 93.075 158.525 93.245 158.715 ;
        RECT 96.755 158.545 96.925 158.735 ;
        RECT 98.595 158.525 98.765 158.715 ;
        RECT 99.510 158.575 99.630 158.685 ;
        RECT 100.435 158.545 100.605 158.735 ;
        RECT 104.115 158.525 104.285 158.715 ;
        RECT 105.955 158.545 106.125 158.735 ;
        RECT 109.635 158.525 109.805 158.715 ;
        RECT 111.475 158.545 111.645 158.735 ;
        RECT 112.390 158.575 112.510 158.685 ;
        RECT 113.325 158.570 113.485 158.680 ;
        RECT 115.155 158.525 115.325 158.735 ;
        RECT 61.195 157.715 62.565 158.525 ;
        RECT 62.575 157.715 68.085 158.525 ;
        RECT 68.095 157.715 73.605 158.525 ;
        RECT 73.615 157.715 79.125 158.525 ;
        RECT 79.135 157.715 84.645 158.525 ;
        RECT 84.655 157.715 86.485 158.525 ;
        RECT 86.965 157.655 87.395 158.440 ;
        RECT 87.415 157.715 92.925 158.525 ;
        RECT 92.935 157.715 98.445 158.525 ;
        RECT 98.455 157.715 103.965 158.525 ;
        RECT 103.975 157.715 109.485 158.525 ;
        RECT 109.495 157.715 112.245 158.525 ;
        RECT 112.725 157.655 113.155 158.440 ;
        RECT 114.095 157.715 115.465 158.525 ;
      LAYER nwell ;
        RECT 61.000 154.495 115.660 157.325 ;
      LAYER pwell ;
        RECT 61.195 153.295 62.565 154.105 ;
        RECT 62.575 153.295 68.085 154.105 ;
        RECT 68.095 153.295 73.605 154.105 ;
        RECT 74.085 153.380 74.515 154.165 ;
        RECT 74.535 153.295 80.045 154.105 ;
        RECT 80.055 153.295 85.565 154.105 ;
        RECT 85.575 153.295 86.945 154.105 ;
        RECT 86.965 153.380 87.395 154.165 ;
        RECT 87.415 153.295 92.925 154.105 ;
        RECT 92.935 153.295 98.445 154.105 ;
        RECT 98.455 153.295 99.825 154.105 ;
        RECT 99.845 153.380 100.275 154.165 ;
        RECT 100.295 153.295 105.805 154.105 ;
        RECT 105.815 153.295 111.325 154.105 ;
        RECT 111.335 153.295 112.705 154.105 ;
        RECT 112.725 153.380 113.155 154.165 ;
        RECT 114.095 153.295 115.465 154.105 ;
        RECT 61.335 153.105 61.505 153.295 ;
        RECT 62.715 153.105 62.885 153.295 ;
        RECT 68.235 153.105 68.405 153.295 ;
        RECT 73.750 153.135 73.870 153.245 ;
        RECT 74.675 153.105 74.845 153.295 ;
        RECT 80.195 153.105 80.365 153.295 ;
        RECT 85.715 153.105 85.885 153.295 ;
        RECT 87.555 153.105 87.725 153.295 ;
        RECT 93.075 153.105 93.245 153.295 ;
        RECT 98.595 153.105 98.765 153.295 ;
        RECT 100.435 153.105 100.605 153.295 ;
        RECT 105.955 153.105 106.125 153.295 ;
        RECT 111.475 153.105 111.645 153.295 ;
        RECT 113.325 153.140 113.485 153.250 ;
        RECT 115.155 153.105 115.325 153.295 ;
        RECT 130.800 94.380 143.260 99.710 ;
        RECT 111.940 88.090 124.400 93.420 ;
        RECT 114.560 48.010 143.540 50.020 ;
        RECT 114.890 15.660 116.900 41.640 ;
        RECT 118.940 15.860 120.950 41.840 ;
        RECT 126.840 34.010 128.850 42.890 ;
        RECT 126.290 22.360 129.390 33.190 ;
      LAYER nwell ;
        RECT 130.890 28.410 134.080 43.820 ;
        RECT 137.240 28.410 140.430 43.820 ;
      LAYER pwell ;
        RECT 131.040 25.560 140.240 28.020 ;
      LAYER nwell ;
        RECT 141.840 26.610 145.030 44.080 ;
      LAYER pwell ;
        RECT 137.840 25.510 138.390 25.560 ;
        RECT 130.340 22.410 141.170 25.510 ;
        RECT 145.840 22.410 148.940 40.110 ;
      LAYER li1 ;
        RECT 61.190 207.505 115.470 207.675 ;
        RECT 61.275 206.755 62.485 207.505 ;
        RECT 62.655 206.960 68.000 207.505 ;
        RECT 61.275 206.215 61.795 206.755 ;
        RECT 61.965 206.045 62.485 206.585 ;
        RECT 64.240 206.130 64.580 206.960 ;
        RECT 68.175 206.735 69.845 207.505 ;
        RECT 61.275 204.955 62.485 206.045 ;
        RECT 66.060 205.390 66.410 206.640 ;
        RECT 68.175 206.215 68.925 206.735 ;
        RECT 70.015 206.685 70.275 207.505 ;
        RECT 70.445 206.685 70.775 207.105 ;
        RECT 70.955 207.020 71.745 207.285 ;
        RECT 70.525 206.595 70.775 206.685 ;
        RECT 69.095 206.045 69.845 206.565 ;
        RECT 62.655 204.955 68.000 205.390 ;
        RECT 68.175 204.955 69.845 206.045 ;
        RECT 70.015 205.635 70.355 206.515 ;
        RECT 70.525 206.345 71.320 206.595 ;
        RECT 70.015 204.955 70.275 205.465 ;
        RECT 70.525 205.125 70.695 206.345 ;
        RECT 71.490 206.165 71.745 207.020 ;
        RECT 71.915 206.865 72.115 207.285 ;
        RECT 72.305 207.045 72.635 207.505 ;
        RECT 71.915 206.345 72.325 206.865 ;
        RECT 72.805 206.855 73.065 207.335 ;
        RECT 72.495 206.165 72.725 206.595 ;
        RECT 70.935 205.995 72.725 206.165 ;
        RECT 70.935 205.630 71.185 205.995 ;
        RECT 71.355 205.635 71.685 205.825 ;
        RECT 71.905 205.700 72.620 205.995 ;
        RECT 72.895 205.825 73.065 206.855 ;
        RECT 74.155 206.780 74.445 207.505 ;
        RECT 74.625 206.780 74.955 207.290 ;
        RECT 75.125 207.105 75.455 207.505 ;
        RECT 76.505 206.935 76.835 207.275 ;
        RECT 77.005 207.105 77.335 207.505 ;
        RECT 77.925 206.955 78.095 207.335 ;
        RECT 78.310 207.125 78.640 207.505 ;
        RECT 71.355 205.460 71.550 205.635 ;
        RECT 70.935 204.955 71.550 205.460 ;
        RECT 71.720 205.125 72.195 205.465 ;
        RECT 72.365 204.955 72.580 205.500 ;
        RECT 72.790 205.125 73.065 205.825 ;
        RECT 74.155 204.955 74.445 206.120 ;
        RECT 74.625 206.015 74.815 206.780 ;
        RECT 75.125 206.765 77.490 206.935 ;
        RECT 77.925 206.785 78.640 206.955 ;
        RECT 75.125 206.595 75.295 206.765 ;
        RECT 74.985 206.265 75.295 206.595 ;
        RECT 75.465 206.265 75.770 206.595 ;
        RECT 74.625 205.165 74.955 206.015 ;
        RECT 75.125 204.955 75.375 206.095 ;
        RECT 75.555 205.935 75.770 206.265 ;
        RECT 75.945 205.935 76.230 206.595 ;
        RECT 76.425 205.935 76.690 206.595 ;
        RECT 76.905 205.935 77.150 206.595 ;
        RECT 77.320 205.765 77.490 206.765 ;
        RECT 77.835 206.235 78.190 206.605 ;
        RECT 78.470 206.595 78.640 206.785 ;
        RECT 78.810 206.760 79.065 207.335 ;
        RECT 78.470 206.265 78.725 206.595 ;
        RECT 78.470 206.055 78.640 206.265 ;
        RECT 75.565 205.595 76.855 205.765 ;
        RECT 75.565 205.175 75.815 205.595 ;
        RECT 76.045 204.955 76.375 205.425 ;
        RECT 76.605 205.175 76.855 205.595 ;
        RECT 77.035 205.595 77.490 205.765 ;
        RECT 77.925 205.885 78.640 206.055 ;
        RECT 78.895 206.030 79.065 206.760 ;
        RECT 79.240 206.665 79.500 207.505 ;
        RECT 79.790 206.875 80.075 207.335 ;
        RECT 80.245 207.045 80.515 207.505 ;
        RECT 79.790 206.705 80.745 206.875 ;
        RECT 77.035 205.165 77.365 205.595 ;
        RECT 77.925 205.125 78.095 205.885 ;
        RECT 78.310 204.955 78.640 205.715 ;
        RECT 78.810 205.125 79.065 206.030 ;
        RECT 79.240 204.955 79.500 206.105 ;
        RECT 79.675 205.975 80.365 206.535 ;
        RECT 80.535 205.805 80.745 206.705 ;
        RECT 79.790 205.585 80.745 205.805 ;
        RECT 80.915 206.535 81.315 207.335 ;
        RECT 81.505 206.875 81.785 207.335 ;
        RECT 82.305 207.045 82.630 207.505 ;
        RECT 81.505 206.705 82.630 206.875 ;
        RECT 82.800 206.765 83.185 207.335 ;
        RECT 82.180 206.595 82.630 206.705 ;
        RECT 80.915 205.975 82.010 206.535 ;
        RECT 82.180 206.265 82.735 206.595 ;
        RECT 79.790 205.125 80.075 205.585 ;
        RECT 80.245 204.955 80.515 205.415 ;
        RECT 80.915 205.125 81.315 205.975 ;
        RECT 82.180 205.805 82.630 206.265 ;
        RECT 82.905 206.095 83.185 206.765 ;
        RECT 81.505 205.585 82.630 205.805 ;
        RECT 81.505 205.125 81.785 205.585 ;
        RECT 82.305 204.955 82.630 205.415 ;
        RECT 82.800 205.125 83.185 206.095 ;
        RECT 83.355 206.560 83.695 207.335 ;
        RECT 83.865 207.045 84.035 207.505 ;
        RECT 84.275 207.070 84.635 207.335 ;
        RECT 84.275 207.065 84.630 207.070 ;
        RECT 84.275 207.055 84.625 207.065 ;
        RECT 84.275 207.050 84.620 207.055 ;
        RECT 84.275 207.040 84.615 207.050 ;
        RECT 85.265 207.045 85.435 207.505 ;
        RECT 84.275 207.035 84.610 207.040 ;
        RECT 84.275 207.025 84.600 207.035 ;
        RECT 84.275 207.015 84.590 207.025 ;
        RECT 84.275 206.875 84.575 207.015 ;
        RECT 83.865 206.685 84.575 206.875 ;
        RECT 84.765 206.875 85.095 206.955 ;
        RECT 85.605 206.875 85.945 207.335 ;
        RECT 84.765 206.685 85.945 206.875 ;
        RECT 87.035 206.780 87.325 207.505 ;
        RECT 83.355 205.125 83.635 206.560 ;
        RECT 83.865 206.115 84.150 206.685 ;
        RECT 88.420 206.665 88.680 207.505 ;
        RECT 88.855 206.760 89.110 207.335 ;
        RECT 89.280 207.125 89.610 207.505 ;
        RECT 89.825 206.955 89.995 207.335 ;
        RECT 89.280 206.785 89.995 206.955 ;
        RECT 84.335 206.285 84.805 206.515 ;
        RECT 84.975 206.495 85.305 206.515 ;
        RECT 84.975 206.315 85.425 206.495 ;
        RECT 85.615 206.315 85.945 206.515 ;
        RECT 83.865 205.900 85.015 206.115 ;
        RECT 83.805 204.955 84.515 205.730 ;
        RECT 84.685 205.125 85.015 205.900 ;
        RECT 85.210 205.200 85.425 206.315 ;
        RECT 85.715 205.975 85.945 206.315 ;
        RECT 85.605 204.955 85.935 205.675 ;
        RECT 87.035 204.955 87.325 206.120 ;
        RECT 88.420 204.955 88.680 206.105 ;
        RECT 88.855 206.030 89.025 206.760 ;
        RECT 89.280 206.595 89.450 206.785 ;
        RECT 90.260 206.665 90.520 207.505 ;
        RECT 90.695 206.760 90.950 207.335 ;
        RECT 91.120 207.125 91.450 207.505 ;
        RECT 91.665 206.955 91.835 207.335 ;
        RECT 92.095 207.125 92.985 207.295 ;
        RECT 91.120 206.785 91.835 206.955 ;
        RECT 89.195 206.265 89.450 206.595 ;
        RECT 89.280 206.055 89.450 206.265 ;
        RECT 89.730 206.235 90.085 206.605 ;
        RECT 88.855 205.125 89.110 206.030 ;
        RECT 89.280 205.885 89.995 206.055 ;
        RECT 89.280 204.955 89.610 205.715 ;
        RECT 89.825 205.125 89.995 205.885 ;
        RECT 90.260 204.955 90.520 206.105 ;
        RECT 90.695 206.030 90.865 206.760 ;
        RECT 91.120 206.595 91.290 206.785 ;
        RECT 91.035 206.265 91.290 206.595 ;
        RECT 91.120 206.055 91.290 206.265 ;
        RECT 91.570 206.235 91.925 206.605 ;
        RECT 92.095 206.570 92.645 206.955 ;
        RECT 92.815 206.400 92.985 207.125 ;
        RECT 92.095 206.330 92.985 206.400 ;
        RECT 93.155 206.825 93.375 207.285 ;
        RECT 93.545 206.965 93.795 207.505 ;
        RECT 93.965 206.855 94.225 207.335 ;
        RECT 94.465 207.105 94.795 207.505 ;
        RECT 94.965 206.935 95.135 207.205 ;
        RECT 95.305 207.105 95.635 207.505 ;
        RECT 95.805 206.935 96.060 207.205 ;
        RECT 93.155 206.800 93.405 206.825 ;
        RECT 93.155 206.375 93.485 206.800 ;
        RECT 92.095 206.305 92.990 206.330 ;
        RECT 92.095 206.290 93.000 206.305 ;
        RECT 92.095 206.275 93.005 206.290 ;
        RECT 92.095 206.270 93.015 206.275 ;
        RECT 92.095 206.260 93.020 206.270 ;
        RECT 92.095 206.250 93.025 206.260 ;
        RECT 92.095 206.245 93.035 206.250 ;
        RECT 92.095 206.235 93.045 206.245 ;
        RECT 92.095 206.230 93.055 206.235 ;
        RECT 90.695 205.125 90.950 206.030 ;
        RECT 91.120 205.885 91.835 206.055 ;
        RECT 91.120 204.955 91.450 205.715 ;
        RECT 91.665 205.125 91.835 205.885 ;
        RECT 92.095 205.780 92.355 206.230 ;
        RECT 92.720 206.225 93.055 206.230 ;
        RECT 92.720 206.220 93.070 206.225 ;
        RECT 92.720 206.210 93.085 206.220 ;
        RECT 92.720 206.205 93.110 206.210 ;
        RECT 93.655 206.205 93.885 206.600 ;
        RECT 92.720 206.200 93.885 206.205 ;
        RECT 92.750 206.165 93.885 206.200 ;
        RECT 92.785 206.140 93.885 206.165 ;
        RECT 92.815 206.110 93.885 206.140 ;
        RECT 92.835 206.080 93.885 206.110 ;
        RECT 92.855 206.050 93.885 206.080 ;
        RECT 92.925 206.040 93.885 206.050 ;
        RECT 92.950 206.030 93.885 206.040 ;
        RECT 92.970 206.015 93.885 206.030 ;
        RECT 92.990 206.000 93.885 206.015 ;
        RECT 92.995 205.990 93.780 206.000 ;
        RECT 93.010 205.955 93.780 205.990 ;
        RECT 92.525 205.635 92.855 205.880 ;
        RECT 93.025 205.705 93.780 205.955 ;
        RECT 94.055 205.825 94.225 206.855 ;
        RECT 94.395 205.925 94.665 206.935 ;
        RECT 94.835 206.765 96.060 206.935 ;
        RECT 94.835 206.095 95.005 206.765 ;
        RECT 96.255 206.695 96.495 207.505 ;
        RECT 96.665 206.695 96.995 207.335 ;
        RECT 97.165 206.695 97.435 207.505 ;
        RECT 97.615 207.045 98.175 207.335 ;
        RECT 98.345 207.045 98.595 207.505 ;
        RECT 95.175 206.265 95.555 206.595 ;
        RECT 95.725 206.265 96.060 206.595 ;
        RECT 96.235 206.265 96.585 206.515 ;
        RECT 94.835 205.925 95.150 206.095 ;
        RECT 92.525 205.610 92.710 205.635 ;
        RECT 92.095 205.510 92.710 205.610 ;
        RECT 92.095 204.955 92.700 205.510 ;
        RECT 92.875 205.125 93.355 205.465 ;
        RECT 93.525 204.955 93.780 205.500 ;
        RECT 93.950 205.125 94.225 205.825 ;
        RECT 94.400 204.955 94.715 205.755 ;
        RECT 94.980 205.310 95.150 205.925 ;
        RECT 95.320 205.585 95.555 206.265 ;
        RECT 96.755 206.095 96.925 206.695 ;
        RECT 97.095 206.265 97.445 206.515 ;
        RECT 95.725 205.310 96.060 206.095 ;
        RECT 94.980 205.140 96.060 205.310 ;
        RECT 96.245 205.925 96.925 206.095 ;
        RECT 96.245 205.140 96.575 205.925 ;
        RECT 97.105 204.955 97.435 206.095 ;
        RECT 97.615 205.675 97.865 207.045 ;
        RECT 99.215 206.875 99.545 207.235 ;
        RECT 98.155 206.685 99.545 206.875 ;
        RECT 99.915 206.780 100.205 207.505 ;
        RECT 100.465 206.955 100.635 207.245 ;
        RECT 100.805 207.125 101.135 207.505 ;
        RECT 100.465 206.785 101.130 206.955 ;
        RECT 98.155 206.595 98.325 206.685 ;
        RECT 98.035 206.265 98.325 206.595 ;
        RECT 98.495 206.265 98.835 206.515 ;
        RECT 99.055 206.265 99.730 206.515 ;
        RECT 98.155 206.015 98.325 206.265 ;
        RECT 98.155 205.845 99.095 206.015 ;
        RECT 99.465 205.905 99.730 206.265 ;
        RECT 97.615 205.125 98.075 205.675 ;
        RECT 98.265 204.955 98.595 205.675 ;
        RECT 98.795 205.295 99.095 205.845 ;
        RECT 99.265 204.955 99.545 205.625 ;
        RECT 99.915 204.955 100.205 206.120 ;
        RECT 100.380 205.965 100.730 206.615 ;
        RECT 100.900 205.795 101.130 206.785 ;
        RECT 100.465 205.625 101.130 205.795 ;
        RECT 100.465 205.125 100.635 205.625 ;
        RECT 100.805 204.955 101.135 205.455 ;
        RECT 101.305 205.125 101.490 207.245 ;
        RECT 101.745 207.045 101.995 207.505 ;
        RECT 102.165 207.055 102.500 207.225 ;
        RECT 102.695 207.055 103.370 207.225 ;
        RECT 102.165 206.915 102.335 207.055 ;
        RECT 101.660 205.925 101.940 206.875 ;
        RECT 102.110 206.785 102.335 206.915 ;
        RECT 102.110 205.680 102.280 206.785 ;
        RECT 102.505 206.635 103.030 206.855 ;
        RECT 102.450 205.870 102.690 206.465 ;
        RECT 102.860 205.935 103.030 206.635 ;
        RECT 103.200 206.275 103.370 207.055 ;
        RECT 103.690 207.005 104.060 207.505 ;
        RECT 104.240 207.055 104.645 207.225 ;
        RECT 104.815 207.055 105.600 207.225 ;
        RECT 104.240 206.825 104.410 207.055 ;
        RECT 103.580 206.525 104.410 206.825 ;
        RECT 104.795 206.555 105.260 206.885 ;
        RECT 103.580 206.495 103.780 206.525 ;
        RECT 103.900 206.275 104.070 206.345 ;
        RECT 103.200 206.105 104.070 206.275 ;
        RECT 103.560 206.015 104.070 206.105 ;
        RECT 102.110 205.550 102.415 205.680 ;
        RECT 102.860 205.570 103.390 205.935 ;
        RECT 101.730 204.955 101.995 205.415 ;
        RECT 102.165 205.125 102.415 205.550 ;
        RECT 103.560 205.400 103.730 206.015 ;
        RECT 102.625 205.230 103.730 205.400 ;
        RECT 103.900 204.955 104.070 205.755 ;
        RECT 104.240 205.455 104.410 206.525 ;
        RECT 104.580 205.625 104.770 206.345 ;
        RECT 104.940 205.595 105.260 206.555 ;
        RECT 105.430 206.595 105.600 207.055 ;
        RECT 105.875 206.975 106.085 207.505 ;
        RECT 106.345 206.765 106.675 207.290 ;
        RECT 106.845 206.895 107.015 207.505 ;
        RECT 107.185 206.850 107.515 207.285 ;
        RECT 107.185 206.765 107.565 206.850 ;
        RECT 106.475 206.595 106.675 206.765 ;
        RECT 107.340 206.725 107.565 206.765 ;
        RECT 105.430 206.265 106.305 206.595 ;
        RECT 106.475 206.265 107.225 206.595 ;
        RECT 104.240 205.125 104.490 205.455 ;
        RECT 105.430 205.425 105.600 206.265 ;
        RECT 106.475 206.060 106.665 206.265 ;
        RECT 107.395 206.145 107.565 206.725 ;
        RECT 107.350 206.095 107.565 206.145 ;
        RECT 105.770 205.685 106.665 206.060 ;
        RECT 107.175 206.015 107.565 206.095 ;
        RECT 107.735 206.765 108.120 207.335 ;
        RECT 108.290 207.045 108.615 207.505 ;
        RECT 109.135 206.875 109.415 207.335 ;
        RECT 107.735 206.095 108.015 206.765 ;
        RECT 108.290 206.705 109.415 206.875 ;
        RECT 108.290 206.595 108.740 206.705 ;
        RECT 108.185 206.265 108.740 206.595 ;
        RECT 109.605 206.535 110.005 207.335 ;
        RECT 110.405 207.045 110.675 207.505 ;
        RECT 110.845 206.875 111.130 207.335 ;
        RECT 104.715 205.255 105.600 205.425 ;
        RECT 105.780 204.955 106.095 205.455 ;
        RECT 106.325 205.125 106.665 205.685 ;
        RECT 106.835 204.955 107.005 205.965 ;
        RECT 107.175 205.170 107.505 206.015 ;
        RECT 107.735 205.125 108.120 206.095 ;
        RECT 108.290 205.805 108.740 206.265 ;
        RECT 108.910 205.975 110.005 206.535 ;
        RECT 108.290 205.585 109.415 205.805 ;
        RECT 108.290 204.955 108.615 205.415 ;
        RECT 109.135 205.125 109.415 205.585 ;
        RECT 109.605 205.125 110.005 205.975 ;
        RECT 110.175 206.705 111.130 206.875 ;
        RECT 111.595 206.845 111.935 207.505 ;
        RECT 110.175 205.805 110.385 206.705 ;
        RECT 110.555 205.975 111.245 206.535 ;
        RECT 110.175 205.585 111.130 205.805 ;
        RECT 110.405 204.955 110.675 205.415 ;
        RECT 110.845 205.125 111.130 205.585 ;
        RECT 111.415 205.125 111.935 206.675 ;
        RECT 112.105 205.850 112.625 207.335 ;
        RECT 112.795 206.780 113.085 207.505 ;
        RECT 114.175 206.755 115.385 207.505 ;
        RECT 112.105 204.955 112.435 205.680 ;
        RECT 112.795 204.955 113.085 206.120 ;
        RECT 114.175 206.045 114.695 206.585 ;
        RECT 114.865 206.215 115.385 206.755 ;
        RECT 114.175 204.955 115.385 206.045 ;
        RECT 61.190 204.785 115.470 204.955 ;
        RECT 61.275 203.695 62.485 204.785 ;
        RECT 62.655 203.695 64.325 204.785 ;
        RECT 61.275 202.985 61.795 203.525 ;
        RECT 61.965 203.155 62.485 203.695 ;
        RECT 62.655 203.005 63.405 203.525 ;
        RECT 63.575 203.175 64.325 203.695 ;
        RECT 64.500 203.635 64.760 204.785 ;
        RECT 64.935 203.710 65.190 204.615 ;
        RECT 65.360 204.025 65.690 204.785 ;
        RECT 65.905 203.855 66.075 204.615 ;
        RECT 61.275 202.235 62.485 202.985 ;
        RECT 62.655 202.235 64.325 203.005 ;
        RECT 64.500 202.235 64.760 203.075 ;
        RECT 64.935 202.980 65.105 203.710 ;
        RECT 65.360 203.685 66.075 203.855 ;
        RECT 65.360 203.475 65.530 203.685 ;
        RECT 66.340 203.635 66.600 204.785 ;
        RECT 66.775 203.710 67.030 204.615 ;
        RECT 67.200 204.025 67.530 204.785 ;
        RECT 67.745 203.855 67.915 204.615 ;
        RECT 68.290 204.155 68.575 204.615 ;
        RECT 68.745 204.325 69.015 204.785 ;
        RECT 68.290 203.935 69.245 204.155 ;
        RECT 65.275 203.145 65.530 203.475 ;
        RECT 64.935 202.405 65.190 202.980 ;
        RECT 65.360 202.955 65.530 203.145 ;
        RECT 65.810 203.135 66.165 203.505 ;
        RECT 65.360 202.785 66.075 202.955 ;
        RECT 65.360 202.235 65.690 202.615 ;
        RECT 65.905 202.405 66.075 202.785 ;
        RECT 66.340 202.235 66.600 203.075 ;
        RECT 66.775 202.980 66.945 203.710 ;
        RECT 67.200 203.685 67.915 203.855 ;
        RECT 67.200 203.475 67.370 203.685 ;
        RECT 67.115 203.145 67.370 203.475 ;
        RECT 66.775 202.405 67.030 202.980 ;
        RECT 67.200 202.955 67.370 203.145 ;
        RECT 67.650 203.135 68.005 203.505 ;
        RECT 68.175 203.205 68.865 203.765 ;
        RECT 69.035 203.035 69.245 203.935 ;
        RECT 67.200 202.785 67.915 202.955 ;
        RECT 67.200 202.235 67.530 202.615 ;
        RECT 67.745 202.405 67.915 202.785 ;
        RECT 68.290 202.865 69.245 203.035 ;
        RECT 69.415 203.765 69.815 204.615 ;
        RECT 70.005 204.155 70.285 204.615 ;
        RECT 70.805 204.325 71.130 204.785 ;
        RECT 70.005 203.935 71.130 204.155 ;
        RECT 69.415 203.205 70.510 203.765 ;
        RECT 70.680 203.475 71.130 203.935 ;
        RECT 71.300 203.645 71.685 204.615 ;
        RECT 68.290 202.405 68.575 202.865 ;
        RECT 68.745 202.235 69.015 202.695 ;
        RECT 69.415 202.405 69.815 203.205 ;
        RECT 70.680 203.145 71.235 203.475 ;
        RECT 70.680 203.035 71.130 203.145 ;
        RECT 70.005 202.865 71.130 203.035 ;
        RECT 71.405 202.975 71.685 203.645 ;
        RECT 72.320 203.635 72.580 204.785 ;
        RECT 72.755 203.710 73.010 204.615 ;
        RECT 73.180 204.025 73.510 204.785 ;
        RECT 73.725 203.855 73.895 204.615 ;
        RECT 70.005 202.405 70.285 202.865 ;
        RECT 70.805 202.235 71.130 202.695 ;
        RECT 71.300 202.405 71.685 202.975 ;
        RECT 72.320 202.235 72.580 203.075 ;
        RECT 72.755 202.980 72.925 203.710 ;
        RECT 73.180 203.685 73.895 203.855 ;
        RECT 73.180 203.475 73.350 203.685 ;
        RECT 74.155 203.620 74.445 204.785 ;
        RECT 74.625 204.175 74.955 204.605 ;
        RECT 75.135 204.345 75.330 204.785 ;
        RECT 75.500 204.175 75.830 204.605 ;
        RECT 74.625 204.005 75.830 204.175 ;
        RECT 74.625 203.675 75.520 204.005 ;
        RECT 76.000 203.835 76.275 204.605 ;
        RECT 75.690 203.645 76.275 203.835 ;
        RECT 76.465 203.725 76.795 204.575 ;
        RECT 73.095 203.145 73.350 203.475 ;
        RECT 72.755 202.405 73.010 202.980 ;
        RECT 73.180 202.955 73.350 203.145 ;
        RECT 73.630 203.135 73.985 203.505 ;
        RECT 74.630 203.145 74.925 203.475 ;
        RECT 75.105 203.145 75.520 203.475 ;
        RECT 73.180 202.785 73.895 202.955 ;
        RECT 73.180 202.235 73.510 202.615 ;
        RECT 73.725 202.405 73.895 202.785 ;
        RECT 74.155 202.235 74.445 202.960 ;
        RECT 74.625 202.235 74.925 202.965 ;
        RECT 75.105 202.525 75.335 203.145 ;
        RECT 75.690 202.975 75.865 203.645 ;
        RECT 75.535 202.795 75.865 202.975 ;
        RECT 76.035 202.825 76.275 203.475 ;
        RECT 76.465 202.960 76.655 203.725 ;
        RECT 76.965 203.645 77.215 204.785 ;
        RECT 77.405 204.145 77.655 204.565 ;
        RECT 77.885 204.315 78.215 204.785 ;
        RECT 78.445 204.145 78.695 204.565 ;
        RECT 77.405 203.975 78.695 204.145 ;
        RECT 78.875 204.145 79.205 204.575 ;
        RECT 78.875 203.975 79.330 204.145 ;
        RECT 77.395 203.475 77.610 203.805 ;
        RECT 76.825 203.145 77.135 203.475 ;
        RECT 77.305 203.145 77.610 203.475 ;
        RECT 77.785 203.145 78.070 203.805 ;
        RECT 78.265 203.145 78.530 203.805 ;
        RECT 78.745 203.145 78.990 203.805 ;
        RECT 76.965 202.975 77.135 203.145 ;
        RECT 79.160 202.975 79.330 203.975 ;
        RECT 75.535 202.415 75.760 202.795 ;
        RECT 75.930 202.235 76.260 202.625 ;
        RECT 76.465 202.450 76.795 202.960 ;
        RECT 76.965 202.805 79.330 202.975 ;
        RECT 79.675 203.645 80.060 204.615 ;
        RECT 80.230 204.325 80.555 204.785 ;
        RECT 81.075 204.155 81.355 204.615 ;
        RECT 80.230 203.935 81.355 204.155 ;
        RECT 79.675 202.975 79.955 203.645 ;
        RECT 80.230 203.475 80.680 203.935 ;
        RECT 81.545 203.765 81.945 204.615 ;
        RECT 82.345 204.325 82.615 204.785 ;
        RECT 82.785 204.155 83.070 204.615 ;
        RECT 80.125 203.145 80.680 203.475 ;
        RECT 80.850 203.205 81.945 203.765 ;
        RECT 80.230 203.035 80.680 203.145 ;
        RECT 76.965 202.235 77.295 202.635 ;
        RECT 78.345 202.465 78.675 202.805 ;
        RECT 78.845 202.235 79.175 202.635 ;
        RECT 79.675 202.405 80.060 202.975 ;
        RECT 80.230 202.865 81.355 203.035 ;
        RECT 80.230 202.235 80.555 202.695 ;
        RECT 81.075 202.405 81.355 202.865 ;
        RECT 81.545 202.405 81.945 203.205 ;
        RECT 82.115 203.935 83.070 204.155 ;
        RECT 82.115 203.035 82.325 203.935 ;
        RECT 82.495 203.205 83.185 203.765 ;
        RECT 83.415 203.645 83.625 204.785 ;
        RECT 83.795 203.635 84.125 204.615 ;
        RECT 84.295 203.645 84.525 204.785 ;
        RECT 84.825 204.115 84.995 204.615 ;
        RECT 85.165 204.285 85.495 204.785 ;
        RECT 84.825 203.945 85.490 204.115 ;
        RECT 82.115 202.865 83.070 203.035 ;
        RECT 82.345 202.235 82.615 202.695 ;
        RECT 82.785 202.405 83.070 202.865 ;
        RECT 83.415 202.235 83.625 203.055 ;
        RECT 83.795 203.035 84.045 203.635 ;
        RECT 84.215 203.225 84.545 203.475 ;
        RECT 84.740 203.125 85.090 203.775 ;
        RECT 83.795 202.405 84.125 203.035 ;
        RECT 84.295 202.235 84.525 203.055 ;
        RECT 85.260 202.955 85.490 203.945 ;
        RECT 84.825 202.785 85.490 202.955 ;
        RECT 84.825 202.495 84.995 202.785 ;
        RECT 85.165 202.235 85.495 202.615 ;
        RECT 85.665 202.495 85.850 204.615 ;
        RECT 86.090 204.325 86.355 204.785 ;
        RECT 86.525 204.190 86.775 204.615 ;
        RECT 86.985 204.340 88.090 204.510 ;
        RECT 86.470 204.060 86.775 204.190 ;
        RECT 86.020 202.865 86.300 203.815 ;
        RECT 86.470 202.955 86.640 204.060 ;
        RECT 86.810 203.275 87.050 203.870 ;
        RECT 87.220 203.805 87.750 204.170 ;
        RECT 87.220 203.105 87.390 203.805 ;
        RECT 87.920 203.725 88.090 204.340 ;
        RECT 88.260 203.985 88.430 204.785 ;
        RECT 88.600 204.285 88.850 204.615 ;
        RECT 89.075 204.315 89.960 204.485 ;
        RECT 87.920 203.635 88.430 203.725 ;
        RECT 86.470 202.825 86.695 202.955 ;
        RECT 86.865 202.885 87.390 203.105 ;
        RECT 87.560 203.465 88.430 203.635 ;
        RECT 86.105 202.235 86.355 202.695 ;
        RECT 86.525 202.685 86.695 202.825 ;
        RECT 87.560 202.685 87.730 203.465 ;
        RECT 88.260 203.395 88.430 203.465 ;
        RECT 87.940 203.215 88.140 203.245 ;
        RECT 88.600 203.215 88.770 204.285 ;
        RECT 88.940 203.395 89.130 204.115 ;
        RECT 87.940 202.915 88.770 203.215 ;
        RECT 89.300 203.185 89.620 204.145 ;
        RECT 86.525 202.515 86.860 202.685 ;
        RECT 87.055 202.515 87.730 202.685 ;
        RECT 88.050 202.235 88.420 202.735 ;
        RECT 88.600 202.685 88.770 202.915 ;
        RECT 89.155 202.855 89.620 203.185 ;
        RECT 89.790 203.475 89.960 204.315 ;
        RECT 90.140 204.285 90.455 204.785 ;
        RECT 90.685 204.055 91.025 204.615 ;
        RECT 90.130 203.680 91.025 204.055 ;
        RECT 91.195 203.775 91.365 204.785 ;
        RECT 90.835 203.475 91.025 203.680 ;
        RECT 91.535 203.725 91.865 204.570 ;
        RECT 91.535 203.645 91.925 203.725 ;
        RECT 91.710 203.595 91.925 203.645 ;
        RECT 89.790 203.145 90.665 203.475 ;
        RECT 90.835 203.145 91.585 203.475 ;
        RECT 89.790 202.685 89.960 203.145 ;
        RECT 90.835 202.975 91.035 203.145 ;
        RECT 91.755 203.015 91.925 203.595 ;
        RECT 91.700 202.975 91.925 203.015 ;
        RECT 88.600 202.515 89.005 202.685 ;
        RECT 89.175 202.515 89.960 202.685 ;
        RECT 90.235 202.235 90.445 202.765 ;
        RECT 90.705 202.450 91.035 202.975 ;
        RECT 91.545 202.890 91.925 202.975 ;
        RECT 92.095 203.645 92.480 204.615 ;
        RECT 92.650 204.325 92.975 204.785 ;
        RECT 93.495 204.155 93.775 204.615 ;
        RECT 92.650 203.935 93.775 204.155 ;
        RECT 92.095 202.975 92.375 203.645 ;
        RECT 92.650 203.475 93.100 203.935 ;
        RECT 93.965 203.765 94.365 204.615 ;
        RECT 94.765 204.325 95.035 204.785 ;
        RECT 95.205 204.155 95.490 204.615 ;
        RECT 92.545 203.145 93.100 203.475 ;
        RECT 93.270 203.205 94.365 203.765 ;
        RECT 92.650 203.035 93.100 203.145 ;
        RECT 91.205 202.235 91.375 202.845 ;
        RECT 91.545 202.455 91.875 202.890 ;
        RECT 92.095 202.405 92.480 202.975 ;
        RECT 92.650 202.865 93.775 203.035 ;
        RECT 92.650 202.235 92.975 202.695 ;
        RECT 93.495 202.405 93.775 202.865 ;
        RECT 93.965 202.405 94.365 203.205 ;
        RECT 94.535 203.935 95.490 204.155 ;
        RECT 95.775 204.065 96.235 204.615 ;
        RECT 96.425 204.065 96.755 204.785 ;
        RECT 94.535 203.035 94.745 203.935 ;
        RECT 94.915 203.205 95.605 203.765 ;
        RECT 94.535 202.865 95.490 203.035 ;
        RECT 94.765 202.235 95.035 202.695 ;
        RECT 95.205 202.405 95.490 202.865 ;
        RECT 95.775 202.695 96.025 204.065 ;
        RECT 96.955 203.895 97.255 204.445 ;
        RECT 97.425 204.115 97.705 204.785 ;
        RECT 98.085 204.175 98.415 204.605 ;
        RECT 98.595 204.345 98.790 204.785 ;
        RECT 98.960 204.175 99.290 204.605 ;
        RECT 96.315 203.725 97.255 203.895 ;
        RECT 98.085 204.005 99.290 204.175 ;
        RECT 96.315 203.475 96.485 203.725 ;
        RECT 97.625 203.475 97.890 203.835 ;
        RECT 98.085 203.675 98.980 204.005 ;
        RECT 99.460 203.835 99.735 204.605 ;
        RECT 99.150 203.645 99.735 203.835 ;
        RECT 96.195 203.145 96.485 203.475 ;
        RECT 96.655 203.225 96.995 203.475 ;
        RECT 97.215 203.225 97.890 203.475 ;
        RECT 98.090 203.145 98.385 203.475 ;
        RECT 98.565 203.145 98.980 203.475 ;
        RECT 96.315 203.055 96.485 203.145 ;
        RECT 96.315 202.865 97.705 203.055 ;
        RECT 95.775 202.405 96.335 202.695 ;
        RECT 96.505 202.235 96.755 202.695 ;
        RECT 97.375 202.505 97.705 202.865 ;
        RECT 98.085 202.235 98.385 202.965 ;
        RECT 98.565 202.525 98.795 203.145 ;
        RECT 99.150 202.975 99.325 203.645 ;
        RECT 99.915 203.620 100.205 204.785 ;
        RECT 100.375 203.645 100.760 204.615 ;
        RECT 100.930 204.325 101.255 204.785 ;
        RECT 101.775 204.155 102.055 204.615 ;
        RECT 100.930 203.935 102.055 204.155 ;
        RECT 98.995 202.795 99.325 202.975 ;
        RECT 99.495 202.825 99.735 203.475 ;
        RECT 100.375 202.975 100.655 203.645 ;
        RECT 100.930 203.475 101.380 203.935 ;
        RECT 102.245 203.765 102.645 204.615 ;
        RECT 103.045 204.325 103.315 204.785 ;
        RECT 103.485 204.155 103.770 204.615 ;
        RECT 100.825 203.145 101.380 203.475 ;
        RECT 101.550 203.205 102.645 203.765 ;
        RECT 100.930 203.035 101.380 203.145 ;
        RECT 98.995 202.415 99.220 202.795 ;
        RECT 99.390 202.235 99.720 202.625 ;
        RECT 99.915 202.235 100.205 202.960 ;
        RECT 100.375 202.405 100.760 202.975 ;
        RECT 100.930 202.865 102.055 203.035 ;
        RECT 100.930 202.235 101.255 202.695 ;
        RECT 101.775 202.405 102.055 202.865 ;
        RECT 102.245 202.405 102.645 203.205 ;
        RECT 102.815 203.935 103.770 204.155 ;
        RECT 102.815 203.035 103.025 203.935 ;
        RECT 103.195 203.205 103.885 203.765 ;
        RECT 104.980 203.595 105.235 204.475 ;
        RECT 105.405 203.645 105.710 204.785 ;
        RECT 106.050 204.405 106.380 204.785 ;
        RECT 106.560 204.235 106.730 204.525 ;
        RECT 106.900 204.325 107.150 204.785 ;
        RECT 105.930 204.065 106.730 204.235 ;
        RECT 107.320 204.275 108.190 204.615 ;
        RECT 102.815 202.865 103.770 203.035 ;
        RECT 103.045 202.235 103.315 202.695 ;
        RECT 103.485 202.405 103.770 202.865 ;
        RECT 104.980 202.945 105.190 203.595 ;
        RECT 105.930 203.475 106.100 204.065 ;
        RECT 107.320 203.895 107.490 204.275 ;
        RECT 108.425 204.155 108.595 204.615 ;
        RECT 108.765 204.325 109.135 204.785 ;
        RECT 109.430 204.185 109.600 204.525 ;
        RECT 109.770 204.355 110.100 204.785 ;
        RECT 110.335 204.185 110.505 204.525 ;
        RECT 106.270 203.725 107.490 203.895 ;
        RECT 107.660 203.815 108.120 204.105 ;
        RECT 108.425 203.985 108.985 204.155 ;
        RECT 109.430 204.015 110.505 204.185 ;
        RECT 110.675 204.285 111.355 204.615 ;
        RECT 111.570 204.285 111.820 204.615 ;
        RECT 111.990 204.325 112.240 204.785 ;
        RECT 108.815 203.845 108.985 203.985 ;
        RECT 107.660 203.805 108.625 203.815 ;
        RECT 107.320 203.635 107.490 203.725 ;
        RECT 107.950 203.645 108.625 203.805 ;
        RECT 105.360 203.445 106.100 203.475 ;
        RECT 105.360 203.145 106.275 203.445 ;
        RECT 105.950 202.970 106.275 203.145 ;
        RECT 104.980 202.415 105.235 202.945 ;
        RECT 105.405 202.235 105.710 202.695 ;
        RECT 105.955 202.615 106.275 202.970 ;
        RECT 106.445 203.185 106.985 203.555 ;
        RECT 107.320 203.465 107.725 203.635 ;
        RECT 106.445 202.785 106.685 203.185 ;
        RECT 107.165 203.015 107.385 203.295 ;
        RECT 106.855 202.845 107.385 203.015 ;
        RECT 106.855 202.615 107.025 202.845 ;
        RECT 107.555 202.685 107.725 203.465 ;
        RECT 107.895 202.855 108.245 203.475 ;
        RECT 108.415 202.855 108.625 203.645 ;
        RECT 108.815 203.675 110.315 203.845 ;
        RECT 108.815 202.985 108.985 203.675 ;
        RECT 110.675 203.505 110.845 204.285 ;
        RECT 111.650 204.155 111.820 204.285 ;
        RECT 109.155 203.335 110.845 203.505 ;
        RECT 111.015 203.725 111.480 204.115 ;
        RECT 111.650 203.985 112.045 204.155 ;
        RECT 109.155 203.155 109.325 203.335 ;
        RECT 105.955 202.445 107.025 202.615 ;
        RECT 107.195 202.235 107.385 202.675 ;
        RECT 107.555 202.405 108.505 202.685 ;
        RECT 108.815 202.595 109.075 202.985 ;
        RECT 109.495 202.915 110.285 203.165 ;
        RECT 108.725 202.425 109.075 202.595 ;
        RECT 109.285 202.235 109.615 202.695 ;
        RECT 110.490 202.625 110.660 203.335 ;
        RECT 111.015 203.135 111.185 203.725 ;
        RECT 110.830 202.915 111.185 203.135 ;
        RECT 111.355 202.915 111.705 203.535 ;
        RECT 111.875 202.625 112.045 203.985 ;
        RECT 112.410 203.815 112.735 204.600 ;
        RECT 112.215 202.765 112.675 203.815 ;
        RECT 110.490 202.455 111.345 202.625 ;
        RECT 111.550 202.455 112.045 202.625 ;
        RECT 112.215 202.235 112.545 202.595 ;
        RECT 112.905 202.495 113.075 204.615 ;
        RECT 113.245 204.285 113.575 204.785 ;
        RECT 113.745 204.115 114.000 204.615 ;
        RECT 113.250 203.945 114.000 204.115 ;
        RECT 113.250 202.955 113.480 203.945 ;
        RECT 113.650 203.125 114.000 203.775 ;
        RECT 114.175 203.695 115.385 204.785 ;
        RECT 114.175 203.155 114.695 203.695 ;
        RECT 114.865 202.985 115.385 203.525 ;
        RECT 113.250 202.785 114.000 202.955 ;
        RECT 113.245 202.235 113.575 202.615 ;
        RECT 113.745 202.495 114.000 202.785 ;
        RECT 114.175 202.235 115.385 202.985 ;
        RECT 61.190 202.065 115.470 202.235 ;
        RECT 61.275 201.315 62.485 202.065 ;
        RECT 61.275 200.775 61.795 201.315 ;
        RECT 63.585 201.255 63.855 202.065 ;
        RECT 64.025 201.255 64.355 201.895 ;
        RECT 64.525 201.255 64.765 202.065 ;
        RECT 64.965 201.335 65.265 202.065 ;
        RECT 61.965 200.605 62.485 201.145 ;
        RECT 63.575 200.825 63.925 201.075 ;
        RECT 64.095 200.655 64.265 201.255 ;
        RECT 65.445 201.155 65.675 201.775 ;
        RECT 65.875 201.505 66.100 201.885 ;
        RECT 66.270 201.675 66.600 202.065 ;
        RECT 65.875 201.325 66.205 201.505 ;
        RECT 64.435 200.825 64.785 201.075 ;
        RECT 64.970 200.825 65.265 201.155 ;
        RECT 65.445 200.825 65.860 201.155 ;
        RECT 66.030 200.655 66.205 201.325 ;
        RECT 66.375 200.825 66.615 201.475 ;
        RECT 66.845 201.410 67.175 201.845 ;
        RECT 67.345 201.455 67.515 202.065 ;
        RECT 66.795 201.325 67.175 201.410 ;
        RECT 67.685 201.325 68.015 201.850 ;
        RECT 68.275 201.535 68.485 202.065 ;
        RECT 68.760 201.615 69.545 201.785 ;
        RECT 69.715 201.615 70.120 201.785 ;
        RECT 66.795 201.285 67.020 201.325 ;
        RECT 66.795 200.705 66.965 201.285 ;
        RECT 67.685 201.155 67.885 201.325 ;
        RECT 68.760 201.155 68.930 201.615 ;
        RECT 67.135 200.825 67.885 201.155 ;
        RECT 68.055 200.825 68.930 201.155 ;
        RECT 66.795 200.655 67.010 200.705 ;
        RECT 61.275 199.515 62.485 200.605 ;
        RECT 63.585 199.515 63.915 200.655 ;
        RECT 64.095 200.485 64.775 200.655 ;
        RECT 64.445 199.700 64.775 200.485 ;
        RECT 64.965 200.295 65.860 200.625 ;
        RECT 66.030 200.465 66.615 200.655 ;
        RECT 66.795 200.575 67.185 200.655 ;
        RECT 64.965 200.125 66.170 200.295 ;
        RECT 64.965 199.695 65.295 200.125 ;
        RECT 65.475 199.515 65.670 199.955 ;
        RECT 65.840 199.695 66.170 200.125 ;
        RECT 66.340 199.695 66.615 200.465 ;
        RECT 66.855 199.730 67.185 200.575 ;
        RECT 67.695 200.620 67.885 200.825 ;
        RECT 67.355 199.515 67.525 200.525 ;
        RECT 67.695 200.245 68.590 200.620 ;
        RECT 67.695 199.685 68.035 200.245 ;
        RECT 68.265 199.515 68.580 200.015 ;
        RECT 68.760 199.985 68.930 200.825 ;
        RECT 69.100 201.115 69.565 201.445 ;
        RECT 69.950 201.385 70.120 201.615 ;
        RECT 70.300 201.565 70.670 202.065 ;
        RECT 70.990 201.615 71.665 201.785 ;
        RECT 71.860 201.615 72.195 201.785 ;
        RECT 69.100 200.155 69.420 201.115 ;
        RECT 69.950 201.085 70.780 201.385 ;
        RECT 69.590 200.185 69.780 200.905 ;
        RECT 69.950 200.015 70.120 201.085 ;
        RECT 70.580 201.055 70.780 201.085 ;
        RECT 70.290 200.835 70.460 200.905 ;
        RECT 70.990 200.835 71.160 201.615 ;
        RECT 72.025 201.475 72.195 201.615 ;
        RECT 72.365 201.605 72.615 202.065 ;
        RECT 70.290 200.665 71.160 200.835 ;
        RECT 71.330 201.195 71.855 201.415 ;
        RECT 72.025 201.345 72.250 201.475 ;
        RECT 70.290 200.575 70.800 200.665 ;
        RECT 68.760 199.815 69.645 199.985 ;
        RECT 69.870 199.685 70.120 200.015 ;
        RECT 70.290 199.515 70.460 200.315 ;
        RECT 70.630 199.960 70.800 200.575 ;
        RECT 71.330 200.495 71.500 201.195 ;
        RECT 70.970 200.130 71.500 200.495 ;
        RECT 71.670 200.430 71.910 201.025 ;
        RECT 72.080 200.240 72.250 201.345 ;
        RECT 72.420 200.485 72.700 201.435 ;
        RECT 71.945 200.110 72.250 200.240 ;
        RECT 70.630 199.790 71.735 199.960 ;
        RECT 71.945 199.685 72.195 200.110 ;
        RECT 72.365 199.515 72.630 199.975 ;
        RECT 72.870 199.685 73.055 201.805 ;
        RECT 73.225 201.685 73.555 202.065 ;
        RECT 73.725 201.515 73.895 201.805 ;
        RECT 73.230 201.345 73.895 201.515 ;
        RECT 73.230 200.355 73.460 201.345 ;
        RECT 74.155 201.265 74.465 202.065 ;
        RECT 74.670 201.265 75.365 201.895 ;
        RECT 75.585 201.410 75.915 201.845 ;
        RECT 76.085 201.455 76.255 202.065 ;
        RECT 75.535 201.325 75.915 201.410 ;
        RECT 76.425 201.325 76.755 201.850 ;
        RECT 77.015 201.535 77.225 202.065 ;
        RECT 77.500 201.615 78.285 201.785 ;
        RECT 78.455 201.615 78.860 201.785 ;
        RECT 75.535 201.285 75.760 201.325 ;
        RECT 73.630 200.525 73.980 201.175 ;
        RECT 74.165 200.825 74.500 201.095 ;
        RECT 74.670 200.665 74.840 201.265 ;
        RECT 75.010 200.825 75.345 201.075 ;
        RECT 75.535 200.705 75.705 201.285 ;
        RECT 76.425 201.155 76.625 201.325 ;
        RECT 77.500 201.155 77.670 201.615 ;
        RECT 75.875 200.825 76.625 201.155 ;
        RECT 76.795 200.825 77.670 201.155 ;
        RECT 73.230 200.185 73.895 200.355 ;
        RECT 73.225 199.515 73.555 200.015 ;
        RECT 73.725 199.685 73.895 200.185 ;
        RECT 74.155 199.515 74.435 200.655 ;
        RECT 74.605 199.685 74.935 200.665 ;
        RECT 75.535 200.655 75.750 200.705 ;
        RECT 75.105 199.515 75.365 200.655 ;
        RECT 75.535 200.575 75.925 200.655 ;
        RECT 75.595 199.730 75.925 200.575 ;
        RECT 76.435 200.620 76.625 200.825 ;
        RECT 76.095 199.515 76.265 200.525 ;
        RECT 76.435 200.245 77.330 200.620 ;
        RECT 76.435 199.685 76.775 200.245 ;
        RECT 77.005 199.515 77.320 200.015 ;
        RECT 77.500 199.985 77.670 200.825 ;
        RECT 77.840 201.115 78.305 201.445 ;
        RECT 78.690 201.385 78.860 201.615 ;
        RECT 79.040 201.565 79.410 202.065 ;
        RECT 79.730 201.615 80.405 201.785 ;
        RECT 80.600 201.615 80.935 201.785 ;
        RECT 77.840 200.155 78.160 201.115 ;
        RECT 78.690 201.085 79.520 201.385 ;
        RECT 78.330 200.185 78.520 200.905 ;
        RECT 78.690 200.015 78.860 201.085 ;
        RECT 79.320 201.055 79.520 201.085 ;
        RECT 79.030 200.835 79.200 200.905 ;
        RECT 79.730 200.835 79.900 201.615 ;
        RECT 80.765 201.475 80.935 201.615 ;
        RECT 81.105 201.605 81.355 202.065 ;
        RECT 79.030 200.665 79.900 200.835 ;
        RECT 80.070 201.195 80.595 201.415 ;
        RECT 80.765 201.345 80.990 201.475 ;
        RECT 79.030 200.575 79.540 200.665 ;
        RECT 77.500 199.815 78.385 199.985 ;
        RECT 78.610 199.685 78.860 200.015 ;
        RECT 79.030 199.515 79.200 200.315 ;
        RECT 79.370 199.960 79.540 200.575 ;
        RECT 80.070 200.495 80.240 201.195 ;
        RECT 79.710 200.130 80.240 200.495 ;
        RECT 80.410 200.430 80.650 201.025 ;
        RECT 80.820 200.240 80.990 201.345 ;
        RECT 81.160 200.485 81.440 201.435 ;
        RECT 80.685 200.110 80.990 200.240 ;
        RECT 79.370 199.790 80.475 199.960 ;
        RECT 80.685 199.685 80.935 200.110 ;
        RECT 81.105 199.515 81.370 199.975 ;
        RECT 81.610 199.685 81.795 201.805 ;
        RECT 81.965 201.685 82.295 202.065 ;
        RECT 82.465 201.515 82.635 201.805 ;
        RECT 81.970 201.345 82.635 201.515 ;
        RECT 81.970 200.355 82.200 201.345 ;
        RECT 82.905 201.255 83.175 202.065 ;
        RECT 83.345 201.255 83.675 201.895 ;
        RECT 83.845 201.255 84.085 202.065 ;
        RECT 82.370 200.525 82.720 201.175 ;
        RECT 82.895 200.825 83.245 201.075 ;
        RECT 83.415 200.655 83.585 201.255 ;
        RECT 84.275 201.120 84.615 201.895 ;
        RECT 84.785 201.605 84.955 202.065 ;
        RECT 85.195 201.630 85.555 201.895 ;
        RECT 85.195 201.625 85.550 201.630 ;
        RECT 85.195 201.615 85.545 201.625 ;
        RECT 85.195 201.610 85.540 201.615 ;
        RECT 85.195 201.600 85.535 201.610 ;
        RECT 86.185 201.605 86.355 202.065 ;
        RECT 85.195 201.595 85.530 201.600 ;
        RECT 85.195 201.585 85.520 201.595 ;
        RECT 85.195 201.575 85.510 201.585 ;
        RECT 85.195 201.435 85.495 201.575 ;
        RECT 84.785 201.245 85.495 201.435 ;
        RECT 85.685 201.435 86.015 201.515 ;
        RECT 86.525 201.435 86.865 201.895 ;
        RECT 85.685 201.245 86.865 201.435 ;
        RECT 87.035 201.340 87.325 202.065 ;
        RECT 83.755 200.825 84.105 201.075 ;
        RECT 81.970 200.185 82.635 200.355 ;
        RECT 81.965 199.515 82.295 200.015 ;
        RECT 82.465 199.685 82.635 200.185 ;
        RECT 82.905 199.515 83.235 200.655 ;
        RECT 83.415 200.485 84.095 200.655 ;
        RECT 83.765 199.700 84.095 200.485 ;
        RECT 84.275 199.685 84.555 201.120 ;
        RECT 84.785 200.675 85.070 201.245 ;
        RECT 87.495 201.120 87.835 201.895 ;
        RECT 88.005 201.605 88.175 202.065 ;
        RECT 88.415 201.630 88.775 201.895 ;
        RECT 88.415 201.625 88.770 201.630 ;
        RECT 88.415 201.615 88.765 201.625 ;
        RECT 88.415 201.610 88.760 201.615 ;
        RECT 88.415 201.600 88.755 201.610 ;
        RECT 89.405 201.605 89.575 202.065 ;
        RECT 88.415 201.595 88.750 201.600 ;
        RECT 88.415 201.585 88.740 201.595 ;
        RECT 88.415 201.575 88.730 201.585 ;
        RECT 88.415 201.435 88.715 201.575 ;
        RECT 88.005 201.245 88.715 201.435 ;
        RECT 88.905 201.435 89.235 201.515 ;
        RECT 89.745 201.435 90.085 201.895 ;
        RECT 88.905 201.245 90.085 201.435 ;
        RECT 90.255 201.325 90.640 201.895 ;
        RECT 90.810 201.605 91.135 202.065 ;
        RECT 91.655 201.435 91.935 201.895 ;
        RECT 85.255 200.845 85.725 201.075 ;
        RECT 85.895 201.055 86.225 201.075 ;
        RECT 85.895 200.875 86.345 201.055 ;
        RECT 86.535 200.875 86.865 201.075 ;
        RECT 84.785 200.460 85.935 200.675 ;
        RECT 84.725 199.515 85.435 200.290 ;
        RECT 85.605 199.685 85.935 200.460 ;
        RECT 86.130 199.760 86.345 200.875 ;
        RECT 86.635 200.535 86.865 200.875 ;
        RECT 86.525 199.515 86.855 200.235 ;
        RECT 87.035 199.515 87.325 200.680 ;
        RECT 87.495 199.685 87.775 201.120 ;
        RECT 88.005 200.675 88.290 201.245 ;
        RECT 88.475 200.845 88.945 201.075 ;
        RECT 89.115 201.055 89.445 201.075 ;
        RECT 89.115 200.875 89.565 201.055 ;
        RECT 89.755 200.875 90.085 201.075 ;
        RECT 88.005 200.460 89.155 200.675 ;
        RECT 87.945 199.515 88.655 200.290 ;
        RECT 88.825 199.685 89.155 200.460 ;
        RECT 89.350 199.760 89.565 200.875 ;
        RECT 89.855 200.535 90.085 200.875 ;
        RECT 90.255 200.655 90.535 201.325 ;
        RECT 90.810 201.265 91.935 201.435 ;
        RECT 90.810 201.155 91.260 201.265 ;
        RECT 90.705 200.825 91.260 201.155 ;
        RECT 92.125 201.095 92.525 201.895 ;
        RECT 92.925 201.605 93.195 202.065 ;
        RECT 93.365 201.435 93.650 201.895 ;
        RECT 89.745 199.515 90.075 200.235 ;
        RECT 90.255 199.685 90.640 200.655 ;
        RECT 90.810 200.365 91.260 200.825 ;
        RECT 91.430 200.535 92.525 201.095 ;
        RECT 90.810 200.145 91.935 200.365 ;
        RECT 90.810 199.515 91.135 199.975 ;
        RECT 91.655 199.685 91.935 200.145 ;
        RECT 92.125 199.685 92.525 200.535 ;
        RECT 92.695 201.265 93.650 201.435 ;
        RECT 94.025 201.515 94.195 201.805 ;
        RECT 94.365 201.685 94.695 202.065 ;
        RECT 94.025 201.345 94.690 201.515 ;
        RECT 92.695 200.365 92.905 201.265 ;
        RECT 93.075 200.535 93.765 201.095 ;
        RECT 93.940 200.525 94.290 201.175 ;
        RECT 92.695 200.145 93.650 200.365 ;
        RECT 94.460 200.355 94.690 201.345 ;
        RECT 92.925 199.515 93.195 199.975 ;
        RECT 93.365 199.685 93.650 200.145 ;
        RECT 94.025 200.185 94.690 200.355 ;
        RECT 94.025 199.685 94.195 200.185 ;
        RECT 94.365 199.515 94.695 200.015 ;
        RECT 94.865 199.685 95.050 201.805 ;
        RECT 95.305 201.605 95.555 202.065 ;
        RECT 95.725 201.615 96.060 201.785 ;
        RECT 96.255 201.615 96.930 201.785 ;
        RECT 95.725 201.475 95.895 201.615 ;
        RECT 95.220 200.485 95.500 201.435 ;
        RECT 95.670 201.345 95.895 201.475 ;
        RECT 95.670 200.240 95.840 201.345 ;
        RECT 96.065 201.195 96.590 201.415 ;
        RECT 96.010 200.430 96.250 201.025 ;
        RECT 96.420 200.495 96.590 201.195 ;
        RECT 96.760 200.835 96.930 201.615 ;
        RECT 97.250 201.565 97.620 202.065 ;
        RECT 97.800 201.615 98.205 201.785 ;
        RECT 98.375 201.615 99.160 201.785 ;
        RECT 97.800 201.385 97.970 201.615 ;
        RECT 97.140 201.085 97.970 201.385 ;
        RECT 98.355 201.115 98.820 201.445 ;
        RECT 97.140 201.055 97.340 201.085 ;
        RECT 97.460 200.835 97.630 200.905 ;
        RECT 96.760 200.665 97.630 200.835 ;
        RECT 97.120 200.575 97.630 200.665 ;
        RECT 95.670 200.110 95.975 200.240 ;
        RECT 96.420 200.130 96.950 200.495 ;
        RECT 95.290 199.515 95.555 199.975 ;
        RECT 95.725 199.685 95.975 200.110 ;
        RECT 97.120 199.960 97.290 200.575 ;
        RECT 96.185 199.790 97.290 199.960 ;
        RECT 97.460 199.515 97.630 200.315 ;
        RECT 97.800 200.015 97.970 201.085 ;
        RECT 98.140 200.185 98.330 200.905 ;
        RECT 98.500 200.155 98.820 201.115 ;
        RECT 98.990 201.155 99.160 201.615 ;
        RECT 99.435 201.535 99.645 202.065 ;
        RECT 99.905 201.325 100.235 201.850 ;
        RECT 100.405 201.455 100.575 202.065 ;
        RECT 100.745 201.410 101.075 201.845 ;
        RECT 100.745 201.325 101.125 201.410 ;
        RECT 100.035 201.155 100.235 201.325 ;
        RECT 100.900 201.285 101.125 201.325 ;
        RECT 98.990 200.825 99.865 201.155 ;
        RECT 100.035 200.825 100.785 201.155 ;
        RECT 97.800 199.685 98.050 200.015 ;
        RECT 98.990 199.985 99.160 200.825 ;
        RECT 100.035 200.620 100.225 200.825 ;
        RECT 100.955 200.705 101.125 201.285 ;
        RECT 100.910 200.655 101.125 200.705 ;
        RECT 99.330 200.245 100.225 200.620 ;
        RECT 100.735 200.575 101.125 200.655 ;
        RECT 101.295 201.325 101.680 201.895 ;
        RECT 101.850 201.605 102.175 202.065 ;
        RECT 102.695 201.435 102.975 201.895 ;
        RECT 101.295 200.655 101.575 201.325 ;
        RECT 101.850 201.265 102.975 201.435 ;
        RECT 101.850 201.155 102.300 201.265 ;
        RECT 101.745 200.825 102.300 201.155 ;
        RECT 103.165 201.095 103.565 201.895 ;
        RECT 103.965 201.605 104.235 202.065 ;
        RECT 104.405 201.435 104.690 201.895 ;
        RECT 98.275 199.815 99.160 199.985 ;
        RECT 99.340 199.515 99.655 200.015 ;
        RECT 99.885 199.685 100.225 200.245 ;
        RECT 100.395 199.515 100.565 200.525 ;
        RECT 100.735 199.730 101.065 200.575 ;
        RECT 101.295 199.685 101.680 200.655 ;
        RECT 101.850 200.365 102.300 200.825 ;
        RECT 102.470 200.535 103.565 201.095 ;
        RECT 101.850 200.145 102.975 200.365 ;
        RECT 101.850 199.515 102.175 199.975 ;
        RECT 102.695 199.685 102.975 200.145 ;
        RECT 103.165 199.685 103.565 200.535 ;
        RECT 103.735 201.265 104.690 201.435 ;
        RECT 105.065 201.515 105.235 201.895 ;
        RECT 105.450 201.685 105.780 202.065 ;
        RECT 105.065 201.345 105.780 201.515 ;
        RECT 103.735 200.365 103.945 201.265 ;
        RECT 104.115 200.535 104.805 201.095 ;
        RECT 104.975 200.795 105.330 201.165 ;
        RECT 105.610 201.155 105.780 201.345 ;
        RECT 105.950 201.320 106.205 201.895 ;
        RECT 105.610 200.825 105.865 201.155 ;
        RECT 105.610 200.615 105.780 200.825 ;
        RECT 105.065 200.445 105.780 200.615 ;
        RECT 106.035 200.590 106.205 201.320 ;
        RECT 106.380 201.225 106.640 202.065 ;
        RECT 106.815 201.325 107.075 201.895 ;
        RECT 107.245 201.665 107.630 202.065 ;
        RECT 107.800 201.495 108.055 201.895 ;
        RECT 107.245 201.325 108.055 201.495 ;
        RECT 108.245 201.325 108.490 201.895 ;
        RECT 108.660 201.665 109.045 202.065 ;
        RECT 109.215 201.495 109.470 201.895 ;
        RECT 108.660 201.325 109.470 201.495 ;
        RECT 109.660 201.325 110.085 201.895 ;
        RECT 110.255 201.665 110.640 202.065 ;
        RECT 110.810 201.495 111.245 201.895 ;
        RECT 110.255 201.325 111.245 201.495 ;
        RECT 103.735 200.145 104.690 200.365 ;
        RECT 103.965 199.515 104.235 199.975 ;
        RECT 104.405 199.685 104.690 200.145 ;
        RECT 105.065 199.685 105.235 200.445 ;
        RECT 105.450 199.515 105.780 200.275 ;
        RECT 105.950 199.685 106.205 200.590 ;
        RECT 106.380 199.515 106.640 200.665 ;
        RECT 106.815 200.655 107.000 201.325 ;
        RECT 107.245 201.155 107.595 201.325 ;
        RECT 108.245 201.155 108.415 201.325 ;
        RECT 108.660 201.155 109.010 201.325 ;
        RECT 109.660 201.155 110.010 201.325 ;
        RECT 110.255 201.155 110.590 201.325 ;
        RECT 111.435 201.255 111.675 202.065 ;
        RECT 111.845 201.255 112.175 201.895 ;
        RECT 112.345 201.255 112.615 202.065 ;
        RECT 112.795 201.340 113.085 202.065 ;
        RECT 114.175 201.315 115.385 202.065 ;
        RECT 107.170 200.825 107.595 201.155 ;
        RECT 106.815 199.685 107.075 200.655 ;
        RECT 107.245 200.305 107.595 200.825 ;
        RECT 107.765 200.655 108.415 201.155 ;
        RECT 108.585 200.825 109.010 201.155 ;
        RECT 107.765 200.475 108.490 200.655 ;
        RECT 107.245 200.110 108.055 200.305 ;
        RECT 107.245 199.515 107.630 199.940 ;
        RECT 107.800 199.685 108.055 200.110 ;
        RECT 108.245 199.685 108.490 200.475 ;
        RECT 108.660 200.305 109.010 200.825 ;
        RECT 109.180 200.655 110.010 201.155 ;
        RECT 110.180 200.825 110.590 201.155 ;
        RECT 109.180 200.475 110.085 200.655 ;
        RECT 108.660 200.110 109.490 200.305 ;
        RECT 108.660 199.515 109.045 199.940 ;
        RECT 109.215 199.685 109.490 200.110 ;
        RECT 109.660 199.685 110.085 200.475 ;
        RECT 110.255 200.280 110.590 200.825 ;
        RECT 110.760 200.450 111.245 201.155 ;
        RECT 111.415 200.825 111.765 201.075 ;
        RECT 111.935 200.655 112.105 201.255 ;
        RECT 112.275 200.825 112.625 201.075 ;
        RECT 111.425 200.485 112.105 200.655 ;
        RECT 110.255 200.110 111.245 200.280 ;
        RECT 110.255 199.515 110.640 199.940 ;
        RECT 110.810 199.685 111.245 200.110 ;
        RECT 111.425 199.700 111.755 200.485 ;
        RECT 112.285 199.515 112.615 200.655 ;
        RECT 112.795 199.515 113.085 200.680 ;
        RECT 114.175 200.605 114.695 201.145 ;
        RECT 114.865 200.775 115.385 201.315 ;
        RECT 114.175 199.515 115.385 200.605 ;
        RECT 61.190 199.345 115.470 199.515 ;
        RECT 61.275 198.255 62.485 199.345 ;
        RECT 61.275 197.545 61.795 198.085 ;
        RECT 61.965 197.715 62.485 198.255 ;
        RECT 63.635 198.205 63.845 199.345 ;
        RECT 64.015 198.195 64.345 199.175 ;
        RECT 64.515 198.205 64.745 199.345 ;
        RECT 65.015 198.285 65.345 199.130 ;
        RECT 65.515 198.335 65.685 199.345 ;
        RECT 65.855 198.615 66.195 199.175 ;
        RECT 66.425 198.845 66.740 199.345 ;
        RECT 66.920 198.875 67.805 199.045 ;
        RECT 64.955 198.205 65.345 198.285 ;
        RECT 65.855 198.240 66.750 198.615 ;
        RECT 61.275 196.795 62.485 197.545 ;
        RECT 63.635 196.795 63.845 197.615 ;
        RECT 64.015 197.595 64.265 198.195 ;
        RECT 64.955 198.155 65.170 198.205 ;
        RECT 64.435 197.785 64.765 198.035 ;
        RECT 64.015 196.965 64.345 197.595 ;
        RECT 64.515 196.795 64.745 197.615 ;
        RECT 64.955 197.575 65.125 198.155 ;
        RECT 65.855 198.035 66.045 198.240 ;
        RECT 66.920 198.035 67.090 198.875 ;
        RECT 68.030 198.845 68.280 199.175 ;
        RECT 65.295 197.705 66.045 198.035 ;
        RECT 66.215 197.705 67.090 198.035 ;
        RECT 64.955 197.535 65.180 197.575 ;
        RECT 65.845 197.535 66.045 197.705 ;
        RECT 64.955 197.450 65.335 197.535 ;
        RECT 65.005 197.015 65.335 197.450 ;
        RECT 65.505 196.795 65.675 197.405 ;
        RECT 65.845 197.010 66.175 197.535 ;
        RECT 66.435 196.795 66.645 197.325 ;
        RECT 66.920 197.245 67.090 197.705 ;
        RECT 67.260 197.745 67.580 198.705 ;
        RECT 67.750 197.955 67.940 198.675 ;
        RECT 68.110 197.775 68.280 198.845 ;
        RECT 68.450 198.545 68.620 199.345 ;
        RECT 68.790 198.900 69.895 199.070 ;
        RECT 68.790 198.285 68.960 198.900 ;
        RECT 70.105 198.750 70.355 199.175 ;
        RECT 70.525 198.885 70.790 199.345 ;
        RECT 69.130 198.365 69.660 198.730 ;
        RECT 70.105 198.620 70.410 198.750 ;
        RECT 68.450 198.195 68.960 198.285 ;
        RECT 68.450 198.025 69.320 198.195 ;
        RECT 68.450 197.955 68.620 198.025 ;
        RECT 68.740 197.775 68.940 197.805 ;
        RECT 67.260 197.415 67.725 197.745 ;
        RECT 68.110 197.475 68.940 197.775 ;
        RECT 68.110 197.245 68.280 197.475 ;
        RECT 66.920 197.075 67.705 197.245 ;
        RECT 67.875 197.075 68.280 197.245 ;
        RECT 68.460 196.795 68.830 197.295 ;
        RECT 69.150 197.245 69.320 198.025 ;
        RECT 69.490 197.665 69.660 198.365 ;
        RECT 69.830 197.835 70.070 198.430 ;
        RECT 69.490 197.445 70.015 197.665 ;
        RECT 70.240 197.515 70.410 198.620 ;
        RECT 70.185 197.385 70.410 197.515 ;
        RECT 70.580 197.425 70.860 198.375 ;
        RECT 70.185 197.245 70.355 197.385 ;
        RECT 69.150 197.075 69.825 197.245 ;
        RECT 70.020 197.075 70.355 197.245 ;
        RECT 70.525 196.795 70.775 197.255 ;
        RECT 71.030 197.055 71.215 199.175 ;
        RECT 71.385 198.845 71.715 199.345 ;
        RECT 71.885 198.675 72.055 199.175 ;
        RECT 71.390 198.505 72.055 198.675 ;
        RECT 71.390 197.515 71.620 198.505 ;
        RECT 71.790 197.685 72.140 198.335 ;
        RECT 72.320 198.195 72.580 199.345 ;
        RECT 72.755 198.270 73.010 199.175 ;
        RECT 73.180 198.585 73.510 199.345 ;
        RECT 73.725 198.415 73.895 199.175 ;
        RECT 71.390 197.345 72.055 197.515 ;
        RECT 71.385 196.795 71.715 197.175 ;
        RECT 71.885 197.055 72.055 197.345 ;
        RECT 72.320 196.795 72.580 197.635 ;
        RECT 72.755 197.540 72.925 198.270 ;
        RECT 73.180 198.245 73.895 198.415 ;
        RECT 73.180 198.035 73.350 198.245 ;
        RECT 74.155 198.180 74.445 199.345 ;
        RECT 75.625 198.675 75.795 199.175 ;
        RECT 75.965 198.845 76.295 199.345 ;
        RECT 75.625 198.505 76.290 198.675 ;
        RECT 73.095 197.705 73.350 198.035 ;
        RECT 72.755 196.965 73.010 197.540 ;
        RECT 73.180 197.515 73.350 197.705 ;
        RECT 73.630 197.695 73.985 198.065 ;
        RECT 75.540 197.685 75.890 198.335 ;
        RECT 73.180 197.345 73.895 197.515 ;
        RECT 73.180 196.795 73.510 197.175 ;
        RECT 73.725 196.965 73.895 197.345 ;
        RECT 74.155 196.795 74.445 197.520 ;
        RECT 76.060 197.515 76.290 198.505 ;
        RECT 75.625 197.345 76.290 197.515 ;
        RECT 75.625 197.055 75.795 197.345 ;
        RECT 75.965 196.795 76.295 197.175 ;
        RECT 76.465 197.055 76.650 199.175 ;
        RECT 76.890 198.885 77.155 199.345 ;
        RECT 77.325 198.750 77.575 199.175 ;
        RECT 77.785 198.900 78.890 199.070 ;
        RECT 77.270 198.620 77.575 198.750 ;
        RECT 76.820 197.425 77.100 198.375 ;
        RECT 77.270 197.515 77.440 198.620 ;
        RECT 77.610 197.835 77.850 198.430 ;
        RECT 78.020 198.365 78.550 198.730 ;
        RECT 78.020 197.665 78.190 198.365 ;
        RECT 78.720 198.285 78.890 198.900 ;
        RECT 79.060 198.545 79.230 199.345 ;
        RECT 79.400 198.845 79.650 199.175 ;
        RECT 79.875 198.875 80.760 199.045 ;
        RECT 78.720 198.195 79.230 198.285 ;
        RECT 77.270 197.385 77.495 197.515 ;
        RECT 77.665 197.445 78.190 197.665 ;
        RECT 78.360 198.025 79.230 198.195 ;
        RECT 76.905 196.795 77.155 197.255 ;
        RECT 77.325 197.245 77.495 197.385 ;
        RECT 78.360 197.245 78.530 198.025 ;
        RECT 79.060 197.955 79.230 198.025 ;
        RECT 78.740 197.775 78.940 197.805 ;
        RECT 79.400 197.775 79.570 198.845 ;
        RECT 79.740 197.955 79.930 198.675 ;
        RECT 78.740 197.475 79.570 197.775 ;
        RECT 80.100 197.745 80.420 198.705 ;
        RECT 77.325 197.075 77.660 197.245 ;
        RECT 77.855 197.075 78.530 197.245 ;
        RECT 78.850 196.795 79.220 197.295 ;
        RECT 79.400 197.245 79.570 197.475 ;
        RECT 79.955 197.415 80.420 197.745 ;
        RECT 80.590 198.035 80.760 198.875 ;
        RECT 80.940 198.845 81.255 199.345 ;
        RECT 81.485 198.615 81.825 199.175 ;
        RECT 80.930 198.240 81.825 198.615 ;
        RECT 81.995 198.335 82.165 199.345 ;
        RECT 81.635 198.035 81.825 198.240 ;
        RECT 82.335 198.285 82.665 199.130 ;
        RECT 82.335 198.205 82.725 198.285 ;
        RECT 82.510 198.155 82.725 198.205 ;
        RECT 82.900 198.195 83.160 199.345 ;
        RECT 83.335 198.270 83.590 199.175 ;
        RECT 83.760 198.585 84.090 199.345 ;
        RECT 84.305 198.415 84.475 199.175 ;
        RECT 80.590 197.705 81.465 198.035 ;
        RECT 81.635 197.705 82.385 198.035 ;
        RECT 80.590 197.245 80.760 197.705 ;
        RECT 81.635 197.535 81.835 197.705 ;
        RECT 82.555 197.575 82.725 198.155 ;
        RECT 82.500 197.535 82.725 197.575 ;
        RECT 79.400 197.075 79.805 197.245 ;
        RECT 79.975 197.075 80.760 197.245 ;
        RECT 81.035 196.795 81.245 197.325 ;
        RECT 81.505 197.010 81.835 197.535 ;
        RECT 82.345 197.450 82.725 197.535 ;
        RECT 82.005 196.795 82.175 197.405 ;
        RECT 82.345 197.015 82.675 197.450 ;
        RECT 82.900 196.795 83.160 197.635 ;
        RECT 83.335 197.540 83.505 198.270 ;
        RECT 83.760 198.245 84.475 198.415 ;
        RECT 84.745 198.395 85.020 199.165 ;
        RECT 85.190 198.735 85.520 199.165 ;
        RECT 85.690 198.905 85.885 199.345 ;
        RECT 86.065 198.735 86.395 199.165 ;
        RECT 85.190 198.565 86.395 198.735 ;
        RECT 83.760 198.035 83.930 198.245 ;
        RECT 84.745 198.205 85.330 198.395 ;
        RECT 85.500 198.235 86.395 198.565 ;
        RECT 86.665 198.675 86.835 199.175 ;
        RECT 87.005 198.845 87.335 199.345 ;
        RECT 86.665 198.505 87.330 198.675 ;
        RECT 83.675 197.705 83.930 198.035 ;
        RECT 83.335 196.965 83.590 197.540 ;
        RECT 83.760 197.515 83.930 197.705 ;
        RECT 84.210 197.695 84.565 198.065 ;
        RECT 83.760 197.345 84.475 197.515 ;
        RECT 84.745 197.385 84.985 198.035 ;
        RECT 85.155 197.535 85.330 198.205 ;
        RECT 85.500 197.705 85.915 198.035 ;
        RECT 86.095 197.705 86.390 198.035 ;
        RECT 85.155 197.355 85.485 197.535 ;
        RECT 83.760 196.795 84.090 197.175 ;
        RECT 84.305 196.965 84.475 197.345 ;
        RECT 84.760 196.795 85.090 197.185 ;
        RECT 85.260 196.975 85.485 197.355 ;
        RECT 85.685 197.085 85.915 197.705 ;
        RECT 86.580 197.685 86.930 198.335 ;
        RECT 86.095 196.795 86.395 197.525 ;
        RECT 87.100 197.515 87.330 198.505 ;
        RECT 86.665 197.345 87.330 197.515 ;
        RECT 86.665 197.055 86.835 197.345 ;
        RECT 87.005 196.795 87.335 197.175 ;
        RECT 87.505 197.055 87.690 199.175 ;
        RECT 87.930 198.885 88.195 199.345 ;
        RECT 88.365 198.750 88.615 199.175 ;
        RECT 88.825 198.900 89.930 199.070 ;
        RECT 88.310 198.620 88.615 198.750 ;
        RECT 87.860 197.425 88.140 198.375 ;
        RECT 88.310 197.515 88.480 198.620 ;
        RECT 88.650 197.835 88.890 198.430 ;
        RECT 89.060 198.365 89.590 198.730 ;
        RECT 89.060 197.665 89.230 198.365 ;
        RECT 89.760 198.285 89.930 198.900 ;
        RECT 90.100 198.545 90.270 199.345 ;
        RECT 90.440 198.845 90.690 199.175 ;
        RECT 90.915 198.875 91.800 199.045 ;
        RECT 89.760 198.195 90.270 198.285 ;
        RECT 88.310 197.385 88.535 197.515 ;
        RECT 88.705 197.445 89.230 197.665 ;
        RECT 89.400 198.025 90.270 198.195 ;
        RECT 87.945 196.795 88.195 197.255 ;
        RECT 88.365 197.245 88.535 197.385 ;
        RECT 89.400 197.245 89.570 198.025 ;
        RECT 90.100 197.955 90.270 198.025 ;
        RECT 89.780 197.775 89.980 197.805 ;
        RECT 90.440 197.775 90.610 198.845 ;
        RECT 90.780 197.955 90.970 198.675 ;
        RECT 89.780 197.475 90.610 197.775 ;
        RECT 91.140 197.745 91.460 198.705 ;
        RECT 88.365 197.075 88.700 197.245 ;
        RECT 88.895 197.075 89.570 197.245 ;
        RECT 89.890 196.795 90.260 197.295 ;
        RECT 90.440 197.245 90.610 197.475 ;
        RECT 90.995 197.415 91.460 197.745 ;
        RECT 91.630 198.035 91.800 198.875 ;
        RECT 91.980 198.845 92.295 199.345 ;
        RECT 92.525 198.615 92.865 199.175 ;
        RECT 91.970 198.240 92.865 198.615 ;
        RECT 93.035 198.335 93.205 199.345 ;
        RECT 92.675 198.035 92.865 198.240 ;
        RECT 93.375 198.285 93.705 199.130 ;
        RECT 93.935 198.915 94.275 199.175 ;
        RECT 93.375 198.205 93.765 198.285 ;
        RECT 93.550 198.155 93.765 198.205 ;
        RECT 91.630 197.705 92.505 198.035 ;
        RECT 92.675 197.705 93.425 198.035 ;
        RECT 91.630 197.245 91.800 197.705 ;
        RECT 92.675 197.535 92.875 197.705 ;
        RECT 93.595 197.575 93.765 198.155 ;
        RECT 93.540 197.535 93.765 197.575 ;
        RECT 90.440 197.075 90.845 197.245 ;
        RECT 91.015 197.075 91.800 197.245 ;
        RECT 92.075 196.795 92.285 197.325 ;
        RECT 92.545 197.010 92.875 197.535 ;
        RECT 93.385 197.450 93.765 197.535 ;
        RECT 93.935 197.515 94.195 198.915 ;
        RECT 94.445 198.545 94.775 199.345 ;
        RECT 95.240 198.375 95.490 199.175 ;
        RECT 95.675 198.625 96.005 199.345 ;
        RECT 96.225 198.375 96.475 199.175 ;
        RECT 96.645 198.965 96.980 199.345 ;
        RECT 94.385 198.205 96.575 198.375 ;
        RECT 94.385 198.035 94.700 198.205 ;
        RECT 94.370 197.785 94.700 198.035 ;
        RECT 93.045 196.795 93.215 197.405 ;
        RECT 93.385 197.015 93.715 197.450 ;
        RECT 93.935 197.005 94.275 197.515 ;
        RECT 94.445 196.795 94.715 197.595 ;
        RECT 94.895 197.065 95.175 198.035 ;
        RECT 95.355 197.065 95.655 198.035 ;
        RECT 95.835 197.070 96.185 198.035 ;
        RECT 96.405 197.295 96.575 198.205 ;
        RECT 96.745 197.475 96.985 198.785 ;
        RECT 97.155 198.475 97.430 199.175 ;
        RECT 97.600 198.800 97.855 199.345 ;
        RECT 98.025 198.835 98.505 199.175 ;
        RECT 98.680 198.790 99.285 199.345 ;
        RECT 98.670 198.690 99.285 198.790 ;
        RECT 98.670 198.665 98.855 198.690 ;
        RECT 97.155 197.445 97.325 198.475 ;
        RECT 97.600 198.345 98.355 198.595 ;
        RECT 98.525 198.420 98.855 198.665 ;
        RECT 97.600 198.310 98.370 198.345 ;
        RECT 97.600 198.300 98.385 198.310 ;
        RECT 97.495 198.285 98.390 198.300 ;
        RECT 97.495 198.270 98.410 198.285 ;
        RECT 97.495 198.260 98.430 198.270 ;
        RECT 97.495 198.250 98.455 198.260 ;
        RECT 97.495 198.220 98.525 198.250 ;
        RECT 97.495 198.190 98.545 198.220 ;
        RECT 97.495 198.160 98.565 198.190 ;
        RECT 97.495 198.135 98.595 198.160 ;
        RECT 97.495 198.100 98.630 198.135 ;
        RECT 97.495 198.095 98.660 198.100 ;
        RECT 97.495 197.700 97.725 198.095 ;
        RECT 98.270 198.090 98.660 198.095 ;
        RECT 98.295 198.080 98.660 198.090 ;
        RECT 98.310 198.075 98.660 198.080 ;
        RECT 98.325 198.070 98.660 198.075 ;
        RECT 99.025 198.070 99.285 198.520 ;
        RECT 99.915 198.180 100.205 199.345 ;
        RECT 100.385 198.625 100.715 199.345 ;
        RECT 98.325 198.065 99.285 198.070 ;
        RECT 98.335 198.055 99.285 198.065 ;
        RECT 98.345 198.050 99.285 198.055 ;
        RECT 98.355 198.040 99.285 198.050 ;
        RECT 98.360 198.030 99.285 198.040 ;
        RECT 98.365 198.025 99.285 198.030 ;
        RECT 98.375 198.010 99.285 198.025 ;
        RECT 98.380 197.995 99.285 198.010 ;
        RECT 98.390 197.970 99.285 197.995 ;
        RECT 97.895 197.500 98.225 197.925 ;
        RECT 96.405 196.965 96.900 197.295 ;
        RECT 97.155 196.965 97.415 197.445 ;
        RECT 97.585 196.795 97.835 197.335 ;
        RECT 98.005 197.015 98.225 197.500 ;
        RECT 98.395 197.900 99.285 197.970 ;
        RECT 100.375 197.985 100.605 198.325 ;
        RECT 100.895 197.985 101.110 199.100 ;
        RECT 101.305 198.400 101.635 199.175 ;
        RECT 101.805 198.570 102.515 199.345 ;
        RECT 101.305 198.185 102.455 198.400 ;
        RECT 98.395 197.175 98.565 197.900 ;
        RECT 100.375 197.785 100.705 197.985 ;
        RECT 100.895 197.805 101.345 197.985 ;
        RECT 101.015 197.785 101.345 197.805 ;
        RECT 101.515 197.785 101.985 198.015 ;
        RECT 98.735 197.345 99.285 197.730 ;
        RECT 102.170 197.615 102.455 198.185 ;
        RECT 102.685 197.740 102.965 199.175 ;
        RECT 103.225 198.675 103.395 199.175 ;
        RECT 103.565 198.845 103.895 199.345 ;
        RECT 103.225 198.505 103.890 198.675 ;
        RECT 98.395 197.005 99.285 197.175 ;
        RECT 99.915 196.795 100.205 197.520 ;
        RECT 100.375 197.425 101.555 197.615 ;
        RECT 100.375 196.965 100.715 197.425 ;
        RECT 101.225 197.345 101.555 197.425 ;
        RECT 101.745 197.425 102.455 197.615 ;
        RECT 101.745 197.285 102.045 197.425 ;
        RECT 101.730 197.275 102.045 197.285 ;
        RECT 101.720 197.265 102.045 197.275 ;
        RECT 101.710 197.260 102.045 197.265 ;
        RECT 100.885 196.795 101.055 197.255 ;
        RECT 101.705 197.250 102.045 197.260 ;
        RECT 101.700 197.245 102.045 197.250 ;
        RECT 101.695 197.235 102.045 197.245 ;
        RECT 101.690 197.230 102.045 197.235 ;
        RECT 101.685 196.965 102.045 197.230 ;
        RECT 102.285 196.795 102.455 197.255 ;
        RECT 102.625 196.965 102.965 197.740 ;
        RECT 103.140 197.685 103.490 198.335 ;
        RECT 103.660 197.515 103.890 198.505 ;
        RECT 103.225 197.345 103.890 197.515 ;
        RECT 103.225 197.055 103.395 197.345 ;
        RECT 103.565 196.795 103.895 197.175 ;
        RECT 104.065 197.055 104.250 199.175 ;
        RECT 104.490 198.885 104.755 199.345 ;
        RECT 104.925 198.750 105.175 199.175 ;
        RECT 105.385 198.900 106.490 199.070 ;
        RECT 104.870 198.620 105.175 198.750 ;
        RECT 104.420 197.425 104.700 198.375 ;
        RECT 104.870 197.515 105.040 198.620 ;
        RECT 105.210 197.835 105.450 198.430 ;
        RECT 105.620 198.365 106.150 198.730 ;
        RECT 105.620 197.665 105.790 198.365 ;
        RECT 106.320 198.285 106.490 198.900 ;
        RECT 106.660 198.545 106.830 199.345 ;
        RECT 107.000 198.845 107.250 199.175 ;
        RECT 107.475 198.875 108.360 199.045 ;
        RECT 106.320 198.195 106.830 198.285 ;
        RECT 104.870 197.385 105.095 197.515 ;
        RECT 105.265 197.445 105.790 197.665 ;
        RECT 105.960 198.025 106.830 198.195 ;
        RECT 104.505 196.795 104.755 197.255 ;
        RECT 104.925 197.245 105.095 197.385 ;
        RECT 105.960 197.245 106.130 198.025 ;
        RECT 106.660 197.955 106.830 198.025 ;
        RECT 106.340 197.775 106.540 197.805 ;
        RECT 107.000 197.775 107.170 198.845 ;
        RECT 107.340 197.955 107.530 198.675 ;
        RECT 106.340 197.475 107.170 197.775 ;
        RECT 107.700 197.745 108.020 198.705 ;
        RECT 104.925 197.075 105.260 197.245 ;
        RECT 105.455 197.075 106.130 197.245 ;
        RECT 106.450 196.795 106.820 197.295 ;
        RECT 107.000 197.245 107.170 197.475 ;
        RECT 107.555 197.415 108.020 197.745 ;
        RECT 108.190 198.035 108.360 198.875 ;
        RECT 108.540 198.845 108.855 199.345 ;
        RECT 109.085 198.615 109.425 199.175 ;
        RECT 108.530 198.240 109.425 198.615 ;
        RECT 109.595 198.335 109.765 199.345 ;
        RECT 109.235 198.035 109.425 198.240 ;
        RECT 109.935 198.285 110.265 199.130 ;
        RECT 109.935 198.205 110.325 198.285 ;
        RECT 110.110 198.155 110.325 198.205 ;
        RECT 108.190 197.705 109.065 198.035 ;
        RECT 109.235 197.705 109.985 198.035 ;
        RECT 108.190 197.245 108.360 197.705 ;
        RECT 109.235 197.535 109.435 197.705 ;
        RECT 110.155 197.575 110.325 198.155 ;
        RECT 110.100 197.535 110.325 197.575 ;
        RECT 107.000 197.075 107.405 197.245 ;
        RECT 107.575 197.075 108.360 197.245 ;
        RECT 108.635 196.795 108.845 197.325 ;
        RECT 109.105 197.010 109.435 197.535 ;
        RECT 109.945 197.450 110.325 197.535 ;
        RECT 110.495 198.205 110.880 199.175 ;
        RECT 111.050 198.885 111.375 199.345 ;
        RECT 111.895 198.715 112.175 199.175 ;
        RECT 111.050 198.495 112.175 198.715 ;
        RECT 110.495 197.535 110.775 198.205 ;
        RECT 111.050 198.035 111.500 198.495 ;
        RECT 112.365 198.325 112.765 199.175 ;
        RECT 113.165 198.885 113.435 199.345 ;
        RECT 113.605 198.715 113.890 199.175 ;
        RECT 110.945 197.705 111.500 198.035 ;
        RECT 111.670 197.765 112.765 198.325 ;
        RECT 111.050 197.595 111.500 197.705 ;
        RECT 109.605 196.795 109.775 197.405 ;
        RECT 109.945 197.015 110.275 197.450 ;
        RECT 110.495 196.965 110.880 197.535 ;
        RECT 111.050 197.425 112.175 197.595 ;
        RECT 111.050 196.795 111.375 197.255 ;
        RECT 111.895 196.965 112.175 197.425 ;
        RECT 112.365 196.965 112.765 197.765 ;
        RECT 112.935 198.495 113.890 198.715 ;
        RECT 112.935 197.595 113.145 198.495 ;
        RECT 113.315 197.765 114.005 198.325 ;
        RECT 114.175 198.255 115.385 199.345 ;
        RECT 114.175 197.715 114.695 198.255 ;
        RECT 112.935 197.425 113.890 197.595 ;
        RECT 114.865 197.545 115.385 198.085 ;
        RECT 113.165 196.795 113.435 197.255 ;
        RECT 113.605 196.965 113.890 197.425 ;
        RECT 114.175 196.795 115.385 197.545 ;
        RECT 61.190 196.625 115.470 196.795 ;
        RECT 61.275 195.875 62.485 196.625 ;
        RECT 62.655 196.080 68.000 196.625 ;
        RECT 61.275 195.335 61.795 195.875 ;
        RECT 61.965 195.165 62.485 195.705 ;
        RECT 64.240 195.250 64.580 196.080 ;
        RECT 68.175 195.855 69.845 196.625 ;
        RECT 70.485 195.900 70.815 196.410 ;
        RECT 70.985 196.225 71.315 196.625 ;
        RECT 72.365 196.055 72.695 196.395 ;
        RECT 72.865 196.225 73.195 196.625 ;
        RECT 61.275 194.075 62.485 195.165 ;
        RECT 66.060 194.510 66.410 195.760 ;
        RECT 68.175 195.335 68.925 195.855 ;
        RECT 69.095 195.165 69.845 195.685 ;
        RECT 62.655 194.075 68.000 194.510 ;
        RECT 68.175 194.075 69.845 195.165 ;
        RECT 70.485 195.135 70.675 195.900 ;
        RECT 70.985 195.885 73.350 196.055 ;
        RECT 70.985 195.715 71.155 195.885 ;
        RECT 70.845 195.385 71.155 195.715 ;
        RECT 71.325 195.385 71.630 195.715 ;
        RECT 70.485 194.285 70.815 195.135 ;
        RECT 70.985 194.075 71.235 195.215 ;
        RECT 71.415 195.055 71.630 195.385 ;
        RECT 71.805 195.055 72.090 195.715 ;
        RECT 72.285 195.055 72.550 195.715 ;
        RECT 72.765 195.055 73.010 195.715 ;
        RECT 73.180 194.885 73.350 195.885 ;
        RECT 71.425 194.715 72.715 194.885 ;
        RECT 71.425 194.295 71.675 194.715 ;
        RECT 71.905 194.075 72.235 194.545 ;
        RECT 72.465 194.295 72.715 194.715 ;
        RECT 72.895 194.715 73.350 194.885 ;
        RECT 74.615 195.975 74.875 196.455 ;
        RECT 75.045 196.085 75.295 196.625 ;
        RECT 74.615 194.945 74.785 195.975 ;
        RECT 75.465 195.920 75.685 196.405 ;
        RECT 74.955 195.325 75.185 195.720 ;
        RECT 75.355 195.495 75.685 195.920 ;
        RECT 75.855 196.245 76.745 196.415 ;
        RECT 75.855 195.520 76.025 196.245 ;
        RECT 77.005 196.145 77.305 196.625 ;
        RECT 76.195 195.690 76.745 196.075 ;
        RECT 77.475 195.975 77.735 196.430 ;
        RECT 77.905 196.145 78.165 196.625 ;
        RECT 78.345 195.975 78.605 196.430 ;
        RECT 78.775 196.145 79.025 196.625 ;
        RECT 79.205 195.975 79.465 196.430 ;
        RECT 79.635 196.145 79.885 196.625 ;
        RECT 80.065 195.975 80.325 196.430 ;
        RECT 80.495 196.145 80.740 196.625 ;
        RECT 80.910 195.975 81.185 196.430 ;
        RECT 81.355 196.145 81.600 196.625 ;
        RECT 81.770 195.975 82.030 196.430 ;
        RECT 82.200 196.145 82.460 196.625 ;
        RECT 82.630 195.975 82.890 196.430 ;
        RECT 83.060 196.145 83.320 196.625 ;
        RECT 83.490 195.975 83.750 196.430 ;
        RECT 83.920 196.065 84.180 196.625 ;
        RECT 77.005 195.805 83.750 195.975 ;
        RECT 75.855 195.450 76.745 195.520 ;
        RECT 75.850 195.425 76.745 195.450 ;
        RECT 75.840 195.410 76.745 195.425 ;
        RECT 75.835 195.395 76.745 195.410 ;
        RECT 75.825 195.390 76.745 195.395 ;
        RECT 75.820 195.380 76.745 195.390 ;
        RECT 75.815 195.370 76.745 195.380 ;
        RECT 75.805 195.365 76.745 195.370 ;
        RECT 75.795 195.355 76.745 195.365 ;
        RECT 75.785 195.350 76.745 195.355 ;
        RECT 75.785 195.345 76.120 195.350 ;
        RECT 75.770 195.340 76.120 195.345 ;
        RECT 75.755 195.330 76.120 195.340 ;
        RECT 75.730 195.325 76.120 195.330 ;
        RECT 74.955 195.320 76.120 195.325 ;
        RECT 74.955 195.285 76.090 195.320 ;
        RECT 74.955 195.260 76.055 195.285 ;
        RECT 74.955 195.230 76.025 195.260 ;
        RECT 74.955 195.200 76.005 195.230 ;
        RECT 74.955 195.170 75.985 195.200 ;
        RECT 74.955 195.160 75.915 195.170 ;
        RECT 74.955 195.150 75.890 195.160 ;
        RECT 74.955 195.135 75.870 195.150 ;
        RECT 74.955 195.120 75.850 195.135 ;
        RECT 75.060 195.110 75.845 195.120 ;
        RECT 75.060 195.075 75.830 195.110 ;
        RECT 72.895 194.285 73.225 194.715 ;
        RECT 74.615 194.245 74.890 194.945 ;
        RECT 75.060 194.825 75.815 195.075 ;
        RECT 75.985 194.755 76.315 195.000 ;
        RECT 76.485 194.900 76.745 195.350 ;
        RECT 77.005 195.265 78.170 195.805 ;
        RECT 84.350 195.635 84.600 196.445 ;
        RECT 84.780 196.100 85.040 196.625 ;
        RECT 85.210 195.635 85.460 196.445 ;
        RECT 85.640 196.115 85.945 196.625 ;
        RECT 78.340 195.385 85.460 195.635 ;
        RECT 85.630 195.385 85.945 195.945 ;
        RECT 87.035 195.900 87.325 196.625 ;
        RECT 87.495 195.950 87.755 196.455 ;
        RECT 87.935 196.245 88.265 196.625 ;
        RECT 88.445 196.075 88.615 196.455 ;
        RECT 88.965 196.145 89.265 196.625 ;
        RECT 76.975 195.215 78.170 195.265 ;
        RECT 76.975 195.095 83.750 195.215 ;
        RECT 77.005 194.990 83.750 195.095 ;
        RECT 76.130 194.730 76.315 194.755 ;
        RECT 76.130 194.630 76.745 194.730 ;
        RECT 75.060 194.075 75.315 194.620 ;
        RECT 75.485 194.245 75.965 194.585 ;
        RECT 76.140 194.075 76.745 194.630 ;
        RECT 77.005 194.075 77.275 194.820 ;
        RECT 77.445 194.250 77.735 194.990 ;
        RECT 78.345 194.975 83.750 194.990 ;
        RECT 77.905 194.080 78.160 194.805 ;
        RECT 78.345 194.250 78.605 194.975 ;
        RECT 78.775 194.080 79.020 194.805 ;
        RECT 79.205 194.250 79.465 194.975 ;
        RECT 79.635 194.080 79.880 194.805 ;
        RECT 80.065 194.250 80.325 194.975 ;
        RECT 80.495 194.080 80.740 194.805 ;
        RECT 80.910 194.250 81.170 194.975 ;
        RECT 81.340 194.080 81.600 194.805 ;
        RECT 81.770 194.250 82.030 194.975 ;
        RECT 82.200 194.080 82.460 194.805 ;
        RECT 82.630 194.250 82.890 194.975 ;
        RECT 83.060 194.080 83.320 194.805 ;
        RECT 83.490 194.250 83.750 194.975 ;
        RECT 83.920 194.080 84.180 194.875 ;
        RECT 84.350 194.250 84.600 195.385 ;
        RECT 77.905 194.075 84.180 194.080 ;
        RECT 84.780 194.075 85.040 194.885 ;
        RECT 85.215 194.245 85.460 195.385 ;
        RECT 85.640 194.075 85.935 194.885 ;
        RECT 87.035 194.075 87.325 195.240 ;
        RECT 87.495 195.150 87.665 195.950 ;
        RECT 87.950 195.905 88.615 196.075 ;
        RECT 89.435 195.975 89.695 196.430 ;
        RECT 89.865 196.145 90.125 196.625 ;
        RECT 90.305 195.975 90.565 196.430 ;
        RECT 90.735 196.145 90.985 196.625 ;
        RECT 91.165 195.975 91.425 196.430 ;
        RECT 91.595 196.145 91.845 196.625 ;
        RECT 92.025 195.975 92.285 196.430 ;
        RECT 92.455 196.145 92.700 196.625 ;
        RECT 92.870 195.975 93.145 196.430 ;
        RECT 93.315 196.145 93.560 196.625 ;
        RECT 93.730 195.975 93.990 196.430 ;
        RECT 94.160 196.145 94.420 196.625 ;
        RECT 94.590 195.975 94.850 196.430 ;
        RECT 95.020 196.145 95.280 196.625 ;
        RECT 95.450 195.975 95.710 196.430 ;
        RECT 95.880 196.065 96.140 196.625 ;
        RECT 87.950 195.650 88.120 195.905 ;
        RECT 88.965 195.805 95.710 195.975 ;
        RECT 87.835 195.320 88.120 195.650 ;
        RECT 88.355 195.355 88.685 195.725 ;
        RECT 87.950 195.175 88.120 195.320 ;
        RECT 88.965 195.215 90.130 195.805 ;
        RECT 96.310 195.635 96.560 196.445 ;
        RECT 96.740 196.100 97.000 196.625 ;
        RECT 97.170 195.635 97.420 196.445 ;
        RECT 97.600 196.115 97.905 196.625 ;
        RECT 90.300 195.385 97.420 195.635 ;
        RECT 97.590 195.385 97.905 195.945 ;
        RECT 98.535 195.680 98.875 196.455 ;
        RECT 99.045 196.165 99.215 196.625 ;
        RECT 99.455 196.190 99.815 196.455 ;
        RECT 99.455 196.185 99.810 196.190 ;
        RECT 99.455 196.175 99.805 196.185 ;
        RECT 99.455 196.170 99.800 196.175 ;
        RECT 99.455 196.160 99.795 196.170 ;
        RECT 100.445 196.165 100.615 196.625 ;
        RECT 99.455 196.155 99.790 196.160 ;
        RECT 99.455 196.145 99.780 196.155 ;
        RECT 99.455 196.135 99.770 196.145 ;
        RECT 99.455 195.995 99.755 196.135 ;
        RECT 99.045 195.805 99.755 195.995 ;
        RECT 99.945 195.995 100.275 196.075 ;
        RECT 100.785 195.995 101.125 196.455 ;
        RECT 101.295 196.115 101.600 196.625 ;
        RECT 99.945 195.805 101.125 195.995 ;
        RECT 87.495 194.245 87.765 195.150 ;
        RECT 87.950 195.005 88.615 195.175 ;
        RECT 87.935 194.075 88.265 194.835 ;
        RECT 88.445 194.245 88.615 195.005 ;
        RECT 88.965 194.990 95.710 195.215 ;
        RECT 88.965 194.075 89.235 194.820 ;
        RECT 89.405 194.250 89.695 194.990 ;
        RECT 90.305 194.975 95.710 194.990 ;
        RECT 89.865 194.080 90.120 194.805 ;
        RECT 90.305 194.250 90.565 194.975 ;
        RECT 90.735 194.080 90.980 194.805 ;
        RECT 91.165 194.250 91.425 194.975 ;
        RECT 91.595 194.080 91.840 194.805 ;
        RECT 92.025 194.250 92.285 194.975 ;
        RECT 92.455 194.080 92.700 194.805 ;
        RECT 92.870 194.250 93.130 194.975 ;
        RECT 93.300 194.080 93.560 194.805 ;
        RECT 93.730 194.250 93.990 194.975 ;
        RECT 94.160 194.080 94.420 194.805 ;
        RECT 94.590 194.250 94.850 194.975 ;
        RECT 95.020 194.080 95.280 194.805 ;
        RECT 95.450 194.250 95.710 194.975 ;
        RECT 95.880 194.080 96.140 194.875 ;
        RECT 96.310 194.250 96.560 195.385 ;
        RECT 89.865 194.075 96.140 194.080 ;
        RECT 96.740 194.075 97.000 194.885 ;
        RECT 97.175 194.245 97.420 195.385 ;
        RECT 97.600 194.075 97.895 194.885 ;
        RECT 98.535 194.245 98.815 195.680 ;
        RECT 99.045 195.235 99.330 195.805 ;
        RECT 99.515 195.405 99.985 195.635 ;
        RECT 100.155 195.615 100.485 195.635 ;
        RECT 100.155 195.435 100.605 195.615 ;
        RECT 100.795 195.435 101.125 195.635 ;
        RECT 99.045 195.020 100.195 195.235 ;
        RECT 98.985 194.075 99.695 194.850 ;
        RECT 99.865 194.245 100.195 195.020 ;
        RECT 100.390 194.320 100.605 195.435 ;
        RECT 100.895 195.095 101.125 195.435 ;
        RECT 101.295 195.385 101.610 195.945 ;
        RECT 101.780 195.635 102.030 196.445 ;
        RECT 102.200 196.100 102.460 196.625 ;
        RECT 102.640 195.635 102.890 196.445 ;
        RECT 103.060 196.065 103.320 196.625 ;
        RECT 103.490 195.975 103.750 196.430 ;
        RECT 103.920 196.145 104.180 196.625 ;
        RECT 104.350 195.975 104.610 196.430 ;
        RECT 104.780 196.145 105.040 196.625 ;
        RECT 105.210 195.975 105.470 196.430 ;
        RECT 105.640 196.145 105.885 196.625 ;
        RECT 106.055 195.975 106.330 196.430 ;
        RECT 106.500 196.145 106.745 196.625 ;
        RECT 106.915 195.975 107.175 196.430 ;
        RECT 107.355 196.145 107.605 196.625 ;
        RECT 107.775 195.975 108.035 196.430 ;
        RECT 108.215 196.145 108.465 196.625 ;
        RECT 108.635 195.975 108.895 196.430 ;
        RECT 109.075 196.145 109.335 196.625 ;
        RECT 109.505 195.975 109.765 196.430 ;
        RECT 109.935 196.145 110.235 196.625 ;
        RECT 110.495 196.165 111.055 196.455 ;
        RECT 111.225 196.165 111.475 196.625 ;
        RECT 103.490 195.945 110.235 195.975 ;
        RECT 103.490 195.805 110.265 195.945 ;
        RECT 109.070 195.775 110.265 195.805 ;
        RECT 101.780 195.385 108.900 195.635 ;
        RECT 100.785 194.075 101.115 194.795 ;
        RECT 101.305 194.075 101.600 194.885 ;
        RECT 101.780 194.245 102.025 195.385 ;
        RECT 102.200 194.075 102.460 194.885 ;
        RECT 102.640 194.250 102.890 195.385 ;
        RECT 109.070 195.215 110.235 195.775 ;
        RECT 103.490 194.990 110.235 195.215 ;
        RECT 103.490 194.975 108.895 194.990 ;
        RECT 103.060 194.080 103.320 194.875 ;
        RECT 103.490 194.250 103.750 194.975 ;
        RECT 103.920 194.080 104.180 194.805 ;
        RECT 104.350 194.250 104.610 194.975 ;
        RECT 104.780 194.080 105.040 194.805 ;
        RECT 105.210 194.250 105.470 194.975 ;
        RECT 105.640 194.080 105.900 194.805 ;
        RECT 106.070 194.250 106.330 194.975 ;
        RECT 106.500 194.080 106.745 194.805 ;
        RECT 106.915 194.250 107.175 194.975 ;
        RECT 107.360 194.080 107.605 194.805 ;
        RECT 107.775 194.250 108.035 194.975 ;
        RECT 108.220 194.080 108.465 194.805 ;
        RECT 108.635 194.250 108.895 194.975 ;
        RECT 109.080 194.080 109.335 194.805 ;
        RECT 109.505 194.250 109.795 194.990 ;
        RECT 103.060 194.075 109.335 194.080 ;
        RECT 109.965 194.075 110.235 194.820 ;
        RECT 110.495 194.795 110.745 196.165 ;
        RECT 112.095 195.995 112.425 196.355 ;
        RECT 111.035 195.805 112.425 195.995 ;
        RECT 112.795 195.900 113.085 196.625 ;
        RECT 114.175 195.875 115.385 196.625 ;
        RECT 111.035 195.715 111.205 195.805 ;
        RECT 110.915 195.385 111.205 195.715 ;
        RECT 111.375 195.385 111.715 195.635 ;
        RECT 111.935 195.385 112.610 195.635 ;
        RECT 111.035 195.135 111.205 195.385 ;
        RECT 111.035 194.965 111.975 195.135 ;
        RECT 112.345 195.025 112.610 195.385 ;
        RECT 110.495 194.245 110.955 194.795 ;
        RECT 111.145 194.075 111.475 194.795 ;
        RECT 111.675 194.415 111.975 194.965 ;
        RECT 112.145 194.075 112.425 194.745 ;
        RECT 112.795 194.075 113.085 195.240 ;
        RECT 114.175 195.165 114.695 195.705 ;
        RECT 114.865 195.335 115.385 195.875 ;
        RECT 114.175 194.075 115.385 195.165 ;
        RECT 61.190 193.905 115.470 194.075 ;
        RECT 61.275 192.815 62.485 193.905 ;
        RECT 62.655 193.470 68.000 193.905 ;
        RECT 61.275 192.105 61.795 192.645 ;
        RECT 61.965 192.275 62.485 192.815 ;
        RECT 61.275 191.355 62.485 192.105 ;
        RECT 64.240 191.900 64.580 192.730 ;
        RECT 66.060 192.220 66.410 193.470 ;
        RECT 68.175 192.815 71.685 193.905 ;
        RECT 68.175 192.125 69.825 192.645 ;
        RECT 69.995 192.295 71.685 192.815 ;
        RECT 72.775 192.830 73.045 193.735 ;
        RECT 73.215 193.145 73.545 193.905 ;
        RECT 73.725 192.975 73.895 193.735 ;
        RECT 62.655 191.355 68.000 191.900 ;
        RECT 68.175 191.355 71.685 192.125 ;
        RECT 72.775 192.030 72.945 192.830 ;
        RECT 73.230 192.805 73.895 192.975 ;
        RECT 73.230 192.660 73.400 192.805 ;
        RECT 74.155 192.740 74.445 193.905 ;
        RECT 74.625 192.765 74.955 193.905 ;
        RECT 75.485 192.935 75.815 193.720 ;
        RECT 76.000 193.105 76.315 193.905 ;
        RECT 76.580 193.550 77.660 193.720 ;
        RECT 76.580 192.935 76.750 193.550 ;
        RECT 75.135 192.765 75.815 192.935 ;
        RECT 73.115 192.330 73.400 192.660 ;
        RECT 73.230 192.075 73.400 192.330 ;
        RECT 73.635 192.255 73.965 192.625 ;
        RECT 74.615 192.345 74.965 192.595 ;
        RECT 75.135 192.165 75.305 192.765 ;
        RECT 75.475 192.345 75.825 192.595 ;
        RECT 72.775 191.525 73.035 192.030 ;
        RECT 73.230 191.905 73.895 192.075 ;
        RECT 73.215 191.355 73.545 191.735 ;
        RECT 73.725 191.525 73.895 191.905 ;
        RECT 74.155 191.355 74.445 192.080 ;
        RECT 74.625 191.355 74.895 192.165 ;
        RECT 75.065 191.525 75.395 192.165 ;
        RECT 75.565 191.355 75.805 192.165 ;
        RECT 75.995 191.925 76.265 192.935 ;
        RECT 76.435 192.765 76.750 192.935 ;
        RECT 76.435 192.095 76.605 192.765 ;
        RECT 76.920 192.595 77.155 193.275 ;
        RECT 77.325 192.765 77.660 193.550 ;
        RECT 77.845 193.295 78.175 193.725 ;
        RECT 78.355 193.465 78.550 193.905 ;
        RECT 78.720 193.295 79.050 193.725 ;
        RECT 77.845 193.125 79.050 193.295 ;
        RECT 77.845 192.795 78.740 193.125 ;
        RECT 79.220 192.955 79.495 193.725 ;
        RECT 78.910 192.765 79.495 192.955 ;
        RECT 79.675 192.765 80.060 193.735 ;
        RECT 80.230 193.445 80.555 193.905 ;
        RECT 81.075 193.275 81.355 193.735 ;
        RECT 80.230 193.055 81.355 193.275 ;
        RECT 76.775 192.265 77.155 192.595 ;
        RECT 77.325 192.265 77.660 192.595 ;
        RECT 77.850 192.265 78.145 192.595 ;
        RECT 78.325 192.265 78.740 192.595 ;
        RECT 76.435 191.925 77.660 192.095 ;
        RECT 76.065 191.355 76.395 191.755 ;
        RECT 76.565 191.655 76.735 191.925 ;
        RECT 76.905 191.355 77.235 191.755 ;
        RECT 77.405 191.655 77.660 191.925 ;
        RECT 77.845 191.355 78.145 192.085 ;
        RECT 78.325 191.645 78.555 192.265 ;
        RECT 78.910 192.095 79.085 192.765 ;
        RECT 78.755 191.915 79.085 192.095 ;
        RECT 79.255 191.945 79.495 192.595 ;
        RECT 79.675 192.095 79.955 192.765 ;
        RECT 80.230 192.595 80.680 193.055 ;
        RECT 81.545 192.885 81.945 193.735 ;
        RECT 82.345 193.445 82.615 193.905 ;
        RECT 82.785 193.275 83.070 193.735 ;
        RECT 83.360 193.525 83.695 193.905 ;
        RECT 80.125 192.265 80.680 192.595 ;
        RECT 80.850 192.325 81.945 192.885 ;
        RECT 80.230 192.155 80.680 192.265 ;
        RECT 78.755 191.535 78.980 191.915 ;
        RECT 79.150 191.355 79.480 191.745 ;
        RECT 79.675 191.525 80.060 192.095 ;
        RECT 80.230 191.985 81.355 192.155 ;
        RECT 80.230 191.355 80.555 191.815 ;
        RECT 81.075 191.525 81.355 191.985 ;
        RECT 81.545 191.525 81.945 192.325 ;
        RECT 82.115 193.055 83.070 193.275 ;
        RECT 82.115 192.155 82.325 193.055 ;
        RECT 82.495 192.325 83.185 192.885 ;
        RECT 82.115 191.985 83.070 192.155 ;
        RECT 83.355 192.035 83.595 193.345 ;
        RECT 83.865 192.935 84.115 193.735 ;
        RECT 84.335 193.185 84.665 193.905 ;
        RECT 84.850 192.935 85.100 193.735 ;
        RECT 85.565 193.105 85.895 193.905 ;
        RECT 86.065 193.475 86.405 193.735 ;
        RECT 86.580 193.480 86.915 193.905 ;
        RECT 83.765 192.765 85.955 192.935 ;
        RECT 82.345 191.355 82.615 191.815 ;
        RECT 82.785 191.525 83.070 191.985 ;
        RECT 83.765 191.855 83.935 192.765 ;
        RECT 85.640 192.595 85.955 192.765 ;
        RECT 83.440 191.525 83.935 191.855 ;
        RECT 84.155 191.630 84.505 192.595 ;
        RECT 84.685 191.625 84.985 192.595 ;
        RECT 85.165 191.625 85.445 192.595 ;
        RECT 85.640 192.345 85.970 192.595 ;
        RECT 85.625 191.355 85.895 192.155 ;
        RECT 86.145 192.075 86.405 193.475 ;
        RECT 87.085 193.300 87.270 193.705 ;
        RECT 86.065 191.565 86.405 192.075 ;
        RECT 86.605 193.125 87.270 193.300 ;
        RECT 87.475 193.125 87.805 193.905 ;
        RECT 86.605 192.095 86.945 193.125 ;
        RECT 87.975 192.935 88.245 193.705 ;
        RECT 87.115 192.765 88.245 192.935 ;
        RECT 87.115 192.265 87.365 192.765 ;
        RECT 86.605 191.925 87.290 192.095 ;
        RECT 87.545 192.015 87.905 192.595 ;
        RECT 86.580 191.355 86.915 191.755 ;
        RECT 87.085 191.525 87.290 191.925 ;
        RECT 88.075 191.855 88.245 192.765 ;
        RECT 87.500 191.355 87.775 191.835 ;
        RECT 87.985 191.525 88.245 191.855 ;
        RECT 88.415 192.300 88.695 193.735 ;
        RECT 88.865 193.130 89.575 193.905 ;
        RECT 89.745 192.960 90.075 193.735 ;
        RECT 88.925 192.745 90.075 192.960 ;
        RECT 88.415 191.525 88.755 192.300 ;
        RECT 88.925 192.175 89.210 192.745 ;
        RECT 89.395 192.345 89.865 192.575 ;
        RECT 90.270 192.545 90.485 193.660 ;
        RECT 90.665 193.185 90.995 193.905 ;
        RECT 90.775 192.545 91.005 192.885 ;
        RECT 90.035 192.365 90.485 192.545 ;
        RECT 90.035 192.345 90.365 192.365 ;
        RECT 90.675 192.345 91.005 192.545 ;
        RECT 91.175 192.715 91.635 193.725 ;
        RECT 92.705 193.395 93.035 193.905 ;
        RECT 94.135 193.235 94.415 193.905 ;
        RECT 91.805 193.055 93.765 193.225 ;
        RECT 91.175 192.205 91.345 192.715 ;
        RECT 91.805 192.515 91.975 193.055 ;
        RECT 91.515 192.345 91.975 192.515 ;
        RECT 92.155 192.265 92.395 192.885 ;
        RECT 92.565 192.265 92.905 192.885 ;
        RECT 93.075 192.265 93.425 192.885 ;
        RECT 88.925 191.985 89.635 192.175 ;
        RECT 89.335 191.845 89.635 191.985 ;
        RECT 89.825 191.985 91.005 192.175 ;
        RECT 89.825 191.905 90.155 191.985 ;
        RECT 89.335 191.835 89.650 191.845 ;
        RECT 89.335 191.825 89.660 191.835 ;
        RECT 89.335 191.820 89.670 191.825 ;
        RECT 88.925 191.355 89.095 191.815 ;
        RECT 89.335 191.810 89.675 191.820 ;
        RECT 89.335 191.805 89.680 191.810 ;
        RECT 89.335 191.795 89.685 191.805 ;
        RECT 89.335 191.790 89.690 191.795 ;
        RECT 89.335 191.525 89.695 191.790 ;
        RECT 90.325 191.355 90.495 191.815 ;
        RECT 90.665 191.525 91.005 191.985 ;
        RECT 91.175 192.095 91.405 192.205 ;
        RECT 93.595 192.095 93.765 193.055 ;
        RECT 94.585 193.015 94.885 193.565 ;
        RECT 95.085 193.185 95.415 193.905 ;
        RECT 95.605 193.185 96.065 193.735 ;
        RECT 93.950 192.595 94.215 192.955 ;
        RECT 94.585 192.845 95.525 193.015 ;
        RECT 95.355 192.595 95.525 192.845 ;
        RECT 93.950 192.345 94.625 192.595 ;
        RECT 94.845 192.345 95.185 192.595 ;
        RECT 95.355 192.265 95.645 192.595 ;
        RECT 95.355 192.175 95.525 192.265 ;
        RECT 91.175 191.925 92.535 192.095 ;
        RECT 91.175 191.525 91.695 191.925 ;
        RECT 91.865 191.355 92.195 191.755 ;
        RECT 92.365 191.580 92.535 191.925 ;
        RECT 92.705 191.355 93.035 192.095 ;
        RECT 93.270 191.925 93.765 192.095 ;
        RECT 94.135 191.985 95.525 192.175 ;
        RECT 93.270 191.675 93.440 191.925 ;
        RECT 94.135 191.625 94.465 191.985 ;
        RECT 95.815 191.815 96.065 193.185 ;
        RECT 95.085 191.355 95.335 191.815 ;
        RECT 95.505 191.525 96.065 191.815 ;
        RECT 97.155 192.300 97.435 193.735 ;
        RECT 97.605 193.130 98.315 193.905 ;
        RECT 98.485 192.960 98.815 193.735 ;
        RECT 97.665 192.745 98.815 192.960 ;
        RECT 97.155 191.525 97.495 192.300 ;
        RECT 97.665 192.175 97.950 192.745 ;
        RECT 98.135 192.345 98.605 192.575 ;
        RECT 99.010 192.545 99.225 193.660 ;
        RECT 99.405 193.185 99.735 193.905 ;
        RECT 99.515 192.545 99.745 192.885 ;
        RECT 99.915 192.740 100.205 193.905 ;
        RECT 98.775 192.365 99.225 192.545 ;
        RECT 98.775 192.345 99.105 192.365 ;
        RECT 99.415 192.345 99.745 192.545 ;
        RECT 100.375 192.300 100.655 193.735 ;
        RECT 100.825 193.130 101.535 193.905 ;
        RECT 101.705 192.960 102.035 193.735 ;
        RECT 100.885 192.745 102.035 192.960 ;
        RECT 97.665 191.985 98.375 192.175 ;
        RECT 98.075 191.845 98.375 191.985 ;
        RECT 98.565 191.985 99.745 192.175 ;
        RECT 98.565 191.905 98.895 191.985 ;
        RECT 98.075 191.835 98.390 191.845 ;
        RECT 98.075 191.825 98.400 191.835 ;
        RECT 98.075 191.820 98.410 191.825 ;
        RECT 97.665 191.355 97.835 191.815 ;
        RECT 98.075 191.810 98.415 191.820 ;
        RECT 98.075 191.805 98.420 191.810 ;
        RECT 98.075 191.795 98.425 191.805 ;
        RECT 98.075 191.790 98.430 191.795 ;
        RECT 98.075 191.525 98.435 191.790 ;
        RECT 99.065 191.355 99.235 191.815 ;
        RECT 99.405 191.525 99.745 191.985 ;
        RECT 99.915 191.355 100.205 192.080 ;
        RECT 100.375 191.525 100.715 192.300 ;
        RECT 100.885 192.175 101.170 192.745 ;
        RECT 101.355 192.345 101.825 192.575 ;
        RECT 102.230 192.545 102.445 193.660 ;
        RECT 102.625 193.185 102.955 193.905 ;
        RECT 103.225 193.235 103.395 193.735 ;
        RECT 103.565 193.405 103.895 193.905 ;
        RECT 103.225 193.065 103.890 193.235 ;
        RECT 102.735 192.545 102.965 192.885 ;
        RECT 101.995 192.365 102.445 192.545 ;
        RECT 101.995 192.345 102.325 192.365 ;
        RECT 102.635 192.345 102.965 192.545 ;
        RECT 103.140 192.245 103.490 192.895 ;
        RECT 100.885 191.985 101.595 192.175 ;
        RECT 101.295 191.845 101.595 191.985 ;
        RECT 101.785 191.985 102.965 192.175 ;
        RECT 103.660 192.075 103.890 193.065 ;
        RECT 101.785 191.905 102.115 191.985 ;
        RECT 101.295 191.835 101.610 191.845 ;
        RECT 101.295 191.825 101.620 191.835 ;
        RECT 101.295 191.820 101.630 191.825 ;
        RECT 100.885 191.355 101.055 191.815 ;
        RECT 101.295 191.810 101.635 191.820 ;
        RECT 101.295 191.805 101.640 191.810 ;
        RECT 101.295 191.795 101.645 191.805 ;
        RECT 101.295 191.790 101.650 191.795 ;
        RECT 101.295 191.525 101.655 191.790 ;
        RECT 102.285 191.355 102.455 191.815 ;
        RECT 102.625 191.525 102.965 191.985 ;
        RECT 103.225 191.905 103.890 192.075 ;
        RECT 103.225 191.615 103.395 191.905 ;
        RECT 103.565 191.355 103.895 191.735 ;
        RECT 104.065 191.615 104.250 193.735 ;
        RECT 104.490 193.445 104.755 193.905 ;
        RECT 104.925 193.310 105.175 193.735 ;
        RECT 105.385 193.460 106.490 193.630 ;
        RECT 104.870 193.180 105.175 193.310 ;
        RECT 104.420 191.985 104.700 192.935 ;
        RECT 104.870 192.075 105.040 193.180 ;
        RECT 105.210 192.395 105.450 192.990 ;
        RECT 105.620 192.925 106.150 193.290 ;
        RECT 105.620 192.225 105.790 192.925 ;
        RECT 106.320 192.845 106.490 193.460 ;
        RECT 106.660 193.105 106.830 193.905 ;
        RECT 107.000 193.405 107.250 193.735 ;
        RECT 107.475 193.435 108.360 193.605 ;
        RECT 106.320 192.755 106.830 192.845 ;
        RECT 104.870 191.945 105.095 192.075 ;
        RECT 105.265 192.005 105.790 192.225 ;
        RECT 105.960 192.585 106.830 192.755 ;
        RECT 104.505 191.355 104.755 191.815 ;
        RECT 104.925 191.805 105.095 191.945 ;
        RECT 105.960 191.805 106.130 192.585 ;
        RECT 106.660 192.515 106.830 192.585 ;
        RECT 106.340 192.335 106.540 192.365 ;
        RECT 107.000 192.335 107.170 193.405 ;
        RECT 107.340 192.515 107.530 193.235 ;
        RECT 106.340 192.035 107.170 192.335 ;
        RECT 107.700 192.305 108.020 193.265 ;
        RECT 104.925 191.635 105.260 191.805 ;
        RECT 105.455 191.635 106.130 191.805 ;
        RECT 106.450 191.355 106.820 191.855 ;
        RECT 107.000 191.805 107.170 192.035 ;
        RECT 107.555 191.975 108.020 192.305 ;
        RECT 108.190 192.595 108.360 193.435 ;
        RECT 108.540 193.405 108.855 193.905 ;
        RECT 109.085 193.175 109.425 193.735 ;
        RECT 108.530 192.800 109.425 193.175 ;
        RECT 109.595 192.895 109.765 193.905 ;
        RECT 109.235 192.595 109.425 192.800 ;
        RECT 109.935 192.845 110.265 193.690 ;
        RECT 109.935 192.765 110.325 192.845 ;
        RECT 110.110 192.715 110.325 192.765 ;
        RECT 108.190 192.265 109.065 192.595 ;
        RECT 109.235 192.265 109.985 192.595 ;
        RECT 108.190 191.805 108.360 192.265 ;
        RECT 109.235 192.095 109.435 192.265 ;
        RECT 110.155 192.135 110.325 192.715 ;
        RECT 110.100 192.095 110.325 192.135 ;
        RECT 107.000 191.635 107.405 191.805 ;
        RECT 107.575 191.635 108.360 191.805 ;
        RECT 108.635 191.355 108.845 191.885 ;
        RECT 109.105 191.570 109.435 192.095 ;
        RECT 109.945 192.010 110.325 192.095 ;
        RECT 110.495 192.765 110.880 193.735 ;
        RECT 111.050 193.445 111.375 193.905 ;
        RECT 111.895 193.275 112.175 193.735 ;
        RECT 111.050 193.055 112.175 193.275 ;
        RECT 110.495 192.095 110.775 192.765 ;
        RECT 111.050 192.595 111.500 193.055 ;
        RECT 112.365 192.885 112.765 193.735 ;
        RECT 113.165 193.445 113.435 193.905 ;
        RECT 113.605 193.275 113.890 193.735 ;
        RECT 110.945 192.265 111.500 192.595 ;
        RECT 111.670 192.325 112.765 192.885 ;
        RECT 111.050 192.155 111.500 192.265 ;
        RECT 109.605 191.355 109.775 191.965 ;
        RECT 109.945 191.575 110.275 192.010 ;
        RECT 110.495 191.525 110.880 192.095 ;
        RECT 111.050 191.985 112.175 192.155 ;
        RECT 111.050 191.355 111.375 191.815 ;
        RECT 111.895 191.525 112.175 191.985 ;
        RECT 112.365 191.525 112.765 192.325 ;
        RECT 112.935 193.055 113.890 193.275 ;
        RECT 112.935 192.155 113.145 193.055 ;
        RECT 113.315 192.325 114.005 192.885 ;
        RECT 114.175 192.815 115.385 193.905 ;
        RECT 114.175 192.275 114.695 192.815 ;
        RECT 112.935 191.985 113.890 192.155 ;
        RECT 114.865 192.105 115.385 192.645 ;
        RECT 113.165 191.355 113.435 191.815 ;
        RECT 113.605 191.525 113.890 191.985 ;
        RECT 114.175 191.355 115.385 192.105 ;
        RECT 61.190 191.185 115.470 191.355 ;
        RECT 61.275 190.435 62.485 191.185 ;
        RECT 62.655 190.640 68.000 191.185 ;
        RECT 61.275 189.895 61.795 190.435 ;
        RECT 61.965 189.725 62.485 190.265 ;
        RECT 64.240 189.810 64.580 190.640 ;
        RECT 68.175 190.415 70.765 191.185 ;
        RECT 61.275 188.635 62.485 189.725 ;
        RECT 66.060 189.070 66.410 190.320 ;
        RECT 68.175 189.895 69.385 190.415 ;
        RECT 69.555 189.725 70.765 190.245 ;
        RECT 62.655 188.635 68.000 189.070 ;
        RECT 68.175 188.635 70.765 189.725 ;
        RECT 71.395 190.240 71.735 191.015 ;
        RECT 71.905 190.725 72.075 191.185 ;
        RECT 72.315 190.750 72.675 191.015 ;
        RECT 72.315 190.745 72.670 190.750 ;
        RECT 72.315 190.735 72.665 190.745 ;
        RECT 72.315 190.730 72.660 190.735 ;
        RECT 72.315 190.720 72.655 190.730 ;
        RECT 73.305 190.725 73.475 191.185 ;
        RECT 72.315 190.715 72.650 190.720 ;
        RECT 72.315 190.705 72.640 190.715 ;
        RECT 72.315 190.695 72.630 190.705 ;
        RECT 72.315 190.555 72.615 190.695 ;
        RECT 71.905 190.365 72.615 190.555 ;
        RECT 72.805 190.555 73.135 190.635 ;
        RECT 73.645 190.555 73.985 191.015 ;
        RECT 72.805 190.365 73.985 190.555 ;
        RECT 74.245 190.635 74.415 190.925 ;
        RECT 74.585 190.805 74.915 191.185 ;
        RECT 74.245 190.465 74.910 190.635 ;
        RECT 71.395 188.805 71.675 190.240 ;
        RECT 71.905 189.795 72.190 190.365 ;
        RECT 72.375 189.965 72.845 190.195 ;
        RECT 73.015 190.175 73.345 190.195 ;
        RECT 73.015 189.995 73.465 190.175 ;
        RECT 73.655 189.995 73.985 190.195 ;
        RECT 71.905 189.580 73.055 189.795 ;
        RECT 71.845 188.635 72.555 189.410 ;
        RECT 72.725 188.805 73.055 189.580 ;
        RECT 73.250 188.880 73.465 189.995 ;
        RECT 73.755 189.655 73.985 189.995 ;
        RECT 74.160 189.645 74.510 190.295 ;
        RECT 74.680 189.475 74.910 190.465 ;
        RECT 73.645 188.635 73.975 189.355 ;
        RECT 74.245 189.305 74.910 189.475 ;
        RECT 74.245 188.805 74.415 189.305 ;
        RECT 74.585 188.635 74.915 189.135 ;
        RECT 75.085 188.805 75.270 190.925 ;
        RECT 75.525 190.725 75.775 191.185 ;
        RECT 75.945 190.735 76.280 190.905 ;
        RECT 76.475 190.735 77.150 190.905 ;
        RECT 75.945 190.595 76.115 190.735 ;
        RECT 75.440 189.605 75.720 190.555 ;
        RECT 75.890 190.465 76.115 190.595 ;
        RECT 75.890 189.360 76.060 190.465 ;
        RECT 76.285 190.315 76.810 190.535 ;
        RECT 76.230 189.550 76.470 190.145 ;
        RECT 76.640 189.615 76.810 190.315 ;
        RECT 76.980 189.955 77.150 190.735 ;
        RECT 77.470 190.685 77.840 191.185 ;
        RECT 78.020 190.735 78.425 190.905 ;
        RECT 78.595 190.735 79.380 190.905 ;
        RECT 78.020 190.505 78.190 190.735 ;
        RECT 77.360 190.205 78.190 190.505 ;
        RECT 78.575 190.235 79.040 190.565 ;
        RECT 77.360 190.175 77.560 190.205 ;
        RECT 77.680 189.955 77.850 190.025 ;
        RECT 76.980 189.785 77.850 189.955 ;
        RECT 77.340 189.695 77.850 189.785 ;
        RECT 75.890 189.230 76.195 189.360 ;
        RECT 76.640 189.250 77.170 189.615 ;
        RECT 75.510 188.635 75.775 189.095 ;
        RECT 75.945 188.805 76.195 189.230 ;
        RECT 77.340 189.080 77.510 189.695 ;
        RECT 76.405 188.910 77.510 189.080 ;
        RECT 77.680 188.635 77.850 189.435 ;
        RECT 78.020 189.135 78.190 190.205 ;
        RECT 78.360 189.305 78.550 190.025 ;
        RECT 78.720 189.275 79.040 190.235 ;
        RECT 79.210 190.275 79.380 190.735 ;
        RECT 79.655 190.655 79.865 191.185 ;
        RECT 80.125 190.445 80.455 190.970 ;
        RECT 80.625 190.575 80.795 191.185 ;
        RECT 80.965 190.530 81.295 190.965 ;
        RECT 80.965 190.445 81.345 190.530 ;
        RECT 80.255 190.275 80.455 190.445 ;
        RECT 81.120 190.405 81.345 190.445 ;
        RECT 79.210 189.945 80.085 190.275 ;
        RECT 80.255 189.945 81.005 190.275 ;
        RECT 78.020 188.805 78.270 189.135 ;
        RECT 79.210 189.105 79.380 189.945 ;
        RECT 80.255 189.740 80.445 189.945 ;
        RECT 81.175 189.825 81.345 190.405 ;
        RECT 81.130 189.775 81.345 189.825 ;
        RECT 79.550 189.365 80.445 189.740 ;
        RECT 80.955 189.695 81.345 189.775 ;
        RECT 82.435 190.445 82.820 191.015 ;
        RECT 82.990 190.725 83.315 191.185 ;
        RECT 83.835 190.555 84.115 191.015 ;
        RECT 82.435 189.775 82.715 190.445 ;
        RECT 82.990 190.385 84.115 190.555 ;
        RECT 82.990 190.275 83.440 190.385 ;
        RECT 82.885 189.945 83.440 190.275 ;
        RECT 84.305 190.215 84.705 191.015 ;
        RECT 85.105 190.725 85.375 191.185 ;
        RECT 85.545 190.555 85.830 191.015 ;
        RECT 78.495 188.935 79.380 189.105 ;
        RECT 79.560 188.635 79.875 189.135 ;
        RECT 80.105 188.805 80.445 189.365 ;
        RECT 80.615 188.635 80.785 189.645 ;
        RECT 80.955 188.850 81.285 189.695 ;
        RECT 82.435 188.805 82.820 189.775 ;
        RECT 82.990 189.485 83.440 189.945 ;
        RECT 83.610 189.655 84.705 190.215 ;
        RECT 82.990 189.265 84.115 189.485 ;
        RECT 82.990 188.635 83.315 189.095 ;
        RECT 83.835 188.805 84.115 189.265 ;
        RECT 84.305 188.805 84.705 189.655 ;
        RECT 84.875 190.385 85.830 190.555 ;
        RECT 87.035 190.460 87.325 191.185 ;
        RECT 87.495 190.445 87.880 191.015 ;
        RECT 88.050 190.725 88.375 191.185 ;
        RECT 88.895 190.555 89.175 191.015 ;
        RECT 84.875 189.485 85.085 190.385 ;
        RECT 85.255 189.655 85.945 190.215 ;
        RECT 84.875 189.265 85.830 189.485 ;
        RECT 85.105 188.635 85.375 189.095 ;
        RECT 85.545 188.805 85.830 189.265 ;
        RECT 87.035 188.635 87.325 189.800 ;
        RECT 87.495 189.775 87.775 190.445 ;
        RECT 88.050 190.385 89.175 190.555 ;
        RECT 88.050 190.275 88.500 190.385 ;
        RECT 87.945 189.945 88.500 190.275 ;
        RECT 89.365 190.215 89.765 191.015 ;
        RECT 90.165 190.725 90.435 191.185 ;
        RECT 90.605 190.555 90.890 191.015 ;
        RECT 87.495 188.805 87.880 189.775 ;
        RECT 88.050 189.485 88.500 189.945 ;
        RECT 88.670 189.655 89.765 190.215 ;
        RECT 88.050 189.265 89.175 189.485 ;
        RECT 88.050 188.635 88.375 189.095 ;
        RECT 88.895 188.805 89.175 189.265 ;
        RECT 89.365 188.805 89.765 189.655 ;
        RECT 89.935 190.385 90.890 190.555 ;
        RECT 92.095 190.445 92.480 191.015 ;
        RECT 92.650 190.725 92.975 191.185 ;
        RECT 93.495 190.555 93.775 191.015 ;
        RECT 89.935 189.485 90.145 190.385 ;
        RECT 90.315 189.655 91.005 190.215 ;
        RECT 92.095 189.775 92.375 190.445 ;
        RECT 92.650 190.385 93.775 190.555 ;
        RECT 92.650 190.275 93.100 190.385 ;
        RECT 92.545 189.945 93.100 190.275 ;
        RECT 93.965 190.215 94.365 191.015 ;
        RECT 94.765 190.725 95.035 191.185 ;
        RECT 95.205 190.555 95.490 191.015 ;
        RECT 89.935 189.265 90.890 189.485 ;
        RECT 90.165 188.635 90.435 189.095 ;
        RECT 90.605 188.805 90.890 189.265 ;
        RECT 92.095 188.805 92.480 189.775 ;
        RECT 92.650 189.485 93.100 189.945 ;
        RECT 93.270 189.655 94.365 190.215 ;
        RECT 92.650 189.265 93.775 189.485 ;
        RECT 92.650 188.635 92.975 189.095 ;
        RECT 93.495 188.805 93.775 189.265 ;
        RECT 93.965 188.805 94.365 189.655 ;
        RECT 94.535 190.385 95.490 190.555 ;
        RECT 95.785 190.460 96.115 190.970 ;
        RECT 96.285 190.785 96.615 191.185 ;
        RECT 97.665 190.615 97.995 190.955 ;
        RECT 98.165 190.785 98.495 191.185 ;
        RECT 99.080 190.685 99.575 191.015 ;
        RECT 94.535 189.485 94.745 190.385 ;
        RECT 94.915 189.655 95.605 190.215 ;
        RECT 95.785 189.695 95.975 190.460 ;
        RECT 96.285 190.445 98.650 190.615 ;
        RECT 96.285 190.275 96.455 190.445 ;
        RECT 96.145 189.945 96.455 190.275 ;
        RECT 96.625 189.945 96.930 190.275 ;
        RECT 94.535 189.265 95.490 189.485 ;
        RECT 94.765 188.635 95.035 189.095 ;
        RECT 95.205 188.805 95.490 189.265 ;
        RECT 95.785 188.845 96.115 189.695 ;
        RECT 96.285 188.635 96.535 189.775 ;
        RECT 96.715 189.615 96.930 189.945 ;
        RECT 97.105 189.615 97.390 190.275 ;
        RECT 97.585 189.615 97.850 190.275 ;
        RECT 98.065 189.615 98.310 190.275 ;
        RECT 98.480 189.445 98.650 190.445 ;
        RECT 96.725 189.275 98.015 189.445 ;
        RECT 96.725 188.855 96.975 189.275 ;
        RECT 97.205 188.635 97.535 189.105 ;
        RECT 97.765 188.855 98.015 189.275 ;
        RECT 98.195 189.275 98.650 189.445 ;
        RECT 98.195 188.845 98.525 189.275 ;
        RECT 98.995 189.195 99.235 190.505 ;
        RECT 99.405 189.775 99.575 190.685 ;
        RECT 99.795 189.945 100.145 190.910 ;
        RECT 100.325 189.945 100.625 190.915 ;
        RECT 100.805 189.945 101.085 190.915 ;
        RECT 101.265 190.385 101.535 191.185 ;
        RECT 101.705 190.465 102.045 190.975 ;
        RECT 101.280 189.945 101.610 190.195 ;
        RECT 101.280 189.775 101.595 189.945 ;
        RECT 99.405 189.605 101.595 189.775 ;
        RECT 99.000 188.635 99.335 189.015 ;
        RECT 99.505 188.805 99.755 189.605 ;
        RECT 99.975 188.635 100.305 189.355 ;
        RECT 100.490 188.805 100.740 189.605 ;
        RECT 101.205 188.635 101.535 189.435 ;
        RECT 101.785 189.065 102.045 190.465 ;
        RECT 101.705 188.805 102.045 189.065 ;
        RECT 103.135 190.445 103.520 191.015 ;
        RECT 103.690 190.725 104.015 191.185 ;
        RECT 104.535 190.555 104.815 191.015 ;
        RECT 103.135 189.775 103.415 190.445 ;
        RECT 103.690 190.385 104.815 190.555 ;
        RECT 103.690 190.275 104.140 190.385 ;
        RECT 103.585 189.945 104.140 190.275 ;
        RECT 105.005 190.215 105.405 191.015 ;
        RECT 105.805 190.725 106.075 191.185 ;
        RECT 106.245 190.555 106.530 191.015 ;
        RECT 103.135 188.805 103.520 189.775 ;
        RECT 103.690 189.485 104.140 189.945 ;
        RECT 104.310 189.655 105.405 190.215 ;
        RECT 103.690 189.265 104.815 189.485 ;
        RECT 103.690 188.635 104.015 189.095 ;
        RECT 104.535 188.805 104.815 189.265 ;
        RECT 105.005 188.805 105.405 189.655 ;
        RECT 105.575 190.385 106.530 190.555 ;
        RECT 105.575 189.485 105.785 190.385 ;
        RECT 106.815 190.240 107.155 191.015 ;
        RECT 107.325 190.725 107.495 191.185 ;
        RECT 107.735 190.750 108.095 191.015 ;
        RECT 107.735 190.745 108.090 190.750 ;
        RECT 107.735 190.735 108.085 190.745 ;
        RECT 107.735 190.730 108.080 190.735 ;
        RECT 107.735 190.720 108.075 190.730 ;
        RECT 108.725 190.725 108.895 191.185 ;
        RECT 107.735 190.715 108.070 190.720 ;
        RECT 107.735 190.705 108.060 190.715 ;
        RECT 107.735 190.695 108.050 190.705 ;
        RECT 107.735 190.555 108.035 190.695 ;
        RECT 107.325 190.365 108.035 190.555 ;
        RECT 108.225 190.555 108.555 190.635 ;
        RECT 109.065 190.555 109.405 191.015 ;
        RECT 108.225 190.365 109.405 190.555 ;
        RECT 109.575 190.465 109.915 190.975 ;
        RECT 105.955 189.655 106.645 190.215 ;
        RECT 105.575 189.265 106.530 189.485 ;
        RECT 105.805 188.635 106.075 189.095 ;
        RECT 106.245 188.805 106.530 189.265 ;
        RECT 106.815 188.805 107.095 190.240 ;
        RECT 107.325 189.795 107.610 190.365 ;
        RECT 107.795 189.965 108.265 190.195 ;
        RECT 108.435 190.175 108.765 190.195 ;
        RECT 108.435 189.995 108.885 190.175 ;
        RECT 109.075 189.995 109.405 190.195 ;
        RECT 107.325 189.580 108.475 189.795 ;
        RECT 107.265 188.635 107.975 189.410 ;
        RECT 108.145 188.805 108.475 189.580 ;
        RECT 108.670 188.880 108.885 189.995 ;
        RECT 109.175 189.655 109.405 189.995 ;
        RECT 109.065 188.635 109.395 189.355 ;
        RECT 109.575 189.065 109.835 190.465 ;
        RECT 110.085 190.385 110.355 191.185 ;
        RECT 110.010 189.945 110.340 190.195 ;
        RECT 110.535 189.945 110.815 190.915 ;
        RECT 110.995 189.945 111.295 190.915 ;
        RECT 111.475 189.945 111.825 190.910 ;
        RECT 112.045 190.685 112.540 191.015 ;
        RECT 110.025 189.775 110.340 189.945 ;
        RECT 112.045 189.775 112.215 190.685 ;
        RECT 110.025 189.605 112.215 189.775 ;
        RECT 109.575 188.805 109.915 189.065 ;
        RECT 110.085 188.635 110.415 189.435 ;
        RECT 110.880 188.805 111.130 189.605 ;
        RECT 111.315 188.635 111.645 189.355 ;
        RECT 111.865 188.805 112.115 189.605 ;
        RECT 112.385 189.195 112.625 190.505 ;
        RECT 112.795 190.460 113.085 191.185 ;
        RECT 114.175 190.435 115.385 191.185 ;
        RECT 112.285 188.635 112.620 189.015 ;
        RECT 112.795 188.635 113.085 189.800 ;
        RECT 114.175 189.725 114.695 190.265 ;
        RECT 114.865 189.895 115.385 190.435 ;
        RECT 114.175 188.635 115.385 189.725 ;
        RECT 61.190 188.465 115.470 188.635 ;
        RECT 61.275 187.375 62.485 188.465 ;
        RECT 62.655 187.375 66.165 188.465 ;
        RECT 66.910 187.835 67.195 188.295 ;
        RECT 67.365 188.005 67.635 188.465 ;
        RECT 66.910 187.615 67.865 187.835 ;
        RECT 61.275 186.665 61.795 187.205 ;
        RECT 61.965 186.835 62.485 187.375 ;
        RECT 62.655 186.685 64.305 187.205 ;
        RECT 64.475 186.855 66.165 187.375 ;
        RECT 66.795 186.885 67.485 187.445 ;
        RECT 67.655 186.715 67.865 187.615 ;
        RECT 61.275 185.915 62.485 186.665 ;
        RECT 62.655 185.915 66.165 186.685 ;
        RECT 66.910 186.545 67.865 186.715 ;
        RECT 68.035 187.445 68.435 188.295 ;
        RECT 68.625 187.835 68.905 188.295 ;
        RECT 69.425 188.005 69.750 188.465 ;
        RECT 68.625 187.615 69.750 187.835 ;
        RECT 68.035 186.885 69.130 187.445 ;
        RECT 69.300 187.155 69.750 187.615 ;
        RECT 69.920 187.325 70.305 188.295 ;
        RECT 66.910 186.085 67.195 186.545 ;
        RECT 67.365 185.915 67.635 186.375 ;
        RECT 68.035 186.085 68.435 186.885 ;
        RECT 69.300 186.825 69.855 187.155 ;
        RECT 69.300 186.715 69.750 186.825 ;
        RECT 68.625 186.545 69.750 186.715 ;
        RECT 70.025 186.655 70.305 187.325 ;
        RECT 68.625 186.085 68.905 186.545 ;
        RECT 69.425 185.915 69.750 186.375 ;
        RECT 69.920 186.085 70.305 186.655 ;
        RECT 70.475 187.325 70.860 188.295 ;
        RECT 71.030 188.005 71.355 188.465 ;
        RECT 71.875 187.835 72.155 188.295 ;
        RECT 71.030 187.615 72.155 187.835 ;
        RECT 70.475 186.655 70.755 187.325 ;
        RECT 71.030 187.155 71.480 187.615 ;
        RECT 72.345 187.445 72.745 188.295 ;
        RECT 73.145 188.005 73.415 188.465 ;
        RECT 73.585 187.835 73.870 188.295 ;
        RECT 70.925 186.825 71.480 187.155 ;
        RECT 71.650 186.885 72.745 187.445 ;
        RECT 71.030 186.715 71.480 186.825 ;
        RECT 70.475 186.085 70.860 186.655 ;
        RECT 71.030 186.545 72.155 186.715 ;
        RECT 71.030 185.915 71.355 186.375 ;
        RECT 71.875 186.085 72.155 186.545 ;
        RECT 72.345 186.085 72.745 186.885 ;
        RECT 72.915 187.615 73.870 187.835 ;
        RECT 72.915 186.715 73.125 187.615 ;
        RECT 73.295 186.885 73.985 187.445 ;
        RECT 74.155 187.300 74.445 188.465 ;
        RECT 74.615 187.910 75.220 188.465 ;
        RECT 75.395 187.955 75.875 188.295 ;
        RECT 76.045 187.920 76.300 188.465 ;
        RECT 74.615 187.810 75.230 187.910 ;
        RECT 75.045 187.785 75.230 187.810 ;
        RECT 74.615 187.190 74.875 187.640 ;
        RECT 75.045 187.540 75.375 187.785 ;
        RECT 75.545 187.465 76.300 187.715 ;
        RECT 76.470 187.595 76.745 188.295 ;
        RECT 77.005 187.795 77.175 188.295 ;
        RECT 77.345 187.965 77.675 188.465 ;
        RECT 77.005 187.625 77.670 187.795 ;
        RECT 75.530 187.430 76.300 187.465 ;
        RECT 75.515 187.420 76.300 187.430 ;
        RECT 75.510 187.405 76.405 187.420 ;
        RECT 75.490 187.390 76.405 187.405 ;
        RECT 75.470 187.380 76.405 187.390 ;
        RECT 75.445 187.370 76.405 187.380 ;
        RECT 75.375 187.340 76.405 187.370 ;
        RECT 75.355 187.310 76.405 187.340 ;
        RECT 75.335 187.280 76.405 187.310 ;
        RECT 75.305 187.255 76.405 187.280 ;
        RECT 75.270 187.220 76.405 187.255 ;
        RECT 75.240 187.215 76.405 187.220 ;
        RECT 75.240 187.210 75.630 187.215 ;
        RECT 75.240 187.200 75.605 187.210 ;
        RECT 75.240 187.195 75.590 187.200 ;
        RECT 75.240 187.190 75.575 187.195 ;
        RECT 74.615 187.185 75.575 187.190 ;
        RECT 74.615 187.175 75.565 187.185 ;
        RECT 74.615 187.170 75.555 187.175 ;
        RECT 74.615 187.160 75.545 187.170 ;
        RECT 74.615 187.150 75.540 187.160 ;
        RECT 74.615 187.145 75.535 187.150 ;
        RECT 74.615 187.130 75.525 187.145 ;
        RECT 74.615 187.115 75.520 187.130 ;
        RECT 74.615 187.090 75.510 187.115 ;
        RECT 74.615 187.020 75.505 187.090 ;
        RECT 72.915 186.545 73.870 186.715 ;
        RECT 73.145 185.915 73.415 186.375 ;
        RECT 73.585 186.085 73.870 186.545 ;
        RECT 74.155 185.915 74.445 186.640 ;
        RECT 74.615 186.465 75.165 186.850 ;
        RECT 75.335 186.295 75.505 187.020 ;
        RECT 74.615 186.125 75.505 186.295 ;
        RECT 75.675 186.620 76.005 187.045 ;
        RECT 76.175 186.820 76.405 187.215 ;
        RECT 75.675 186.595 75.925 186.620 ;
        RECT 75.675 186.135 75.895 186.595 ;
        RECT 76.575 186.565 76.745 187.595 ;
        RECT 76.920 186.805 77.270 187.455 ;
        RECT 77.440 186.635 77.670 187.625 ;
        RECT 76.065 185.915 76.315 186.455 ;
        RECT 76.485 186.085 76.745 186.565 ;
        RECT 77.005 186.465 77.670 186.635 ;
        RECT 77.005 186.175 77.175 186.465 ;
        RECT 77.345 185.915 77.675 186.295 ;
        RECT 77.845 186.175 78.030 188.295 ;
        RECT 78.270 188.005 78.535 188.465 ;
        RECT 78.705 187.870 78.955 188.295 ;
        RECT 79.165 188.020 80.270 188.190 ;
        RECT 78.650 187.740 78.955 187.870 ;
        RECT 78.200 186.545 78.480 187.495 ;
        RECT 78.650 186.635 78.820 187.740 ;
        RECT 78.990 186.955 79.230 187.550 ;
        RECT 79.400 187.485 79.930 187.850 ;
        RECT 79.400 186.785 79.570 187.485 ;
        RECT 80.100 187.405 80.270 188.020 ;
        RECT 80.440 187.665 80.610 188.465 ;
        RECT 80.780 187.965 81.030 188.295 ;
        RECT 81.255 187.995 82.140 188.165 ;
        RECT 80.100 187.315 80.610 187.405 ;
        RECT 78.650 186.505 78.875 186.635 ;
        RECT 79.045 186.565 79.570 186.785 ;
        RECT 79.740 187.145 80.610 187.315 ;
        RECT 78.285 185.915 78.535 186.375 ;
        RECT 78.705 186.365 78.875 186.505 ;
        RECT 79.740 186.365 79.910 187.145 ;
        RECT 80.440 187.075 80.610 187.145 ;
        RECT 80.120 186.895 80.320 186.925 ;
        RECT 80.780 186.895 80.950 187.965 ;
        RECT 81.120 187.075 81.310 187.795 ;
        RECT 80.120 186.595 80.950 186.895 ;
        RECT 81.480 186.865 81.800 187.825 ;
        RECT 78.705 186.195 79.040 186.365 ;
        RECT 79.235 186.195 79.910 186.365 ;
        RECT 80.230 185.915 80.600 186.415 ;
        RECT 80.780 186.365 80.950 186.595 ;
        RECT 81.335 186.535 81.800 186.865 ;
        RECT 81.970 187.155 82.140 187.995 ;
        RECT 82.320 187.965 82.635 188.465 ;
        RECT 82.865 187.735 83.205 188.295 ;
        RECT 82.310 187.360 83.205 187.735 ;
        RECT 83.375 187.455 83.545 188.465 ;
        RECT 83.015 187.155 83.205 187.360 ;
        RECT 83.715 187.405 84.045 188.250 ;
        RECT 84.285 187.855 84.615 188.285 ;
        RECT 84.795 188.025 84.990 188.465 ;
        RECT 85.160 187.855 85.490 188.285 ;
        RECT 84.285 187.685 85.490 187.855 ;
        RECT 83.715 187.325 84.105 187.405 ;
        RECT 84.285 187.355 85.180 187.685 ;
        RECT 85.660 187.515 85.935 188.285 ;
        RECT 86.665 187.795 86.835 188.295 ;
        RECT 87.005 187.965 87.335 188.465 ;
        RECT 86.665 187.625 87.330 187.795 ;
        RECT 83.890 187.275 84.105 187.325 ;
        RECT 81.970 186.825 82.845 187.155 ;
        RECT 83.015 186.825 83.765 187.155 ;
        RECT 81.970 186.365 82.140 186.825 ;
        RECT 83.015 186.655 83.215 186.825 ;
        RECT 83.935 186.695 84.105 187.275 ;
        RECT 85.350 187.325 85.935 187.515 ;
        RECT 84.290 186.825 84.585 187.155 ;
        RECT 84.765 186.825 85.180 187.155 ;
        RECT 83.880 186.655 84.105 186.695 ;
        RECT 80.780 186.195 81.185 186.365 ;
        RECT 81.355 186.195 82.140 186.365 ;
        RECT 82.415 185.915 82.625 186.445 ;
        RECT 82.885 186.130 83.215 186.655 ;
        RECT 83.725 186.570 84.105 186.655 ;
        RECT 83.385 185.915 83.555 186.525 ;
        RECT 83.725 186.135 84.055 186.570 ;
        RECT 84.285 185.915 84.585 186.645 ;
        RECT 84.765 186.205 84.995 186.825 ;
        RECT 85.350 186.655 85.525 187.325 ;
        RECT 85.195 186.475 85.525 186.655 ;
        RECT 85.695 186.505 85.935 187.155 ;
        RECT 86.580 186.805 86.930 187.455 ;
        RECT 87.100 186.635 87.330 187.625 ;
        RECT 85.195 186.095 85.420 186.475 ;
        RECT 86.665 186.465 87.330 186.635 ;
        RECT 85.590 185.915 85.920 186.305 ;
        RECT 86.665 186.175 86.835 186.465 ;
        RECT 87.005 185.915 87.335 186.295 ;
        RECT 87.505 186.175 87.690 188.295 ;
        RECT 87.930 188.005 88.195 188.465 ;
        RECT 88.365 187.870 88.615 188.295 ;
        RECT 88.825 188.020 89.930 188.190 ;
        RECT 88.310 187.740 88.615 187.870 ;
        RECT 87.860 186.545 88.140 187.495 ;
        RECT 88.310 186.635 88.480 187.740 ;
        RECT 88.650 186.955 88.890 187.550 ;
        RECT 89.060 187.485 89.590 187.850 ;
        RECT 89.060 186.785 89.230 187.485 ;
        RECT 89.760 187.405 89.930 188.020 ;
        RECT 90.100 187.665 90.270 188.465 ;
        RECT 90.440 187.965 90.690 188.295 ;
        RECT 90.915 187.995 91.800 188.165 ;
        RECT 89.760 187.315 90.270 187.405 ;
        RECT 88.310 186.505 88.535 186.635 ;
        RECT 88.705 186.565 89.230 186.785 ;
        RECT 89.400 187.145 90.270 187.315 ;
        RECT 87.945 185.915 88.195 186.375 ;
        RECT 88.365 186.365 88.535 186.505 ;
        RECT 89.400 186.365 89.570 187.145 ;
        RECT 90.100 187.075 90.270 187.145 ;
        RECT 89.780 186.895 89.980 186.925 ;
        RECT 90.440 186.895 90.610 187.965 ;
        RECT 90.780 187.075 90.970 187.795 ;
        RECT 89.780 186.595 90.610 186.895 ;
        RECT 91.140 186.865 91.460 187.825 ;
        RECT 88.365 186.195 88.700 186.365 ;
        RECT 88.895 186.195 89.570 186.365 ;
        RECT 89.890 185.915 90.260 186.415 ;
        RECT 90.440 186.365 90.610 186.595 ;
        RECT 90.995 186.535 91.460 186.865 ;
        RECT 91.630 187.155 91.800 187.995 ;
        RECT 91.980 187.965 92.295 188.465 ;
        RECT 92.525 187.735 92.865 188.295 ;
        RECT 91.970 187.360 92.865 187.735 ;
        RECT 93.035 187.455 93.205 188.465 ;
        RECT 92.675 187.155 92.865 187.360 ;
        RECT 93.375 187.405 93.705 188.250 ;
        RECT 93.945 187.855 94.275 188.285 ;
        RECT 94.455 188.025 94.650 188.465 ;
        RECT 94.820 187.855 95.150 188.285 ;
        RECT 93.945 187.685 95.150 187.855 ;
        RECT 93.375 187.325 93.765 187.405 ;
        RECT 93.945 187.355 94.840 187.685 ;
        RECT 95.320 187.515 95.595 188.285 ;
        RECT 96.350 187.835 96.635 188.295 ;
        RECT 96.805 188.005 97.075 188.465 ;
        RECT 96.350 187.615 97.305 187.835 ;
        RECT 93.550 187.275 93.765 187.325 ;
        RECT 91.630 186.825 92.505 187.155 ;
        RECT 92.675 186.825 93.425 187.155 ;
        RECT 91.630 186.365 91.800 186.825 ;
        RECT 92.675 186.655 92.875 186.825 ;
        RECT 93.595 186.695 93.765 187.275 ;
        RECT 95.010 187.325 95.595 187.515 ;
        RECT 93.950 186.825 94.245 187.155 ;
        RECT 94.425 186.825 94.840 187.155 ;
        RECT 93.540 186.655 93.765 186.695 ;
        RECT 90.440 186.195 90.845 186.365 ;
        RECT 91.015 186.195 91.800 186.365 ;
        RECT 92.075 185.915 92.285 186.445 ;
        RECT 92.545 186.130 92.875 186.655 ;
        RECT 93.385 186.570 93.765 186.655 ;
        RECT 93.045 185.915 93.215 186.525 ;
        RECT 93.385 186.135 93.715 186.570 ;
        RECT 93.945 185.915 94.245 186.645 ;
        RECT 94.425 186.205 94.655 186.825 ;
        RECT 95.010 186.655 95.185 187.325 ;
        RECT 94.855 186.475 95.185 186.655 ;
        RECT 95.355 186.505 95.595 187.155 ;
        RECT 96.235 186.885 96.925 187.445 ;
        RECT 97.095 186.715 97.305 187.615 ;
        RECT 96.350 186.545 97.305 186.715 ;
        RECT 97.475 187.445 97.875 188.295 ;
        RECT 98.065 187.835 98.345 188.295 ;
        RECT 98.865 188.005 99.190 188.465 ;
        RECT 98.065 187.615 99.190 187.835 ;
        RECT 97.475 186.885 98.570 187.445 ;
        RECT 98.740 187.155 99.190 187.615 ;
        RECT 99.360 187.325 99.745 188.295 ;
        RECT 94.855 186.095 95.080 186.475 ;
        RECT 95.250 185.915 95.580 186.305 ;
        RECT 96.350 186.085 96.635 186.545 ;
        RECT 96.805 185.915 97.075 186.375 ;
        RECT 97.475 186.085 97.875 186.885 ;
        RECT 98.740 186.825 99.295 187.155 ;
        RECT 98.740 186.715 99.190 186.825 ;
        RECT 98.065 186.545 99.190 186.715 ;
        RECT 99.465 186.655 99.745 187.325 ;
        RECT 99.915 187.300 100.205 188.465 ;
        RECT 100.375 187.325 100.635 188.295 ;
        RECT 100.805 188.040 101.190 188.465 ;
        RECT 101.360 187.870 101.615 188.295 ;
        RECT 100.805 187.675 101.615 187.870 ;
        RECT 98.065 186.085 98.345 186.545 ;
        RECT 98.865 185.915 99.190 186.375 ;
        RECT 99.360 186.085 99.745 186.655 ;
        RECT 100.375 186.655 100.560 187.325 ;
        RECT 100.805 187.155 101.155 187.675 ;
        RECT 101.805 187.505 102.050 188.295 ;
        RECT 102.220 188.040 102.605 188.465 ;
        RECT 102.775 187.870 103.050 188.295 ;
        RECT 100.730 186.825 101.155 187.155 ;
        RECT 101.325 187.325 102.050 187.505 ;
        RECT 102.220 187.675 103.050 187.870 ;
        RECT 101.325 186.825 101.975 187.325 ;
        RECT 102.220 187.155 102.570 187.675 ;
        RECT 103.220 187.505 103.645 188.295 ;
        RECT 103.815 188.040 104.200 188.465 ;
        RECT 104.370 187.870 104.805 188.295 ;
        RECT 102.145 186.825 102.570 187.155 ;
        RECT 102.740 187.325 103.645 187.505 ;
        RECT 103.815 187.700 104.805 187.870 ;
        RECT 102.740 186.825 103.570 187.325 ;
        RECT 103.815 187.155 104.150 187.700 ;
        RECT 103.740 186.825 104.150 187.155 ;
        RECT 104.320 186.825 104.805 187.530 ;
        RECT 104.985 187.495 105.315 188.280 ;
        RECT 104.985 187.325 105.665 187.495 ;
        RECT 105.845 187.325 106.175 188.465 ;
        RECT 106.355 187.325 106.740 188.295 ;
        RECT 106.910 188.005 107.235 188.465 ;
        RECT 107.755 187.835 108.035 188.295 ;
        RECT 106.910 187.615 108.035 187.835 ;
        RECT 104.975 186.905 105.325 187.155 ;
        RECT 100.805 186.655 101.155 186.825 ;
        RECT 101.805 186.655 101.975 186.825 ;
        RECT 102.220 186.655 102.570 186.825 ;
        RECT 103.220 186.655 103.570 186.825 ;
        RECT 103.815 186.655 104.150 186.825 ;
        RECT 105.495 186.725 105.665 187.325 ;
        RECT 105.835 186.905 106.185 187.155 ;
        RECT 99.915 185.915 100.205 186.640 ;
        RECT 100.375 186.085 100.635 186.655 ;
        RECT 100.805 186.485 101.615 186.655 ;
        RECT 100.805 185.915 101.190 186.315 ;
        RECT 101.360 186.085 101.615 186.485 ;
        RECT 101.805 186.085 102.050 186.655 ;
        RECT 102.220 186.485 103.030 186.655 ;
        RECT 102.220 185.915 102.605 186.315 ;
        RECT 102.775 186.085 103.030 186.485 ;
        RECT 103.220 186.085 103.645 186.655 ;
        RECT 103.815 186.485 104.805 186.655 ;
        RECT 103.815 185.915 104.200 186.315 ;
        RECT 104.370 186.085 104.805 186.485 ;
        RECT 104.995 185.915 105.235 186.725 ;
        RECT 105.405 186.085 105.735 186.725 ;
        RECT 105.905 185.915 106.175 186.725 ;
        RECT 106.355 186.655 106.635 187.325 ;
        RECT 106.910 187.155 107.360 187.615 ;
        RECT 108.225 187.445 108.625 188.295 ;
        RECT 109.025 188.005 109.295 188.465 ;
        RECT 109.465 187.835 109.750 188.295 ;
        RECT 106.805 186.825 107.360 187.155 ;
        RECT 107.530 186.885 108.625 187.445 ;
        RECT 106.910 186.715 107.360 186.825 ;
        RECT 106.355 186.085 106.740 186.655 ;
        RECT 106.910 186.545 108.035 186.715 ;
        RECT 106.910 185.915 107.235 186.375 ;
        RECT 107.755 186.085 108.035 186.545 ;
        RECT 108.225 186.085 108.625 186.885 ;
        RECT 108.795 187.615 109.750 187.835 ;
        RECT 110.150 187.835 110.435 188.295 ;
        RECT 110.605 188.005 110.875 188.465 ;
        RECT 110.150 187.615 111.105 187.835 ;
        RECT 108.795 186.715 109.005 187.615 ;
        RECT 109.175 186.885 109.865 187.445 ;
        RECT 110.035 186.885 110.725 187.445 ;
        RECT 110.895 186.715 111.105 187.615 ;
        RECT 108.795 186.545 109.750 186.715 ;
        RECT 109.025 185.915 109.295 186.375 ;
        RECT 109.465 186.085 109.750 186.545 ;
        RECT 110.150 186.545 111.105 186.715 ;
        RECT 111.275 187.445 111.675 188.295 ;
        RECT 111.865 187.835 112.145 188.295 ;
        RECT 112.665 188.005 112.990 188.465 ;
        RECT 111.865 187.615 112.990 187.835 ;
        RECT 111.275 186.885 112.370 187.445 ;
        RECT 112.540 187.155 112.990 187.615 ;
        RECT 113.160 187.325 113.545 188.295 ;
        RECT 110.150 186.085 110.435 186.545 ;
        RECT 110.605 185.915 110.875 186.375 ;
        RECT 111.275 186.085 111.675 186.885 ;
        RECT 112.540 186.825 113.095 187.155 ;
        RECT 112.540 186.715 112.990 186.825 ;
        RECT 111.865 186.545 112.990 186.715 ;
        RECT 113.265 186.655 113.545 187.325 ;
        RECT 114.175 187.375 115.385 188.465 ;
        RECT 114.175 186.835 114.695 187.375 ;
        RECT 114.865 186.665 115.385 187.205 ;
        RECT 111.865 186.085 112.145 186.545 ;
        RECT 112.665 185.915 112.990 186.375 ;
        RECT 113.160 186.085 113.545 186.655 ;
        RECT 114.175 185.915 115.385 186.665 ;
        RECT 61.190 185.745 115.470 185.915 ;
        RECT 61.275 184.995 62.485 185.745 ;
        RECT 62.655 185.200 68.000 185.745 ;
        RECT 61.275 184.455 61.795 184.995 ;
        RECT 61.965 184.285 62.485 184.825 ;
        RECT 64.240 184.370 64.580 185.200 ;
        RECT 68.175 184.995 69.385 185.745 ;
        RECT 69.645 185.195 69.815 185.485 ;
        RECT 69.985 185.365 70.315 185.745 ;
        RECT 69.645 185.025 70.310 185.195 ;
        RECT 61.275 183.195 62.485 184.285 ;
        RECT 66.060 183.630 66.410 184.880 ;
        RECT 68.175 184.455 68.695 184.995 ;
        RECT 68.865 184.285 69.385 184.825 ;
        RECT 62.655 183.195 68.000 183.630 ;
        RECT 68.175 183.195 69.385 184.285 ;
        RECT 69.560 184.205 69.910 184.855 ;
        RECT 70.080 184.035 70.310 185.025 ;
        RECT 69.645 183.865 70.310 184.035 ;
        RECT 69.645 183.365 69.815 183.865 ;
        RECT 69.985 183.195 70.315 183.695 ;
        RECT 70.485 183.365 70.670 185.485 ;
        RECT 70.925 185.285 71.175 185.745 ;
        RECT 71.345 185.295 71.680 185.465 ;
        RECT 71.875 185.295 72.550 185.465 ;
        RECT 71.345 185.155 71.515 185.295 ;
        RECT 70.840 184.165 71.120 185.115 ;
        RECT 71.290 185.025 71.515 185.155 ;
        RECT 71.290 183.920 71.460 185.025 ;
        RECT 71.685 184.875 72.210 185.095 ;
        RECT 71.630 184.110 71.870 184.705 ;
        RECT 72.040 184.175 72.210 184.875 ;
        RECT 72.380 184.515 72.550 185.295 ;
        RECT 72.870 185.245 73.240 185.745 ;
        RECT 73.420 185.295 73.825 185.465 ;
        RECT 73.995 185.295 74.780 185.465 ;
        RECT 73.420 185.065 73.590 185.295 ;
        RECT 72.760 184.765 73.590 185.065 ;
        RECT 73.975 184.795 74.440 185.125 ;
        RECT 72.760 184.735 72.960 184.765 ;
        RECT 73.080 184.515 73.250 184.585 ;
        RECT 72.380 184.345 73.250 184.515 ;
        RECT 72.740 184.255 73.250 184.345 ;
        RECT 71.290 183.790 71.595 183.920 ;
        RECT 72.040 183.810 72.570 184.175 ;
        RECT 70.910 183.195 71.175 183.655 ;
        RECT 71.345 183.365 71.595 183.790 ;
        RECT 72.740 183.640 72.910 184.255 ;
        RECT 71.805 183.470 72.910 183.640 ;
        RECT 73.080 183.195 73.250 183.995 ;
        RECT 73.420 183.695 73.590 184.765 ;
        RECT 73.760 183.865 73.950 184.585 ;
        RECT 74.120 183.835 74.440 184.795 ;
        RECT 74.610 184.835 74.780 185.295 ;
        RECT 75.055 185.215 75.265 185.745 ;
        RECT 75.525 185.005 75.855 185.530 ;
        RECT 76.025 185.135 76.195 185.745 ;
        RECT 76.365 185.090 76.695 185.525 ;
        RECT 77.005 185.195 77.175 185.485 ;
        RECT 77.345 185.365 77.675 185.745 ;
        RECT 76.365 185.005 76.745 185.090 ;
        RECT 77.005 185.025 77.670 185.195 ;
        RECT 75.655 184.835 75.855 185.005 ;
        RECT 76.520 184.965 76.745 185.005 ;
        RECT 74.610 184.505 75.485 184.835 ;
        RECT 75.655 184.505 76.405 184.835 ;
        RECT 73.420 183.365 73.670 183.695 ;
        RECT 74.610 183.665 74.780 184.505 ;
        RECT 75.655 184.300 75.845 184.505 ;
        RECT 76.575 184.385 76.745 184.965 ;
        RECT 76.530 184.335 76.745 184.385 ;
        RECT 74.950 183.925 75.845 184.300 ;
        RECT 76.355 184.255 76.745 184.335 ;
        RECT 73.895 183.495 74.780 183.665 ;
        RECT 74.960 183.195 75.275 183.695 ;
        RECT 75.505 183.365 75.845 183.925 ;
        RECT 76.015 183.195 76.185 184.205 ;
        RECT 76.355 183.410 76.685 184.255 ;
        RECT 76.920 184.205 77.270 184.855 ;
        RECT 77.440 184.035 77.670 185.025 ;
        RECT 77.005 183.865 77.670 184.035 ;
        RECT 77.005 183.365 77.175 183.865 ;
        RECT 77.345 183.195 77.675 183.695 ;
        RECT 77.845 183.365 78.030 185.485 ;
        RECT 78.285 185.285 78.535 185.745 ;
        RECT 78.705 185.295 79.040 185.465 ;
        RECT 79.235 185.295 79.910 185.465 ;
        RECT 78.705 185.155 78.875 185.295 ;
        RECT 78.200 184.165 78.480 185.115 ;
        RECT 78.650 185.025 78.875 185.155 ;
        RECT 78.650 183.920 78.820 185.025 ;
        RECT 79.045 184.875 79.570 185.095 ;
        RECT 78.990 184.110 79.230 184.705 ;
        RECT 79.400 184.175 79.570 184.875 ;
        RECT 79.740 184.515 79.910 185.295 ;
        RECT 80.230 185.245 80.600 185.745 ;
        RECT 80.780 185.295 81.185 185.465 ;
        RECT 81.355 185.295 82.140 185.465 ;
        RECT 80.780 185.065 80.950 185.295 ;
        RECT 80.120 184.765 80.950 185.065 ;
        RECT 81.335 184.795 81.800 185.125 ;
        RECT 80.120 184.735 80.320 184.765 ;
        RECT 80.440 184.515 80.610 184.585 ;
        RECT 79.740 184.345 80.610 184.515 ;
        RECT 80.100 184.255 80.610 184.345 ;
        RECT 78.650 183.790 78.955 183.920 ;
        RECT 79.400 183.810 79.930 184.175 ;
        RECT 78.270 183.195 78.535 183.655 ;
        RECT 78.705 183.365 78.955 183.790 ;
        RECT 80.100 183.640 80.270 184.255 ;
        RECT 79.165 183.470 80.270 183.640 ;
        RECT 80.440 183.195 80.610 183.995 ;
        RECT 80.780 183.695 80.950 184.765 ;
        RECT 81.120 183.865 81.310 184.585 ;
        RECT 81.480 183.835 81.800 184.795 ;
        RECT 81.970 184.835 82.140 185.295 ;
        RECT 82.415 185.215 82.625 185.745 ;
        RECT 82.885 185.005 83.215 185.530 ;
        RECT 83.385 185.135 83.555 185.745 ;
        RECT 83.725 185.090 84.055 185.525 ;
        RECT 83.725 185.005 84.105 185.090 ;
        RECT 83.015 184.835 83.215 185.005 ;
        RECT 83.880 184.965 84.105 185.005 ;
        RECT 81.970 184.505 82.845 184.835 ;
        RECT 83.015 184.505 83.765 184.835 ;
        RECT 80.780 183.365 81.030 183.695 ;
        RECT 81.970 183.665 82.140 184.505 ;
        RECT 83.015 184.300 83.205 184.505 ;
        RECT 83.935 184.385 84.105 184.965 ;
        RECT 84.285 184.935 84.555 185.745 ;
        RECT 84.725 184.935 85.055 185.575 ;
        RECT 85.225 184.935 85.465 185.745 ;
        RECT 85.655 184.995 86.865 185.745 ;
        RECT 87.035 185.020 87.325 185.745 ;
        RECT 87.495 184.995 88.705 185.745 ;
        RECT 84.275 184.505 84.625 184.755 ;
        RECT 83.890 184.335 84.105 184.385 ;
        RECT 84.795 184.335 84.965 184.935 ;
        RECT 85.135 184.505 85.485 184.755 ;
        RECT 85.655 184.455 86.175 184.995 ;
        RECT 82.310 183.925 83.205 184.300 ;
        RECT 83.715 184.255 84.105 184.335 ;
        RECT 81.255 183.495 82.140 183.665 ;
        RECT 82.320 183.195 82.635 183.695 ;
        RECT 82.865 183.365 83.205 183.925 ;
        RECT 83.375 183.195 83.545 184.205 ;
        RECT 83.715 183.410 84.045 184.255 ;
        RECT 84.285 183.195 84.615 184.335 ;
        RECT 84.795 184.165 85.475 184.335 ;
        RECT 86.345 184.285 86.865 184.825 ;
        RECT 87.495 184.455 88.015 184.995 ;
        RECT 88.885 184.935 89.155 185.745 ;
        RECT 89.325 184.935 89.655 185.575 ;
        RECT 89.825 184.935 90.065 185.745 ;
        RECT 90.345 185.195 90.515 185.485 ;
        RECT 90.685 185.365 91.015 185.745 ;
        RECT 90.345 185.025 91.010 185.195 ;
        RECT 85.145 183.380 85.475 184.165 ;
        RECT 85.655 183.195 86.865 184.285 ;
        RECT 87.035 183.195 87.325 184.360 ;
        RECT 88.185 184.285 88.705 184.825 ;
        RECT 88.875 184.505 89.225 184.755 ;
        RECT 89.395 184.335 89.565 184.935 ;
        RECT 89.735 184.505 90.085 184.755 ;
        RECT 87.495 183.195 88.705 184.285 ;
        RECT 88.885 183.195 89.215 184.335 ;
        RECT 89.395 184.165 90.075 184.335 ;
        RECT 90.260 184.205 90.610 184.855 ;
        RECT 89.745 183.380 90.075 184.165 ;
        RECT 90.780 184.035 91.010 185.025 ;
        RECT 90.345 183.865 91.010 184.035 ;
        RECT 90.345 183.365 90.515 183.865 ;
        RECT 90.685 183.195 91.015 183.695 ;
        RECT 91.185 183.365 91.370 185.485 ;
        RECT 91.625 185.285 91.875 185.745 ;
        RECT 92.045 185.295 92.380 185.465 ;
        RECT 92.575 185.295 93.250 185.465 ;
        RECT 92.045 185.155 92.215 185.295 ;
        RECT 91.540 184.165 91.820 185.115 ;
        RECT 91.990 185.025 92.215 185.155 ;
        RECT 91.990 183.920 92.160 185.025 ;
        RECT 92.385 184.875 92.910 185.095 ;
        RECT 92.330 184.110 92.570 184.705 ;
        RECT 92.740 184.175 92.910 184.875 ;
        RECT 93.080 184.515 93.250 185.295 ;
        RECT 93.570 185.245 93.940 185.745 ;
        RECT 94.120 185.295 94.525 185.465 ;
        RECT 94.695 185.295 95.480 185.465 ;
        RECT 94.120 185.065 94.290 185.295 ;
        RECT 93.460 184.765 94.290 185.065 ;
        RECT 94.675 184.795 95.140 185.125 ;
        RECT 93.460 184.735 93.660 184.765 ;
        RECT 93.780 184.515 93.950 184.585 ;
        RECT 93.080 184.345 93.950 184.515 ;
        RECT 93.440 184.255 93.950 184.345 ;
        RECT 91.990 183.790 92.295 183.920 ;
        RECT 92.740 183.810 93.270 184.175 ;
        RECT 91.610 183.195 91.875 183.655 ;
        RECT 92.045 183.365 92.295 183.790 ;
        RECT 93.440 183.640 93.610 184.255 ;
        RECT 92.505 183.470 93.610 183.640 ;
        RECT 93.780 183.195 93.950 183.995 ;
        RECT 94.120 183.695 94.290 184.765 ;
        RECT 94.460 183.865 94.650 184.585 ;
        RECT 94.820 183.835 95.140 184.795 ;
        RECT 95.310 184.835 95.480 185.295 ;
        RECT 95.755 185.215 95.965 185.745 ;
        RECT 96.225 185.005 96.555 185.530 ;
        RECT 96.725 185.135 96.895 185.745 ;
        RECT 97.065 185.090 97.395 185.525 ;
        RECT 97.705 185.195 97.875 185.485 ;
        RECT 98.045 185.365 98.375 185.745 ;
        RECT 97.065 185.005 97.445 185.090 ;
        RECT 97.705 185.025 98.370 185.195 ;
        RECT 96.355 184.835 96.555 185.005 ;
        RECT 97.220 184.965 97.445 185.005 ;
        RECT 95.310 184.505 96.185 184.835 ;
        RECT 96.355 184.505 97.105 184.835 ;
        RECT 94.120 183.365 94.370 183.695 ;
        RECT 95.310 183.665 95.480 184.505 ;
        RECT 96.355 184.300 96.545 184.505 ;
        RECT 97.275 184.385 97.445 184.965 ;
        RECT 97.230 184.335 97.445 184.385 ;
        RECT 95.650 183.925 96.545 184.300 ;
        RECT 97.055 184.255 97.445 184.335 ;
        RECT 94.595 183.495 95.480 183.665 ;
        RECT 95.660 183.195 95.975 183.695 ;
        RECT 96.205 183.365 96.545 183.925 ;
        RECT 96.715 183.195 96.885 184.205 ;
        RECT 97.055 183.410 97.385 184.255 ;
        RECT 97.620 184.205 97.970 184.855 ;
        RECT 98.140 184.035 98.370 185.025 ;
        RECT 97.705 183.865 98.370 184.035 ;
        RECT 97.705 183.365 97.875 183.865 ;
        RECT 98.045 183.195 98.375 183.695 ;
        RECT 98.545 183.365 98.730 185.485 ;
        RECT 98.985 185.285 99.235 185.745 ;
        RECT 99.405 185.295 99.740 185.465 ;
        RECT 99.935 185.295 100.610 185.465 ;
        RECT 99.405 185.155 99.575 185.295 ;
        RECT 98.900 184.165 99.180 185.115 ;
        RECT 99.350 185.025 99.575 185.155 ;
        RECT 99.350 183.920 99.520 185.025 ;
        RECT 99.745 184.875 100.270 185.095 ;
        RECT 99.690 184.110 99.930 184.705 ;
        RECT 100.100 184.175 100.270 184.875 ;
        RECT 100.440 184.515 100.610 185.295 ;
        RECT 100.930 185.245 101.300 185.745 ;
        RECT 101.480 185.295 101.885 185.465 ;
        RECT 102.055 185.295 102.840 185.465 ;
        RECT 101.480 185.065 101.650 185.295 ;
        RECT 100.820 184.765 101.650 185.065 ;
        RECT 102.035 184.795 102.500 185.125 ;
        RECT 100.820 184.735 101.020 184.765 ;
        RECT 101.140 184.515 101.310 184.585 ;
        RECT 100.440 184.345 101.310 184.515 ;
        RECT 100.800 184.255 101.310 184.345 ;
        RECT 99.350 183.790 99.655 183.920 ;
        RECT 100.100 183.810 100.630 184.175 ;
        RECT 98.970 183.195 99.235 183.655 ;
        RECT 99.405 183.365 99.655 183.790 ;
        RECT 100.800 183.640 100.970 184.255 ;
        RECT 99.865 183.470 100.970 183.640 ;
        RECT 101.140 183.195 101.310 183.995 ;
        RECT 101.480 183.695 101.650 184.765 ;
        RECT 101.820 183.865 102.010 184.585 ;
        RECT 102.180 183.835 102.500 184.795 ;
        RECT 102.670 184.835 102.840 185.295 ;
        RECT 103.115 185.215 103.325 185.745 ;
        RECT 103.585 185.005 103.915 185.530 ;
        RECT 104.085 185.135 104.255 185.745 ;
        RECT 104.425 185.090 104.755 185.525 ;
        RECT 105.065 185.195 105.235 185.485 ;
        RECT 105.405 185.365 105.735 185.745 ;
        RECT 104.425 185.005 104.805 185.090 ;
        RECT 105.065 185.025 105.730 185.195 ;
        RECT 103.715 184.835 103.915 185.005 ;
        RECT 104.580 184.965 104.805 185.005 ;
        RECT 102.670 184.505 103.545 184.835 ;
        RECT 103.715 184.505 104.465 184.835 ;
        RECT 101.480 183.365 101.730 183.695 ;
        RECT 102.670 183.665 102.840 184.505 ;
        RECT 103.715 184.300 103.905 184.505 ;
        RECT 104.635 184.385 104.805 184.965 ;
        RECT 104.590 184.335 104.805 184.385 ;
        RECT 103.010 183.925 103.905 184.300 ;
        RECT 104.415 184.255 104.805 184.335 ;
        RECT 101.955 183.495 102.840 183.665 ;
        RECT 103.020 183.195 103.335 183.695 ;
        RECT 103.565 183.365 103.905 183.925 ;
        RECT 104.075 183.195 104.245 184.205 ;
        RECT 104.415 183.410 104.745 184.255 ;
        RECT 104.980 184.205 105.330 184.855 ;
        RECT 105.500 184.035 105.730 185.025 ;
        RECT 105.065 183.865 105.730 184.035 ;
        RECT 105.065 183.365 105.235 183.865 ;
        RECT 105.405 183.195 105.735 183.695 ;
        RECT 105.905 183.365 106.090 185.485 ;
        RECT 106.345 185.285 106.595 185.745 ;
        RECT 106.765 185.295 107.100 185.465 ;
        RECT 107.295 185.295 107.970 185.465 ;
        RECT 106.765 185.155 106.935 185.295 ;
        RECT 106.260 184.165 106.540 185.115 ;
        RECT 106.710 185.025 106.935 185.155 ;
        RECT 106.710 183.920 106.880 185.025 ;
        RECT 107.105 184.875 107.630 185.095 ;
        RECT 107.050 184.110 107.290 184.705 ;
        RECT 107.460 184.175 107.630 184.875 ;
        RECT 107.800 184.515 107.970 185.295 ;
        RECT 108.290 185.245 108.660 185.745 ;
        RECT 108.840 185.295 109.245 185.465 ;
        RECT 109.415 185.295 110.200 185.465 ;
        RECT 108.840 185.065 109.010 185.295 ;
        RECT 108.180 184.765 109.010 185.065 ;
        RECT 109.395 184.795 109.860 185.125 ;
        RECT 108.180 184.735 108.380 184.765 ;
        RECT 108.500 184.515 108.670 184.585 ;
        RECT 107.800 184.345 108.670 184.515 ;
        RECT 108.160 184.255 108.670 184.345 ;
        RECT 106.710 183.790 107.015 183.920 ;
        RECT 107.460 183.810 107.990 184.175 ;
        RECT 106.330 183.195 106.595 183.655 ;
        RECT 106.765 183.365 107.015 183.790 ;
        RECT 108.160 183.640 108.330 184.255 ;
        RECT 107.225 183.470 108.330 183.640 ;
        RECT 108.500 183.195 108.670 183.995 ;
        RECT 108.840 183.695 109.010 184.765 ;
        RECT 109.180 183.865 109.370 184.585 ;
        RECT 109.540 183.835 109.860 184.795 ;
        RECT 110.030 184.835 110.200 185.295 ;
        RECT 110.475 185.215 110.685 185.745 ;
        RECT 110.945 185.005 111.275 185.530 ;
        RECT 111.445 185.135 111.615 185.745 ;
        RECT 111.785 185.090 112.115 185.525 ;
        RECT 111.785 185.005 112.165 185.090 ;
        RECT 112.795 185.020 113.085 185.745 ;
        RECT 111.075 184.835 111.275 185.005 ;
        RECT 111.940 184.965 112.165 185.005 ;
        RECT 114.175 184.995 115.385 185.745 ;
        RECT 110.030 184.505 110.905 184.835 ;
        RECT 111.075 184.505 111.825 184.835 ;
        RECT 108.840 183.365 109.090 183.695 ;
        RECT 110.030 183.665 110.200 184.505 ;
        RECT 111.075 184.300 111.265 184.505 ;
        RECT 111.995 184.385 112.165 184.965 ;
        RECT 111.950 184.335 112.165 184.385 ;
        RECT 110.370 183.925 111.265 184.300 ;
        RECT 111.775 184.255 112.165 184.335 ;
        RECT 109.315 183.495 110.200 183.665 ;
        RECT 110.380 183.195 110.695 183.695 ;
        RECT 110.925 183.365 111.265 183.925 ;
        RECT 111.435 183.195 111.605 184.205 ;
        RECT 111.775 183.410 112.105 184.255 ;
        RECT 112.795 183.195 113.085 184.360 ;
        RECT 114.175 184.285 114.695 184.825 ;
        RECT 114.865 184.455 115.385 184.995 ;
        RECT 114.175 183.195 115.385 184.285 ;
        RECT 61.190 183.025 115.470 183.195 ;
        RECT 61.275 181.935 62.485 183.025 ;
        RECT 62.655 182.590 68.000 183.025 ;
        RECT 68.175 182.590 73.520 183.025 ;
        RECT 61.275 181.225 61.795 181.765 ;
        RECT 61.965 181.395 62.485 181.935 ;
        RECT 61.275 180.475 62.485 181.225 ;
        RECT 64.240 181.020 64.580 181.850 ;
        RECT 66.060 181.340 66.410 182.590 ;
        RECT 69.760 181.020 70.100 181.850 ;
        RECT 71.580 181.340 71.930 182.590 ;
        RECT 74.155 181.860 74.445 183.025 ;
        RECT 74.615 181.935 76.285 183.025 ;
        RECT 74.615 181.245 75.365 181.765 ;
        RECT 75.535 181.415 76.285 181.935 ;
        RECT 76.925 182.075 77.200 182.845 ;
        RECT 77.370 182.415 77.700 182.845 ;
        RECT 77.870 182.585 78.065 183.025 ;
        RECT 78.245 182.415 78.575 182.845 ;
        RECT 77.370 182.245 78.575 182.415 ;
        RECT 76.925 181.885 77.510 182.075 ;
        RECT 77.680 181.915 78.575 182.245 ;
        RECT 62.655 180.475 68.000 181.020 ;
        RECT 68.175 180.475 73.520 181.020 ;
        RECT 74.155 180.475 74.445 181.200 ;
        RECT 74.615 180.475 76.285 181.245 ;
        RECT 76.925 181.065 77.165 181.715 ;
        RECT 77.335 181.215 77.510 181.885 ;
        RECT 77.680 181.385 78.095 181.715 ;
        RECT 78.275 181.385 78.570 181.715 ;
        RECT 79.215 181.420 79.495 182.855 ;
        RECT 79.665 182.250 80.375 183.025 ;
        RECT 80.545 182.080 80.875 182.855 ;
        RECT 79.725 181.865 80.875 182.080 ;
        RECT 77.335 181.035 77.665 181.215 ;
        RECT 76.940 180.475 77.270 180.865 ;
        RECT 77.440 180.655 77.665 181.035 ;
        RECT 77.865 180.765 78.095 181.385 ;
        RECT 78.275 180.475 78.575 181.205 ;
        RECT 79.215 180.645 79.555 181.420 ;
        RECT 79.725 181.295 80.010 181.865 ;
        RECT 80.195 181.465 80.665 181.695 ;
        RECT 81.070 181.665 81.285 182.780 ;
        RECT 81.465 182.305 81.795 183.025 ;
        RECT 81.575 181.665 81.805 182.005 ;
        RECT 80.835 181.485 81.285 181.665 ;
        RECT 80.835 181.465 81.165 181.485 ;
        RECT 81.475 181.465 81.805 181.665 ;
        RECT 82.895 181.885 83.280 182.855 ;
        RECT 83.450 182.565 83.775 183.025 ;
        RECT 84.295 182.395 84.575 182.855 ;
        RECT 83.450 182.175 84.575 182.395 ;
        RECT 79.725 181.105 80.435 181.295 ;
        RECT 80.135 180.965 80.435 181.105 ;
        RECT 80.625 181.105 81.805 181.295 ;
        RECT 80.625 181.025 80.955 181.105 ;
        RECT 80.135 180.955 80.450 180.965 ;
        RECT 80.135 180.945 80.460 180.955 ;
        RECT 80.135 180.940 80.470 180.945 ;
        RECT 79.725 180.475 79.895 180.935 ;
        RECT 80.135 180.930 80.475 180.940 ;
        RECT 80.135 180.925 80.480 180.930 ;
        RECT 80.135 180.915 80.485 180.925 ;
        RECT 80.135 180.910 80.490 180.915 ;
        RECT 80.135 180.645 80.495 180.910 ;
        RECT 81.125 180.475 81.295 180.935 ;
        RECT 81.465 180.645 81.805 181.105 ;
        RECT 82.895 181.215 83.175 181.885 ;
        RECT 83.450 181.715 83.900 182.175 ;
        RECT 84.765 182.005 85.165 182.855 ;
        RECT 85.565 182.565 85.835 183.025 ;
        RECT 86.005 182.395 86.290 182.855 ;
        RECT 83.345 181.385 83.900 181.715 ;
        RECT 84.070 181.445 85.165 182.005 ;
        RECT 83.450 181.275 83.900 181.385 ;
        RECT 82.895 180.645 83.280 181.215 ;
        RECT 83.450 181.105 84.575 181.275 ;
        RECT 83.450 180.475 83.775 180.935 ;
        RECT 84.295 180.645 84.575 181.105 ;
        RECT 84.765 180.645 85.165 181.445 ;
        RECT 85.335 182.175 86.290 182.395 ;
        RECT 87.585 182.355 87.755 182.855 ;
        RECT 87.925 182.525 88.255 183.025 ;
        RECT 87.585 182.185 88.250 182.355 ;
        RECT 85.335 181.275 85.545 182.175 ;
        RECT 85.715 181.445 86.405 182.005 ;
        RECT 87.500 181.365 87.850 182.015 ;
        RECT 85.335 181.105 86.290 181.275 ;
        RECT 88.020 181.195 88.250 182.185 ;
        RECT 85.565 180.475 85.835 180.935 ;
        RECT 86.005 180.645 86.290 181.105 ;
        RECT 87.585 181.025 88.250 181.195 ;
        RECT 87.585 180.735 87.755 181.025 ;
        RECT 87.925 180.475 88.255 180.855 ;
        RECT 88.425 180.735 88.610 182.855 ;
        RECT 88.850 182.565 89.115 183.025 ;
        RECT 89.285 182.430 89.535 182.855 ;
        RECT 89.745 182.580 90.850 182.750 ;
        RECT 89.230 182.300 89.535 182.430 ;
        RECT 88.780 181.105 89.060 182.055 ;
        RECT 89.230 181.195 89.400 182.300 ;
        RECT 89.570 181.515 89.810 182.110 ;
        RECT 89.980 182.045 90.510 182.410 ;
        RECT 89.980 181.345 90.150 182.045 ;
        RECT 90.680 181.965 90.850 182.580 ;
        RECT 91.020 182.225 91.190 183.025 ;
        RECT 91.360 182.525 91.610 182.855 ;
        RECT 91.835 182.555 92.720 182.725 ;
        RECT 90.680 181.875 91.190 181.965 ;
        RECT 89.230 181.065 89.455 181.195 ;
        RECT 89.625 181.125 90.150 181.345 ;
        RECT 90.320 181.705 91.190 181.875 ;
        RECT 88.865 180.475 89.115 180.935 ;
        RECT 89.285 180.925 89.455 181.065 ;
        RECT 90.320 180.925 90.490 181.705 ;
        RECT 91.020 181.635 91.190 181.705 ;
        RECT 90.700 181.455 90.900 181.485 ;
        RECT 91.360 181.455 91.530 182.525 ;
        RECT 91.700 181.635 91.890 182.355 ;
        RECT 90.700 181.155 91.530 181.455 ;
        RECT 92.060 181.425 92.380 182.385 ;
        RECT 89.285 180.755 89.620 180.925 ;
        RECT 89.815 180.755 90.490 180.925 ;
        RECT 90.810 180.475 91.180 180.975 ;
        RECT 91.360 180.925 91.530 181.155 ;
        RECT 91.915 181.095 92.380 181.425 ;
        RECT 92.550 181.715 92.720 182.555 ;
        RECT 92.900 182.525 93.215 183.025 ;
        RECT 93.445 182.295 93.785 182.855 ;
        RECT 92.890 181.920 93.785 182.295 ;
        RECT 93.955 182.015 94.125 183.025 ;
        RECT 93.595 181.715 93.785 181.920 ;
        RECT 94.295 181.965 94.625 182.810 ;
        RECT 95.890 182.395 96.175 182.855 ;
        RECT 96.345 182.565 96.615 183.025 ;
        RECT 95.890 182.175 96.845 182.395 ;
        RECT 94.295 181.885 94.685 181.965 ;
        RECT 94.470 181.835 94.685 181.885 ;
        RECT 92.550 181.385 93.425 181.715 ;
        RECT 93.595 181.385 94.345 181.715 ;
        RECT 92.550 180.925 92.720 181.385 ;
        RECT 93.595 181.215 93.795 181.385 ;
        RECT 94.515 181.255 94.685 181.835 ;
        RECT 95.775 181.445 96.465 182.005 ;
        RECT 96.635 181.275 96.845 182.175 ;
        RECT 94.460 181.215 94.685 181.255 ;
        RECT 91.360 180.755 91.765 180.925 ;
        RECT 91.935 180.755 92.720 180.925 ;
        RECT 92.995 180.475 93.205 181.005 ;
        RECT 93.465 180.690 93.795 181.215 ;
        RECT 94.305 181.130 94.685 181.215 ;
        RECT 93.965 180.475 94.135 181.085 ;
        RECT 94.305 180.695 94.635 181.130 ;
        RECT 95.890 181.105 96.845 181.275 ;
        RECT 97.015 182.005 97.415 182.855 ;
        RECT 97.605 182.395 97.885 182.855 ;
        RECT 98.405 182.565 98.730 183.025 ;
        RECT 97.605 182.175 98.730 182.395 ;
        RECT 97.015 181.445 98.110 182.005 ;
        RECT 98.280 181.715 98.730 182.175 ;
        RECT 98.900 181.885 99.285 182.855 ;
        RECT 95.890 180.645 96.175 181.105 ;
        RECT 96.345 180.475 96.615 180.935 ;
        RECT 97.015 180.645 97.415 181.445 ;
        RECT 98.280 181.385 98.835 181.715 ;
        RECT 98.280 181.275 98.730 181.385 ;
        RECT 97.605 181.105 98.730 181.275 ;
        RECT 99.005 181.215 99.285 181.885 ;
        RECT 99.915 181.860 100.205 183.025 ;
        RECT 101.300 181.875 101.560 183.025 ;
        RECT 101.735 181.950 101.990 182.855 ;
        RECT 102.160 182.265 102.490 183.025 ;
        RECT 102.705 182.095 102.875 182.855 ;
        RECT 97.605 180.645 97.885 181.105 ;
        RECT 98.405 180.475 98.730 180.935 ;
        RECT 98.900 180.645 99.285 181.215 ;
        RECT 99.915 180.475 100.205 181.200 ;
        RECT 101.300 180.475 101.560 181.315 ;
        RECT 101.735 181.220 101.905 181.950 ;
        RECT 102.160 181.925 102.875 182.095 ;
        RECT 102.160 181.715 102.330 181.925 ;
        RECT 102.075 181.385 102.330 181.715 ;
        RECT 101.735 180.645 101.990 181.220 ;
        RECT 102.160 181.195 102.330 181.385 ;
        RECT 102.610 181.375 102.965 181.745 ;
        RECT 103.135 181.420 103.415 182.855 ;
        RECT 103.585 182.250 104.295 183.025 ;
        RECT 104.465 182.080 104.795 182.855 ;
        RECT 103.645 181.865 104.795 182.080 ;
        RECT 102.160 181.025 102.875 181.195 ;
        RECT 102.160 180.475 102.490 180.855 ;
        RECT 102.705 180.645 102.875 181.025 ;
        RECT 103.135 180.645 103.475 181.420 ;
        RECT 103.645 181.295 103.930 181.865 ;
        RECT 104.115 181.465 104.585 181.695 ;
        RECT 104.990 181.665 105.205 182.780 ;
        RECT 105.385 182.305 105.715 183.025 ;
        RECT 105.495 181.665 105.725 182.005 ;
        RECT 105.955 181.965 106.285 182.810 ;
        RECT 106.455 182.015 106.625 183.025 ;
        RECT 106.795 182.295 107.135 182.855 ;
        RECT 107.365 182.525 107.680 183.025 ;
        RECT 107.860 182.555 108.745 182.725 ;
        RECT 104.755 181.485 105.205 181.665 ;
        RECT 104.755 181.465 105.085 181.485 ;
        RECT 105.395 181.465 105.725 181.665 ;
        RECT 105.895 181.885 106.285 181.965 ;
        RECT 106.795 181.920 107.690 182.295 ;
        RECT 105.895 181.835 106.110 181.885 ;
        RECT 103.645 181.105 104.355 181.295 ;
        RECT 104.055 180.965 104.355 181.105 ;
        RECT 104.545 181.105 105.725 181.295 ;
        RECT 105.895 181.255 106.065 181.835 ;
        RECT 106.795 181.715 106.985 181.920 ;
        RECT 107.860 181.715 108.030 182.555 ;
        RECT 108.970 182.525 109.220 182.855 ;
        RECT 106.235 181.385 106.985 181.715 ;
        RECT 107.155 181.385 108.030 181.715 ;
        RECT 105.895 181.215 106.120 181.255 ;
        RECT 106.785 181.215 106.985 181.385 ;
        RECT 105.895 181.130 106.275 181.215 ;
        RECT 104.545 181.025 104.875 181.105 ;
        RECT 104.055 180.955 104.370 180.965 ;
        RECT 104.055 180.945 104.380 180.955 ;
        RECT 104.055 180.940 104.390 180.945 ;
        RECT 103.645 180.475 103.815 180.935 ;
        RECT 104.055 180.930 104.395 180.940 ;
        RECT 104.055 180.925 104.400 180.930 ;
        RECT 104.055 180.915 104.405 180.925 ;
        RECT 104.055 180.910 104.410 180.915 ;
        RECT 104.055 180.645 104.415 180.910 ;
        RECT 105.045 180.475 105.215 180.935 ;
        RECT 105.385 180.645 105.725 181.105 ;
        RECT 105.945 180.695 106.275 181.130 ;
        RECT 106.445 180.475 106.615 181.085 ;
        RECT 106.785 180.690 107.115 181.215 ;
        RECT 107.375 180.475 107.585 181.005 ;
        RECT 107.860 180.925 108.030 181.385 ;
        RECT 108.200 181.425 108.520 182.385 ;
        RECT 108.690 181.635 108.880 182.355 ;
        RECT 109.050 181.455 109.220 182.525 ;
        RECT 109.390 182.225 109.560 183.025 ;
        RECT 109.730 182.580 110.835 182.750 ;
        RECT 109.730 181.965 109.900 182.580 ;
        RECT 111.045 182.430 111.295 182.855 ;
        RECT 111.465 182.565 111.730 183.025 ;
        RECT 110.070 182.045 110.600 182.410 ;
        RECT 111.045 182.300 111.350 182.430 ;
        RECT 109.390 181.875 109.900 181.965 ;
        RECT 109.390 181.705 110.260 181.875 ;
        RECT 109.390 181.635 109.560 181.705 ;
        RECT 109.680 181.455 109.880 181.485 ;
        RECT 108.200 181.095 108.665 181.425 ;
        RECT 109.050 181.155 109.880 181.455 ;
        RECT 109.050 180.925 109.220 181.155 ;
        RECT 107.860 180.755 108.645 180.925 ;
        RECT 108.815 180.755 109.220 180.925 ;
        RECT 109.400 180.475 109.770 180.975 ;
        RECT 110.090 180.925 110.260 181.705 ;
        RECT 110.430 181.345 110.600 182.045 ;
        RECT 110.770 181.515 111.010 182.110 ;
        RECT 110.430 181.125 110.955 181.345 ;
        RECT 111.180 181.195 111.350 182.300 ;
        RECT 111.125 181.065 111.350 181.195 ;
        RECT 111.520 181.105 111.800 182.055 ;
        RECT 111.125 180.925 111.295 181.065 ;
        RECT 110.090 180.755 110.765 180.925 ;
        RECT 110.960 180.755 111.295 180.925 ;
        RECT 111.465 180.475 111.715 180.935 ;
        RECT 111.970 180.735 112.155 182.855 ;
        RECT 112.325 182.525 112.655 183.025 ;
        RECT 112.825 182.355 112.995 182.855 ;
        RECT 112.330 182.185 112.995 182.355 ;
        RECT 112.330 181.195 112.560 182.185 ;
        RECT 112.730 181.365 113.080 182.015 ;
        RECT 114.175 181.935 115.385 183.025 ;
        RECT 114.175 181.395 114.695 181.935 ;
        RECT 114.865 181.225 115.385 181.765 ;
        RECT 112.330 181.025 112.995 181.195 ;
        RECT 112.325 180.475 112.655 180.855 ;
        RECT 112.825 180.735 112.995 181.025 ;
        RECT 114.175 180.475 115.385 181.225 ;
        RECT 61.190 180.305 115.470 180.475 ;
        RECT 61.275 179.555 62.485 180.305 ;
        RECT 62.655 179.760 68.000 180.305 ;
        RECT 68.175 179.760 73.520 180.305 ;
        RECT 73.695 179.760 79.040 180.305 ;
        RECT 79.215 179.760 84.560 180.305 ;
        RECT 61.275 179.015 61.795 179.555 ;
        RECT 61.965 178.845 62.485 179.385 ;
        RECT 64.240 178.930 64.580 179.760 ;
        RECT 61.275 177.755 62.485 178.845 ;
        RECT 66.060 178.190 66.410 179.440 ;
        RECT 69.760 178.930 70.100 179.760 ;
        RECT 71.580 178.190 71.930 179.440 ;
        RECT 75.280 178.930 75.620 179.760 ;
        RECT 77.100 178.190 77.450 179.440 ;
        RECT 80.800 178.930 81.140 179.760 ;
        RECT 84.735 179.535 86.405 180.305 ;
        RECT 87.035 179.580 87.325 180.305 ;
        RECT 87.495 179.760 92.840 180.305 ;
        RECT 82.620 178.190 82.970 179.440 ;
        RECT 84.735 179.015 85.485 179.535 ;
        RECT 85.655 178.845 86.405 179.365 ;
        RECT 89.080 178.930 89.420 179.760 ;
        RECT 93.015 179.535 94.685 180.305 ;
        RECT 95.055 179.675 95.385 180.035 ;
        RECT 96.005 179.845 96.255 180.305 ;
        RECT 96.425 179.845 96.985 180.135 ;
        RECT 62.655 177.755 68.000 178.190 ;
        RECT 68.175 177.755 73.520 178.190 ;
        RECT 73.695 177.755 79.040 178.190 ;
        RECT 79.215 177.755 84.560 178.190 ;
        RECT 84.735 177.755 86.405 178.845 ;
        RECT 87.035 177.755 87.325 178.920 ;
        RECT 90.900 178.190 91.250 179.440 ;
        RECT 93.015 179.015 93.765 179.535 ;
        RECT 95.055 179.485 96.445 179.675 ;
        RECT 96.275 179.395 96.445 179.485 ;
        RECT 93.935 178.845 94.685 179.365 ;
        RECT 87.495 177.755 92.840 178.190 ;
        RECT 93.015 177.755 94.685 178.845 ;
        RECT 94.870 179.065 95.545 179.315 ;
        RECT 95.765 179.065 96.105 179.315 ;
        RECT 96.275 179.065 96.565 179.395 ;
        RECT 94.870 178.705 95.135 179.065 ;
        RECT 96.275 178.815 96.445 179.065 ;
        RECT 95.505 178.645 96.445 178.815 ;
        RECT 95.055 177.755 95.335 178.425 ;
        RECT 95.505 178.095 95.805 178.645 ;
        RECT 96.735 178.475 96.985 179.845 ;
        RECT 97.155 179.535 100.665 180.305 ;
        RECT 97.155 179.015 98.805 179.535 ;
        RECT 101.765 179.495 102.035 180.305 ;
        RECT 102.205 179.495 102.535 180.135 ;
        RECT 102.705 179.495 102.945 180.305 ;
        RECT 104.065 179.575 104.365 180.305 ;
        RECT 98.975 178.845 100.665 179.365 ;
        RECT 101.755 179.065 102.105 179.315 ;
        RECT 102.275 178.895 102.445 179.495 ;
        RECT 104.545 179.395 104.775 180.015 ;
        RECT 104.975 179.745 105.200 180.125 ;
        RECT 105.370 179.915 105.700 180.305 ;
        RECT 104.975 179.565 105.305 179.745 ;
        RECT 102.615 179.065 102.965 179.315 ;
        RECT 104.070 179.065 104.365 179.395 ;
        RECT 104.545 179.065 104.960 179.395 ;
        RECT 105.130 178.895 105.305 179.565 ;
        RECT 105.475 179.065 105.715 179.715 ;
        RECT 105.895 179.555 107.105 180.305 ;
        RECT 107.390 179.675 107.675 180.135 ;
        RECT 107.845 179.845 108.115 180.305 ;
        RECT 105.895 179.015 106.415 179.555 ;
        RECT 107.390 179.505 108.345 179.675 ;
        RECT 96.005 177.755 96.335 178.475 ;
        RECT 96.525 177.925 96.985 178.475 ;
        RECT 97.155 177.755 100.665 178.845 ;
        RECT 101.765 177.755 102.095 178.895 ;
        RECT 102.275 178.725 102.955 178.895 ;
        RECT 102.625 177.940 102.955 178.725 ;
        RECT 104.065 178.535 104.960 178.865 ;
        RECT 105.130 178.705 105.715 178.895 ;
        RECT 106.585 178.845 107.105 179.385 ;
        RECT 104.065 178.365 105.270 178.535 ;
        RECT 104.065 177.935 104.395 178.365 ;
        RECT 104.575 177.755 104.770 178.195 ;
        RECT 104.940 177.935 105.270 178.365 ;
        RECT 105.440 177.935 105.715 178.705 ;
        RECT 105.895 177.755 107.105 178.845 ;
        RECT 107.275 178.775 107.965 179.335 ;
        RECT 108.135 178.605 108.345 179.505 ;
        RECT 107.390 178.385 108.345 178.605 ;
        RECT 108.515 179.335 108.915 180.135 ;
        RECT 109.105 179.675 109.385 180.135 ;
        RECT 109.905 179.845 110.230 180.305 ;
        RECT 109.105 179.505 110.230 179.675 ;
        RECT 110.400 179.565 110.785 180.135 ;
        RECT 110.980 179.915 111.310 180.305 ;
        RECT 111.480 179.745 111.705 180.125 ;
        RECT 109.780 179.395 110.230 179.505 ;
        RECT 108.515 178.775 109.610 179.335 ;
        RECT 109.780 179.065 110.335 179.395 ;
        RECT 107.390 177.925 107.675 178.385 ;
        RECT 107.845 177.755 108.115 178.215 ;
        RECT 108.515 177.925 108.915 178.775 ;
        RECT 109.780 178.605 110.230 179.065 ;
        RECT 110.505 178.895 110.785 179.565 ;
        RECT 110.965 179.065 111.205 179.715 ;
        RECT 111.375 179.565 111.705 179.745 ;
        RECT 111.375 178.895 111.550 179.565 ;
        RECT 111.905 179.395 112.135 180.015 ;
        RECT 112.315 179.575 112.615 180.305 ;
        RECT 112.795 179.580 113.085 180.305 ;
        RECT 114.175 179.555 115.385 180.305 ;
        RECT 111.720 179.065 112.135 179.395 ;
        RECT 112.315 179.065 112.610 179.395 ;
        RECT 109.105 178.385 110.230 178.605 ;
        RECT 109.105 177.925 109.385 178.385 ;
        RECT 109.905 177.755 110.230 178.215 ;
        RECT 110.400 177.925 110.785 178.895 ;
        RECT 110.965 178.705 111.550 178.895 ;
        RECT 110.965 177.935 111.240 178.705 ;
        RECT 111.720 178.535 112.615 178.865 ;
        RECT 111.410 178.365 112.615 178.535 ;
        RECT 111.410 177.935 111.740 178.365 ;
        RECT 111.910 177.755 112.105 178.195 ;
        RECT 112.285 177.935 112.615 178.365 ;
        RECT 112.795 177.755 113.085 178.920 ;
        RECT 114.175 178.845 114.695 179.385 ;
        RECT 114.865 179.015 115.385 179.555 ;
        RECT 114.175 177.755 115.385 178.845 ;
        RECT 61.190 177.585 115.470 177.755 ;
        RECT 61.275 176.495 62.485 177.585 ;
        RECT 62.655 177.150 68.000 177.585 ;
        RECT 68.175 177.150 73.520 177.585 ;
        RECT 61.275 175.785 61.795 176.325 ;
        RECT 61.965 175.955 62.485 176.495 ;
        RECT 61.275 175.035 62.485 175.785 ;
        RECT 64.240 175.580 64.580 176.410 ;
        RECT 66.060 175.900 66.410 177.150 ;
        RECT 69.760 175.580 70.100 176.410 ;
        RECT 71.580 175.900 71.930 177.150 ;
        RECT 74.155 176.420 74.445 177.585 ;
        RECT 74.615 177.150 79.960 177.585 ;
        RECT 80.135 177.150 85.480 177.585 ;
        RECT 85.655 177.150 91.000 177.585 ;
        RECT 91.175 177.150 96.520 177.585 ;
        RECT 62.655 175.035 68.000 175.580 ;
        RECT 68.175 175.035 73.520 175.580 ;
        RECT 74.155 175.035 74.445 175.760 ;
        RECT 76.200 175.580 76.540 176.410 ;
        RECT 78.020 175.900 78.370 177.150 ;
        RECT 81.720 175.580 82.060 176.410 ;
        RECT 83.540 175.900 83.890 177.150 ;
        RECT 87.240 175.580 87.580 176.410 ;
        RECT 89.060 175.900 89.410 177.150 ;
        RECT 92.760 175.580 93.100 176.410 ;
        RECT 94.580 175.900 94.930 177.150 ;
        RECT 96.695 176.495 99.285 177.585 ;
        RECT 96.695 175.805 97.905 176.325 ;
        RECT 98.075 175.975 99.285 176.495 ;
        RECT 99.915 176.420 100.205 177.585 ;
        RECT 100.375 177.150 105.720 177.585 ;
        RECT 74.615 175.035 79.960 175.580 ;
        RECT 80.135 175.035 85.480 175.580 ;
        RECT 85.655 175.035 91.000 175.580 ;
        RECT 91.175 175.035 96.520 175.580 ;
        RECT 96.695 175.035 99.285 175.805 ;
        RECT 99.915 175.035 100.205 175.760 ;
        RECT 101.960 175.580 102.300 176.410 ;
        RECT 103.780 175.900 104.130 177.150 ;
        RECT 105.895 176.495 107.565 177.585 ;
        RECT 108.395 176.915 108.675 177.585 ;
        RECT 108.845 176.695 109.145 177.245 ;
        RECT 109.345 176.865 109.675 177.585 ;
        RECT 109.865 176.865 110.325 177.415 ;
        RECT 105.895 175.805 106.645 176.325 ;
        RECT 106.815 175.975 107.565 176.495 ;
        RECT 108.210 176.275 108.475 176.635 ;
        RECT 108.845 176.525 109.785 176.695 ;
        RECT 109.615 176.275 109.785 176.525 ;
        RECT 108.210 176.025 108.885 176.275 ;
        RECT 109.105 176.025 109.445 176.275 ;
        RECT 109.615 175.945 109.905 176.275 ;
        RECT 109.615 175.855 109.785 175.945 ;
        RECT 100.375 175.035 105.720 175.580 ;
        RECT 105.895 175.035 107.565 175.805 ;
        RECT 108.395 175.665 109.785 175.855 ;
        RECT 108.395 175.305 108.725 175.665 ;
        RECT 110.075 175.495 110.325 176.865 ;
        RECT 109.345 175.035 109.595 175.495 ;
        RECT 109.765 175.205 110.325 175.495 ;
        RECT 110.495 176.715 110.770 177.415 ;
        RECT 110.940 177.040 111.195 177.585 ;
        RECT 111.365 177.075 111.845 177.415 ;
        RECT 112.020 177.030 112.625 177.585 ;
        RECT 112.010 176.930 112.625 177.030 ;
        RECT 112.010 176.905 112.195 176.930 ;
        RECT 110.495 175.685 110.665 176.715 ;
        RECT 110.940 176.585 111.695 176.835 ;
        RECT 111.865 176.660 112.195 176.905 ;
        RECT 110.940 176.550 111.710 176.585 ;
        RECT 110.940 176.540 111.725 176.550 ;
        RECT 110.835 176.525 111.730 176.540 ;
        RECT 110.835 176.510 111.750 176.525 ;
        RECT 110.835 176.500 111.770 176.510 ;
        RECT 110.835 176.490 111.795 176.500 ;
        RECT 110.835 176.460 111.865 176.490 ;
        RECT 110.835 176.430 111.885 176.460 ;
        RECT 110.835 176.400 111.905 176.430 ;
        RECT 110.835 176.375 111.935 176.400 ;
        RECT 110.835 176.340 111.970 176.375 ;
        RECT 110.835 176.335 112.000 176.340 ;
        RECT 110.835 175.940 111.065 176.335 ;
        RECT 111.610 176.330 112.000 176.335 ;
        RECT 111.635 176.320 112.000 176.330 ;
        RECT 111.650 176.315 112.000 176.320 ;
        RECT 111.665 176.310 112.000 176.315 ;
        RECT 112.365 176.310 112.625 176.760 ;
        RECT 112.795 176.495 114.005 177.585 ;
        RECT 111.665 176.305 112.625 176.310 ;
        RECT 111.675 176.295 112.625 176.305 ;
        RECT 111.685 176.290 112.625 176.295 ;
        RECT 111.695 176.280 112.625 176.290 ;
        RECT 111.700 176.270 112.625 176.280 ;
        RECT 111.705 176.265 112.625 176.270 ;
        RECT 111.715 176.250 112.625 176.265 ;
        RECT 111.720 176.235 112.625 176.250 ;
        RECT 111.730 176.210 112.625 176.235 ;
        RECT 111.235 175.740 111.565 176.165 ;
        RECT 111.315 175.715 111.565 175.740 ;
        RECT 110.495 175.205 110.755 175.685 ;
        RECT 110.925 175.035 111.175 175.575 ;
        RECT 111.345 175.255 111.565 175.715 ;
        RECT 111.735 176.140 112.625 176.210 ;
        RECT 111.735 175.415 111.905 176.140 ;
        RECT 112.075 175.585 112.625 175.970 ;
        RECT 112.795 175.785 113.315 176.325 ;
        RECT 113.485 175.955 114.005 176.495 ;
        RECT 114.175 176.495 115.385 177.585 ;
        RECT 114.175 175.955 114.695 176.495 ;
        RECT 114.865 175.785 115.385 176.325 ;
        RECT 111.735 175.245 112.625 175.415 ;
        RECT 112.795 175.035 114.005 175.785 ;
        RECT 114.175 175.035 115.385 175.785 ;
        RECT 61.190 174.865 115.470 175.035 ;
        RECT 61.275 174.115 62.485 174.865 ;
        RECT 62.655 174.320 68.000 174.865 ;
        RECT 68.175 174.320 73.520 174.865 ;
        RECT 73.695 174.320 79.040 174.865 ;
        RECT 79.215 174.320 84.560 174.865 ;
        RECT 61.275 173.575 61.795 174.115 ;
        RECT 61.965 173.405 62.485 173.945 ;
        RECT 64.240 173.490 64.580 174.320 ;
        RECT 61.275 172.315 62.485 173.405 ;
        RECT 66.060 172.750 66.410 174.000 ;
        RECT 69.760 173.490 70.100 174.320 ;
        RECT 71.580 172.750 71.930 174.000 ;
        RECT 75.280 173.490 75.620 174.320 ;
        RECT 77.100 172.750 77.450 174.000 ;
        RECT 80.800 173.490 81.140 174.320 ;
        RECT 84.735 174.095 86.405 174.865 ;
        RECT 87.035 174.140 87.325 174.865 ;
        RECT 87.495 174.320 92.840 174.865 ;
        RECT 93.015 174.320 98.360 174.865 ;
        RECT 98.535 174.320 103.880 174.865 ;
        RECT 104.055 174.320 109.400 174.865 ;
        RECT 82.620 172.750 82.970 174.000 ;
        RECT 84.735 173.575 85.485 174.095 ;
        RECT 85.655 173.405 86.405 173.925 ;
        RECT 89.080 173.490 89.420 174.320 ;
        RECT 62.655 172.315 68.000 172.750 ;
        RECT 68.175 172.315 73.520 172.750 ;
        RECT 73.695 172.315 79.040 172.750 ;
        RECT 79.215 172.315 84.560 172.750 ;
        RECT 84.735 172.315 86.405 173.405 ;
        RECT 87.035 172.315 87.325 173.480 ;
        RECT 90.900 172.750 91.250 174.000 ;
        RECT 94.600 173.490 94.940 174.320 ;
        RECT 96.420 172.750 96.770 174.000 ;
        RECT 100.120 173.490 100.460 174.320 ;
        RECT 101.940 172.750 102.290 174.000 ;
        RECT 105.640 173.490 105.980 174.320 ;
        RECT 109.575 174.115 110.785 174.865 ;
        RECT 111.025 174.465 111.355 174.865 ;
        RECT 111.525 174.295 111.695 174.565 ;
        RECT 111.865 174.465 112.195 174.865 ;
        RECT 112.365 174.295 112.620 174.565 ;
        RECT 107.460 172.750 107.810 174.000 ;
        RECT 109.575 173.575 110.095 174.115 ;
        RECT 110.265 173.405 110.785 173.945 ;
        RECT 87.495 172.315 92.840 172.750 ;
        RECT 93.015 172.315 98.360 172.750 ;
        RECT 98.535 172.315 103.880 172.750 ;
        RECT 104.055 172.315 109.400 172.750 ;
        RECT 109.575 172.315 110.785 173.405 ;
        RECT 110.955 173.285 111.225 174.295 ;
        RECT 111.395 174.125 112.620 174.295 ;
        RECT 112.795 174.140 113.085 174.865 ;
        RECT 111.395 173.455 111.565 174.125 ;
        RECT 114.175 174.115 115.385 174.865 ;
        RECT 111.735 173.625 112.115 173.955 ;
        RECT 112.285 173.625 112.620 173.955 ;
        RECT 111.395 173.285 111.710 173.455 ;
        RECT 110.960 172.315 111.275 173.115 ;
        RECT 111.540 172.670 111.710 173.285 ;
        RECT 111.880 172.945 112.115 173.625 ;
        RECT 112.285 172.670 112.620 173.455 ;
        RECT 111.540 172.500 112.620 172.670 ;
        RECT 112.795 172.315 113.085 173.480 ;
        RECT 114.175 173.405 114.695 173.945 ;
        RECT 114.865 173.575 115.385 174.115 ;
        RECT 114.175 172.315 115.385 173.405 ;
        RECT 61.190 172.145 115.470 172.315 ;
        RECT 61.275 171.055 62.485 172.145 ;
        RECT 62.655 171.710 68.000 172.145 ;
        RECT 68.175 171.710 73.520 172.145 ;
        RECT 61.275 170.345 61.795 170.885 ;
        RECT 61.965 170.515 62.485 171.055 ;
        RECT 61.275 169.595 62.485 170.345 ;
        RECT 64.240 170.140 64.580 170.970 ;
        RECT 66.060 170.460 66.410 171.710 ;
        RECT 69.760 170.140 70.100 170.970 ;
        RECT 71.580 170.460 71.930 171.710 ;
        RECT 74.155 170.980 74.445 172.145 ;
        RECT 74.615 171.710 79.960 172.145 ;
        RECT 80.135 171.710 85.480 172.145 ;
        RECT 85.655 171.710 91.000 172.145 ;
        RECT 91.175 171.710 96.520 172.145 ;
        RECT 62.655 169.595 68.000 170.140 ;
        RECT 68.175 169.595 73.520 170.140 ;
        RECT 74.155 169.595 74.445 170.320 ;
        RECT 76.200 170.140 76.540 170.970 ;
        RECT 78.020 170.460 78.370 171.710 ;
        RECT 81.720 170.140 82.060 170.970 ;
        RECT 83.540 170.460 83.890 171.710 ;
        RECT 87.240 170.140 87.580 170.970 ;
        RECT 89.060 170.460 89.410 171.710 ;
        RECT 92.760 170.140 93.100 170.970 ;
        RECT 94.580 170.460 94.930 171.710 ;
        RECT 96.695 171.055 99.285 172.145 ;
        RECT 96.695 170.365 97.905 170.885 ;
        RECT 98.075 170.535 99.285 171.055 ;
        RECT 99.915 170.980 100.205 172.145 ;
        RECT 100.375 171.710 105.720 172.145 ;
        RECT 105.895 171.710 111.240 172.145 ;
        RECT 74.615 169.595 79.960 170.140 ;
        RECT 80.135 169.595 85.480 170.140 ;
        RECT 85.655 169.595 91.000 170.140 ;
        RECT 91.175 169.595 96.520 170.140 ;
        RECT 96.695 169.595 99.285 170.365 ;
        RECT 99.915 169.595 100.205 170.320 ;
        RECT 101.960 170.140 102.300 170.970 ;
        RECT 103.780 170.460 104.130 171.710 ;
        RECT 107.480 170.140 107.820 170.970 ;
        RECT 109.300 170.460 109.650 171.710 ;
        RECT 111.415 171.055 114.005 172.145 ;
        RECT 111.415 170.365 112.625 170.885 ;
        RECT 112.795 170.535 114.005 171.055 ;
        RECT 114.175 171.055 115.385 172.145 ;
        RECT 114.175 170.515 114.695 171.055 ;
        RECT 100.375 169.595 105.720 170.140 ;
        RECT 105.895 169.595 111.240 170.140 ;
        RECT 111.415 169.595 114.005 170.365 ;
        RECT 114.865 170.345 115.385 170.885 ;
        RECT 114.175 169.595 115.385 170.345 ;
        RECT 61.190 169.425 115.470 169.595 ;
        RECT 61.275 168.675 62.485 169.425 ;
        RECT 62.655 168.880 68.000 169.425 ;
        RECT 68.175 168.880 73.520 169.425 ;
        RECT 73.695 168.880 79.040 169.425 ;
        RECT 79.215 168.880 84.560 169.425 ;
        RECT 61.275 168.135 61.795 168.675 ;
        RECT 61.965 167.965 62.485 168.505 ;
        RECT 64.240 168.050 64.580 168.880 ;
        RECT 61.275 166.875 62.485 167.965 ;
        RECT 66.060 167.310 66.410 168.560 ;
        RECT 69.760 168.050 70.100 168.880 ;
        RECT 71.580 167.310 71.930 168.560 ;
        RECT 75.280 168.050 75.620 168.880 ;
        RECT 77.100 167.310 77.450 168.560 ;
        RECT 80.800 168.050 81.140 168.880 ;
        RECT 84.735 168.655 86.405 169.425 ;
        RECT 87.035 168.700 87.325 169.425 ;
        RECT 87.495 168.880 92.840 169.425 ;
        RECT 93.015 168.880 98.360 169.425 ;
        RECT 98.535 168.880 103.880 169.425 ;
        RECT 104.055 168.880 109.400 169.425 ;
        RECT 82.620 167.310 82.970 168.560 ;
        RECT 84.735 168.135 85.485 168.655 ;
        RECT 85.655 167.965 86.405 168.485 ;
        RECT 89.080 168.050 89.420 168.880 ;
        RECT 62.655 166.875 68.000 167.310 ;
        RECT 68.175 166.875 73.520 167.310 ;
        RECT 73.695 166.875 79.040 167.310 ;
        RECT 79.215 166.875 84.560 167.310 ;
        RECT 84.735 166.875 86.405 167.965 ;
        RECT 87.035 166.875 87.325 168.040 ;
        RECT 90.900 167.310 91.250 168.560 ;
        RECT 94.600 168.050 94.940 168.880 ;
        RECT 96.420 167.310 96.770 168.560 ;
        RECT 100.120 168.050 100.460 168.880 ;
        RECT 101.940 167.310 102.290 168.560 ;
        RECT 105.640 168.050 105.980 168.880 ;
        RECT 109.575 168.655 112.165 169.425 ;
        RECT 112.795 168.700 113.085 169.425 ;
        RECT 114.175 168.675 115.385 169.425 ;
        RECT 107.460 167.310 107.810 168.560 ;
        RECT 109.575 168.135 110.785 168.655 ;
        RECT 110.955 167.965 112.165 168.485 ;
        RECT 87.495 166.875 92.840 167.310 ;
        RECT 93.015 166.875 98.360 167.310 ;
        RECT 98.535 166.875 103.880 167.310 ;
        RECT 104.055 166.875 109.400 167.310 ;
        RECT 109.575 166.875 112.165 167.965 ;
        RECT 112.795 166.875 113.085 168.040 ;
        RECT 114.175 167.965 114.695 168.505 ;
        RECT 114.865 168.135 115.385 168.675 ;
        RECT 114.175 166.875 115.385 167.965 ;
        RECT 61.190 166.705 115.470 166.875 ;
        RECT 61.275 165.615 62.485 166.705 ;
        RECT 62.655 166.270 68.000 166.705 ;
        RECT 68.175 166.270 73.520 166.705 ;
        RECT 61.275 164.905 61.795 165.445 ;
        RECT 61.965 165.075 62.485 165.615 ;
        RECT 61.275 164.155 62.485 164.905 ;
        RECT 64.240 164.700 64.580 165.530 ;
        RECT 66.060 165.020 66.410 166.270 ;
        RECT 69.760 164.700 70.100 165.530 ;
        RECT 71.580 165.020 71.930 166.270 ;
        RECT 74.155 165.540 74.445 166.705 ;
        RECT 74.615 166.270 79.960 166.705 ;
        RECT 80.135 166.270 85.480 166.705 ;
        RECT 85.655 166.270 91.000 166.705 ;
        RECT 91.175 166.270 96.520 166.705 ;
        RECT 62.655 164.155 68.000 164.700 ;
        RECT 68.175 164.155 73.520 164.700 ;
        RECT 74.155 164.155 74.445 164.880 ;
        RECT 76.200 164.700 76.540 165.530 ;
        RECT 78.020 165.020 78.370 166.270 ;
        RECT 81.720 164.700 82.060 165.530 ;
        RECT 83.540 165.020 83.890 166.270 ;
        RECT 87.240 164.700 87.580 165.530 ;
        RECT 89.060 165.020 89.410 166.270 ;
        RECT 92.760 164.700 93.100 165.530 ;
        RECT 94.580 165.020 94.930 166.270 ;
        RECT 96.695 165.615 99.285 166.705 ;
        RECT 96.695 164.925 97.905 165.445 ;
        RECT 98.075 165.095 99.285 165.615 ;
        RECT 99.915 165.540 100.205 166.705 ;
        RECT 100.375 166.270 105.720 166.705 ;
        RECT 105.895 166.270 111.240 166.705 ;
        RECT 74.615 164.155 79.960 164.700 ;
        RECT 80.135 164.155 85.480 164.700 ;
        RECT 85.655 164.155 91.000 164.700 ;
        RECT 91.175 164.155 96.520 164.700 ;
        RECT 96.695 164.155 99.285 164.925 ;
        RECT 99.915 164.155 100.205 164.880 ;
        RECT 101.960 164.700 102.300 165.530 ;
        RECT 103.780 165.020 104.130 166.270 ;
        RECT 107.480 164.700 107.820 165.530 ;
        RECT 109.300 165.020 109.650 166.270 ;
        RECT 111.415 165.615 114.005 166.705 ;
        RECT 111.415 164.925 112.625 165.445 ;
        RECT 112.795 165.095 114.005 165.615 ;
        RECT 114.175 165.615 115.385 166.705 ;
        RECT 114.175 165.075 114.695 165.615 ;
        RECT 100.375 164.155 105.720 164.700 ;
        RECT 105.895 164.155 111.240 164.700 ;
        RECT 111.415 164.155 114.005 164.925 ;
        RECT 114.865 164.905 115.385 165.445 ;
        RECT 114.175 164.155 115.385 164.905 ;
        RECT 61.190 163.985 115.470 164.155 ;
        RECT 61.275 163.235 62.485 163.985 ;
        RECT 62.655 163.440 68.000 163.985 ;
        RECT 68.175 163.440 73.520 163.985 ;
        RECT 73.695 163.440 79.040 163.985 ;
        RECT 79.215 163.440 84.560 163.985 ;
        RECT 61.275 162.695 61.795 163.235 ;
        RECT 61.965 162.525 62.485 163.065 ;
        RECT 64.240 162.610 64.580 163.440 ;
        RECT 61.275 161.435 62.485 162.525 ;
        RECT 66.060 161.870 66.410 163.120 ;
        RECT 69.760 162.610 70.100 163.440 ;
        RECT 71.580 161.870 71.930 163.120 ;
        RECT 75.280 162.610 75.620 163.440 ;
        RECT 77.100 161.870 77.450 163.120 ;
        RECT 80.800 162.610 81.140 163.440 ;
        RECT 84.735 163.215 86.405 163.985 ;
        RECT 87.035 163.260 87.325 163.985 ;
        RECT 87.495 163.440 92.840 163.985 ;
        RECT 93.015 163.440 98.360 163.985 ;
        RECT 98.535 163.440 103.880 163.985 ;
        RECT 104.055 163.440 109.400 163.985 ;
        RECT 82.620 161.870 82.970 163.120 ;
        RECT 84.735 162.695 85.485 163.215 ;
        RECT 85.655 162.525 86.405 163.045 ;
        RECT 89.080 162.610 89.420 163.440 ;
        RECT 62.655 161.435 68.000 161.870 ;
        RECT 68.175 161.435 73.520 161.870 ;
        RECT 73.695 161.435 79.040 161.870 ;
        RECT 79.215 161.435 84.560 161.870 ;
        RECT 84.735 161.435 86.405 162.525 ;
        RECT 87.035 161.435 87.325 162.600 ;
        RECT 90.900 161.870 91.250 163.120 ;
        RECT 94.600 162.610 94.940 163.440 ;
        RECT 96.420 161.870 96.770 163.120 ;
        RECT 100.120 162.610 100.460 163.440 ;
        RECT 101.940 161.870 102.290 163.120 ;
        RECT 105.640 162.610 105.980 163.440 ;
        RECT 109.575 163.215 112.165 163.985 ;
        RECT 112.795 163.260 113.085 163.985 ;
        RECT 114.175 163.235 115.385 163.985 ;
        RECT 107.460 161.870 107.810 163.120 ;
        RECT 109.575 162.695 110.785 163.215 ;
        RECT 110.955 162.525 112.165 163.045 ;
        RECT 87.495 161.435 92.840 161.870 ;
        RECT 93.015 161.435 98.360 161.870 ;
        RECT 98.535 161.435 103.880 161.870 ;
        RECT 104.055 161.435 109.400 161.870 ;
        RECT 109.575 161.435 112.165 162.525 ;
        RECT 112.795 161.435 113.085 162.600 ;
        RECT 114.175 162.525 114.695 163.065 ;
        RECT 114.865 162.695 115.385 163.235 ;
        RECT 114.175 161.435 115.385 162.525 ;
        RECT 61.190 161.265 115.470 161.435 ;
        RECT 61.275 160.175 62.485 161.265 ;
        RECT 62.655 160.830 68.000 161.265 ;
        RECT 68.175 160.830 73.520 161.265 ;
        RECT 61.275 159.465 61.795 160.005 ;
        RECT 61.965 159.635 62.485 160.175 ;
        RECT 61.275 158.715 62.485 159.465 ;
        RECT 64.240 159.260 64.580 160.090 ;
        RECT 66.060 159.580 66.410 160.830 ;
        RECT 69.760 159.260 70.100 160.090 ;
        RECT 71.580 159.580 71.930 160.830 ;
        RECT 74.155 160.100 74.445 161.265 ;
        RECT 74.615 160.830 79.960 161.265 ;
        RECT 80.135 160.830 85.480 161.265 ;
        RECT 85.655 160.830 91.000 161.265 ;
        RECT 91.175 160.830 96.520 161.265 ;
        RECT 62.655 158.715 68.000 159.260 ;
        RECT 68.175 158.715 73.520 159.260 ;
        RECT 74.155 158.715 74.445 159.440 ;
        RECT 76.200 159.260 76.540 160.090 ;
        RECT 78.020 159.580 78.370 160.830 ;
        RECT 81.720 159.260 82.060 160.090 ;
        RECT 83.540 159.580 83.890 160.830 ;
        RECT 87.240 159.260 87.580 160.090 ;
        RECT 89.060 159.580 89.410 160.830 ;
        RECT 92.760 159.260 93.100 160.090 ;
        RECT 94.580 159.580 94.930 160.830 ;
        RECT 96.695 160.175 99.285 161.265 ;
        RECT 96.695 159.485 97.905 160.005 ;
        RECT 98.075 159.655 99.285 160.175 ;
        RECT 99.915 160.100 100.205 161.265 ;
        RECT 100.375 160.830 105.720 161.265 ;
        RECT 105.895 160.830 111.240 161.265 ;
        RECT 74.615 158.715 79.960 159.260 ;
        RECT 80.135 158.715 85.480 159.260 ;
        RECT 85.655 158.715 91.000 159.260 ;
        RECT 91.175 158.715 96.520 159.260 ;
        RECT 96.695 158.715 99.285 159.485 ;
        RECT 99.915 158.715 100.205 159.440 ;
        RECT 101.960 159.260 102.300 160.090 ;
        RECT 103.780 159.580 104.130 160.830 ;
        RECT 107.480 159.260 107.820 160.090 ;
        RECT 109.300 159.580 109.650 160.830 ;
        RECT 111.415 160.175 114.005 161.265 ;
        RECT 111.415 159.485 112.625 160.005 ;
        RECT 112.795 159.655 114.005 160.175 ;
        RECT 114.175 160.175 115.385 161.265 ;
        RECT 114.175 159.635 114.695 160.175 ;
        RECT 100.375 158.715 105.720 159.260 ;
        RECT 105.895 158.715 111.240 159.260 ;
        RECT 111.415 158.715 114.005 159.485 ;
        RECT 114.865 159.465 115.385 160.005 ;
        RECT 114.175 158.715 115.385 159.465 ;
        RECT 61.190 158.545 115.470 158.715 ;
        RECT 61.275 157.795 62.485 158.545 ;
        RECT 62.655 158.000 68.000 158.545 ;
        RECT 68.175 158.000 73.520 158.545 ;
        RECT 73.695 158.000 79.040 158.545 ;
        RECT 79.215 158.000 84.560 158.545 ;
        RECT 61.275 157.255 61.795 157.795 ;
        RECT 61.965 157.085 62.485 157.625 ;
        RECT 64.240 157.170 64.580 158.000 ;
        RECT 61.275 155.995 62.485 157.085 ;
        RECT 66.060 156.430 66.410 157.680 ;
        RECT 69.760 157.170 70.100 158.000 ;
        RECT 71.580 156.430 71.930 157.680 ;
        RECT 75.280 157.170 75.620 158.000 ;
        RECT 77.100 156.430 77.450 157.680 ;
        RECT 80.800 157.170 81.140 158.000 ;
        RECT 84.735 157.775 86.405 158.545 ;
        RECT 87.035 157.820 87.325 158.545 ;
        RECT 87.495 158.000 92.840 158.545 ;
        RECT 93.015 158.000 98.360 158.545 ;
        RECT 98.535 158.000 103.880 158.545 ;
        RECT 104.055 158.000 109.400 158.545 ;
        RECT 82.620 156.430 82.970 157.680 ;
        RECT 84.735 157.255 85.485 157.775 ;
        RECT 85.655 157.085 86.405 157.605 ;
        RECT 89.080 157.170 89.420 158.000 ;
        RECT 62.655 155.995 68.000 156.430 ;
        RECT 68.175 155.995 73.520 156.430 ;
        RECT 73.695 155.995 79.040 156.430 ;
        RECT 79.215 155.995 84.560 156.430 ;
        RECT 84.735 155.995 86.405 157.085 ;
        RECT 87.035 155.995 87.325 157.160 ;
        RECT 90.900 156.430 91.250 157.680 ;
        RECT 94.600 157.170 94.940 158.000 ;
        RECT 96.420 156.430 96.770 157.680 ;
        RECT 100.120 157.170 100.460 158.000 ;
        RECT 101.940 156.430 102.290 157.680 ;
        RECT 105.640 157.170 105.980 158.000 ;
        RECT 109.575 157.775 112.165 158.545 ;
        RECT 112.795 157.820 113.085 158.545 ;
        RECT 114.175 157.795 115.385 158.545 ;
        RECT 107.460 156.430 107.810 157.680 ;
        RECT 109.575 157.255 110.785 157.775 ;
        RECT 110.955 157.085 112.165 157.605 ;
        RECT 87.495 155.995 92.840 156.430 ;
        RECT 93.015 155.995 98.360 156.430 ;
        RECT 98.535 155.995 103.880 156.430 ;
        RECT 104.055 155.995 109.400 156.430 ;
        RECT 109.575 155.995 112.165 157.085 ;
        RECT 112.795 155.995 113.085 157.160 ;
        RECT 114.175 157.085 114.695 157.625 ;
        RECT 114.865 157.255 115.385 157.795 ;
        RECT 114.175 155.995 115.385 157.085 ;
        RECT 61.190 155.825 115.470 155.995 ;
        RECT 61.275 154.735 62.485 155.825 ;
        RECT 62.655 155.390 68.000 155.825 ;
        RECT 68.175 155.390 73.520 155.825 ;
        RECT 61.275 154.025 61.795 154.565 ;
        RECT 61.965 154.195 62.485 154.735 ;
        RECT 61.275 153.275 62.485 154.025 ;
        RECT 64.240 153.820 64.580 154.650 ;
        RECT 66.060 154.140 66.410 155.390 ;
        RECT 69.760 153.820 70.100 154.650 ;
        RECT 71.580 154.140 71.930 155.390 ;
        RECT 74.155 154.660 74.445 155.825 ;
        RECT 74.615 155.390 79.960 155.825 ;
        RECT 80.135 155.390 85.480 155.825 ;
        RECT 62.655 153.275 68.000 153.820 ;
        RECT 68.175 153.275 73.520 153.820 ;
        RECT 74.155 153.275 74.445 154.000 ;
        RECT 76.200 153.820 76.540 154.650 ;
        RECT 78.020 154.140 78.370 155.390 ;
        RECT 81.720 153.820 82.060 154.650 ;
        RECT 83.540 154.140 83.890 155.390 ;
        RECT 85.655 154.735 86.865 155.825 ;
        RECT 85.655 154.025 86.175 154.565 ;
        RECT 86.345 154.195 86.865 154.735 ;
        RECT 87.035 154.660 87.325 155.825 ;
        RECT 87.495 155.390 92.840 155.825 ;
        RECT 93.015 155.390 98.360 155.825 ;
        RECT 74.615 153.275 79.960 153.820 ;
        RECT 80.135 153.275 85.480 153.820 ;
        RECT 85.655 153.275 86.865 154.025 ;
        RECT 87.035 153.275 87.325 154.000 ;
        RECT 89.080 153.820 89.420 154.650 ;
        RECT 90.900 154.140 91.250 155.390 ;
        RECT 94.600 153.820 94.940 154.650 ;
        RECT 96.420 154.140 96.770 155.390 ;
        RECT 98.535 154.735 99.745 155.825 ;
        RECT 98.535 154.025 99.055 154.565 ;
        RECT 99.225 154.195 99.745 154.735 ;
        RECT 99.915 154.660 100.205 155.825 ;
        RECT 100.375 155.390 105.720 155.825 ;
        RECT 105.895 155.390 111.240 155.825 ;
        RECT 87.495 153.275 92.840 153.820 ;
        RECT 93.015 153.275 98.360 153.820 ;
        RECT 98.535 153.275 99.745 154.025 ;
        RECT 99.915 153.275 100.205 154.000 ;
        RECT 101.960 153.820 102.300 154.650 ;
        RECT 103.780 154.140 104.130 155.390 ;
        RECT 107.480 153.820 107.820 154.650 ;
        RECT 109.300 154.140 109.650 155.390 ;
        RECT 111.415 154.735 112.625 155.825 ;
        RECT 111.415 154.025 111.935 154.565 ;
        RECT 112.105 154.195 112.625 154.735 ;
        RECT 112.795 154.660 113.085 155.825 ;
        RECT 114.175 154.735 115.385 155.825 ;
        RECT 114.175 154.195 114.695 154.735 ;
        RECT 114.865 154.025 115.385 154.565 ;
        RECT 100.375 153.275 105.720 153.820 ;
        RECT 105.895 153.275 111.240 153.820 ;
        RECT 111.415 153.275 112.625 154.025 ;
        RECT 112.795 153.275 113.085 154.000 ;
        RECT 114.175 153.275 115.385 154.025 ;
        RECT 61.190 153.105 115.470 153.275 ;
        RECT 130.980 99.360 143.080 99.530 ;
        RECT 130.980 94.730 131.150 99.360 ;
        RECT 131.630 98.530 133.790 98.880 ;
        RECT 140.270 95.210 142.430 95.560 ;
        RECT 142.910 94.730 143.080 99.360 ;
        RECT 130.980 94.560 143.080 94.730 ;
        RECT 112.120 93.070 124.220 93.240 ;
        RECT 112.120 88.440 112.290 93.070 ;
        RECT 112.770 92.240 114.930 92.590 ;
        RECT 121.410 88.920 123.570 89.270 ;
        RECT 124.050 88.440 124.220 93.070 ;
        RECT 112.120 88.270 124.220 88.440 ;
        RECT 106.000 83.700 108.290 86.550 ;
        RECT 114.740 49.670 143.360 49.840 ;
        RECT 114.740 48.360 114.910 49.670 ;
        RECT 115.390 48.840 117.550 49.190 ;
        RECT 140.550 48.840 142.710 49.190 ;
        RECT 143.190 48.360 143.360 49.670 ;
        RECT 114.740 48.190 143.360 48.360 ;
        RECT 142.020 43.730 144.850 43.900 ;
        RECT 131.070 43.470 133.900 43.640 ;
        RECT 131.070 43.110 131.240 43.470 ;
        RECT 127.020 42.540 128.670 42.710 ;
        RECT 127.020 42.410 127.190 42.540 ;
        RECT 119.120 41.490 120.770 41.660 ;
        RECT 115.070 41.290 116.720 41.460 ;
        RECT 115.070 16.010 115.240 41.290 ;
        RECT 115.720 38.650 116.070 40.810 ;
        RECT 115.720 16.490 116.070 18.650 ;
        RECT 116.550 16.010 116.720 41.290 ;
        RECT 119.120 16.210 119.290 41.490 ;
        RECT 119.770 38.850 120.120 41.010 ;
        RECT 119.770 16.690 120.120 18.850 ;
        RECT 120.600 16.210 120.770 41.490 ;
        RECT 125.190 34.360 127.190 42.410 ;
        RECT 127.670 39.900 128.020 42.060 ;
        RECT 127.670 34.840 128.020 37.000 ;
        RECT 128.500 34.360 128.670 42.540 ;
        RECT 125.190 34.190 128.670 34.360 ;
        RECT 125.190 33.010 128.340 34.190 ;
        RECT 125.190 32.840 129.210 33.010 ;
        RECT 125.190 22.710 126.640 32.840 ;
        RECT 127.320 32.270 128.360 32.440 ;
        RECT 126.980 30.210 127.150 32.210 ;
        RECT 128.530 30.210 128.700 32.210 ;
        RECT 127.320 29.980 128.360 30.150 ;
        RECT 126.980 27.920 127.150 29.920 ;
        RECT 128.530 27.920 128.700 29.920 ;
        RECT 127.320 27.690 128.360 27.860 ;
        RECT 126.980 25.630 127.150 27.630 ;
        RECT 128.530 25.630 128.700 27.630 ;
        RECT 127.320 25.400 128.360 25.570 ;
        RECT 126.980 23.340 127.150 25.340 ;
        RECT 128.530 23.340 128.700 25.340 ;
        RECT 129.040 25.010 129.210 32.840 ;
        RECT 130.940 31.210 131.240 43.110 ;
        RECT 131.965 42.900 133.005 43.070 ;
        RECT 131.580 40.840 131.750 42.840 ;
        RECT 133.220 40.840 133.390 42.840 ;
        RECT 131.965 40.610 133.005 40.780 ;
        RECT 131.580 38.550 131.750 40.550 ;
        RECT 133.220 38.550 133.390 40.550 ;
        RECT 131.965 38.320 133.005 38.490 ;
        RECT 131.580 36.260 131.750 38.260 ;
        RECT 133.220 36.260 133.390 38.260 ;
        RECT 131.965 36.030 133.005 36.200 ;
        RECT 131.580 33.970 131.750 35.970 ;
        RECT 133.220 33.970 133.390 35.970 ;
        RECT 131.965 33.740 133.005 33.910 ;
        RECT 131.580 31.680 131.750 33.680 ;
        RECT 133.220 31.680 133.390 33.680 ;
        RECT 131.965 31.450 133.005 31.620 ;
        RECT 131.070 28.760 131.240 31.210 ;
        RECT 131.580 29.390 131.750 31.390 ;
        RECT 133.220 29.390 133.390 31.390 ;
        RECT 131.965 29.160 133.005 29.330 ;
        RECT 133.730 28.760 133.900 43.470 ;
        RECT 131.070 28.590 133.900 28.760 ;
        RECT 137.420 43.470 140.250 43.640 ;
        RECT 137.420 28.760 137.590 43.470 ;
        RECT 140.080 43.110 140.250 43.470 ;
        RECT 142.020 43.360 142.190 43.730 ;
        RECT 138.315 42.900 139.355 43.070 ;
        RECT 137.930 40.840 138.100 42.840 ;
        RECT 139.570 40.840 139.740 42.840 ;
        RECT 138.315 40.610 139.355 40.780 ;
        RECT 137.930 38.550 138.100 40.550 ;
        RECT 139.570 38.550 139.740 40.550 ;
        RECT 138.315 38.320 139.355 38.490 ;
        RECT 137.930 36.260 138.100 38.260 ;
        RECT 139.570 36.260 139.740 38.260 ;
        RECT 138.315 36.030 139.355 36.200 ;
        RECT 137.930 33.970 138.100 35.970 ;
        RECT 139.570 33.970 139.740 35.970 ;
        RECT 138.315 33.740 139.355 33.910 ;
        RECT 137.930 31.680 138.100 33.680 ;
        RECT 139.570 31.680 139.740 33.680 ;
        RECT 138.315 31.450 139.355 31.620 ;
        RECT 137.930 29.390 138.100 31.390 ;
        RECT 139.570 29.390 139.740 31.390 ;
        RECT 140.080 31.210 140.390 43.110 ;
        RECT 138.315 29.160 139.355 29.330 ;
        RECT 140.080 28.760 140.250 31.210 ;
        RECT 137.420 28.590 140.250 28.760 ;
        RECT 131.220 27.670 135.460 27.840 ;
        RECT 131.220 25.910 131.390 27.670 ;
        RECT 132.070 27.100 134.610 27.270 ;
        RECT 131.730 26.540 131.900 27.040 ;
        RECT 134.780 26.540 134.950 27.040 ;
        RECT 132.070 26.310 134.610 26.480 ;
        RECT 135.290 25.910 135.460 27.670 ;
        RECT 131.220 25.740 135.460 25.910 ;
        RECT 135.820 27.670 140.060 27.840 ;
        RECT 141.990 27.810 142.190 43.360 ;
        RECT 142.915 43.160 143.955 43.330 ;
        RECT 142.530 42.600 142.700 43.100 ;
        RECT 144.170 42.600 144.340 43.100 ;
        RECT 142.915 42.370 143.955 42.540 ;
        RECT 142.530 41.810 142.700 42.310 ;
        RECT 144.170 41.810 144.340 42.310 ;
        RECT 142.915 41.580 143.955 41.750 ;
        RECT 142.530 41.020 142.700 41.520 ;
        RECT 144.170 41.020 144.340 41.520 ;
        RECT 142.915 40.790 143.955 40.960 ;
        RECT 142.530 40.230 142.700 40.730 ;
        RECT 144.170 40.230 144.340 40.730 ;
        RECT 142.915 40.000 143.955 40.170 ;
        RECT 142.530 39.440 142.700 39.940 ;
        RECT 144.170 39.440 144.340 39.940 ;
        RECT 142.915 39.210 143.955 39.380 ;
        RECT 142.530 38.650 142.700 39.150 ;
        RECT 144.170 38.650 144.340 39.150 ;
        RECT 142.915 38.420 143.955 38.590 ;
        RECT 142.530 37.860 142.700 38.360 ;
        RECT 144.170 37.860 144.340 38.360 ;
        RECT 142.915 37.630 143.955 37.800 ;
        RECT 142.530 37.070 142.700 37.570 ;
        RECT 144.170 37.070 144.340 37.570 ;
        RECT 142.915 36.840 143.955 37.010 ;
        RECT 142.530 36.280 142.700 36.780 ;
        RECT 144.170 36.280 144.340 36.780 ;
        RECT 142.915 36.050 143.955 36.220 ;
        RECT 142.530 35.490 142.700 35.990 ;
        RECT 144.170 35.490 144.340 35.990 ;
        RECT 142.915 35.260 143.955 35.430 ;
        RECT 142.530 34.700 142.700 35.200 ;
        RECT 144.170 34.700 144.340 35.200 ;
        RECT 142.915 34.470 143.955 34.640 ;
        RECT 142.530 33.910 142.700 34.410 ;
        RECT 144.170 33.910 144.340 34.410 ;
        RECT 142.915 33.680 143.955 33.850 ;
        RECT 142.530 33.120 142.700 33.620 ;
        RECT 144.170 33.120 144.340 33.620 ;
        RECT 142.915 32.890 143.955 33.060 ;
        RECT 142.530 32.330 142.700 32.830 ;
        RECT 144.170 32.330 144.340 32.830 ;
        RECT 142.915 32.100 143.955 32.270 ;
        RECT 142.530 31.540 142.700 32.040 ;
        RECT 144.170 31.540 144.340 32.040 ;
        RECT 142.915 31.310 143.955 31.480 ;
        RECT 142.530 30.750 142.700 31.250 ;
        RECT 144.170 30.750 144.340 31.250 ;
        RECT 142.915 30.520 143.955 30.690 ;
        RECT 142.530 29.960 142.700 30.460 ;
        RECT 144.170 29.960 144.340 30.460 ;
        RECT 142.915 29.730 143.955 29.900 ;
        RECT 142.530 29.170 142.700 29.670 ;
        RECT 144.170 29.170 144.340 29.670 ;
        RECT 142.915 28.940 143.955 29.110 ;
        RECT 142.530 28.380 142.700 28.880 ;
        RECT 144.170 28.380 144.340 28.880 ;
        RECT 142.915 28.150 143.955 28.320 ;
        RECT 135.820 25.910 135.990 27.670 ;
        RECT 136.670 27.100 139.210 27.270 ;
        RECT 136.330 26.540 136.500 27.040 ;
        RECT 139.380 26.540 139.550 27.040 ;
        RECT 136.670 26.310 139.210 26.480 ;
        RECT 139.890 25.910 140.060 27.670 ;
        RECT 142.020 26.960 142.190 27.810 ;
        RECT 142.530 27.590 142.700 28.090 ;
        RECT 144.170 27.590 144.340 28.090 ;
        RECT 142.915 27.360 143.955 27.530 ;
        RECT 144.680 26.960 144.850 43.730 ;
        RECT 142.020 26.790 144.850 26.960 ;
        RECT 146.020 39.760 148.760 39.930 ;
        RECT 135.820 25.740 140.190 25.910 ;
        RECT 131.240 25.710 132.040 25.740 ;
        RECT 139.390 25.710 140.190 25.740 ;
        RECT 130.520 25.260 140.990 25.330 ;
        RECT 146.020 25.260 146.190 39.760 ;
        RECT 146.870 39.190 147.910 39.360 ;
        RECT 146.530 37.130 146.700 39.130 ;
        RECT 148.080 37.130 148.250 39.130 ;
        RECT 146.870 36.900 147.910 37.070 ;
        RECT 148.590 37.060 148.760 39.760 ;
        RECT 146.530 34.840 146.700 36.840 ;
        RECT 148.080 34.840 148.250 36.840 ;
        RECT 146.870 34.610 147.910 34.780 ;
        RECT 146.530 32.550 146.700 34.550 ;
        RECT 148.080 32.550 148.250 34.550 ;
        RECT 146.870 32.320 147.910 32.490 ;
        RECT 146.530 30.260 146.700 32.260 ;
        RECT 148.080 30.260 148.250 32.260 ;
        RECT 146.870 30.030 147.910 30.200 ;
        RECT 146.530 27.970 146.700 29.970 ;
        RECT 148.080 27.970 148.250 29.970 ;
        RECT 146.870 27.740 147.910 27.910 ;
        RECT 146.530 25.680 146.700 27.680 ;
        RECT 148.080 25.680 148.250 27.680 ;
        RECT 146.870 25.450 147.910 25.620 ;
        RECT 130.520 25.160 146.190 25.260 ;
        RECT 130.520 25.010 130.690 25.160 ;
        RECT 127.320 23.110 128.360 23.280 ;
        RECT 129.040 22.760 130.690 25.010 ;
        RECT 131.320 24.650 133.320 24.820 ;
        RECT 133.610 24.650 135.610 24.820 ;
        RECT 135.900 24.650 137.900 24.820 ;
        RECT 138.190 24.650 140.190 24.820 ;
        RECT 140.820 24.660 146.190 25.160 ;
        RECT 131.090 23.440 131.260 24.480 ;
        RECT 133.380 23.440 133.550 24.480 ;
        RECT 135.670 23.440 135.840 24.480 ;
        RECT 137.960 23.440 138.130 24.480 ;
        RECT 140.250 23.440 140.420 24.480 ;
        RECT 131.320 23.100 133.320 23.270 ;
        RECT 133.610 23.100 135.610 23.270 ;
        RECT 135.900 23.100 137.900 23.270 ;
        RECT 138.190 23.100 140.190 23.270 ;
        RECT 140.790 23.060 146.190 24.660 ;
        RECT 146.530 23.390 146.700 25.390 ;
        RECT 148.080 23.390 148.250 25.390 ;
        RECT 146.870 23.160 147.910 23.330 ;
        RECT 140.820 22.760 146.190 23.060 ;
        RECT 148.590 22.760 149.340 37.060 ;
        RECT 126.890 22.710 128.790 22.760 ;
        RECT 129.040 22.710 149.340 22.760 ;
        RECT 125.190 20.510 149.340 22.710 ;
        RECT 119.120 16.040 120.770 16.210 ;
        RECT 115.070 15.840 116.720 16.010 ;
      LAYER mcon ;
        RECT 61.335 207.505 61.505 207.675 ;
        RECT 61.795 207.505 61.965 207.675 ;
        RECT 62.255 207.505 62.425 207.675 ;
        RECT 62.715 207.505 62.885 207.675 ;
        RECT 63.175 207.505 63.345 207.675 ;
        RECT 63.635 207.505 63.805 207.675 ;
        RECT 64.095 207.505 64.265 207.675 ;
        RECT 64.555 207.505 64.725 207.675 ;
        RECT 65.015 207.505 65.185 207.675 ;
        RECT 65.475 207.505 65.645 207.675 ;
        RECT 65.935 207.505 66.105 207.675 ;
        RECT 66.395 207.505 66.565 207.675 ;
        RECT 66.855 207.505 67.025 207.675 ;
        RECT 67.315 207.505 67.485 207.675 ;
        RECT 67.775 207.505 67.945 207.675 ;
        RECT 68.235 207.505 68.405 207.675 ;
        RECT 68.695 207.505 68.865 207.675 ;
        RECT 69.155 207.505 69.325 207.675 ;
        RECT 69.615 207.505 69.785 207.675 ;
        RECT 70.075 207.505 70.245 207.675 ;
        RECT 70.535 207.505 70.705 207.675 ;
        RECT 70.995 207.505 71.165 207.675 ;
        RECT 71.455 207.505 71.625 207.675 ;
        RECT 71.915 207.505 72.085 207.675 ;
        RECT 72.375 207.505 72.545 207.675 ;
        RECT 72.835 207.505 73.005 207.675 ;
        RECT 73.295 207.505 73.465 207.675 ;
        RECT 73.755 207.505 73.925 207.675 ;
        RECT 74.215 207.505 74.385 207.675 ;
        RECT 74.675 207.505 74.845 207.675 ;
        RECT 75.135 207.505 75.305 207.675 ;
        RECT 75.595 207.505 75.765 207.675 ;
        RECT 76.055 207.505 76.225 207.675 ;
        RECT 76.515 207.505 76.685 207.675 ;
        RECT 76.975 207.505 77.145 207.675 ;
        RECT 77.435 207.505 77.605 207.675 ;
        RECT 77.895 207.505 78.065 207.675 ;
        RECT 78.355 207.505 78.525 207.675 ;
        RECT 78.815 207.505 78.985 207.675 ;
        RECT 79.275 207.505 79.445 207.675 ;
        RECT 79.735 207.505 79.905 207.675 ;
        RECT 80.195 207.505 80.365 207.675 ;
        RECT 80.655 207.505 80.825 207.675 ;
        RECT 81.115 207.505 81.285 207.675 ;
        RECT 81.575 207.505 81.745 207.675 ;
        RECT 82.035 207.505 82.205 207.675 ;
        RECT 82.495 207.505 82.665 207.675 ;
        RECT 82.955 207.505 83.125 207.675 ;
        RECT 83.415 207.505 83.585 207.675 ;
        RECT 83.875 207.505 84.045 207.675 ;
        RECT 84.335 207.505 84.505 207.675 ;
        RECT 84.795 207.505 84.965 207.675 ;
        RECT 85.255 207.505 85.425 207.675 ;
        RECT 85.715 207.505 85.885 207.675 ;
        RECT 86.175 207.505 86.345 207.675 ;
        RECT 86.635 207.505 86.805 207.675 ;
        RECT 87.095 207.505 87.265 207.675 ;
        RECT 87.555 207.505 87.725 207.675 ;
        RECT 88.015 207.505 88.185 207.675 ;
        RECT 88.475 207.505 88.645 207.675 ;
        RECT 88.935 207.505 89.105 207.675 ;
        RECT 89.395 207.505 89.565 207.675 ;
        RECT 89.855 207.505 90.025 207.675 ;
        RECT 90.315 207.505 90.485 207.675 ;
        RECT 90.775 207.505 90.945 207.675 ;
        RECT 91.235 207.505 91.405 207.675 ;
        RECT 91.695 207.505 91.865 207.675 ;
        RECT 92.155 207.505 92.325 207.675 ;
        RECT 92.615 207.505 92.785 207.675 ;
        RECT 93.075 207.505 93.245 207.675 ;
        RECT 93.535 207.505 93.705 207.675 ;
        RECT 93.995 207.505 94.165 207.675 ;
        RECT 94.455 207.505 94.625 207.675 ;
        RECT 94.915 207.505 95.085 207.675 ;
        RECT 95.375 207.505 95.545 207.675 ;
        RECT 95.835 207.505 96.005 207.675 ;
        RECT 96.295 207.505 96.465 207.675 ;
        RECT 96.755 207.505 96.925 207.675 ;
        RECT 97.215 207.505 97.385 207.675 ;
        RECT 97.675 207.505 97.845 207.675 ;
        RECT 98.135 207.505 98.305 207.675 ;
        RECT 98.595 207.505 98.765 207.675 ;
        RECT 99.055 207.505 99.225 207.675 ;
        RECT 99.515 207.505 99.685 207.675 ;
        RECT 99.975 207.505 100.145 207.675 ;
        RECT 100.435 207.505 100.605 207.675 ;
        RECT 100.895 207.505 101.065 207.675 ;
        RECT 101.355 207.505 101.525 207.675 ;
        RECT 101.815 207.505 101.985 207.675 ;
        RECT 102.275 207.505 102.445 207.675 ;
        RECT 102.735 207.505 102.905 207.675 ;
        RECT 103.195 207.505 103.365 207.675 ;
        RECT 103.655 207.505 103.825 207.675 ;
        RECT 104.115 207.505 104.285 207.675 ;
        RECT 104.575 207.505 104.745 207.675 ;
        RECT 105.035 207.505 105.205 207.675 ;
        RECT 105.495 207.505 105.665 207.675 ;
        RECT 105.955 207.505 106.125 207.675 ;
        RECT 106.415 207.505 106.585 207.675 ;
        RECT 106.875 207.505 107.045 207.675 ;
        RECT 107.335 207.505 107.505 207.675 ;
        RECT 107.795 207.505 107.965 207.675 ;
        RECT 108.255 207.505 108.425 207.675 ;
        RECT 108.715 207.505 108.885 207.675 ;
        RECT 109.175 207.505 109.345 207.675 ;
        RECT 109.635 207.505 109.805 207.675 ;
        RECT 110.095 207.505 110.265 207.675 ;
        RECT 110.555 207.505 110.725 207.675 ;
        RECT 111.015 207.505 111.185 207.675 ;
        RECT 111.475 207.505 111.645 207.675 ;
        RECT 111.935 207.505 112.105 207.675 ;
        RECT 112.395 207.505 112.565 207.675 ;
        RECT 112.855 207.505 113.025 207.675 ;
        RECT 113.315 207.505 113.485 207.675 ;
        RECT 113.775 207.505 113.945 207.675 ;
        RECT 114.235 207.505 114.405 207.675 ;
        RECT 114.695 207.505 114.865 207.675 ;
        RECT 115.155 207.505 115.325 207.675 ;
        RECT 70.075 206.315 70.245 206.485 ;
        RECT 71.915 206.655 72.085 206.825 ;
        RECT 78.815 206.995 78.985 207.165 ;
        RECT 71.915 205.295 72.085 205.465 ;
        RECT 72.835 205.295 73.005 205.465 ;
        RECT 74.675 205.635 74.845 205.805 ;
        RECT 75.595 205.975 75.765 206.145 ;
        RECT 76.055 206.315 76.225 206.485 ;
        RECT 76.515 205.975 76.685 206.145 ;
        RECT 76.975 205.975 77.145 206.145 ;
        RECT 77.895 206.315 78.065 206.485 ;
        RECT 79.735 206.315 79.905 206.485 ;
        RECT 82.955 205.975 83.125 206.145 ;
        RECT 88.935 206.995 89.105 207.165 ;
        RECT 84.335 206.315 84.505 206.485 ;
        RECT 83.415 205.295 83.585 205.465 ;
        RECT 85.255 205.635 85.425 205.805 ;
        RECT 90.775 206.995 90.945 207.165 ;
        RECT 89.855 206.315 90.025 206.485 ;
        RECT 92.155 206.655 92.325 206.825 ;
        RECT 91.695 206.315 91.865 206.485 ;
        RECT 93.235 206.655 93.405 206.825 ;
        RECT 94.455 205.975 94.625 206.145 ;
        RECT 95.835 206.315 96.005 206.485 ;
        RECT 96.295 206.315 96.465 206.485 ;
        RECT 93.995 205.635 94.165 205.805 ;
        RECT 93.075 205.295 93.245 205.465 ;
        RECT 95.375 205.975 95.545 206.145 ;
        RECT 97.215 206.315 97.385 206.485 ;
        RECT 95.835 205.635 96.005 205.805 ;
        RECT 96.295 205.295 96.465 205.465 ;
        RECT 98.595 206.315 98.765 206.485 ;
        RECT 99.515 205.975 99.685 206.145 ;
        RECT 100.435 206.315 100.605 206.485 ;
        RECT 97.675 205.295 97.845 205.465 ;
        RECT 100.920 205.635 101.090 205.805 ;
        RECT 101.315 205.975 101.485 206.145 ;
        RECT 101.770 206.315 101.940 206.485 ;
        RECT 102.505 205.975 102.675 206.145 ;
        RECT 103.020 205.635 103.190 205.805 ;
        RECT 104.590 205.635 104.760 205.805 ;
        RECT 105.025 205.975 105.195 206.145 ;
        RECT 107.335 205.295 107.505 205.465 ;
        RECT 107.795 205.295 107.965 205.465 ;
        RECT 112.395 205.975 112.565 206.145 ;
        RECT 61.335 204.785 61.505 204.955 ;
        RECT 61.795 204.785 61.965 204.955 ;
        RECT 62.255 204.785 62.425 204.955 ;
        RECT 62.715 204.785 62.885 204.955 ;
        RECT 63.175 204.785 63.345 204.955 ;
        RECT 63.635 204.785 63.805 204.955 ;
        RECT 64.095 204.785 64.265 204.955 ;
        RECT 64.555 204.785 64.725 204.955 ;
        RECT 65.015 204.785 65.185 204.955 ;
        RECT 65.475 204.785 65.645 204.955 ;
        RECT 65.935 204.785 66.105 204.955 ;
        RECT 66.395 204.785 66.565 204.955 ;
        RECT 66.855 204.785 67.025 204.955 ;
        RECT 67.315 204.785 67.485 204.955 ;
        RECT 67.775 204.785 67.945 204.955 ;
        RECT 68.235 204.785 68.405 204.955 ;
        RECT 68.695 204.785 68.865 204.955 ;
        RECT 69.155 204.785 69.325 204.955 ;
        RECT 69.615 204.785 69.785 204.955 ;
        RECT 70.075 204.785 70.245 204.955 ;
        RECT 70.535 204.785 70.705 204.955 ;
        RECT 70.995 204.785 71.165 204.955 ;
        RECT 71.455 204.785 71.625 204.955 ;
        RECT 71.915 204.785 72.085 204.955 ;
        RECT 72.375 204.785 72.545 204.955 ;
        RECT 72.835 204.785 73.005 204.955 ;
        RECT 73.295 204.785 73.465 204.955 ;
        RECT 73.755 204.785 73.925 204.955 ;
        RECT 74.215 204.785 74.385 204.955 ;
        RECT 74.675 204.785 74.845 204.955 ;
        RECT 75.135 204.785 75.305 204.955 ;
        RECT 75.595 204.785 75.765 204.955 ;
        RECT 76.055 204.785 76.225 204.955 ;
        RECT 76.515 204.785 76.685 204.955 ;
        RECT 76.975 204.785 77.145 204.955 ;
        RECT 77.435 204.785 77.605 204.955 ;
        RECT 77.895 204.785 78.065 204.955 ;
        RECT 78.355 204.785 78.525 204.955 ;
        RECT 78.815 204.785 78.985 204.955 ;
        RECT 79.275 204.785 79.445 204.955 ;
        RECT 79.735 204.785 79.905 204.955 ;
        RECT 80.195 204.785 80.365 204.955 ;
        RECT 80.655 204.785 80.825 204.955 ;
        RECT 81.115 204.785 81.285 204.955 ;
        RECT 81.575 204.785 81.745 204.955 ;
        RECT 82.035 204.785 82.205 204.955 ;
        RECT 82.495 204.785 82.665 204.955 ;
        RECT 82.955 204.785 83.125 204.955 ;
        RECT 83.415 204.785 83.585 204.955 ;
        RECT 83.875 204.785 84.045 204.955 ;
        RECT 84.335 204.785 84.505 204.955 ;
        RECT 84.795 204.785 84.965 204.955 ;
        RECT 85.255 204.785 85.425 204.955 ;
        RECT 85.715 204.785 85.885 204.955 ;
        RECT 86.175 204.785 86.345 204.955 ;
        RECT 86.635 204.785 86.805 204.955 ;
        RECT 87.095 204.785 87.265 204.955 ;
        RECT 87.555 204.785 87.725 204.955 ;
        RECT 88.015 204.785 88.185 204.955 ;
        RECT 88.475 204.785 88.645 204.955 ;
        RECT 88.935 204.785 89.105 204.955 ;
        RECT 89.395 204.785 89.565 204.955 ;
        RECT 89.855 204.785 90.025 204.955 ;
        RECT 90.315 204.785 90.485 204.955 ;
        RECT 90.775 204.785 90.945 204.955 ;
        RECT 91.235 204.785 91.405 204.955 ;
        RECT 91.695 204.785 91.865 204.955 ;
        RECT 92.155 204.785 92.325 204.955 ;
        RECT 92.615 204.785 92.785 204.955 ;
        RECT 93.075 204.785 93.245 204.955 ;
        RECT 93.535 204.785 93.705 204.955 ;
        RECT 93.995 204.785 94.165 204.955 ;
        RECT 94.455 204.785 94.625 204.955 ;
        RECT 94.915 204.785 95.085 204.955 ;
        RECT 95.375 204.785 95.545 204.955 ;
        RECT 95.835 204.785 96.005 204.955 ;
        RECT 96.295 204.785 96.465 204.955 ;
        RECT 96.755 204.785 96.925 204.955 ;
        RECT 97.215 204.785 97.385 204.955 ;
        RECT 97.675 204.785 97.845 204.955 ;
        RECT 98.135 204.785 98.305 204.955 ;
        RECT 98.595 204.785 98.765 204.955 ;
        RECT 99.055 204.785 99.225 204.955 ;
        RECT 99.515 204.785 99.685 204.955 ;
        RECT 99.975 204.785 100.145 204.955 ;
        RECT 100.435 204.785 100.605 204.955 ;
        RECT 100.895 204.785 101.065 204.955 ;
        RECT 101.355 204.785 101.525 204.955 ;
        RECT 101.815 204.785 101.985 204.955 ;
        RECT 102.275 204.785 102.445 204.955 ;
        RECT 102.735 204.785 102.905 204.955 ;
        RECT 103.195 204.785 103.365 204.955 ;
        RECT 103.655 204.785 103.825 204.955 ;
        RECT 104.115 204.785 104.285 204.955 ;
        RECT 104.575 204.785 104.745 204.955 ;
        RECT 105.035 204.785 105.205 204.955 ;
        RECT 105.495 204.785 105.665 204.955 ;
        RECT 105.955 204.785 106.125 204.955 ;
        RECT 106.415 204.785 106.585 204.955 ;
        RECT 106.875 204.785 107.045 204.955 ;
        RECT 107.335 204.785 107.505 204.955 ;
        RECT 107.795 204.785 107.965 204.955 ;
        RECT 108.255 204.785 108.425 204.955 ;
        RECT 108.715 204.785 108.885 204.955 ;
        RECT 109.175 204.785 109.345 204.955 ;
        RECT 109.635 204.785 109.805 204.955 ;
        RECT 110.095 204.785 110.265 204.955 ;
        RECT 110.555 204.785 110.725 204.955 ;
        RECT 111.015 204.785 111.185 204.955 ;
        RECT 111.475 204.785 111.645 204.955 ;
        RECT 111.935 204.785 112.105 204.955 ;
        RECT 112.395 204.785 112.565 204.955 ;
        RECT 112.855 204.785 113.025 204.955 ;
        RECT 113.315 204.785 113.485 204.955 ;
        RECT 113.775 204.785 113.945 204.955 ;
        RECT 114.235 204.785 114.405 204.955 ;
        RECT 114.695 204.785 114.865 204.955 ;
        RECT 115.155 204.785 115.325 204.955 ;
        RECT 65.015 204.275 65.185 204.445 ;
        RECT 66.855 204.275 67.025 204.445 ;
        RECT 65.935 203.255 66.105 203.425 ;
        RECT 68.235 203.595 68.405 203.765 ;
        RECT 67.775 203.255 67.945 203.425 ;
        RECT 72.835 204.275 73.005 204.445 ;
        RECT 71.455 202.575 71.625 202.745 ;
        RECT 76.055 203.935 76.225 204.105 ;
        RECT 73.755 203.255 73.925 203.425 ;
        RECT 74.675 203.255 74.845 203.425 ;
        RECT 75.135 203.255 75.305 203.425 ;
        RECT 76.055 202.915 76.225 203.085 ;
        RECT 77.435 203.255 77.605 203.425 ;
        RECT 77.895 203.595 78.065 203.765 ;
        RECT 78.355 203.255 78.525 203.425 ;
        RECT 78.815 203.255 78.985 203.425 ;
        RECT 79.735 202.915 79.905 203.085 ;
        RECT 76.515 202.575 76.685 202.745 ;
        RECT 82.495 203.595 82.665 203.765 ;
        RECT 85.280 203.935 85.450 204.105 ;
        RECT 84.335 203.255 84.505 203.425 ;
        RECT 84.795 203.255 84.965 203.425 ;
        RECT 83.875 202.575 84.045 202.745 ;
        RECT 85.675 203.595 85.845 203.765 ;
        RECT 86.020 202.915 86.190 203.085 ;
        RECT 87.380 203.935 87.550 204.105 ;
        RECT 86.865 203.595 87.035 203.765 ;
        RECT 88.950 203.935 89.120 204.105 ;
        RECT 89.385 203.595 89.555 203.765 ;
        RECT 91.695 203.935 91.865 204.105 ;
        RECT 92.155 202.575 92.325 202.745 ;
        RECT 95.375 203.255 95.545 203.425 ;
        RECT 97.675 203.595 97.845 203.765 ;
        RECT 99.515 203.935 99.685 204.105 ;
        RECT 96.755 203.255 96.925 203.425 ;
        RECT 98.135 203.255 98.305 203.425 ;
        RECT 95.835 202.575 96.005 202.745 ;
        RECT 98.595 202.575 98.765 202.745 ;
        RECT 99.515 202.915 99.685 203.085 ;
        RECT 100.435 202.915 100.605 203.085 ;
        RECT 103.195 203.595 103.365 203.765 ;
        RECT 107.895 203.935 108.065 204.105 ;
        RECT 105.035 202.575 105.205 202.745 ;
        RECT 106.815 203.230 106.985 203.400 ;
        RECT 106.515 202.915 106.685 203.085 ;
        RECT 107.895 203.255 108.065 203.425 ;
        RECT 111.015 203.935 111.185 204.105 ;
        RECT 109.755 202.915 109.925 203.085 ;
        RECT 110.115 202.915 110.285 203.085 ;
        RECT 111.475 203.255 111.645 203.425 ;
        RECT 112.905 203.935 113.075 204.105 ;
        RECT 112.395 203.595 112.565 203.765 ;
        RECT 113.310 203.255 113.480 203.425 ;
        RECT 113.775 203.255 113.945 203.425 ;
        RECT 61.335 202.065 61.505 202.235 ;
        RECT 61.795 202.065 61.965 202.235 ;
        RECT 62.255 202.065 62.425 202.235 ;
        RECT 62.715 202.065 62.885 202.235 ;
        RECT 63.175 202.065 63.345 202.235 ;
        RECT 63.635 202.065 63.805 202.235 ;
        RECT 64.095 202.065 64.265 202.235 ;
        RECT 64.555 202.065 64.725 202.235 ;
        RECT 65.015 202.065 65.185 202.235 ;
        RECT 65.475 202.065 65.645 202.235 ;
        RECT 65.935 202.065 66.105 202.235 ;
        RECT 66.395 202.065 66.565 202.235 ;
        RECT 66.855 202.065 67.025 202.235 ;
        RECT 67.315 202.065 67.485 202.235 ;
        RECT 67.775 202.065 67.945 202.235 ;
        RECT 68.235 202.065 68.405 202.235 ;
        RECT 68.695 202.065 68.865 202.235 ;
        RECT 69.155 202.065 69.325 202.235 ;
        RECT 69.615 202.065 69.785 202.235 ;
        RECT 70.075 202.065 70.245 202.235 ;
        RECT 70.535 202.065 70.705 202.235 ;
        RECT 70.995 202.065 71.165 202.235 ;
        RECT 71.455 202.065 71.625 202.235 ;
        RECT 71.915 202.065 72.085 202.235 ;
        RECT 72.375 202.065 72.545 202.235 ;
        RECT 72.835 202.065 73.005 202.235 ;
        RECT 73.295 202.065 73.465 202.235 ;
        RECT 73.755 202.065 73.925 202.235 ;
        RECT 74.215 202.065 74.385 202.235 ;
        RECT 74.675 202.065 74.845 202.235 ;
        RECT 75.135 202.065 75.305 202.235 ;
        RECT 75.595 202.065 75.765 202.235 ;
        RECT 76.055 202.065 76.225 202.235 ;
        RECT 76.515 202.065 76.685 202.235 ;
        RECT 76.975 202.065 77.145 202.235 ;
        RECT 77.435 202.065 77.605 202.235 ;
        RECT 77.895 202.065 78.065 202.235 ;
        RECT 78.355 202.065 78.525 202.235 ;
        RECT 78.815 202.065 78.985 202.235 ;
        RECT 79.275 202.065 79.445 202.235 ;
        RECT 79.735 202.065 79.905 202.235 ;
        RECT 80.195 202.065 80.365 202.235 ;
        RECT 80.655 202.065 80.825 202.235 ;
        RECT 81.115 202.065 81.285 202.235 ;
        RECT 81.575 202.065 81.745 202.235 ;
        RECT 82.035 202.065 82.205 202.235 ;
        RECT 82.495 202.065 82.665 202.235 ;
        RECT 82.955 202.065 83.125 202.235 ;
        RECT 83.415 202.065 83.585 202.235 ;
        RECT 83.875 202.065 84.045 202.235 ;
        RECT 84.335 202.065 84.505 202.235 ;
        RECT 84.795 202.065 84.965 202.235 ;
        RECT 85.255 202.065 85.425 202.235 ;
        RECT 85.715 202.065 85.885 202.235 ;
        RECT 86.175 202.065 86.345 202.235 ;
        RECT 86.635 202.065 86.805 202.235 ;
        RECT 87.095 202.065 87.265 202.235 ;
        RECT 87.555 202.065 87.725 202.235 ;
        RECT 88.015 202.065 88.185 202.235 ;
        RECT 88.475 202.065 88.645 202.235 ;
        RECT 88.935 202.065 89.105 202.235 ;
        RECT 89.395 202.065 89.565 202.235 ;
        RECT 89.855 202.065 90.025 202.235 ;
        RECT 90.315 202.065 90.485 202.235 ;
        RECT 90.775 202.065 90.945 202.235 ;
        RECT 91.235 202.065 91.405 202.235 ;
        RECT 91.695 202.065 91.865 202.235 ;
        RECT 92.155 202.065 92.325 202.235 ;
        RECT 92.615 202.065 92.785 202.235 ;
        RECT 93.075 202.065 93.245 202.235 ;
        RECT 93.535 202.065 93.705 202.235 ;
        RECT 93.995 202.065 94.165 202.235 ;
        RECT 94.455 202.065 94.625 202.235 ;
        RECT 94.915 202.065 95.085 202.235 ;
        RECT 95.375 202.065 95.545 202.235 ;
        RECT 95.835 202.065 96.005 202.235 ;
        RECT 96.295 202.065 96.465 202.235 ;
        RECT 96.755 202.065 96.925 202.235 ;
        RECT 97.215 202.065 97.385 202.235 ;
        RECT 97.675 202.065 97.845 202.235 ;
        RECT 98.135 202.065 98.305 202.235 ;
        RECT 98.595 202.065 98.765 202.235 ;
        RECT 99.055 202.065 99.225 202.235 ;
        RECT 99.515 202.065 99.685 202.235 ;
        RECT 99.975 202.065 100.145 202.235 ;
        RECT 100.435 202.065 100.605 202.235 ;
        RECT 100.895 202.065 101.065 202.235 ;
        RECT 101.355 202.065 101.525 202.235 ;
        RECT 101.815 202.065 101.985 202.235 ;
        RECT 102.275 202.065 102.445 202.235 ;
        RECT 102.735 202.065 102.905 202.235 ;
        RECT 103.195 202.065 103.365 202.235 ;
        RECT 103.655 202.065 103.825 202.235 ;
        RECT 104.115 202.065 104.285 202.235 ;
        RECT 104.575 202.065 104.745 202.235 ;
        RECT 105.035 202.065 105.205 202.235 ;
        RECT 105.495 202.065 105.665 202.235 ;
        RECT 105.955 202.065 106.125 202.235 ;
        RECT 106.415 202.065 106.585 202.235 ;
        RECT 106.875 202.065 107.045 202.235 ;
        RECT 107.335 202.065 107.505 202.235 ;
        RECT 107.795 202.065 107.965 202.235 ;
        RECT 108.255 202.065 108.425 202.235 ;
        RECT 108.715 202.065 108.885 202.235 ;
        RECT 109.175 202.065 109.345 202.235 ;
        RECT 109.635 202.065 109.805 202.235 ;
        RECT 110.095 202.065 110.265 202.235 ;
        RECT 110.555 202.065 110.725 202.235 ;
        RECT 111.015 202.065 111.185 202.235 ;
        RECT 111.475 202.065 111.645 202.235 ;
        RECT 111.935 202.065 112.105 202.235 ;
        RECT 112.395 202.065 112.565 202.235 ;
        RECT 112.855 202.065 113.025 202.235 ;
        RECT 113.315 202.065 113.485 202.235 ;
        RECT 113.775 202.065 113.945 202.235 ;
        RECT 114.235 202.065 114.405 202.235 ;
        RECT 114.695 202.065 114.865 202.235 ;
        RECT 115.155 202.065 115.325 202.235 ;
        RECT 63.635 200.875 63.805 201.045 ;
        RECT 65.475 201.215 65.645 201.385 ;
        RECT 64.555 200.875 64.725 201.045 ;
        RECT 65.015 200.875 65.185 201.045 ;
        RECT 66.395 200.875 66.565 201.045 ;
        RECT 64.555 199.855 64.725 200.025 ;
        RECT 66.395 199.855 66.565 200.025 ;
        RECT 66.855 200.195 67.025 200.365 ;
        RECT 69.165 200.535 69.335 200.705 ;
        RECT 69.600 200.195 69.770 200.365 ;
        RECT 71.685 200.535 71.855 200.705 ;
        RECT 71.170 200.195 71.340 200.365 ;
        RECT 72.420 200.875 72.590 201.045 ;
        RECT 72.875 200.535 73.045 200.705 ;
        RECT 74.675 201.555 74.845 201.725 ;
        RECT 74.215 200.875 74.385 201.045 ;
        RECT 73.755 200.535 73.925 200.705 ;
        RECT 75.135 200.875 75.305 201.045 ;
        RECT 73.270 200.195 73.440 200.365 ;
        RECT 75.595 199.855 75.765 200.025 ;
        RECT 77.905 200.535 78.075 200.705 ;
        RECT 78.340 200.195 78.510 200.365 ;
        RECT 80.425 200.535 80.595 200.705 ;
        RECT 79.910 200.195 80.080 200.365 ;
        RECT 81.270 201.215 81.440 201.385 ;
        RECT 81.615 200.535 81.785 200.705 ;
        RECT 84.335 201.555 84.505 201.725 ;
        RECT 82.955 200.875 83.125 201.045 ;
        RECT 82.495 200.535 82.665 200.705 ;
        RECT 83.875 200.875 84.045 201.045 ;
        RECT 82.010 200.195 82.180 200.365 ;
        RECT 83.415 200.535 83.585 200.705 ;
        RECT 85.255 200.875 85.425 201.045 ;
        RECT 86.175 200.875 86.345 201.045 ;
        RECT 86.635 200.875 86.805 201.045 ;
        RECT 88.475 200.875 88.645 201.045 ;
        RECT 87.555 199.855 87.725 200.025 ;
        RECT 90.315 200.535 90.485 200.705 ;
        RECT 89.395 200.195 89.565 200.365 ;
        RECT 93.535 200.875 93.705 201.045 ;
        RECT 93.995 200.875 94.165 201.045 ;
        RECT 94.480 200.195 94.650 200.365 ;
        RECT 94.875 200.535 95.045 200.705 ;
        RECT 95.330 200.875 95.500 201.045 ;
        RECT 96.065 200.535 96.235 200.705 ;
        RECT 96.580 200.195 96.750 200.365 ;
        RECT 98.150 200.195 98.320 200.365 ;
        RECT 98.585 200.535 98.755 200.705 ;
        RECT 101.355 201.555 101.525 201.725 ;
        RECT 100.895 199.855 101.065 200.025 ;
        RECT 105.955 201.555 106.125 201.725 ;
        RECT 104.115 200.875 104.285 201.045 ;
        RECT 105.035 200.875 105.205 201.045 ;
        RECT 109.635 200.535 109.805 200.705 ;
        RECT 111.475 200.875 111.645 201.045 ;
        RECT 111.015 200.535 111.185 200.705 ;
        RECT 112.395 200.875 112.565 201.045 ;
        RECT 111.475 199.855 111.645 200.025 ;
        RECT 61.335 199.345 61.505 199.515 ;
        RECT 61.795 199.345 61.965 199.515 ;
        RECT 62.255 199.345 62.425 199.515 ;
        RECT 62.715 199.345 62.885 199.515 ;
        RECT 63.175 199.345 63.345 199.515 ;
        RECT 63.635 199.345 63.805 199.515 ;
        RECT 64.095 199.345 64.265 199.515 ;
        RECT 64.555 199.345 64.725 199.515 ;
        RECT 65.015 199.345 65.185 199.515 ;
        RECT 65.475 199.345 65.645 199.515 ;
        RECT 65.935 199.345 66.105 199.515 ;
        RECT 66.395 199.345 66.565 199.515 ;
        RECT 66.855 199.345 67.025 199.515 ;
        RECT 67.315 199.345 67.485 199.515 ;
        RECT 67.775 199.345 67.945 199.515 ;
        RECT 68.235 199.345 68.405 199.515 ;
        RECT 68.695 199.345 68.865 199.515 ;
        RECT 69.155 199.345 69.325 199.515 ;
        RECT 69.615 199.345 69.785 199.515 ;
        RECT 70.075 199.345 70.245 199.515 ;
        RECT 70.535 199.345 70.705 199.515 ;
        RECT 70.995 199.345 71.165 199.515 ;
        RECT 71.455 199.345 71.625 199.515 ;
        RECT 71.915 199.345 72.085 199.515 ;
        RECT 72.375 199.345 72.545 199.515 ;
        RECT 72.835 199.345 73.005 199.515 ;
        RECT 73.295 199.345 73.465 199.515 ;
        RECT 73.755 199.345 73.925 199.515 ;
        RECT 74.215 199.345 74.385 199.515 ;
        RECT 74.675 199.345 74.845 199.515 ;
        RECT 75.135 199.345 75.305 199.515 ;
        RECT 75.595 199.345 75.765 199.515 ;
        RECT 76.055 199.345 76.225 199.515 ;
        RECT 76.515 199.345 76.685 199.515 ;
        RECT 76.975 199.345 77.145 199.515 ;
        RECT 77.435 199.345 77.605 199.515 ;
        RECT 77.895 199.345 78.065 199.515 ;
        RECT 78.355 199.345 78.525 199.515 ;
        RECT 78.815 199.345 78.985 199.515 ;
        RECT 79.275 199.345 79.445 199.515 ;
        RECT 79.735 199.345 79.905 199.515 ;
        RECT 80.195 199.345 80.365 199.515 ;
        RECT 80.655 199.345 80.825 199.515 ;
        RECT 81.115 199.345 81.285 199.515 ;
        RECT 81.575 199.345 81.745 199.515 ;
        RECT 82.035 199.345 82.205 199.515 ;
        RECT 82.495 199.345 82.665 199.515 ;
        RECT 82.955 199.345 83.125 199.515 ;
        RECT 83.415 199.345 83.585 199.515 ;
        RECT 83.875 199.345 84.045 199.515 ;
        RECT 84.335 199.345 84.505 199.515 ;
        RECT 84.795 199.345 84.965 199.515 ;
        RECT 85.255 199.345 85.425 199.515 ;
        RECT 85.715 199.345 85.885 199.515 ;
        RECT 86.175 199.345 86.345 199.515 ;
        RECT 86.635 199.345 86.805 199.515 ;
        RECT 87.095 199.345 87.265 199.515 ;
        RECT 87.555 199.345 87.725 199.515 ;
        RECT 88.015 199.345 88.185 199.515 ;
        RECT 88.475 199.345 88.645 199.515 ;
        RECT 88.935 199.345 89.105 199.515 ;
        RECT 89.395 199.345 89.565 199.515 ;
        RECT 89.855 199.345 90.025 199.515 ;
        RECT 90.315 199.345 90.485 199.515 ;
        RECT 90.775 199.345 90.945 199.515 ;
        RECT 91.235 199.345 91.405 199.515 ;
        RECT 91.695 199.345 91.865 199.515 ;
        RECT 92.155 199.345 92.325 199.515 ;
        RECT 92.615 199.345 92.785 199.515 ;
        RECT 93.075 199.345 93.245 199.515 ;
        RECT 93.535 199.345 93.705 199.515 ;
        RECT 93.995 199.345 94.165 199.515 ;
        RECT 94.455 199.345 94.625 199.515 ;
        RECT 94.915 199.345 95.085 199.515 ;
        RECT 95.375 199.345 95.545 199.515 ;
        RECT 95.835 199.345 96.005 199.515 ;
        RECT 96.295 199.345 96.465 199.515 ;
        RECT 96.755 199.345 96.925 199.515 ;
        RECT 97.215 199.345 97.385 199.515 ;
        RECT 97.675 199.345 97.845 199.515 ;
        RECT 98.135 199.345 98.305 199.515 ;
        RECT 98.595 199.345 98.765 199.515 ;
        RECT 99.055 199.345 99.225 199.515 ;
        RECT 99.515 199.345 99.685 199.515 ;
        RECT 99.975 199.345 100.145 199.515 ;
        RECT 100.435 199.345 100.605 199.515 ;
        RECT 100.895 199.345 101.065 199.515 ;
        RECT 101.355 199.345 101.525 199.515 ;
        RECT 101.815 199.345 101.985 199.515 ;
        RECT 102.275 199.345 102.445 199.515 ;
        RECT 102.735 199.345 102.905 199.515 ;
        RECT 103.195 199.345 103.365 199.515 ;
        RECT 103.655 199.345 103.825 199.515 ;
        RECT 104.115 199.345 104.285 199.515 ;
        RECT 104.575 199.345 104.745 199.515 ;
        RECT 105.035 199.345 105.205 199.515 ;
        RECT 105.495 199.345 105.665 199.515 ;
        RECT 105.955 199.345 106.125 199.515 ;
        RECT 106.415 199.345 106.585 199.515 ;
        RECT 106.875 199.345 107.045 199.515 ;
        RECT 107.335 199.345 107.505 199.515 ;
        RECT 107.795 199.345 107.965 199.515 ;
        RECT 108.255 199.345 108.425 199.515 ;
        RECT 108.715 199.345 108.885 199.515 ;
        RECT 109.175 199.345 109.345 199.515 ;
        RECT 109.635 199.345 109.805 199.515 ;
        RECT 110.095 199.345 110.265 199.515 ;
        RECT 110.555 199.345 110.725 199.515 ;
        RECT 111.015 199.345 111.185 199.515 ;
        RECT 111.475 199.345 111.645 199.515 ;
        RECT 111.935 199.345 112.105 199.515 ;
        RECT 112.395 199.345 112.565 199.515 ;
        RECT 112.855 199.345 113.025 199.515 ;
        RECT 113.315 199.345 113.485 199.515 ;
        RECT 113.775 199.345 113.945 199.515 ;
        RECT 114.235 199.345 114.405 199.515 ;
        RECT 114.695 199.345 114.865 199.515 ;
        RECT 115.155 199.345 115.325 199.515 ;
        RECT 64.095 198.495 64.265 198.665 ;
        RECT 65.015 198.835 65.185 199.005 ;
        RECT 64.555 197.815 64.725 197.985 ;
        RECT 67.325 198.155 67.495 198.325 ;
        RECT 67.760 198.495 67.930 198.665 ;
        RECT 69.330 198.495 69.500 198.665 ;
        RECT 69.845 198.155 70.015 198.325 ;
        RECT 70.580 197.815 70.750 197.985 ;
        RECT 71.035 198.155 71.205 198.325 ;
        RECT 71.430 198.495 71.600 198.665 ;
        RECT 71.915 198.155 72.085 198.325 ;
        RECT 72.835 198.495 73.005 198.665 ;
        RECT 76.080 198.495 76.250 198.665 ;
        RECT 73.755 197.815 73.925 197.985 ;
        RECT 75.595 197.815 75.765 197.985 ;
        RECT 76.475 198.155 76.645 198.325 ;
        RECT 76.820 197.475 76.990 197.645 ;
        RECT 78.180 198.495 78.350 198.665 ;
        RECT 77.665 198.155 77.835 198.325 ;
        RECT 79.750 198.495 79.920 198.665 ;
        RECT 80.185 198.155 80.355 198.325 ;
        RECT 83.415 198.495 83.585 198.665 ;
        RECT 82.495 197.135 82.665 197.305 ;
        RECT 84.795 198.835 84.965 199.005 ;
        RECT 87.120 198.495 87.290 198.665 ;
        RECT 84.335 197.815 84.505 197.985 ;
        RECT 84.795 197.475 84.965 197.645 ;
        RECT 86.635 198.155 86.805 198.325 ;
        RECT 86.175 197.815 86.345 197.985 ;
        RECT 85.715 197.135 85.885 197.305 ;
        RECT 87.515 198.155 87.685 198.325 ;
        RECT 87.970 197.475 88.140 197.645 ;
        RECT 89.220 198.495 89.390 198.665 ;
        RECT 88.705 198.155 88.875 198.325 ;
        RECT 90.790 198.495 90.960 198.665 ;
        RECT 91.225 198.155 91.395 198.325 ;
        RECT 93.535 198.835 93.705 199.005 ;
        RECT 96.755 198.495 96.925 198.665 ;
        RECT 93.995 197.135 94.165 197.305 ;
        RECT 94.915 197.135 95.085 197.305 ;
        RECT 95.375 197.815 95.545 197.985 ;
        RECT 95.835 197.475 96.005 197.645 ;
        RECT 98.135 198.835 98.305 199.005 ;
        RECT 100.895 198.495 101.065 198.665 ;
        RECT 97.215 197.135 97.385 197.305 ;
        RECT 98.055 197.135 98.225 197.305 ;
        RECT 102.735 198.835 102.905 199.005 ;
        RECT 100.435 197.815 100.605 197.985 ;
        RECT 101.815 197.815 101.985 197.985 ;
        RECT 99.055 197.475 99.225 197.645 ;
        RECT 103.680 198.495 103.850 198.665 ;
        RECT 103.195 197.815 103.365 197.985 ;
        RECT 104.075 198.155 104.245 198.325 ;
        RECT 104.420 197.475 104.590 197.645 ;
        RECT 105.780 198.495 105.950 198.665 ;
        RECT 105.265 198.155 105.435 198.325 ;
        RECT 107.350 198.495 107.520 198.665 ;
        RECT 107.785 198.155 107.955 198.325 ;
        RECT 110.095 198.495 110.265 198.665 ;
        RECT 110.555 197.135 110.725 197.305 ;
        RECT 113.315 198.155 113.485 198.325 ;
        RECT 61.335 196.625 61.505 196.795 ;
        RECT 61.795 196.625 61.965 196.795 ;
        RECT 62.255 196.625 62.425 196.795 ;
        RECT 62.715 196.625 62.885 196.795 ;
        RECT 63.175 196.625 63.345 196.795 ;
        RECT 63.635 196.625 63.805 196.795 ;
        RECT 64.095 196.625 64.265 196.795 ;
        RECT 64.555 196.625 64.725 196.795 ;
        RECT 65.015 196.625 65.185 196.795 ;
        RECT 65.475 196.625 65.645 196.795 ;
        RECT 65.935 196.625 66.105 196.795 ;
        RECT 66.395 196.625 66.565 196.795 ;
        RECT 66.855 196.625 67.025 196.795 ;
        RECT 67.315 196.625 67.485 196.795 ;
        RECT 67.775 196.625 67.945 196.795 ;
        RECT 68.235 196.625 68.405 196.795 ;
        RECT 68.695 196.625 68.865 196.795 ;
        RECT 69.155 196.625 69.325 196.795 ;
        RECT 69.615 196.625 69.785 196.795 ;
        RECT 70.075 196.625 70.245 196.795 ;
        RECT 70.535 196.625 70.705 196.795 ;
        RECT 70.995 196.625 71.165 196.795 ;
        RECT 71.455 196.625 71.625 196.795 ;
        RECT 71.915 196.625 72.085 196.795 ;
        RECT 72.375 196.625 72.545 196.795 ;
        RECT 72.835 196.625 73.005 196.795 ;
        RECT 73.295 196.625 73.465 196.795 ;
        RECT 73.755 196.625 73.925 196.795 ;
        RECT 74.215 196.625 74.385 196.795 ;
        RECT 74.675 196.625 74.845 196.795 ;
        RECT 75.135 196.625 75.305 196.795 ;
        RECT 75.595 196.625 75.765 196.795 ;
        RECT 76.055 196.625 76.225 196.795 ;
        RECT 76.515 196.625 76.685 196.795 ;
        RECT 76.975 196.625 77.145 196.795 ;
        RECT 77.435 196.625 77.605 196.795 ;
        RECT 77.895 196.625 78.065 196.795 ;
        RECT 78.355 196.625 78.525 196.795 ;
        RECT 78.815 196.625 78.985 196.795 ;
        RECT 79.275 196.625 79.445 196.795 ;
        RECT 79.735 196.625 79.905 196.795 ;
        RECT 80.195 196.625 80.365 196.795 ;
        RECT 80.655 196.625 80.825 196.795 ;
        RECT 81.115 196.625 81.285 196.795 ;
        RECT 81.575 196.625 81.745 196.795 ;
        RECT 82.035 196.625 82.205 196.795 ;
        RECT 82.495 196.625 82.665 196.795 ;
        RECT 82.955 196.625 83.125 196.795 ;
        RECT 83.415 196.625 83.585 196.795 ;
        RECT 83.875 196.625 84.045 196.795 ;
        RECT 84.335 196.625 84.505 196.795 ;
        RECT 84.795 196.625 84.965 196.795 ;
        RECT 85.255 196.625 85.425 196.795 ;
        RECT 85.715 196.625 85.885 196.795 ;
        RECT 86.175 196.625 86.345 196.795 ;
        RECT 86.635 196.625 86.805 196.795 ;
        RECT 87.095 196.625 87.265 196.795 ;
        RECT 87.555 196.625 87.725 196.795 ;
        RECT 88.015 196.625 88.185 196.795 ;
        RECT 88.475 196.625 88.645 196.795 ;
        RECT 88.935 196.625 89.105 196.795 ;
        RECT 89.395 196.625 89.565 196.795 ;
        RECT 89.855 196.625 90.025 196.795 ;
        RECT 90.315 196.625 90.485 196.795 ;
        RECT 90.775 196.625 90.945 196.795 ;
        RECT 91.235 196.625 91.405 196.795 ;
        RECT 91.695 196.625 91.865 196.795 ;
        RECT 92.155 196.625 92.325 196.795 ;
        RECT 92.615 196.625 92.785 196.795 ;
        RECT 93.075 196.625 93.245 196.795 ;
        RECT 93.535 196.625 93.705 196.795 ;
        RECT 93.995 196.625 94.165 196.795 ;
        RECT 94.455 196.625 94.625 196.795 ;
        RECT 94.915 196.625 95.085 196.795 ;
        RECT 95.375 196.625 95.545 196.795 ;
        RECT 95.835 196.625 96.005 196.795 ;
        RECT 96.295 196.625 96.465 196.795 ;
        RECT 96.755 196.625 96.925 196.795 ;
        RECT 97.215 196.625 97.385 196.795 ;
        RECT 97.675 196.625 97.845 196.795 ;
        RECT 98.135 196.625 98.305 196.795 ;
        RECT 98.595 196.625 98.765 196.795 ;
        RECT 99.055 196.625 99.225 196.795 ;
        RECT 99.515 196.625 99.685 196.795 ;
        RECT 99.975 196.625 100.145 196.795 ;
        RECT 100.435 196.625 100.605 196.795 ;
        RECT 100.895 196.625 101.065 196.795 ;
        RECT 101.355 196.625 101.525 196.795 ;
        RECT 101.815 196.625 101.985 196.795 ;
        RECT 102.275 196.625 102.445 196.795 ;
        RECT 102.735 196.625 102.905 196.795 ;
        RECT 103.195 196.625 103.365 196.795 ;
        RECT 103.655 196.625 103.825 196.795 ;
        RECT 104.115 196.625 104.285 196.795 ;
        RECT 104.575 196.625 104.745 196.795 ;
        RECT 105.035 196.625 105.205 196.795 ;
        RECT 105.495 196.625 105.665 196.795 ;
        RECT 105.955 196.625 106.125 196.795 ;
        RECT 106.415 196.625 106.585 196.795 ;
        RECT 106.875 196.625 107.045 196.795 ;
        RECT 107.335 196.625 107.505 196.795 ;
        RECT 107.795 196.625 107.965 196.795 ;
        RECT 108.255 196.625 108.425 196.795 ;
        RECT 108.715 196.625 108.885 196.795 ;
        RECT 109.175 196.625 109.345 196.795 ;
        RECT 109.635 196.625 109.805 196.795 ;
        RECT 110.095 196.625 110.265 196.795 ;
        RECT 110.555 196.625 110.725 196.795 ;
        RECT 111.015 196.625 111.185 196.795 ;
        RECT 111.475 196.625 111.645 196.795 ;
        RECT 111.935 196.625 112.105 196.795 ;
        RECT 112.395 196.625 112.565 196.795 ;
        RECT 112.855 196.625 113.025 196.795 ;
        RECT 113.315 196.625 113.485 196.795 ;
        RECT 113.775 196.625 113.945 196.795 ;
        RECT 114.235 196.625 114.405 196.795 ;
        RECT 114.695 196.625 114.865 196.795 ;
        RECT 115.155 196.625 115.325 196.795 ;
        RECT 70.535 196.115 70.705 196.285 ;
        RECT 74.675 196.115 74.845 196.285 ;
        RECT 71.455 195.435 71.625 195.605 ;
        RECT 71.915 195.095 72.085 195.265 ;
        RECT 72.375 195.095 72.545 195.265 ;
        RECT 72.835 195.435 73.005 195.605 ;
        RECT 75.515 196.115 75.685 196.285 ;
        RECT 76.515 195.775 76.685 195.945 ;
        RECT 85.715 195.775 85.885 195.945 ;
        RECT 87.555 196.115 87.725 196.285 ;
        RECT 75.595 194.415 75.765 194.585 ;
        RECT 91.235 196.115 91.405 196.285 ;
        RECT 88.475 195.435 88.645 195.605 ;
        RECT 98.595 196.115 98.765 196.285 ;
        RECT 97.675 195.435 97.845 195.605 ;
        RECT 101.355 195.775 101.525 195.945 ;
        RECT 99.515 195.435 99.685 195.605 ;
        RECT 100.895 195.435 101.065 195.605 ;
        RECT 110.095 195.775 110.265 195.945 ;
        RECT 100.435 194.415 100.605 194.585 ;
        RECT 111.475 195.435 111.645 195.605 ;
        RECT 112.395 195.095 112.565 195.265 ;
        RECT 110.555 194.415 110.725 194.585 ;
        RECT 61.335 193.905 61.505 194.075 ;
        RECT 61.795 193.905 61.965 194.075 ;
        RECT 62.255 193.905 62.425 194.075 ;
        RECT 62.715 193.905 62.885 194.075 ;
        RECT 63.175 193.905 63.345 194.075 ;
        RECT 63.635 193.905 63.805 194.075 ;
        RECT 64.095 193.905 64.265 194.075 ;
        RECT 64.555 193.905 64.725 194.075 ;
        RECT 65.015 193.905 65.185 194.075 ;
        RECT 65.475 193.905 65.645 194.075 ;
        RECT 65.935 193.905 66.105 194.075 ;
        RECT 66.395 193.905 66.565 194.075 ;
        RECT 66.855 193.905 67.025 194.075 ;
        RECT 67.315 193.905 67.485 194.075 ;
        RECT 67.775 193.905 67.945 194.075 ;
        RECT 68.235 193.905 68.405 194.075 ;
        RECT 68.695 193.905 68.865 194.075 ;
        RECT 69.155 193.905 69.325 194.075 ;
        RECT 69.615 193.905 69.785 194.075 ;
        RECT 70.075 193.905 70.245 194.075 ;
        RECT 70.535 193.905 70.705 194.075 ;
        RECT 70.995 193.905 71.165 194.075 ;
        RECT 71.455 193.905 71.625 194.075 ;
        RECT 71.915 193.905 72.085 194.075 ;
        RECT 72.375 193.905 72.545 194.075 ;
        RECT 72.835 193.905 73.005 194.075 ;
        RECT 73.295 193.905 73.465 194.075 ;
        RECT 73.755 193.905 73.925 194.075 ;
        RECT 74.215 193.905 74.385 194.075 ;
        RECT 74.675 193.905 74.845 194.075 ;
        RECT 75.135 193.905 75.305 194.075 ;
        RECT 75.595 193.905 75.765 194.075 ;
        RECT 76.055 193.905 76.225 194.075 ;
        RECT 76.515 193.905 76.685 194.075 ;
        RECT 76.975 193.905 77.145 194.075 ;
        RECT 77.435 193.905 77.605 194.075 ;
        RECT 77.895 193.905 78.065 194.075 ;
        RECT 78.355 193.905 78.525 194.075 ;
        RECT 78.815 193.905 78.985 194.075 ;
        RECT 79.275 193.905 79.445 194.075 ;
        RECT 79.735 193.905 79.905 194.075 ;
        RECT 80.195 193.905 80.365 194.075 ;
        RECT 80.655 193.905 80.825 194.075 ;
        RECT 81.115 193.905 81.285 194.075 ;
        RECT 81.575 193.905 81.745 194.075 ;
        RECT 82.035 193.905 82.205 194.075 ;
        RECT 82.495 193.905 82.665 194.075 ;
        RECT 82.955 193.905 83.125 194.075 ;
        RECT 83.415 193.905 83.585 194.075 ;
        RECT 83.875 193.905 84.045 194.075 ;
        RECT 84.335 193.905 84.505 194.075 ;
        RECT 84.795 193.905 84.965 194.075 ;
        RECT 85.255 193.905 85.425 194.075 ;
        RECT 85.715 193.905 85.885 194.075 ;
        RECT 86.175 193.905 86.345 194.075 ;
        RECT 86.635 193.905 86.805 194.075 ;
        RECT 87.095 193.905 87.265 194.075 ;
        RECT 87.555 193.905 87.725 194.075 ;
        RECT 88.015 193.905 88.185 194.075 ;
        RECT 88.475 193.905 88.645 194.075 ;
        RECT 88.935 193.905 89.105 194.075 ;
        RECT 89.395 193.905 89.565 194.075 ;
        RECT 89.855 193.905 90.025 194.075 ;
        RECT 90.315 193.905 90.485 194.075 ;
        RECT 90.775 193.905 90.945 194.075 ;
        RECT 91.235 193.905 91.405 194.075 ;
        RECT 91.695 193.905 91.865 194.075 ;
        RECT 92.155 193.905 92.325 194.075 ;
        RECT 92.615 193.905 92.785 194.075 ;
        RECT 93.075 193.905 93.245 194.075 ;
        RECT 93.535 193.905 93.705 194.075 ;
        RECT 93.995 193.905 94.165 194.075 ;
        RECT 94.455 193.905 94.625 194.075 ;
        RECT 94.915 193.905 95.085 194.075 ;
        RECT 95.375 193.905 95.545 194.075 ;
        RECT 95.835 193.905 96.005 194.075 ;
        RECT 96.295 193.905 96.465 194.075 ;
        RECT 96.755 193.905 96.925 194.075 ;
        RECT 97.215 193.905 97.385 194.075 ;
        RECT 97.675 193.905 97.845 194.075 ;
        RECT 98.135 193.905 98.305 194.075 ;
        RECT 98.595 193.905 98.765 194.075 ;
        RECT 99.055 193.905 99.225 194.075 ;
        RECT 99.515 193.905 99.685 194.075 ;
        RECT 99.975 193.905 100.145 194.075 ;
        RECT 100.435 193.905 100.605 194.075 ;
        RECT 100.895 193.905 101.065 194.075 ;
        RECT 101.355 193.905 101.525 194.075 ;
        RECT 101.815 193.905 101.985 194.075 ;
        RECT 102.275 193.905 102.445 194.075 ;
        RECT 102.735 193.905 102.905 194.075 ;
        RECT 103.195 193.905 103.365 194.075 ;
        RECT 103.655 193.905 103.825 194.075 ;
        RECT 104.115 193.905 104.285 194.075 ;
        RECT 104.575 193.905 104.745 194.075 ;
        RECT 105.035 193.905 105.205 194.075 ;
        RECT 105.495 193.905 105.665 194.075 ;
        RECT 105.955 193.905 106.125 194.075 ;
        RECT 106.415 193.905 106.585 194.075 ;
        RECT 106.875 193.905 107.045 194.075 ;
        RECT 107.335 193.905 107.505 194.075 ;
        RECT 107.795 193.905 107.965 194.075 ;
        RECT 108.255 193.905 108.425 194.075 ;
        RECT 108.715 193.905 108.885 194.075 ;
        RECT 109.175 193.905 109.345 194.075 ;
        RECT 109.635 193.905 109.805 194.075 ;
        RECT 110.095 193.905 110.265 194.075 ;
        RECT 110.555 193.905 110.725 194.075 ;
        RECT 111.015 193.905 111.185 194.075 ;
        RECT 111.475 193.905 111.645 194.075 ;
        RECT 111.935 193.905 112.105 194.075 ;
        RECT 112.395 193.905 112.565 194.075 ;
        RECT 112.855 193.905 113.025 194.075 ;
        RECT 113.315 193.905 113.485 194.075 ;
        RECT 113.775 193.905 113.945 194.075 ;
        RECT 114.235 193.905 114.405 194.075 ;
        RECT 114.695 193.905 114.865 194.075 ;
        RECT 115.155 193.905 115.325 194.075 ;
        RECT 72.835 193.395 73.005 193.565 ;
        RECT 75.595 193.055 75.765 193.225 ;
        RECT 73.755 192.375 73.925 192.545 ;
        RECT 74.675 192.375 74.845 192.545 ;
        RECT 75.595 192.375 75.765 192.545 ;
        RECT 76.055 192.375 76.225 192.545 ;
        RECT 79.275 193.055 79.445 193.225 ;
        RECT 79.735 193.395 79.905 193.565 ;
        RECT 76.975 192.375 77.145 192.545 ;
        RECT 77.435 192.375 77.605 192.545 ;
        RECT 77.895 192.375 78.065 192.545 ;
        RECT 78.355 192.375 78.525 192.545 ;
        RECT 77.435 191.695 77.605 191.865 ;
        RECT 79.275 192.035 79.445 192.205 ;
        RECT 82.955 192.375 83.125 192.545 ;
        RECT 83.415 192.035 83.585 192.205 ;
        RECT 84.335 191.695 84.505 191.865 ;
        RECT 84.795 191.695 84.965 191.865 ;
        RECT 86.175 192.375 86.345 192.545 ;
        RECT 85.255 192.035 85.425 192.205 ;
        RECT 86.635 192.715 86.805 192.885 ;
        RECT 87.555 192.375 87.725 192.545 ;
        RECT 90.315 193.055 90.485 193.225 ;
        RECT 89.395 192.375 89.565 192.545 ;
        RECT 90.775 192.375 90.945 192.545 ;
        RECT 92.155 192.375 92.325 192.545 ;
        RECT 92.615 192.375 92.785 192.545 ;
        RECT 93.075 192.375 93.245 192.545 ;
        RECT 88.475 191.695 88.645 191.865 ;
        RECT 91.235 192.035 91.405 192.205 ;
        RECT 95.835 193.395 96.005 193.565 ;
        RECT 94.455 192.375 94.625 192.545 ;
        RECT 94.915 192.375 95.085 192.545 ;
        RECT 99.055 193.055 99.225 193.225 ;
        RECT 98.135 192.375 98.305 192.545 ;
        RECT 99.515 192.375 99.685 192.545 ;
        RECT 102.275 193.395 102.445 193.565 ;
        RECT 97.215 191.695 97.385 191.865 ;
        RECT 100.435 192.035 100.605 192.205 ;
        RECT 103.680 193.055 103.850 193.225 ;
        RECT 101.355 192.375 101.525 192.545 ;
        RECT 102.735 192.375 102.905 192.545 ;
        RECT 103.195 192.375 103.365 192.545 ;
        RECT 104.075 192.715 104.245 192.885 ;
        RECT 104.420 192.035 104.590 192.205 ;
        RECT 105.780 193.055 105.950 193.225 ;
        RECT 105.265 192.715 105.435 192.885 ;
        RECT 107.350 193.055 107.520 193.225 ;
        RECT 107.785 192.715 107.955 192.885 ;
        RECT 110.555 192.035 110.725 192.205 ;
        RECT 110.095 191.695 110.265 191.865 ;
        RECT 113.315 192.375 113.485 192.545 ;
        RECT 61.335 191.185 61.505 191.355 ;
        RECT 61.795 191.185 61.965 191.355 ;
        RECT 62.255 191.185 62.425 191.355 ;
        RECT 62.715 191.185 62.885 191.355 ;
        RECT 63.175 191.185 63.345 191.355 ;
        RECT 63.635 191.185 63.805 191.355 ;
        RECT 64.095 191.185 64.265 191.355 ;
        RECT 64.555 191.185 64.725 191.355 ;
        RECT 65.015 191.185 65.185 191.355 ;
        RECT 65.475 191.185 65.645 191.355 ;
        RECT 65.935 191.185 66.105 191.355 ;
        RECT 66.395 191.185 66.565 191.355 ;
        RECT 66.855 191.185 67.025 191.355 ;
        RECT 67.315 191.185 67.485 191.355 ;
        RECT 67.775 191.185 67.945 191.355 ;
        RECT 68.235 191.185 68.405 191.355 ;
        RECT 68.695 191.185 68.865 191.355 ;
        RECT 69.155 191.185 69.325 191.355 ;
        RECT 69.615 191.185 69.785 191.355 ;
        RECT 70.075 191.185 70.245 191.355 ;
        RECT 70.535 191.185 70.705 191.355 ;
        RECT 70.995 191.185 71.165 191.355 ;
        RECT 71.455 191.185 71.625 191.355 ;
        RECT 71.915 191.185 72.085 191.355 ;
        RECT 72.375 191.185 72.545 191.355 ;
        RECT 72.835 191.185 73.005 191.355 ;
        RECT 73.295 191.185 73.465 191.355 ;
        RECT 73.755 191.185 73.925 191.355 ;
        RECT 74.215 191.185 74.385 191.355 ;
        RECT 74.675 191.185 74.845 191.355 ;
        RECT 75.135 191.185 75.305 191.355 ;
        RECT 75.595 191.185 75.765 191.355 ;
        RECT 76.055 191.185 76.225 191.355 ;
        RECT 76.515 191.185 76.685 191.355 ;
        RECT 76.975 191.185 77.145 191.355 ;
        RECT 77.435 191.185 77.605 191.355 ;
        RECT 77.895 191.185 78.065 191.355 ;
        RECT 78.355 191.185 78.525 191.355 ;
        RECT 78.815 191.185 78.985 191.355 ;
        RECT 79.275 191.185 79.445 191.355 ;
        RECT 79.735 191.185 79.905 191.355 ;
        RECT 80.195 191.185 80.365 191.355 ;
        RECT 80.655 191.185 80.825 191.355 ;
        RECT 81.115 191.185 81.285 191.355 ;
        RECT 81.575 191.185 81.745 191.355 ;
        RECT 82.035 191.185 82.205 191.355 ;
        RECT 82.495 191.185 82.665 191.355 ;
        RECT 82.955 191.185 83.125 191.355 ;
        RECT 83.415 191.185 83.585 191.355 ;
        RECT 83.875 191.185 84.045 191.355 ;
        RECT 84.335 191.185 84.505 191.355 ;
        RECT 84.795 191.185 84.965 191.355 ;
        RECT 85.255 191.185 85.425 191.355 ;
        RECT 85.715 191.185 85.885 191.355 ;
        RECT 86.175 191.185 86.345 191.355 ;
        RECT 86.635 191.185 86.805 191.355 ;
        RECT 87.095 191.185 87.265 191.355 ;
        RECT 87.555 191.185 87.725 191.355 ;
        RECT 88.015 191.185 88.185 191.355 ;
        RECT 88.475 191.185 88.645 191.355 ;
        RECT 88.935 191.185 89.105 191.355 ;
        RECT 89.395 191.185 89.565 191.355 ;
        RECT 89.855 191.185 90.025 191.355 ;
        RECT 90.315 191.185 90.485 191.355 ;
        RECT 90.775 191.185 90.945 191.355 ;
        RECT 91.235 191.185 91.405 191.355 ;
        RECT 91.695 191.185 91.865 191.355 ;
        RECT 92.155 191.185 92.325 191.355 ;
        RECT 92.615 191.185 92.785 191.355 ;
        RECT 93.075 191.185 93.245 191.355 ;
        RECT 93.535 191.185 93.705 191.355 ;
        RECT 93.995 191.185 94.165 191.355 ;
        RECT 94.455 191.185 94.625 191.355 ;
        RECT 94.915 191.185 95.085 191.355 ;
        RECT 95.375 191.185 95.545 191.355 ;
        RECT 95.835 191.185 96.005 191.355 ;
        RECT 96.295 191.185 96.465 191.355 ;
        RECT 96.755 191.185 96.925 191.355 ;
        RECT 97.215 191.185 97.385 191.355 ;
        RECT 97.675 191.185 97.845 191.355 ;
        RECT 98.135 191.185 98.305 191.355 ;
        RECT 98.595 191.185 98.765 191.355 ;
        RECT 99.055 191.185 99.225 191.355 ;
        RECT 99.515 191.185 99.685 191.355 ;
        RECT 99.975 191.185 100.145 191.355 ;
        RECT 100.435 191.185 100.605 191.355 ;
        RECT 100.895 191.185 101.065 191.355 ;
        RECT 101.355 191.185 101.525 191.355 ;
        RECT 101.815 191.185 101.985 191.355 ;
        RECT 102.275 191.185 102.445 191.355 ;
        RECT 102.735 191.185 102.905 191.355 ;
        RECT 103.195 191.185 103.365 191.355 ;
        RECT 103.655 191.185 103.825 191.355 ;
        RECT 104.115 191.185 104.285 191.355 ;
        RECT 104.575 191.185 104.745 191.355 ;
        RECT 105.035 191.185 105.205 191.355 ;
        RECT 105.495 191.185 105.665 191.355 ;
        RECT 105.955 191.185 106.125 191.355 ;
        RECT 106.415 191.185 106.585 191.355 ;
        RECT 106.875 191.185 107.045 191.355 ;
        RECT 107.335 191.185 107.505 191.355 ;
        RECT 107.795 191.185 107.965 191.355 ;
        RECT 108.255 191.185 108.425 191.355 ;
        RECT 108.715 191.185 108.885 191.355 ;
        RECT 109.175 191.185 109.345 191.355 ;
        RECT 109.635 191.185 109.805 191.355 ;
        RECT 110.095 191.185 110.265 191.355 ;
        RECT 110.555 191.185 110.725 191.355 ;
        RECT 111.015 191.185 111.185 191.355 ;
        RECT 111.475 191.185 111.645 191.355 ;
        RECT 111.935 191.185 112.105 191.355 ;
        RECT 112.395 191.185 112.565 191.355 ;
        RECT 112.855 191.185 113.025 191.355 ;
        RECT 113.315 191.185 113.485 191.355 ;
        RECT 113.775 191.185 113.945 191.355 ;
        RECT 114.235 191.185 114.405 191.355 ;
        RECT 114.695 191.185 114.865 191.355 ;
        RECT 115.155 191.185 115.325 191.355 ;
        RECT 72.375 189.995 72.545 190.165 ;
        RECT 73.755 189.995 73.925 190.165 ;
        RECT 71.455 188.975 71.625 189.145 ;
        RECT 74.215 189.995 74.385 190.165 ;
        RECT 73.295 188.975 73.465 189.145 ;
        RECT 74.700 189.315 74.870 189.485 ;
        RECT 75.095 189.655 75.265 189.825 ;
        RECT 75.550 189.995 75.720 190.165 ;
        RECT 76.285 189.655 76.455 189.825 ;
        RECT 76.800 189.315 76.970 189.485 ;
        RECT 78.370 189.315 78.540 189.485 ;
        RECT 78.805 189.655 78.975 189.825 ;
        RECT 82.495 190.675 82.665 190.845 ;
        RECT 81.115 188.975 81.285 189.145 ;
        RECT 85.715 189.655 85.885 189.825 ;
        RECT 87.555 188.975 87.725 189.145 ;
        RECT 92.155 190.675 92.325 190.845 ;
        RECT 90.315 189.995 90.485 190.165 ;
        RECT 95.835 190.675 96.005 190.845 ;
        RECT 95.375 189.655 95.545 189.825 ;
        RECT 96.755 189.655 96.925 189.825 ;
        RECT 97.215 189.995 97.385 190.165 ;
        RECT 97.675 189.995 97.845 190.165 ;
        RECT 98.135 189.655 98.305 189.825 ;
        RECT 99.055 189.995 99.225 190.165 ;
        RECT 99.975 189.995 100.145 190.165 ;
        RECT 100.435 190.675 100.605 190.845 ;
        RECT 100.895 190.335 101.065 190.505 ;
        RECT 101.815 188.975 101.985 189.145 ;
        RECT 103.195 190.675 103.365 190.845 ;
        RECT 109.635 190.675 109.805 190.845 ;
        RECT 107.795 189.995 107.965 190.165 ;
        RECT 108.715 189.995 108.885 190.165 ;
        RECT 106.875 188.975 107.045 189.145 ;
        RECT 110.555 190.335 110.725 190.505 ;
        RECT 111.015 189.995 111.185 190.165 ;
        RECT 111.475 190.675 111.645 190.845 ;
        RECT 112.395 189.315 112.565 189.485 ;
        RECT 61.335 188.465 61.505 188.635 ;
        RECT 61.795 188.465 61.965 188.635 ;
        RECT 62.255 188.465 62.425 188.635 ;
        RECT 62.715 188.465 62.885 188.635 ;
        RECT 63.175 188.465 63.345 188.635 ;
        RECT 63.635 188.465 63.805 188.635 ;
        RECT 64.095 188.465 64.265 188.635 ;
        RECT 64.555 188.465 64.725 188.635 ;
        RECT 65.015 188.465 65.185 188.635 ;
        RECT 65.475 188.465 65.645 188.635 ;
        RECT 65.935 188.465 66.105 188.635 ;
        RECT 66.395 188.465 66.565 188.635 ;
        RECT 66.855 188.465 67.025 188.635 ;
        RECT 67.315 188.465 67.485 188.635 ;
        RECT 67.775 188.465 67.945 188.635 ;
        RECT 68.235 188.465 68.405 188.635 ;
        RECT 68.695 188.465 68.865 188.635 ;
        RECT 69.155 188.465 69.325 188.635 ;
        RECT 69.615 188.465 69.785 188.635 ;
        RECT 70.075 188.465 70.245 188.635 ;
        RECT 70.535 188.465 70.705 188.635 ;
        RECT 70.995 188.465 71.165 188.635 ;
        RECT 71.455 188.465 71.625 188.635 ;
        RECT 71.915 188.465 72.085 188.635 ;
        RECT 72.375 188.465 72.545 188.635 ;
        RECT 72.835 188.465 73.005 188.635 ;
        RECT 73.295 188.465 73.465 188.635 ;
        RECT 73.755 188.465 73.925 188.635 ;
        RECT 74.215 188.465 74.385 188.635 ;
        RECT 74.675 188.465 74.845 188.635 ;
        RECT 75.135 188.465 75.305 188.635 ;
        RECT 75.595 188.465 75.765 188.635 ;
        RECT 76.055 188.465 76.225 188.635 ;
        RECT 76.515 188.465 76.685 188.635 ;
        RECT 76.975 188.465 77.145 188.635 ;
        RECT 77.435 188.465 77.605 188.635 ;
        RECT 77.895 188.465 78.065 188.635 ;
        RECT 78.355 188.465 78.525 188.635 ;
        RECT 78.815 188.465 78.985 188.635 ;
        RECT 79.275 188.465 79.445 188.635 ;
        RECT 79.735 188.465 79.905 188.635 ;
        RECT 80.195 188.465 80.365 188.635 ;
        RECT 80.655 188.465 80.825 188.635 ;
        RECT 81.115 188.465 81.285 188.635 ;
        RECT 81.575 188.465 81.745 188.635 ;
        RECT 82.035 188.465 82.205 188.635 ;
        RECT 82.495 188.465 82.665 188.635 ;
        RECT 82.955 188.465 83.125 188.635 ;
        RECT 83.415 188.465 83.585 188.635 ;
        RECT 83.875 188.465 84.045 188.635 ;
        RECT 84.335 188.465 84.505 188.635 ;
        RECT 84.795 188.465 84.965 188.635 ;
        RECT 85.255 188.465 85.425 188.635 ;
        RECT 85.715 188.465 85.885 188.635 ;
        RECT 86.175 188.465 86.345 188.635 ;
        RECT 86.635 188.465 86.805 188.635 ;
        RECT 87.095 188.465 87.265 188.635 ;
        RECT 87.555 188.465 87.725 188.635 ;
        RECT 88.015 188.465 88.185 188.635 ;
        RECT 88.475 188.465 88.645 188.635 ;
        RECT 88.935 188.465 89.105 188.635 ;
        RECT 89.395 188.465 89.565 188.635 ;
        RECT 89.855 188.465 90.025 188.635 ;
        RECT 90.315 188.465 90.485 188.635 ;
        RECT 90.775 188.465 90.945 188.635 ;
        RECT 91.235 188.465 91.405 188.635 ;
        RECT 91.695 188.465 91.865 188.635 ;
        RECT 92.155 188.465 92.325 188.635 ;
        RECT 92.615 188.465 92.785 188.635 ;
        RECT 93.075 188.465 93.245 188.635 ;
        RECT 93.535 188.465 93.705 188.635 ;
        RECT 93.995 188.465 94.165 188.635 ;
        RECT 94.455 188.465 94.625 188.635 ;
        RECT 94.915 188.465 95.085 188.635 ;
        RECT 95.375 188.465 95.545 188.635 ;
        RECT 95.835 188.465 96.005 188.635 ;
        RECT 96.295 188.465 96.465 188.635 ;
        RECT 96.755 188.465 96.925 188.635 ;
        RECT 97.215 188.465 97.385 188.635 ;
        RECT 97.675 188.465 97.845 188.635 ;
        RECT 98.135 188.465 98.305 188.635 ;
        RECT 98.595 188.465 98.765 188.635 ;
        RECT 99.055 188.465 99.225 188.635 ;
        RECT 99.515 188.465 99.685 188.635 ;
        RECT 99.975 188.465 100.145 188.635 ;
        RECT 100.435 188.465 100.605 188.635 ;
        RECT 100.895 188.465 101.065 188.635 ;
        RECT 101.355 188.465 101.525 188.635 ;
        RECT 101.815 188.465 101.985 188.635 ;
        RECT 102.275 188.465 102.445 188.635 ;
        RECT 102.735 188.465 102.905 188.635 ;
        RECT 103.195 188.465 103.365 188.635 ;
        RECT 103.655 188.465 103.825 188.635 ;
        RECT 104.115 188.465 104.285 188.635 ;
        RECT 104.575 188.465 104.745 188.635 ;
        RECT 105.035 188.465 105.205 188.635 ;
        RECT 105.495 188.465 105.665 188.635 ;
        RECT 105.955 188.465 106.125 188.635 ;
        RECT 106.415 188.465 106.585 188.635 ;
        RECT 106.875 188.465 107.045 188.635 ;
        RECT 107.335 188.465 107.505 188.635 ;
        RECT 107.795 188.465 107.965 188.635 ;
        RECT 108.255 188.465 108.425 188.635 ;
        RECT 108.715 188.465 108.885 188.635 ;
        RECT 109.175 188.465 109.345 188.635 ;
        RECT 109.635 188.465 109.805 188.635 ;
        RECT 110.095 188.465 110.265 188.635 ;
        RECT 110.555 188.465 110.725 188.635 ;
        RECT 111.015 188.465 111.185 188.635 ;
        RECT 111.475 188.465 111.645 188.635 ;
        RECT 111.935 188.465 112.105 188.635 ;
        RECT 112.395 188.465 112.565 188.635 ;
        RECT 112.855 188.465 113.025 188.635 ;
        RECT 113.315 188.465 113.485 188.635 ;
        RECT 113.775 188.465 113.945 188.635 ;
        RECT 114.235 188.465 114.405 188.635 ;
        RECT 114.695 188.465 114.865 188.635 ;
        RECT 115.155 188.465 115.325 188.635 ;
        RECT 67.315 187.275 67.485 187.445 ;
        RECT 70.075 186.595 70.245 186.765 ;
        RECT 70.535 187.955 70.705 188.125 ;
        RECT 73.755 187.275 73.925 187.445 ;
        RECT 75.595 187.955 75.765 188.125 ;
        RECT 74.675 186.595 74.845 186.765 ;
        RECT 75.755 186.595 75.925 186.765 ;
        RECT 77.460 187.615 77.630 187.785 ;
        RECT 76.975 186.935 77.145 187.105 ;
        RECT 76.515 186.255 76.685 186.425 ;
        RECT 77.855 187.275 78.025 187.445 ;
        RECT 78.255 186.935 78.425 187.105 ;
        RECT 79.560 187.615 79.730 187.785 ;
        RECT 79.045 187.275 79.215 187.445 ;
        RECT 81.130 187.615 81.300 187.785 ;
        RECT 81.565 187.275 81.735 187.445 ;
        RECT 85.715 187.955 85.885 188.125 ;
        RECT 87.120 187.615 87.290 187.785 ;
        RECT 84.335 186.935 84.505 187.105 ;
        RECT 83.875 186.255 84.045 186.425 ;
        RECT 84.795 186.255 84.965 186.425 ;
        RECT 85.715 186.935 85.885 187.105 ;
        RECT 86.635 186.935 86.805 187.105 ;
        RECT 87.515 187.275 87.685 187.445 ;
        RECT 87.970 186.935 88.140 187.105 ;
        RECT 89.220 187.615 89.390 187.785 ;
        RECT 88.705 187.275 88.875 187.445 ;
        RECT 90.790 187.615 90.960 187.785 ;
        RECT 91.225 187.275 91.395 187.445 ;
        RECT 93.535 187.955 93.705 188.125 ;
        RECT 95.375 187.955 95.545 188.125 ;
        RECT 93.995 186.935 94.165 187.105 ;
        RECT 94.455 186.255 94.625 186.425 ;
        RECT 96.755 186.935 96.925 187.105 ;
        RECT 95.375 186.595 95.545 186.765 ;
        RECT 99.515 187.955 99.685 188.125 ;
        RECT 105.035 187.955 105.205 188.125 ;
        RECT 103.195 186.935 103.365 187.105 ;
        RECT 104.575 187.275 104.745 187.445 ;
        RECT 105.035 186.935 105.205 187.105 ;
        RECT 105.955 186.935 106.125 187.105 ;
        RECT 106.415 186.255 106.585 186.425 ;
        RECT 109.635 187.275 109.805 187.445 ;
        RECT 110.555 186.935 110.725 187.105 ;
        RECT 113.315 186.255 113.485 186.425 ;
        RECT 61.335 185.745 61.505 185.915 ;
        RECT 61.795 185.745 61.965 185.915 ;
        RECT 62.255 185.745 62.425 185.915 ;
        RECT 62.715 185.745 62.885 185.915 ;
        RECT 63.175 185.745 63.345 185.915 ;
        RECT 63.635 185.745 63.805 185.915 ;
        RECT 64.095 185.745 64.265 185.915 ;
        RECT 64.555 185.745 64.725 185.915 ;
        RECT 65.015 185.745 65.185 185.915 ;
        RECT 65.475 185.745 65.645 185.915 ;
        RECT 65.935 185.745 66.105 185.915 ;
        RECT 66.395 185.745 66.565 185.915 ;
        RECT 66.855 185.745 67.025 185.915 ;
        RECT 67.315 185.745 67.485 185.915 ;
        RECT 67.775 185.745 67.945 185.915 ;
        RECT 68.235 185.745 68.405 185.915 ;
        RECT 68.695 185.745 68.865 185.915 ;
        RECT 69.155 185.745 69.325 185.915 ;
        RECT 69.615 185.745 69.785 185.915 ;
        RECT 70.075 185.745 70.245 185.915 ;
        RECT 70.535 185.745 70.705 185.915 ;
        RECT 70.995 185.745 71.165 185.915 ;
        RECT 71.455 185.745 71.625 185.915 ;
        RECT 71.915 185.745 72.085 185.915 ;
        RECT 72.375 185.745 72.545 185.915 ;
        RECT 72.835 185.745 73.005 185.915 ;
        RECT 73.295 185.745 73.465 185.915 ;
        RECT 73.755 185.745 73.925 185.915 ;
        RECT 74.215 185.745 74.385 185.915 ;
        RECT 74.675 185.745 74.845 185.915 ;
        RECT 75.135 185.745 75.305 185.915 ;
        RECT 75.595 185.745 75.765 185.915 ;
        RECT 76.055 185.745 76.225 185.915 ;
        RECT 76.515 185.745 76.685 185.915 ;
        RECT 76.975 185.745 77.145 185.915 ;
        RECT 77.435 185.745 77.605 185.915 ;
        RECT 77.895 185.745 78.065 185.915 ;
        RECT 78.355 185.745 78.525 185.915 ;
        RECT 78.815 185.745 78.985 185.915 ;
        RECT 79.275 185.745 79.445 185.915 ;
        RECT 79.735 185.745 79.905 185.915 ;
        RECT 80.195 185.745 80.365 185.915 ;
        RECT 80.655 185.745 80.825 185.915 ;
        RECT 81.115 185.745 81.285 185.915 ;
        RECT 81.575 185.745 81.745 185.915 ;
        RECT 82.035 185.745 82.205 185.915 ;
        RECT 82.495 185.745 82.665 185.915 ;
        RECT 82.955 185.745 83.125 185.915 ;
        RECT 83.415 185.745 83.585 185.915 ;
        RECT 83.875 185.745 84.045 185.915 ;
        RECT 84.335 185.745 84.505 185.915 ;
        RECT 84.795 185.745 84.965 185.915 ;
        RECT 85.255 185.745 85.425 185.915 ;
        RECT 85.715 185.745 85.885 185.915 ;
        RECT 86.175 185.745 86.345 185.915 ;
        RECT 86.635 185.745 86.805 185.915 ;
        RECT 87.095 185.745 87.265 185.915 ;
        RECT 87.555 185.745 87.725 185.915 ;
        RECT 88.015 185.745 88.185 185.915 ;
        RECT 88.475 185.745 88.645 185.915 ;
        RECT 88.935 185.745 89.105 185.915 ;
        RECT 89.395 185.745 89.565 185.915 ;
        RECT 89.855 185.745 90.025 185.915 ;
        RECT 90.315 185.745 90.485 185.915 ;
        RECT 90.775 185.745 90.945 185.915 ;
        RECT 91.235 185.745 91.405 185.915 ;
        RECT 91.695 185.745 91.865 185.915 ;
        RECT 92.155 185.745 92.325 185.915 ;
        RECT 92.615 185.745 92.785 185.915 ;
        RECT 93.075 185.745 93.245 185.915 ;
        RECT 93.535 185.745 93.705 185.915 ;
        RECT 93.995 185.745 94.165 185.915 ;
        RECT 94.455 185.745 94.625 185.915 ;
        RECT 94.915 185.745 95.085 185.915 ;
        RECT 95.375 185.745 95.545 185.915 ;
        RECT 95.835 185.745 96.005 185.915 ;
        RECT 96.295 185.745 96.465 185.915 ;
        RECT 96.755 185.745 96.925 185.915 ;
        RECT 97.215 185.745 97.385 185.915 ;
        RECT 97.675 185.745 97.845 185.915 ;
        RECT 98.135 185.745 98.305 185.915 ;
        RECT 98.595 185.745 98.765 185.915 ;
        RECT 99.055 185.745 99.225 185.915 ;
        RECT 99.515 185.745 99.685 185.915 ;
        RECT 99.975 185.745 100.145 185.915 ;
        RECT 100.435 185.745 100.605 185.915 ;
        RECT 100.895 185.745 101.065 185.915 ;
        RECT 101.355 185.745 101.525 185.915 ;
        RECT 101.815 185.745 101.985 185.915 ;
        RECT 102.275 185.745 102.445 185.915 ;
        RECT 102.735 185.745 102.905 185.915 ;
        RECT 103.195 185.745 103.365 185.915 ;
        RECT 103.655 185.745 103.825 185.915 ;
        RECT 104.115 185.745 104.285 185.915 ;
        RECT 104.575 185.745 104.745 185.915 ;
        RECT 105.035 185.745 105.205 185.915 ;
        RECT 105.495 185.745 105.665 185.915 ;
        RECT 105.955 185.745 106.125 185.915 ;
        RECT 106.415 185.745 106.585 185.915 ;
        RECT 106.875 185.745 107.045 185.915 ;
        RECT 107.335 185.745 107.505 185.915 ;
        RECT 107.795 185.745 107.965 185.915 ;
        RECT 108.255 185.745 108.425 185.915 ;
        RECT 108.715 185.745 108.885 185.915 ;
        RECT 109.175 185.745 109.345 185.915 ;
        RECT 109.635 185.745 109.805 185.915 ;
        RECT 110.095 185.745 110.265 185.915 ;
        RECT 110.555 185.745 110.725 185.915 ;
        RECT 111.015 185.745 111.185 185.915 ;
        RECT 111.475 185.745 111.645 185.915 ;
        RECT 111.935 185.745 112.105 185.915 ;
        RECT 112.395 185.745 112.565 185.915 ;
        RECT 112.855 185.745 113.025 185.915 ;
        RECT 113.315 185.745 113.485 185.915 ;
        RECT 113.775 185.745 113.945 185.915 ;
        RECT 114.235 185.745 114.405 185.915 ;
        RECT 114.695 185.745 114.865 185.915 ;
        RECT 115.155 185.745 115.325 185.915 ;
        RECT 69.615 184.555 69.785 184.725 ;
        RECT 70.100 183.875 70.270 184.045 ;
        RECT 70.495 184.215 70.665 184.385 ;
        RECT 70.950 184.555 71.120 184.725 ;
        RECT 71.685 184.215 71.855 184.385 ;
        RECT 72.200 183.875 72.370 184.045 ;
        RECT 73.770 183.875 73.940 184.045 ;
        RECT 74.205 184.215 74.375 184.385 ;
        RECT 76.515 185.235 76.685 185.405 ;
        RECT 76.975 184.215 77.145 184.385 ;
        RECT 77.460 183.875 77.630 184.045 ;
        RECT 77.855 184.215 78.025 184.385 ;
        RECT 78.310 184.555 78.480 184.725 ;
        RECT 79.045 184.215 79.215 184.385 ;
        RECT 79.560 183.875 79.730 184.045 ;
        RECT 81.130 183.875 81.300 184.045 ;
        RECT 81.565 184.215 81.735 184.385 ;
        RECT 84.335 184.555 84.505 184.725 ;
        RECT 85.255 184.555 85.425 184.725 ;
        RECT 83.875 183.875 84.045 184.045 ;
        RECT 85.255 183.535 85.425 183.705 ;
        RECT 88.935 184.555 89.105 184.725 ;
        RECT 89.855 184.555 90.025 184.725 ;
        RECT 90.315 184.215 90.485 184.385 ;
        RECT 89.855 183.875 90.025 184.045 ;
        RECT 90.800 183.875 90.970 184.045 ;
        RECT 91.195 184.215 91.365 184.385 ;
        RECT 91.650 184.555 91.820 184.725 ;
        RECT 92.385 184.215 92.555 184.385 ;
        RECT 92.900 183.875 93.070 184.045 ;
        RECT 94.470 183.875 94.640 184.045 ;
        RECT 94.905 184.215 95.075 184.385 ;
        RECT 97.675 184.215 97.845 184.385 ;
        RECT 97.215 183.535 97.385 183.705 ;
        RECT 98.160 183.875 98.330 184.045 ;
        RECT 98.555 184.215 98.725 184.385 ;
        RECT 99.010 184.555 99.180 184.725 ;
        RECT 99.745 184.215 99.915 184.385 ;
        RECT 100.260 183.875 100.430 184.045 ;
        RECT 101.830 183.875 102.000 184.045 ;
        RECT 102.265 184.215 102.435 184.385 ;
        RECT 104.575 185.235 104.745 185.405 ;
        RECT 105.035 184.215 105.205 184.385 ;
        RECT 105.520 183.875 105.690 184.045 ;
        RECT 105.915 184.215 106.085 184.385 ;
        RECT 106.370 184.555 106.540 184.725 ;
        RECT 107.105 184.215 107.275 184.385 ;
        RECT 107.620 183.875 107.790 184.045 ;
        RECT 109.190 183.875 109.360 184.045 ;
        RECT 109.625 184.215 109.795 184.385 ;
        RECT 111.935 185.235 112.105 185.405 ;
        RECT 61.335 183.025 61.505 183.195 ;
        RECT 61.795 183.025 61.965 183.195 ;
        RECT 62.255 183.025 62.425 183.195 ;
        RECT 62.715 183.025 62.885 183.195 ;
        RECT 63.175 183.025 63.345 183.195 ;
        RECT 63.635 183.025 63.805 183.195 ;
        RECT 64.095 183.025 64.265 183.195 ;
        RECT 64.555 183.025 64.725 183.195 ;
        RECT 65.015 183.025 65.185 183.195 ;
        RECT 65.475 183.025 65.645 183.195 ;
        RECT 65.935 183.025 66.105 183.195 ;
        RECT 66.395 183.025 66.565 183.195 ;
        RECT 66.855 183.025 67.025 183.195 ;
        RECT 67.315 183.025 67.485 183.195 ;
        RECT 67.775 183.025 67.945 183.195 ;
        RECT 68.235 183.025 68.405 183.195 ;
        RECT 68.695 183.025 68.865 183.195 ;
        RECT 69.155 183.025 69.325 183.195 ;
        RECT 69.615 183.025 69.785 183.195 ;
        RECT 70.075 183.025 70.245 183.195 ;
        RECT 70.535 183.025 70.705 183.195 ;
        RECT 70.995 183.025 71.165 183.195 ;
        RECT 71.455 183.025 71.625 183.195 ;
        RECT 71.915 183.025 72.085 183.195 ;
        RECT 72.375 183.025 72.545 183.195 ;
        RECT 72.835 183.025 73.005 183.195 ;
        RECT 73.295 183.025 73.465 183.195 ;
        RECT 73.755 183.025 73.925 183.195 ;
        RECT 74.215 183.025 74.385 183.195 ;
        RECT 74.675 183.025 74.845 183.195 ;
        RECT 75.135 183.025 75.305 183.195 ;
        RECT 75.595 183.025 75.765 183.195 ;
        RECT 76.055 183.025 76.225 183.195 ;
        RECT 76.515 183.025 76.685 183.195 ;
        RECT 76.975 183.025 77.145 183.195 ;
        RECT 77.435 183.025 77.605 183.195 ;
        RECT 77.895 183.025 78.065 183.195 ;
        RECT 78.355 183.025 78.525 183.195 ;
        RECT 78.815 183.025 78.985 183.195 ;
        RECT 79.275 183.025 79.445 183.195 ;
        RECT 79.735 183.025 79.905 183.195 ;
        RECT 80.195 183.025 80.365 183.195 ;
        RECT 80.655 183.025 80.825 183.195 ;
        RECT 81.115 183.025 81.285 183.195 ;
        RECT 81.575 183.025 81.745 183.195 ;
        RECT 82.035 183.025 82.205 183.195 ;
        RECT 82.495 183.025 82.665 183.195 ;
        RECT 82.955 183.025 83.125 183.195 ;
        RECT 83.415 183.025 83.585 183.195 ;
        RECT 83.875 183.025 84.045 183.195 ;
        RECT 84.335 183.025 84.505 183.195 ;
        RECT 84.795 183.025 84.965 183.195 ;
        RECT 85.255 183.025 85.425 183.195 ;
        RECT 85.715 183.025 85.885 183.195 ;
        RECT 86.175 183.025 86.345 183.195 ;
        RECT 86.635 183.025 86.805 183.195 ;
        RECT 87.095 183.025 87.265 183.195 ;
        RECT 87.555 183.025 87.725 183.195 ;
        RECT 88.015 183.025 88.185 183.195 ;
        RECT 88.475 183.025 88.645 183.195 ;
        RECT 88.935 183.025 89.105 183.195 ;
        RECT 89.395 183.025 89.565 183.195 ;
        RECT 89.855 183.025 90.025 183.195 ;
        RECT 90.315 183.025 90.485 183.195 ;
        RECT 90.775 183.025 90.945 183.195 ;
        RECT 91.235 183.025 91.405 183.195 ;
        RECT 91.695 183.025 91.865 183.195 ;
        RECT 92.155 183.025 92.325 183.195 ;
        RECT 92.615 183.025 92.785 183.195 ;
        RECT 93.075 183.025 93.245 183.195 ;
        RECT 93.535 183.025 93.705 183.195 ;
        RECT 93.995 183.025 94.165 183.195 ;
        RECT 94.455 183.025 94.625 183.195 ;
        RECT 94.915 183.025 95.085 183.195 ;
        RECT 95.375 183.025 95.545 183.195 ;
        RECT 95.835 183.025 96.005 183.195 ;
        RECT 96.295 183.025 96.465 183.195 ;
        RECT 96.755 183.025 96.925 183.195 ;
        RECT 97.215 183.025 97.385 183.195 ;
        RECT 97.675 183.025 97.845 183.195 ;
        RECT 98.135 183.025 98.305 183.195 ;
        RECT 98.595 183.025 98.765 183.195 ;
        RECT 99.055 183.025 99.225 183.195 ;
        RECT 99.515 183.025 99.685 183.195 ;
        RECT 99.975 183.025 100.145 183.195 ;
        RECT 100.435 183.025 100.605 183.195 ;
        RECT 100.895 183.025 101.065 183.195 ;
        RECT 101.355 183.025 101.525 183.195 ;
        RECT 101.815 183.025 101.985 183.195 ;
        RECT 102.275 183.025 102.445 183.195 ;
        RECT 102.735 183.025 102.905 183.195 ;
        RECT 103.195 183.025 103.365 183.195 ;
        RECT 103.655 183.025 103.825 183.195 ;
        RECT 104.115 183.025 104.285 183.195 ;
        RECT 104.575 183.025 104.745 183.195 ;
        RECT 105.035 183.025 105.205 183.195 ;
        RECT 105.495 183.025 105.665 183.195 ;
        RECT 105.955 183.025 106.125 183.195 ;
        RECT 106.415 183.025 106.585 183.195 ;
        RECT 106.875 183.025 107.045 183.195 ;
        RECT 107.335 183.025 107.505 183.195 ;
        RECT 107.795 183.025 107.965 183.195 ;
        RECT 108.255 183.025 108.425 183.195 ;
        RECT 108.715 183.025 108.885 183.195 ;
        RECT 109.175 183.025 109.345 183.195 ;
        RECT 109.635 183.025 109.805 183.195 ;
        RECT 110.095 183.025 110.265 183.195 ;
        RECT 110.555 183.025 110.725 183.195 ;
        RECT 111.015 183.025 111.185 183.195 ;
        RECT 111.475 183.025 111.645 183.195 ;
        RECT 111.935 183.025 112.105 183.195 ;
        RECT 112.395 183.025 112.565 183.195 ;
        RECT 112.855 183.025 113.025 183.195 ;
        RECT 113.315 183.025 113.485 183.195 ;
        RECT 113.775 183.025 113.945 183.195 ;
        RECT 114.235 183.025 114.405 183.195 ;
        RECT 114.695 183.025 114.865 183.195 ;
        RECT 115.155 183.025 115.325 183.195 ;
        RECT 76.975 182.515 77.145 182.685 ;
        RECT 79.275 182.515 79.445 182.685 ;
        RECT 76.975 181.155 77.145 181.325 ;
        RECT 78.355 181.495 78.525 181.665 ;
        RECT 81.115 182.175 81.285 182.345 ;
        RECT 77.895 180.815 78.065 180.985 ;
        RECT 80.195 181.495 80.365 181.665 ;
        RECT 81.575 181.495 81.745 181.665 ;
        RECT 82.955 181.495 83.125 181.665 ;
        RECT 88.040 182.175 88.210 182.345 ;
        RECT 85.715 181.495 85.885 181.665 ;
        RECT 87.555 181.835 87.725 182.005 ;
        RECT 88.435 181.835 88.605 182.005 ;
        RECT 88.890 181.495 89.060 181.665 ;
        RECT 90.140 182.175 90.310 182.345 ;
        RECT 89.625 181.835 89.795 182.005 ;
        RECT 91.710 182.175 91.880 182.345 ;
        RECT 92.145 181.835 92.315 182.005 ;
        RECT 94.455 182.175 94.625 182.345 ;
        RECT 96.295 181.835 96.465 182.005 ;
        RECT 99.055 182.515 99.225 182.685 ;
        RECT 101.815 182.175 101.985 182.345 ;
        RECT 103.195 182.515 103.365 182.685 ;
        RECT 102.735 181.495 102.905 181.665 ;
        RECT 105.955 182.515 106.125 182.685 ;
        RECT 105.495 181.835 105.665 182.005 ;
        RECT 104.115 181.495 104.285 181.665 ;
        RECT 105.035 181.495 105.205 181.665 ;
        RECT 108.265 181.835 108.435 182.005 ;
        RECT 108.700 182.175 108.870 182.345 ;
        RECT 110.270 182.175 110.440 182.345 ;
        RECT 110.785 181.835 110.955 182.005 ;
        RECT 111.630 181.155 111.800 181.325 ;
        RECT 111.975 181.835 112.145 182.005 ;
        RECT 112.370 182.175 112.540 182.345 ;
        RECT 112.855 181.495 113.025 181.665 ;
        RECT 61.335 180.305 61.505 180.475 ;
        RECT 61.795 180.305 61.965 180.475 ;
        RECT 62.255 180.305 62.425 180.475 ;
        RECT 62.715 180.305 62.885 180.475 ;
        RECT 63.175 180.305 63.345 180.475 ;
        RECT 63.635 180.305 63.805 180.475 ;
        RECT 64.095 180.305 64.265 180.475 ;
        RECT 64.555 180.305 64.725 180.475 ;
        RECT 65.015 180.305 65.185 180.475 ;
        RECT 65.475 180.305 65.645 180.475 ;
        RECT 65.935 180.305 66.105 180.475 ;
        RECT 66.395 180.305 66.565 180.475 ;
        RECT 66.855 180.305 67.025 180.475 ;
        RECT 67.315 180.305 67.485 180.475 ;
        RECT 67.775 180.305 67.945 180.475 ;
        RECT 68.235 180.305 68.405 180.475 ;
        RECT 68.695 180.305 68.865 180.475 ;
        RECT 69.155 180.305 69.325 180.475 ;
        RECT 69.615 180.305 69.785 180.475 ;
        RECT 70.075 180.305 70.245 180.475 ;
        RECT 70.535 180.305 70.705 180.475 ;
        RECT 70.995 180.305 71.165 180.475 ;
        RECT 71.455 180.305 71.625 180.475 ;
        RECT 71.915 180.305 72.085 180.475 ;
        RECT 72.375 180.305 72.545 180.475 ;
        RECT 72.835 180.305 73.005 180.475 ;
        RECT 73.295 180.305 73.465 180.475 ;
        RECT 73.755 180.305 73.925 180.475 ;
        RECT 74.215 180.305 74.385 180.475 ;
        RECT 74.675 180.305 74.845 180.475 ;
        RECT 75.135 180.305 75.305 180.475 ;
        RECT 75.595 180.305 75.765 180.475 ;
        RECT 76.055 180.305 76.225 180.475 ;
        RECT 76.515 180.305 76.685 180.475 ;
        RECT 76.975 180.305 77.145 180.475 ;
        RECT 77.435 180.305 77.605 180.475 ;
        RECT 77.895 180.305 78.065 180.475 ;
        RECT 78.355 180.305 78.525 180.475 ;
        RECT 78.815 180.305 78.985 180.475 ;
        RECT 79.275 180.305 79.445 180.475 ;
        RECT 79.735 180.305 79.905 180.475 ;
        RECT 80.195 180.305 80.365 180.475 ;
        RECT 80.655 180.305 80.825 180.475 ;
        RECT 81.115 180.305 81.285 180.475 ;
        RECT 81.575 180.305 81.745 180.475 ;
        RECT 82.035 180.305 82.205 180.475 ;
        RECT 82.495 180.305 82.665 180.475 ;
        RECT 82.955 180.305 83.125 180.475 ;
        RECT 83.415 180.305 83.585 180.475 ;
        RECT 83.875 180.305 84.045 180.475 ;
        RECT 84.335 180.305 84.505 180.475 ;
        RECT 84.795 180.305 84.965 180.475 ;
        RECT 85.255 180.305 85.425 180.475 ;
        RECT 85.715 180.305 85.885 180.475 ;
        RECT 86.175 180.305 86.345 180.475 ;
        RECT 86.635 180.305 86.805 180.475 ;
        RECT 87.095 180.305 87.265 180.475 ;
        RECT 87.555 180.305 87.725 180.475 ;
        RECT 88.015 180.305 88.185 180.475 ;
        RECT 88.475 180.305 88.645 180.475 ;
        RECT 88.935 180.305 89.105 180.475 ;
        RECT 89.395 180.305 89.565 180.475 ;
        RECT 89.855 180.305 90.025 180.475 ;
        RECT 90.315 180.305 90.485 180.475 ;
        RECT 90.775 180.305 90.945 180.475 ;
        RECT 91.235 180.305 91.405 180.475 ;
        RECT 91.695 180.305 91.865 180.475 ;
        RECT 92.155 180.305 92.325 180.475 ;
        RECT 92.615 180.305 92.785 180.475 ;
        RECT 93.075 180.305 93.245 180.475 ;
        RECT 93.535 180.305 93.705 180.475 ;
        RECT 93.995 180.305 94.165 180.475 ;
        RECT 94.455 180.305 94.625 180.475 ;
        RECT 94.915 180.305 95.085 180.475 ;
        RECT 95.375 180.305 95.545 180.475 ;
        RECT 95.835 180.305 96.005 180.475 ;
        RECT 96.295 180.305 96.465 180.475 ;
        RECT 96.755 180.305 96.925 180.475 ;
        RECT 97.215 180.305 97.385 180.475 ;
        RECT 97.675 180.305 97.845 180.475 ;
        RECT 98.135 180.305 98.305 180.475 ;
        RECT 98.595 180.305 98.765 180.475 ;
        RECT 99.055 180.305 99.225 180.475 ;
        RECT 99.515 180.305 99.685 180.475 ;
        RECT 99.975 180.305 100.145 180.475 ;
        RECT 100.435 180.305 100.605 180.475 ;
        RECT 100.895 180.305 101.065 180.475 ;
        RECT 101.355 180.305 101.525 180.475 ;
        RECT 101.815 180.305 101.985 180.475 ;
        RECT 102.275 180.305 102.445 180.475 ;
        RECT 102.735 180.305 102.905 180.475 ;
        RECT 103.195 180.305 103.365 180.475 ;
        RECT 103.655 180.305 103.825 180.475 ;
        RECT 104.115 180.305 104.285 180.475 ;
        RECT 104.575 180.305 104.745 180.475 ;
        RECT 105.035 180.305 105.205 180.475 ;
        RECT 105.495 180.305 105.665 180.475 ;
        RECT 105.955 180.305 106.125 180.475 ;
        RECT 106.415 180.305 106.585 180.475 ;
        RECT 106.875 180.305 107.045 180.475 ;
        RECT 107.335 180.305 107.505 180.475 ;
        RECT 107.795 180.305 107.965 180.475 ;
        RECT 108.255 180.305 108.425 180.475 ;
        RECT 108.715 180.305 108.885 180.475 ;
        RECT 109.175 180.305 109.345 180.475 ;
        RECT 109.635 180.305 109.805 180.475 ;
        RECT 110.095 180.305 110.265 180.475 ;
        RECT 110.555 180.305 110.725 180.475 ;
        RECT 111.015 180.305 111.185 180.475 ;
        RECT 111.475 180.305 111.645 180.475 ;
        RECT 111.935 180.305 112.105 180.475 ;
        RECT 112.395 180.305 112.565 180.475 ;
        RECT 112.855 180.305 113.025 180.475 ;
        RECT 113.315 180.305 113.485 180.475 ;
        RECT 113.775 180.305 113.945 180.475 ;
        RECT 114.235 180.305 114.405 180.475 ;
        RECT 114.695 180.305 114.865 180.475 ;
        RECT 115.155 180.305 115.325 180.475 ;
        RECT 96.755 179.795 96.925 179.965 ;
        RECT 95.375 179.115 95.545 179.285 ;
        RECT 95.835 179.115 96.005 179.285 ;
        RECT 102.275 179.795 102.445 179.965 ;
        RECT 104.575 179.795 104.745 179.965 ;
        RECT 101.815 179.115 101.985 179.285 ;
        RECT 102.735 179.115 102.905 179.285 ;
        RECT 104.115 179.115 104.285 179.285 ;
        RECT 105.495 179.115 105.665 179.285 ;
        RECT 105.495 178.435 105.665 178.605 ;
        RECT 107.795 179.115 107.965 179.285 ;
        RECT 110.555 179.115 110.725 179.285 ;
        RECT 111.015 179.115 111.185 179.285 ;
        RECT 111.935 179.795 112.105 179.965 ;
        RECT 112.395 179.115 112.565 179.285 ;
        RECT 111.015 178.435 111.185 178.605 ;
        RECT 61.335 177.585 61.505 177.755 ;
        RECT 61.795 177.585 61.965 177.755 ;
        RECT 62.255 177.585 62.425 177.755 ;
        RECT 62.715 177.585 62.885 177.755 ;
        RECT 63.175 177.585 63.345 177.755 ;
        RECT 63.635 177.585 63.805 177.755 ;
        RECT 64.095 177.585 64.265 177.755 ;
        RECT 64.555 177.585 64.725 177.755 ;
        RECT 65.015 177.585 65.185 177.755 ;
        RECT 65.475 177.585 65.645 177.755 ;
        RECT 65.935 177.585 66.105 177.755 ;
        RECT 66.395 177.585 66.565 177.755 ;
        RECT 66.855 177.585 67.025 177.755 ;
        RECT 67.315 177.585 67.485 177.755 ;
        RECT 67.775 177.585 67.945 177.755 ;
        RECT 68.235 177.585 68.405 177.755 ;
        RECT 68.695 177.585 68.865 177.755 ;
        RECT 69.155 177.585 69.325 177.755 ;
        RECT 69.615 177.585 69.785 177.755 ;
        RECT 70.075 177.585 70.245 177.755 ;
        RECT 70.535 177.585 70.705 177.755 ;
        RECT 70.995 177.585 71.165 177.755 ;
        RECT 71.455 177.585 71.625 177.755 ;
        RECT 71.915 177.585 72.085 177.755 ;
        RECT 72.375 177.585 72.545 177.755 ;
        RECT 72.835 177.585 73.005 177.755 ;
        RECT 73.295 177.585 73.465 177.755 ;
        RECT 73.755 177.585 73.925 177.755 ;
        RECT 74.215 177.585 74.385 177.755 ;
        RECT 74.675 177.585 74.845 177.755 ;
        RECT 75.135 177.585 75.305 177.755 ;
        RECT 75.595 177.585 75.765 177.755 ;
        RECT 76.055 177.585 76.225 177.755 ;
        RECT 76.515 177.585 76.685 177.755 ;
        RECT 76.975 177.585 77.145 177.755 ;
        RECT 77.435 177.585 77.605 177.755 ;
        RECT 77.895 177.585 78.065 177.755 ;
        RECT 78.355 177.585 78.525 177.755 ;
        RECT 78.815 177.585 78.985 177.755 ;
        RECT 79.275 177.585 79.445 177.755 ;
        RECT 79.735 177.585 79.905 177.755 ;
        RECT 80.195 177.585 80.365 177.755 ;
        RECT 80.655 177.585 80.825 177.755 ;
        RECT 81.115 177.585 81.285 177.755 ;
        RECT 81.575 177.585 81.745 177.755 ;
        RECT 82.035 177.585 82.205 177.755 ;
        RECT 82.495 177.585 82.665 177.755 ;
        RECT 82.955 177.585 83.125 177.755 ;
        RECT 83.415 177.585 83.585 177.755 ;
        RECT 83.875 177.585 84.045 177.755 ;
        RECT 84.335 177.585 84.505 177.755 ;
        RECT 84.795 177.585 84.965 177.755 ;
        RECT 85.255 177.585 85.425 177.755 ;
        RECT 85.715 177.585 85.885 177.755 ;
        RECT 86.175 177.585 86.345 177.755 ;
        RECT 86.635 177.585 86.805 177.755 ;
        RECT 87.095 177.585 87.265 177.755 ;
        RECT 87.555 177.585 87.725 177.755 ;
        RECT 88.015 177.585 88.185 177.755 ;
        RECT 88.475 177.585 88.645 177.755 ;
        RECT 88.935 177.585 89.105 177.755 ;
        RECT 89.395 177.585 89.565 177.755 ;
        RECT 89.855 177.585 90.025 177.755 ;
        RECT 90.315 177.585 90.485 177.755 ;
        RECT 90.775 177.585 90.945 177.755 ;
        RECT 91.235 177.585 91.405 177.755 ;
        RECT 91.695 177.585 91.865 177.755 ;
        RECT 92.155 177.585 92.325 177.755 ;
        RECT 92.615 177.585 92.785 177.755 ;
        RECT 93.075 177.585 93.245 177.755 ;
        RECT 93.535 177.585 93.705 177.755 ;
        RECT 93.995 177.585 94.165 177.755 ;
        RECT 94.455 177.585 94.625 177.755 ;
        RECT 94.915 177.585 95.085 177.755 ;
        RECT 95.375 177.585 95.545 177.755 ;
        RECT 95.835 177.585 96.005 177.755 ;
        RECT 96.295 177.585 96.465 177.755 ;
        RECT 96.755 177.585 96.925 177.755 ;
        RECT 97.215 177.585 97.385 177.755 ;
        RECT 97.675 177.585 97.845 177.755 ;
        RECT 98.135 177.585 98.305 177.755 ;
        RECT 98.595 177.585 98.765 177.755 ;
        RECT 99.055 177.585 99.225 177.755 ;
        RECT 99.515 177.585 99.685 177.755 ;
        RECT 99.975 177.585 100.145 177.755 ;
        RECT 100.435 177.585 100.605 177.755 ;
        RECT 100.895 177.585 101.065 177.755 ;
        RECT 101.355 177.585 101.525 177.755 ;
        RECT 101.815 177.585 101.985 177.755 ;
        RECT 102.275 177.585 102.445 177.755 ;
        RECT 102.735 177.585 102.905 177.755 ;
        RECT 103.195 177.585 103.365 177.755 ;
        RECT 103.655 177.585 103.825 177.755 ;
        RECT 104.115 177.585 104.285 177.755 ;
        RECT 104.575 177.585 104.745 177.755 ;
        RECT 105.035 177.585 105.205 177.755 ;
        RECT 105.495 177.585 105.665 177.755 ;
        RECT 105.955 177.585 106.125 177.755 ;
        RECT 106.415 177.585 106.585 177.755 ;
        RECT 106.875 177.585 107.045 177.755 ;
        RECT 107.335 177.585 107.505 177.755 ;
        RECT 107.795 177.585 107.965 177.755 ;
        RECT 108.255 177.585 108.425 177.755 ;
        RECT 108.715 177.585 108.885 177.755 ;
        RECT 109.175 177.585 109.345 177.755 ;
        RECT 109.635 177.585 109.805 177.755 ;
        RECT 110.095 177.585 110.265 177.755 ;
        RECT 110.555 177.585 110.725 177.755 ;
        RECT 111.015 177.585 111.185 177.755 ;
        RECT 111.475 177.585 111.645 177.755 ;
        RECT 111.935 177.585 112.105 177.755 ;
        RECT 112.395 177.585 112.565 177.755 ;
        RECT 112.855 177.585 113.025 177.755 ;
        RECT 113.315 177.585 113.485 177.755 ;
        RECT 113.775 177.585 113.945 177.755 ;
        RECT 114.235 177.585 114.405 177.755 ;
        RECT 114.695 177.585 114.865 177.755 ;
        RECT 115.155 177.585 115.325 177.755 ;
        RECT 110.095 177.075 110.265 177.245 ;
        RECT 108.255 176.395 108.425 176.565 ;
        RECT 109.175 176.055 109.345 176.225 ;
        RECT 111.475 177.075 111.645 177.245 ;
        RECT 110.555 176.735 110.725 176.905 ;
        RECT 112.395 175.715 112.565 175.885 ;
        RECT 61.335 174.865 61.505 175.035 ;
        RECT 61.795 174.865 61.965 175.035 ;
        RECT 62.255 174.865 62.425 175.035 ;
        RECT 62.715 174.865 62.885 175.035 ;
        RECT 63.175 174.865 63.345 175.035 ;
        RECT 63.635 174.865 63.805 175.035 ;
        RECT 64.095 174.865 64.265 175.035 ;
        RECT 64.555 174.865 64.725 175.035 ;
        RECT 65.015 174.865 65.185 175.035 ;
        RECT 65.475 174.865 65.645 175.035 ;
        RECT 65.935 174.865 66.105 175.035 ;
        RECT 66.395 174.865 66.565 175.035 ;
        RECT 66.855 174.865 67.025 175.035 ;
        RECT 67.315 174.865 67.485 175.035 ;
        RECT 67.775 174.865 67.945 175.035 ;
        RECT 68.235 174.865 68.405 175.035 ;
        RECT 68.695 174.865 68.865 175.035 ;
        RECT 69.155 174.865 69.325 175.035 ;
        RECT 69.615 174.865 69.785 175.035 ;
        RECT 70.075 174.865 70.245 175.035 ;
        RECT 70.535 174.865 70.705 175.035 ;
        RECT 70.995 174.865 71.165 175.035 ;
        RECT 71.455 174.865 71.625 175.035 ;
        RECT 71.915 174.865 72.085 175.035 ;
        RECT 72.375 174.865 72.545 175.035 ;
        RECT 72.835 174.865 73.005 175.035 ;
        RECT 73.295 174.865 73.465 175.035 ;
        RECT 73.755 174.865 73.925 175.035 ;
        RECT 74.215 174.865 74.385 175.035 ;
        RECT 74.675 174.865 74.845 175.035 ;
        RECT 75.135 174.865 75.305 175.035 ;
        RECT 75.595 174.865 75.765 175.035 ;
        RECT 76.055 174.865 76.225 175.035 ;
        RECT 76.515 174.865 76.685 175.035 ;
        RECT 76.975 174.865 77.145 175.035 ;
        RECT 77.435 174.865 77.605 175.035 ;
        RECT 77.895 174.865 78.065 175.035 ;
        RECT 78.355 174.865 78.525 175.035 ;
        RECT 78.815 174.865 78.985 175.035 ;
        RECT 79.275 174.865 79.445 175.035 ;
        RECT 79.735 174.865 79.905 175.035 ;
        RECT 80.195 174.865 80.365 175.035 ;
        RECT 80.655 174.865 80.825 175.035 ;
        RECT 81.115 174.865 81.285 175.035 ;
        RECT 81.575 174.865 81.745 175.035 ;
        RECT 82.035 174.865 82.205 175.035 ;
        RECT 82.495 174.865 82.665 175.035 ;
        RECT 82.955 174.865 83.125 175.035 ;
        RECT 83.415 174.865 83.585 175.035 ;
        RECT 83.875 174.865 84.045 175.035 ;
        RECT 84.335 174.865 84.505 175.035 ;
        RECT 84.795 174.865 84.965 175.035 ;
        RECT 85.255 174.865 85.425 175.035 ;
        RECT 85.715 174.865 85.885 175.035 ;
        RECT 86.175 174.865 86.345 175.035 ;
        RECT 86.635 174.865 86.805 175.035 ;
        RECT 87.095 174.865 87.265 175.035 ;
        RECT 87.555 174.865 87.725 175.035 ;
        RECT 88.015 174.865 88.185 175.035 ;
        RECT 88.475 174.865 88.645 175.035 ;
        RECT 88.935 174.865 89.105 175.035 ;
        RECT 89.395 174.865 89.565 175.035 ;
        RECT 89.855 174.865 90.025 175.035 ;
        RECT 90.315 174.865 90.485 175.035 ;
        RECT 90.775 174.865 90.945 175.035 ;
        RECT 91.235 174.865 91.405 175.035 ;
        RECT 91.695 174.865 91.865 175.035 ;
        RECT 92.155 174.865 92.325 175.035 ;
        RECT 92.615 174.865 92.785 175.035 ;
        RECT 93.075 174.865 93.245 175.035 ;
        RECT 93.535 174.865 93.705 175.035 ;
        RECT 93.995 174.865 94.165 175.035 ;
        RECT 94.455 174.865 94.625 175.035 ;
        RECT 94.915 174.865 95.085 175.035 ;
        RECT 95.375 174.865 95.545 175.035 ;
        RECT 95.835 174.865 96.005 175.035 ;
        RECT 96.295 174.865 96.465 175.035 ;
        RECT 96.755 174.865 96.925 175.035 ;
        RECT 97.215 174.865 97.385 175.035 ;
        RECT 97.675 174.865 97.845 175.035 ;
        RECT 98.135 174.865 98.305 175.035 ;
        RECT 98.595 174.865 98.765 175.035 ;
        RECT 99.055 174.865 99.225 175.035 ;
        RECT 99.515 174.865 99.685 175.035 ;
        RECT 99.975 174.865 100.145 175.035 ;
        RECT 100.435 174.865 100.605 175.035 ;
        RECT 100.895 174.865 101.065 175.035 ;
        RECT 101.355 174.865 101.525 175.035 ;
        RECT 101.815 174.865 101.985 175.035 ;
        RECT 102.275 174.865 102.445 175.035 ;
        RECT 102.735 174.865 102.905 175.035 ;
        RECT 103.195 174.865 103.365 175.035 ;
        RECT 103.655 174.865 103.825 175.035 ;
        RECT 104.115 174.865 104.285 175.035 ;
        RECT 104.575 174.865 104.745 175.035 ;
        RECT 105.035 174.865 105.205 175.035 ;
        RECT 105.495 174.865 105.665 175.035 ;
        RECT 105.955 174.865 106.125 175.035 ;
        RECT 106.415 174.865 106.585 175.035 ;
        RECT 106.875 174.865 107.045 175.035 ;
        RECT 107.335 174.865 107.505 175.035 ;
        RECT 107.795 174.865 107.965 175.035 ;
        RECT 108.255 174.865 108.425 175.035 ;
        RECT 108.715 174.865 108.885 175.035 ;
        RECT 109.175 174.865 109.345 175.035 ;
        RECT 109.635 174.865 109.805 175.035 ;
        RECT 110.095 174.865 110.265 175.035 ;
        RECT 110.555 174.865 110.725 175.035 ;
        RECT 111.015 174.865 111.185 175.035 ;
        RECT 111.475 174.865 111.645 175.035 ;
        RECT 111.935 174.865 112.105 175.035 ;
        RECT 112.395 174.865 112.565 175.035 ;
        RECT 112.855 174.865 113.025 175.035 ;
        RECT 113.315 174.865 113.485 175.035 ;
        RECT 113.775 174.865 113.945 175.035 ;
        RECT 114.235 174.865 114.405 175.035 ;
        RECT 114.695 174.865 114.865 175.035 ;
        RECT 115.155 174.865 115.325 175.035 ;
        RECT 112.395 174.355 112.565 174.525 ;
        RECT 111.015 173.675 111.185 173.845 ;
        RECT 111.935 173.675 112.105 173.845 ;
        RECT 112.395 173.675 112.565 173.845 ;
        RECT 61.335 172.145 61.505 172.315 ;
        RECT 61.795 172.145 61.965 172.315 ;
        RECT 62.255 172.145 62.425 172.315 ;
        RECT 62.715 172.145 62.885 172.315 ;
        RECT 63.175 172.145 63.345 172.315 ;
        RECT 63.635 172.145 63.805 172.315 ;
        RECT 64.095 172.145 64.265 172.315 ;
        RECT 64.555 172.145 64.725 172.315 ;
        RECT 65.015 172.145 65.185 172.315 ;
        RECT 65.475 172.145 65.645 172.315 ;
        RECT 65.935 172.145 66.105 172.315 ;
        RECT 66.395 172.145 66.565 172.315 ;
        RECT 66.855 172.145 67.025 172.315 ;
        RECT 67.315 172.145 67.485 172.315 ;
        RECT 67.775 172.145 67.945 172.315 ;
        RECT 68.235 172.145 68.405 172.315 ;
        RECT 68.695 172.145 68.865 172.315 ;
        RECT 69.155 172.145 69.325 172.315 ;
        RECT 69.615 172.145 69.785 172.315 ;
        RECT 70.075 172.145 70.245 172.315 ;
        RECT 70.535 172.145 70.705 172.315 ;
        RECT 70.995 172.145 71.165 172.315 ;
        RECT 71.455 172.145 71.625 172.315 ;
        RECT 71.915 172.145 72.085 172.315 ;
        RECT 72.375 172.145 72.545 172.315 ;
        RECT 72.835 172.145 73.005 172.315 ;
        RECT 73.295 172.145 73.465 172.315 ;
        RECT 73.755 172.145 73.925 172.315 ;
        RECT 74.215 172.145 74.385 172.315 ;
        RECT 74.675 172.145 74.845 172.315 ;
        RECT 75.135 172.145 75.305 172.315 ;
        RECT 75.595 172.145 75.765 172.315 ;
        RECT 76.055 172.145 76.225 172.315 ;
        RECT 76.515 172.145 76.685 172.315 ;
        RECT 76.975 172.145 77.145 172.315 ;
        RECT 77.435 172.145 77.605 172.315 ;
        RECT 77.895 172.145 78.065 172.315 ;
        RECT 78.355 172.145 78.525 172.315 ;
        RECT 78.815 172.145 78.985 172.315 ;
        RECT 79.275 172.145 79.445 172.315 ;
        RECT 79.735 172.145 79.905 172.315 ;
        RECT 80.195 172.145 80.365 172.315 ;
        RECT 80.655 172.145 80.825 172.315 ;
        RECT 81.115 172.145 81.285 172.315 ;
        RECT 81.575 172.145 81.745 172.315 ;
        RECT 82.035 172.145 82.205 172.315 ;
        RECT 82.495 172.145 82.665 172.315 ;
        RECT 82.955 172.145 83.125 172.315 ;
        RECT 83.415 172.145 83.585 172.315 ;
        RECT 83.875 172.145 84.045 172.315 ;
        RECT 84.335 172.145 84.505 172.315 ;
        RECT 84.795 172.145 84.965 172.315 ;
        RECT 85.255 172.145 85.425 172.315 ;
        RECT 85.715 172.145 85.885 172.315 ;
        RECT 86.175 172.145 86.345 172.315 ;
        RECT 86.635 172.145 86.805 172.315 ;
        RECT 87.095 172.145 87.265 172.315 ;
        RECT 87.555 172.145 87.725 172.315 ;
        RECT 88.015 172.145 88.185 172.315 ;
        RECT 88.475 172.145 88.645 172.315 ;
        RECT 88.935 172.145 89.105 172.315 ;
        RECT 89.395 172.145 89.565 172.315 ;
        RECT 89.855 172.145 90.025 172.315 ;
        RECT 90.315 172.145 90.485 172.315 ;
        RECT 90.775 172.145 90.945 172.315 ;
        RECT 91.235 172.145 91.405 172.315 ;
        RECT 91.695 172.145 91.865 172.315 ;
        RECT 92.155 172.145 92.325 172.315 ;
        RECT 92.615 172.145 92.785 172.315 ;
        RECT 93.075 172.145 93.245 172.315 ;
        RECT 93.535 172.145 93.705 172.315 ;
        RECT 93.995 172.145 94.165 172.315 ;
        RECT 94.455 172.145 94.625 172.315 ;
        RECT 94.915 172.145 95.085 172.315 ;
        RECT 95.375 172.145 95.545 172.315 ;
        RECT 95.835 172.145 96.005 172.315 ;
        RECT 96.295 172.145 96.465 172.315 ;
        RECT 96.755 172.145 96.925 172.315 ;
        RECT 97.215 172.145 97.385 172.315 ;
        RECT 97.675 172.145 97.845 172.315 ;
        RECT 98.135 172.145 98.305 172.315 ;
        RECT 98.595 172.145 98.765 172.315 ;
        RECT 99.055 172.145 99.225 172.315 ;
        RECT 99.515 172.145 99.685 172.315 ;
        RECT 99.975 172.145 100.145 172.315 ;
        RECT 100.435 172.145 100.605 172.315 ;
        RECT 100.895 172.145 101.065 172.315 ;
        RECT 101.355 172.145 101.525 172.315 ;
        RECT 101.815 172.145 101.985 172.315 ;
        RECT 102.275 172.145 102.445 172.315 ;
        RECT 102.735 172.145 102.905 172.315 ;
        RECT 103.195 172.145 103.365 172.315 ;
        RECT 103.655 172.145 103.825 172.315 ;
        RECT 104.115 172.145 104.285 172.315 ;
        RECT 104.575 172.145 104.745 172.315 ;
        RECT 105.035 172.145 105.205 172.315 ;
        RECT 105.495 172.145 105.665 172.315 ;
        RECT 105.955 172.145 106.125 172.315 ;
        RECT 106.415 172.145 106.585 172.315 ;
        RECT 106.875 172.145 107.045 172.315 ;
        RECT 107.335 172.145 107.505 172.315 ;
        RECT 107.795 172.145 107.965 172.315 ;
        RECT 108.255 172.145 108.425 172.315 ;
        RECT 108.715 172.145 108.885 172.315 ;
        RECT 109.175 172.145 109.345 172.315 ;
        RECT 109.635 172.145 109.805 172.315 ;
        RECT 110.095 172.145 110.265 172.315 ;
        RECT 110.555 172.145 110.725 172.315 ;
        RECT 111.015 172.145 111.185 172.315 ;
        RECT 111.475 172.145 111.645 172.315 ;
        RECT 111.935 172.145 112.105 172.315 ;
        RECT 112.395 172.145 112.565 172.315 ;
        RECT 112.855 172.145 113.025 172.315 ;
        RECT 113.315 172.145 113.485 172.315 ;
        RECT 113.775 172.145 113.945 172.315 ;
        RECT 114.235 172.145 114.405 172.315 ;
        RECT 114.695 172.145 114.865 172.315 ;
        RECT 115.155 172.145 115.325 172.315 ;
        RECT 61.335 169.425 61.505 169.595 ;
        RECT 61.795 169.425 61.965 169.595 ;
        RECT 62.255 169.425 62.425 169.595 ;
        RECT 62.715 169.425 62.885 169.595 ;
        RECT 63.175 169.425 63.345 169.595 ;
        RECT 63.635 169.425 63.805 169.595 ;
        RECT 64.095 169.425 64.265 169.595 ;
        RECT 64.555 169.425 64.725 169.595 ;
        RECT 65.015 169.425 65.185 169.595 ;
        RECT 65.475 169.425 65.645 169.595 ;
        RECT 65.935 169.425 66.105 169.595 ;
        RECT 66.395 169.425 66.565 169.595 ;
        RECT 66.855 169.425 67.025 169.595 ;
        RECT 67.315 169.425 67.485 169.595 ;
        RECT 67.775 169.425 67.945 169.595 ;
        RECT 68.235 169.425 68.405 169.595 ;
        RECT 68.695 169.425 68.865 169.595 ;
        RECT 69.155 169.425 69.325 169.595 ;
        RECT 69.615 169.425 69.785 169.595 ;
        RECT 70.075 169.425 70.245 169.595 ;
        RECT 70.535 169.425 70.705 169.595 ;
        RECT 70.995 169.425 71.165 169.595 ;
        RECT 71.455 169.425 71.625 169.595 ;
        RECT 71.915 169.425 72.085 169.595 ;
        RECT 72.375 169.425 72.545 169.595 ;
        RECT 72.835 169.425 73.005 169.595 ;
        RECT 73.295 169.425 73.465 169.595 ;
        RECT 73.755 169.425 73.925 169.595 ;
        RECT 74.215 169.425 74.385 169.595 ;
        RECT 74.675 169.425 74.845 169.595 ;
        RECT 75.135 169.425 75.305 169.595 ;
        RECT 75.595 169.425 75.765 169.595 ;
        RECT 76.055 169.425 76.225 169.595 ;
        RECT 76.515 169.425 76.685 169.595 ;
        RECT 76.975 169.425 77.145 169.595 ;
        RECT 77.435 169.425 77.605 169.595 ;
        RECT 77.895 169.425 78.065 169.595 ;
        RECT 78.355 169.425 78.525 169.595 ;
        RECT 78.815 169.425 78.985 169.595 ;
        RECT 79.275 169.425 79.445 169.595 ;
        RECT 79.735 169.425 79.905 169.595 ;
        RECT 80.195 169.425 80.365 169.595 ;
        RECT 80.655 169.425 80.825 169.595 ;
        RECT 81.115 169.425 81.285 169.595 ;
        RECT 81.575 169.425 81.745 169.595 ;
        RECT 82.035 169.425 82.205 169.595 ;
        RECT 82.495 169.425 82.665 169.595 ;
        RECT 82.955 169.425 83.125 169.595 ;
        RECT 83.415 169.425 83.585 169.595 ;
        RECT 83.875 169.425 84.045 169.595 ;
        RECT 84.335 169.425 84.505 169.595 ;
        RECT 84.795 169.425 84.965 169.595 ;
        RECT 85.255 169.425 85.425 169.595 ;
        RECT 85.715 169.425 85.885 169.595 ;
        RECT 86.175 169.425 86.345 169.595 ;
        RECT 86.635 169.425 86.805 169.595 ;
        RECT 87.095 169.425 87.265 169.595 ;
        RECT 87.555 169.425 87.725 169.595 ;
        RECT 88.015 169.425 88.185 169.595 ;
        RECT 88.475 169.425 88.645 169.595 ;
        RECT 88.935 169.425 89.105 169.595 ;
        RECT 89.395 169.425 89.565 169.595 ;
        RECT 89.855 169.425 90.025 169.595 ;
        RECT 90.315 169.425 90.485 169.595 ;
        RECT 90.775 169.425 90.945 169.595 ;
        RECT 91.235 169.425 91.405 169.595 ;
        RECT 91.695 169.425 91.865 169.595 ;
        RECT 92.155 169.425 92.325 169.595 ;
        RECT 92.615 169.425 92.785 169.595 ;
        RECT 93.075 169.425 93.245 169.595 ;
        RECT 93.535 169.425 93.705 169.595 ;
        RECT 93.995 169.425 94.165 169.595 ;
        RECT 94.455 169.425 94.625 169.595 ;
        RECT 94.915 169.425 95.085 169.595 ;
        RECT 95.375 169.425 95.545 169.595 ;
        RECT 95.835 169.425 96.005 169.595 ;
        RECT 96.295 169.425 96.465 169.595 ;
        RECT 96.755 169.425 96.925 169.595 ;
        RECT 97.215 169.425 97.385 169.595 ;
        RECT 97.675 169.425 97.845 169.595 ;
        RECT 98.135 169.425 98.305 169.595 ;
        RECT 98.595 169.425 98.765 169.595 ;
        RECT 99.055 169.425 99.225 169.595 ;
        RECT 99.515 169.425 99.685 169.595 ;
        RECT 99.975 169.425 100.145 169.595 ;
        RECT 100.435 169.425 100.605 169.595 ;
        RECT 100.895 169.425 101.065 169.595 ;
        RECT 101.355 169.425 101.525 169.595 ;
        RECT 101.815 169.425 101.985 169.595 ;
        RECT 102.275 169.425 102.445 169.595 ;
        RECT 102.735 169.425 102.905 169.595 ;
        RECT 103.195 169.425 103.365 169.595 ;
        RECT 103.655 169.425 103.825 169.595 ;
        RECT 104.115 169.425 104.285 169.595 ;
        RECT 104.575 169.425 104.745 169.595 ;
        RECT 105.035 169.425 105.205 169.595 ;
        RECT 105.495 169.425 105.665 169.595 ;
        RECT 105.955 169.425 106.125 169.595 ;
        RECT 106.415 169.425 106.585 169.595 ;
        RECT 106.875 169.425 107.045 169.595 ;
        RECT 107.335 169.425 107.505 169.595 ;
        RECT 107.795 169.425 107.965 169.595 ;
        RECT 108.255 169.425 108.425 169.595 ;
        RECT 108.715 169.425 108.885 169.595 ;
        RECT 109.175 169.425 109.345 169.595 ;
        RECT 109.635 169.425 109.805 169.595 ;
        RECT 110.095 169.425 110.265 169.595 ;
        RECT 110.555 169.425 110.725 169.595 ;
        RECT 111.015 169.425 111.185 169.595 ;
        RECT 111.475 169.425 111.645 169.595 ;
        RECT 111.935 169.425 112.105 169.595 ;
        RECT 112.395 169.425 112.565 169.595 ;
        RECT 112.855 169.425 113.025 169.595 ;
        RECT 113.315 169.425 113.485 169.595 ;
        RECT 113.775 169.425 113.945 169.595 ;
        RECT 114.235 169.425 114.405 169.595 ;
        RECT 114.695 169.425 114.865 169.595 ;
        RECT 115.155 169.425 115.325 169.595 ;
        RECT 61.335 166.705 61.505 166.875 ;
        RECT 61.795 166.705 61.965 166.875 ;
        RECT 62.255 166.705 62.425 166.875 ;
        RECT 62.715 166.705 62.885 166.875 ;
        RECT 63.175 166.705 63.345 166.875 ;
        RECT 63.635 166.705 63.805 166.875 ;
        RECT 64.095 166.705 64.265 166.875 ;
        RECT 64.555 166.705 64.725 166.875 ;
        RECT 65.015 166.705 65.185 166.875 ;
        RECT 65.475 166.705 65.645 166.875 ;
        RECT 65.935 166.705 66.105 166.875 ;
        RECT 66.395 166.705 66.565 166.875 ;
        RECT 66.855 166.705 67.025 166.875 ;
        RECT 67.315 166.705 67.485 166.875 ;
        RECT 67.775 166.705 67.945 166.875 ;
        RECT 68.235 166.705 68.405 166.875 ;
        RECT 68.695 166.705 68.865 166.875 ;
        RECT 69.155 166.705 69.325 166.875 ;
        RECT 69.615 166.705 69.785 166.875 ;
        RECT 70.075 166.705 70.245 166.875 ;
        RECT 70.535 166.705 70.705 166.875 ;
        RECT 70.995 166.705 71.165 166.875 ;
        RECT 71.455 166.705 71.625 166.875 ;
        RECT 71.915 166.705 72.085 166.875 ;
        RECT 72.375 166.705 72.545 166.875 ;
        RECT 72.835 166.705 73.005 166.875 ;
        RECT 73.295 166.705 73.465 166.875 ;
        RECT 73.755 166.705 73.925 166.875 ;
        RECT 74.215 166.705 74.385 166.875 ;
        RECT 74.675 166.705 74.845 166.875 ;
        RECT 75.135 166.705 75.305 166.875 ;
        RECT 75.595 166.705 75.765 166.875 ;
        RECT 76.055 166.705 76.225 166.875 ;
        RECT 76.515 166.705 76.685 166.875 ;
        RECT 76.975 166.705 77.145 166.875 ;
        RECT 77.435 166.705 77.605 166.875 ;
        RECT 77.895 166.705 78.065 166.875 ;
        RECT 78.355 166.705 78.525 166.875 ;
        RECT 78.815 166.705 78.985 166.875 ;
        RECT 79.275 166.705 79.445 166.875 ;
        RECT 79.735 166.705 79.905 166.875 ;
        RECT 80.195 166.705 80.365 166.875 ;
        RECT 80.655 166.705 80.825 166.875 ;
        RECT 81.115 166.705 81.285 166.875 ;
        RECT 81.575 166.705 81.745 166.875 ;
        RECT 82.035 166.705 82.205 166.875 ;
        RECT 82.495 166.705 82.665 166.875 ;
        RECT 82.955 166.705 83.125 166.875 ;
        RECT 83.415 166.705 83.585 166.875 ;
        RECT 83.875 166.705 84.045 166.875 ;
        RECT 84.335 166.705 84.505 166.875 ;
        RECT 84.795 166.705 84.965 166.875 ;
        RECT 85.255 166.705 85.425 166.875 ;
        RECT 85.715 166.705 85.885 166.875 ;
        RECT 86.175 166.705 86.345 166.875 ;
        RECT 86.635 166.705 86.805 166.875 ;
        RECT 87.095 166.705 87.265 166.875 ;
        RECT 87.555 166.705 87.725 166.875 ;
        RECT 88.015 166.705 88.185 166.875 ;
        RECT 88.475 166.705 88.645 166.875 ;
        RECT 88.935 166.705 89.105 166.875 ;
        RECT 89.395 166.705 89.565 166.875 ;
        RECT 89.855 166.705 90.025 166.875 ;
        RECT 90.315 166.705 90.485 166.875 ;
        RECT 90.775 166.705 90.945 166.875 ;
        RECT 91.235 166.705 91.405 166.875 ;
        RECT 91.695 166.705 91.865 166.875 ;
        RECT 92.155 166.705 92.325 166.875 ;
        RECT 92.615 166.705 92.785 166.875 ;
        RECT 93.075 166.705 93.245 166.875 ;
        RECT 93.535 166.705 93.705 166.875 ;
        RECT 93.995 166.705 94.165 166.875 ;
        RECT 94.455 166.705 94.625 166.875 ;
        RECT 94.915 166.705 95.085 166.875 ;
        RECT 95.375 166.705 95.545 166.875 ;
        RECT 95.835 166.705 96.005 166.875 ;
        RECT 96.295 166.705 96.465 166.875 ;
        RECT 96.755 166.705 96.925 166.875 ;
        RECT 97.215 166.705 97.385 166.875 ;
        RECT 97.675 166.705 97.845 166.875 ;
        RECT 98.135 166.705 98.305 166.875 ;
        RECT 98.595 166.705 98.765 166.875 ;
        RECT 99.055 166.705 99.225 166.875 ;
        RECT 99.515 166.705 99.685 166.875 ;
        RECT 99.975 166.705 100.145 166.875 ;
        RECT 100.435 166.705 100.605 166.875 ;
        RECT 100.895 166.705 101.065 166.875 ;
        RECT 101.355 166.705 101.525 166.875 ;
        RECT 101.815 166.705 101.985 166.875 ;
        RECT 102.275 166.705 102.445 166.875 ;
        RECT 102.735 166.705 102.905 166.875 ;
        RECT 103.195 166.705 103.365 166.875 ;
        RECT 103.655 166.705 103.825 166.875 ;
        RECT 104.115 166.705 104.285 166.875 ;
        RECT 104.575 166.705 104.745 166.875 ;
        RECT 105.035 166.705 105.205 166.875 ;
        RECT 105.495 166.705 105.665 166.875 ;
        RECT 105.955 166.705 106.125 166.875 ;
        RECT 106.415 166.705 106.585 166.875 ;
        RECT 106.875 166.705 107.045 166.875 ;
        RECT 107.335 166.705 107.505 166.875 ;
        RECT 107.795 166.705 107.965 166.875 ;
        RECT 108.255 166.705 108.425 166.875 ;
        RECT 108.715 166.705 108.885 166.875 ;
        RECT 109.175 166.705 109.345 166.875 ;
        RECT 109.635 166.705 109.805 166.875 ;
        RECT 110.095 166.705 110.265 166.875 ;
        RECT 110.555 166.705 110.725 166.875 ;
        RECT 111.015 166.705 111.185 166.875 ;
        RECT 111.475 166.705 111.645 166.875 ;
        RECT 111.935 166.705 112.105 166.875 ;
        RECT 112.395 166.705 112.565 166.875 ;
        RECT 112.855 166.705 113.025 166.875 ;
        RECT 113.315 166.705 113.485 166.875 ;
        RECT 113.775 166.705 113.945 166.875 ;
        RECT 114.235 166.705 114.405 166.875 ;
        RECT 114.695 166.705 114.865 166.875 ;
        RECT 115.155 166.705 115.325 166.875 ;
        RECT 61.335 163.985 61.505 164.155 ;
        RECT 61.795 163.985 61.965 164.155 ;
        RECT 62.255 163.985 62.425 164.155 ;
        RECT 62.715 163.985 62.885 164.155 ;
        RECT 63.175 163.985 63.345 164.155 ;
        RECT 63.635 163.985 63.805 164.155 ;
        RECT 64.095 163.985 64.265 164.155 ;
        RECT 64.555 163.985 64.725 164.155 ;
        RECT 65.015 163.985 65.185 164.155 ;
        RECT 65.475 163.985 65.645 164.155 ;
        RECT 65.935 163.985 66.105 164.155 ;
        RECT 66.395 163.985 66.565 164.155 ;
        RECT 66.855 163.985 67.025 164.155 ;
        RECT 67.315 163.985 67.485 164.155 ;
        RECT 67.775 163.985 67.945 164.155 ;
        RECT 68.235 163.985 68.405 164.155 ;
        RECT 68.695 163.985 68.865 164.155 ;
        RECT 69.155 163.985 69.325 164.155 ;
        RECT 69.615 163.985 69.785 164.155 ;
        RECT 70.075 163.985 70.245 164.155 ;
        RECT 70.535 163.985 70.705 164.155 ;
        RECT 70.995 163.985 71.165 164.155 ;
        RECT 71.455 163.985 71.625 164.155 ;
        RECT 71.915 163.985 72.085 164.155 ;
        RECT 72.375 163.985 72.545 164.155 ;
        RECT 72.835 163.985 73.005 164.155 ;
        RECT 73.295 163.985 73.465 164.155 ;
        RECT 73.755 163.985 73.925 164.155 ;
        RECT 74.215 163.985 74.385 164.155 ;
        RECT 74.675 163.985 74.845 164.155 ;
        RECT 75.135 163.985 75.305 164.155 ;
        RECT 75.595 163.985 75.765 164.155 ;
        RECT 76.055 163.985 76.225 164.155 ;
        RECT 76.515 163.985 76.685 164.155 ;
        RECT 76.975 163.985 77.145 164.155 ;
        RECT 77.435 163.985 77.605 164.155 ;
        RECT 77.895 163.985 78.065 164.155 ;
        RECT 78.355 163.985 78.525 164.155 ;
        RECT 78.815 163.985 78.985 164.155 ;
        RECT 79.275 163.985 79.445 164.155 ;
        RECT 79.735 163.985 79.905 164.155 ;
        RECT 80.195 163.985 80.365 164.155 ;
        RECT 80.655 163.985 80.825 164.155 ;
        RECT 81.115 163.985 81.285 164.155 ;
        RECT 81.575 163.985 81.745 164.155 ;
        RECT 82.035 163.985 82.205 164.155 ;
        RECT 82.495 163.985 82.665 164.155 ;
        RECT 82.955 163.985 83.125 164.155 ;
        RECT 83.415 163.985 83.585 164.155 ;
        RECT 83.875 163.985 84.045 164.155 ;
        RECT 84.335 163.985 84.505 164.155 ;
        RECT 84.795 163.985 84.965 164.155 ;
        RECT 85.255 163.985 85.425 164.155 ;
        RECT 85.715 163.985 85.885 164.155 ;
        RECT 86.175 163.985 86.345 164.155 ;
        RECT 86.635 163.985 86.805 164.155 ;
        RECT 87.095 163.985 87.265 164.155 ;
        RECT 87.555 163.985 87.725 164.155 ;
        RECT 88.015 163.985 88.185 164.155 ;
        RECT 88.475 163.985 88.645 164.155 ;
        RECT 88.935 163.985 89.105 164.155 ;
        RECT 89.395 163.985 89.565 164.155 ;
        RECT 89.855 163.985 90.025 164.155 ;
        RECT 90.315 163.985 90.485 164.155 ;
        RECT 90.775 163.985 90.945 164.155 ;
        RECT 91.235 163.985 91.405 164.155 ;
        RECT 91.695 163.985 91.865 164.155 ;
        RECT 92.155 163.985 92.325 164.155 ;
        RECT 92.615 163.985 92.785 164.155 ;
        RECT 93.075 163.985 93.245 164.155 ;
        RECT 93.535 163.985 93.705 164.155 ;
        RECT 93.995 163.985 94.165 164.155 ;
        RECT 94.455 163.985 94.625 164.155 ;
        RECT 94.915 163.985 95.085 164.155 ;
        RECT 95.375 163.985 95.545 164.155 ;
        RECT 95.835 163.985 96.005 164.155 ;
        RECT 96.295 163.985 96.465 164.155 ;
        RECT 96.755 163.985 96.925 164.155 ;
        RECT 97.215 163.985 97.385 164.155 ;
        RECT 97.675 163.985 97.845 164.155 ;
        RECT 98.135 163.985 98.305 164.155 ;
        RECT 98.595 163.985 98.765 164.155 ;
        RECT 99.055 163.985 99.225 164.155 ;
        RECT 99.515 163.985 99.685 164.155 ;
        RECT 99.975 163.985 100.145 164.155 ;
        RECT 100.435 163.985 100.605 164.155 ;
        RECT 100.895 163.985 101.065 164.155 ;
        RECT 101.355 163.985 101.525 164.155 ;
        RECT 101.815 163.985 101.985 164.155 ;
        RECT 102.275 163.985 102.445 164.155 ;
        RECT 102.735 163.985 102.905 164.155 ;
        RECT 103.195 163.985 103.365 164.155 ;
        RECT 103.655 163.985 103.825 164.155 ;
        RECT 104.115 163.985 104.285 164.155 ;
        RECT 104.575 163.985 104.745 164.155 ;
        RECT 105.035 163.985 105.205 164.155 ;
        RECT 105.495 163.985 105.665 164.155 ;
        RECT 105.955 163.985 106.125 164.155 ;
        RECT 106.415 163.985 106.585 164.155 ;
        RECT 106.875 163.985 107.045 164.155 ;
        RECT 107.335 163.985 107.505 164.155 ;
        RECT 107.795 163.985 107.965 164.155 ;
        RECT 108.255 163.985 108.425 164.155 ;
        RECT 108.715 163.985 108.885 164.155 ;
        RECT 109.175 163.985 109.345 164.155 ;
        RECT 109.635 163.985 109.805 164.155 ;
        RECT 110.095 163.985 110.265 164.155 ;
        RECT 110.555 163.985 110.725 164.155 ;
        RECT 111.015 163.985 111.185 164.155 ;
        RECT 111.475 163.985 111.645 164.155 ;
        RECT 111.935 163.985 112.105 164.155 ;
        RECT 112.395 163.985 112.565 164.155 ;
        RECT 112.855 163.985 113.025 164.155 ;
        RECT 113.315 163.985 113.485 164.155 ;
        RECT 113.775 163.985 113.945 164.155 ;
        RECT 114.235 163.985 114.405 164.155 ;
        RECT 114.695 163.985 114.865 164.155 ;
        RECT 115.155 163.985 115.325 164.155 ;
        RECT 61.335 161.265 61.505 161.435 ;
        RECT 61.795 161.265 61.965 161.435 ;
        RECT 62.255 161.265 62.425 161.435 ;
        RECT 62.715 161.265 62.885 161.435 ;
        RECT 63.175 161.265 63.345 161.435 ;
        RECT 63.635 161.265 63.805 161.435 ;
        RECT 64.095 161.265 64.265 161.435 ;
        RECT 64.555 161.265 64.725 161.435 ;
        RECT 65.015 161.265 65.185 161.435 ;
        RECT 65.475 161.265 65.645 161.435 ;
        RECT 65.935 161.265 66.105 161.435 ;
        RECT 66.395 161.265 66.565 161.435 ;
        RECT 66.855 161.265 67.025 161.435 ;
        RECT 67.315 161.265 67.485 161.435 ;
        RECT 67.775 161.265 67.945 161.435 ;
        RECT 68.235 161.265 68.405 161.435 ;
        RECT 68.695 161.265 68.865 161.435 ;
        RECT 69.155 161.265 69.325 161.435 ;
        RECT 69.615 161.265 69.785 161.435 ;
        RECT 70.075 161.265 70.245 161.435 ;
        RECT 70.535 161.265 70.705 161.435 ;
        RECT 70.995 161.265 71.165 161.435 ;
        RECT 71.455 161.265 71.625 161.435 ;
        RECT 71.915 161.265 72.085 161.435 ;
        RECT 72.375 161.265 72.545 161.435 ;
        RECT 72.835 161.265 73.005 161.435 ;
        RECT 73.295 161.265 73.465 161.435 ;
        RECT 73.755 161.265 73.925 161.435 ;
        RECT 74.215 161.265 74.385 161.435 ;
        RECT 74.675 161.265 74.845 161.435 ;
        RECT 75.135 161.265 75.305 161.435 ;
        RECT 75.595 161.265 75.765 161.435 ;
        RECT 76.055 161.265 76.225 161.435 ;
        RECT 76.515 161.265 76.685 161.435 ;
        RECT 76.975 161.265 77.145 161.435 ;
        RECT 77.435 161.265 77.605 161.435 ;
        RECT 77.895 161.265 78.065 161.435 ;
        RECT 78.355 161.265 78.525 161.435 ;
        RECT 78.815 161.265 78.985 161.435 ;
        RECT 79.275 161.265 79.445 161.435 ;
        RECT 79.735 161.265 79.905 161.435 ;
        RECT 80.195 161.265 80.365 161.435 ;
        RECT 80.655 161.265 80.825 161.435 ;
        RECT 81.115 161.265 81.285 161.435 ;
        RECT 81.575 161.265 81.745 161.435 ;
        RECT 82.035 161.265 82.205 161.435 ;
        RECT 82.495 161.265 82.665 161.435 ;
        RECT 82.955 161.265 83.125 161.435 ;
        RECT 83.415 161.265 83.585 161.435 ;
        RECT 83.875 161.265 84.045 161.435 ;
        RECT 84.335 161.265 84.505 161.435 ;
        RECT 84.795 161.265 84.965 161.435 ;
        RECT 85.255 161.265 85.425 161.435 ;
        RECT 85.715 161.265 85.885 161.435 ;
        RECT 86.175 161.265 86.345 161.435 ;
        RECT 86.635 161.265 86.805 161.435 ;
        RECT 87.095 161.265 87.265 161.435 ;
        RECT 87.555 161.265 87.725 161.435 ;
        RECT 88.015 161.265 88.185 161.435 ;
        RECT 88.475 161.265 88.645 161.435 ;
        RECT 88.935 161.265 89.105 161.435 ;
        RECT 89.395 161.265 89.565 161.435 ;
        RECT 89.855 161.265 90.025 161.435 ;
        RECT 90.315 161.265 90.485 161.435 ;
        RECT 90.775 161.265 90.945 161.435 ;
        RECT 91.235 161.265 91.405 161.435 ;
        RECT 91.695 161.265 91.865 161.435 ;
        RECT 92.155 161.265 92.325 161.435 ;
        RECT 92.615 161.265 92.785 161.435 ;
        RECT 93.075 161.265 93.245 161.435 ;
        RECT 93.535 161.265 93.705 161.435 ;
        RECT 93.995 161.265 94.165 161.435 ;
        RECT 94.455 161.265 94.625 161.435 ;
        RECT 94.915 161.265 95.085 161.435 ;
        RECT 95.375 161.265 95.545 161.435 ;
        RECT 95.835 161.265 96.005 161.435 ;
        RECT 96.295 161.265 96.465 161.435 ;
        RECT 96.755 161.265 96.925 161.435 ;
        RECT 97.215 161.265 97.385 161.435 ;
        RECT 97.675 161.265 97.845 161.435 ;
        RECT 98.135 161.265 98.305 161.435 ;
        RECT 98.595 161.265 98.765 161.435 ;
        RECT 99.055 161.265 99.225 161.435 ;
        RECT 99.515 161.265 99.685 161.435 ;
        RECT 99.975 161.265 100.145 161.435 ;
        RECT 100.435 161.265 100.605 161.435 ;
        RECT 100.895 161.265 101.065 161.435 ;
        RECT 101.355 161.265 101.525 161.435 ;
        RECT 101.815 161.265 101.985 161.435 ;
        RECT 102.275 161.265 102.445 161.435 ;
        RECT 102.735 161.265 102.905 161.435 ;
        RECT 103.195 161.265 103.365 161.435 ;
        RECT 103.655 161.265 103.825 161.435 ;
        RECT 104.115 161.265 104.285 161.435 ;
        RECT 104.575 161.265 104.745 161.435 ;
        RECT 105.035 161.265 105.205 161.435 ;
        RECT 105.495 161.265 105.665 161.435 ;
        RECT 105.955 161.265 106.125 161.435 ;
        RECT 106.415 161.265 106.585 161.435 ;
        RECT 106.875 161.265 107.045 161.435 ;
        RECT 107.335 161.265 107.505 161.435 ;
        RECT 107.795 161.265 107.965 161.435 ;
        RECT 108.255 161.265 108.425 161.435 ;
        RECT 108.715 161.265 108.885 161.435 ;
        RECT 109.175 161.265 109.345 161.435 ;
        RECT 109.635 161.265 109.805 161.435 ;
        RECT 110.095 161.265 110.265 161.435 ;
        RECT 110.555 161.265 110.725 161.435 ;
        RECT 111.015 161.265 111.185 161.435 ;
        RECT 111.475 161.265 111.645 161.435 ;
        RECT 111.935 161.265 112.105 161.435 ;
        RECT 112.395 161.265 112.565 161.435 ;
        RECT 112.855 161.265 113.025 161.435 ;
        RECT 113.315 161.265 113.485 161.435 ;
        RECT 113.775 161.265 113.945 161.435 ;
        RECT 114.235 161.265 114.405 161.435 ;
        RECT 114.695 161.265 114.865 161.435 ;
        RECT 115.155 161.265 115.325 161.435 ;
        RECT 61.335 158.545 61.505 158.715 ;
        RECT 61.795 158.545 61.965 158.715 ;
        RECT 62.255 158.545 62.425 158.715 ;
        RECT 62.715 158.545 62.885 158.715 ;
        RECT 63.175 158.545 63.345 158.715 ;
        RECT 63.635 158.545 63.805 158.715 ;
        RECT 64.095 158.545 64.265 158.715 ;
        RECT 64.555 158.545 64.725 158.715 ;
        RECT 65.015 158.545 65.185 158.715 ;
        RECT 65.475 158.545 65.645 158.715 ;
        RECT 65.935 158.545 66.105 158.715 ;
        RECT 66.395 158.545 66.565 158.715 ;
        RECT 66.855 158.545 67.025 158.715 ;
        RECT 67.315 158.545 67.485 158.715 ;
        RECT 67.775 158.545 67.945 158.715 ;
        RECT 68.235 158.545 68.405 158.715 ;
        RECT 68.695 158.545 68.865 158.715 ;
        RECT 69.155 158.545 69.325 158.715 ;
        RECT 69.615 158.545 69.785 158.715 ;
        RECT 70.075 158.545 70.245 158.715 ;
        RECT 70.535 158.545 70.705 158.715 ;
        RECT 70.995 158.545 71.165 158.715 ;
        RECT 71.455 158.545 71.625 158.715 ;
        RECT 71.915 158.545 72.085 158.715 ;
        RECT 72.375 158.545 72.545 158.715 ;
        RECT 72.835 158.545 73.005 158.715 ;
        RECT 73.295 158.545 73.465 158.715 ;
        RECT 73.755 158.545 73.925 158.715 ;
        RECT 74.215 158.545 74.385 158.715 ;
        RECT 74.675 158.545 74.845 158.715 ;
        RECT 75.135 158.545 75.305 158.715 ;
        RECT 75.595 158.545 75.765 158.715 ;
        RECT 76.055 158.545 76.225 158.715 ;
        RECT 76.515 158.545 76.685 158.715 ;
        RECT 76.975 158.545 77.145 158.715 ;
        RECT 77.435 158.545 77.605 158.715 ;
        RECT 77.895 158.545 78.065 158.715 ;
        RECT 78.355 158.545 78.525 158.715 ;
        RECT 78.815 158.545 78.985 158.715 ;
        RECT 79.275 158.545 79.445 158.715 ;
        RECT 79.735 158.545 79.905 158.715 ;
        RECT 80.195 158.545 80.365 158.715 ;
        RECT 80.655 158.545 80.825 158.715 ;
        RECT 81.115 158.545 81.285 158.715 ;
        RECT 81.575 158.545 81.745 158.715 ;
        RECT 82.035 158.545 82.205 158.715 ;
        RECT 82.495 158.545 82.665 158.715 ;
        RECT 82.955 158.545 83.125 158.715 ;
        RECT 83.415 158.545 83.585 158.715 ;
        RECT 83.875 158.545 84.045 158.715 ;
        RECT 84.335 158.545 84.505 158.715 ;
        RECT 84.795 158.545 84.965 158.715 ;
        RECT 85.255 158.545 85.425 158.715 ;
        RECT 85.715 158.545 85.885 158.715 ;
        RECT 86.175 158.545 86.345 158.715 ;
        RECT 86.635 158.545 86.805 158.715 ;
        RECT 87.095 158.545 87.265 158.715 ;
        RECT 87.555 158.545 87.725 158.715 ;
        RECT 88.015 158.545 88.185 158.715 ;
        RECT 88.475 158.545 88.645 158.715 ;
        RECT 88.935 158.545 89.105 158.715 ;
        RECT 89.395 158.545 89.565 158.715 ;
        RECT 89.855 158.545 90.025 158.715 ;
        RECT 90.315 158.545 90.485 158.715 ;
        RECT 90.775 158.545 90.945 158.715 ;
        RECT 91.235 158.545 91.405 158.715 ;
        RECT 91.695 158.545 91.865 158.715 ;
        RECT 92.155 158.545 92.325 158.715 ;
        RECT 92.615 158.545 92.785 158.715 ;
        RECT 93.075 158.545 93.245 158.715 ;
        RECT 93.535 158.545 93.705 158.715 ;
        RECT 93.995 158.545 94.165 158.715 ;
        RECT 94.455 158.545 94.625 158.715 ;
        RECT 94.915 158.545 95.085 158.715 ;
        RECT 95.375 158.545 95.545 158.715 ;
        RECT 95.835 158.545 96.005 158.715 ;
        RECT 96.295 158.545 96.465 158.715 ;
        RECT 96.755 158.545 96.925 158.715 ;
        RECT 97.215 158.545 97.385 158.715 ;
        RECT 97.675 158.545 97.845 158.715 ;
        RECT 98.135 158.545 98.305 158.715 ;
        RECT 98.595 158.545 98.765 158.715 ;
        RECT 99.055 158.545 99.225 158.715 ;
        RECT 99.515 158.545 99.685 158.715 ;
        RECT 99.975 158.545 100.145 158.715 ;
        RECT 100.435 158.545 100.605 158.715 ;
        RECT 100.895 158.545 101.065 158.715 ;
        RECT 101.355 158.545 101.525 158.715 ;
        RECT 101.815 158.545 101.985 158.715 ;
        RECT 102.275 158.545 102.445 158.715 ;
        RECT 102.735 158.545 102.905 158.715 ;
        RECT 103.195 158.545 103.365 158.715 ;
        RECT 103.655 158.545 103.825 158.715 ;
        RECT 104.115 158.545 104.285 158.715 ;
        RECT 104.575 158.545 104.745 158.715 ;
        RECT 105.035 158.545 105.205 158.715 ;
        RECT 105.495 158.545 105.665 158.715 ;
        RECT 105.955 158.545 106.125 158.715 ;
        RECT 106.415 158.545 106.585 158.715 ;
        RECT 106.875 158.545 107.045 158.715 ;
        RECT 107.335 158.545 107.505 158.715 ;
        RECT 107.795 158.545 107.965 158.715 ;
        RECT 108.255 158.545 108.425 158.715 ;
        RECT 108.715 158.545 108.885 158.715 ;
        RECT 109.175 158.545 109.345 158.715 ;
        RECT 109.635 158.545 109.805 158.715 ;
        RECT 110.095 158.545 110.265 158.715 ;
        RECT 110.555 158.545 110.725 158.715 ;
        RECT 111.015 158.545 111.185 158.715 ;
        RECT 111.475 158.545 111.645 158.715 ;
        RECT 111.935 158.545 112.105 158.715 ;
        RECT 112.395 158.545 112.565 158.715 ;
        RECT 112.855 158.545 113.025 158.715 ;
        RECT 113.315 158.545 113.485 158.715 ;
        RECT 113.775 158.545 113.945 158.715 ;
        RECT 114.235 158.545 114.405 158.715 ;
        RECT 114.695 158.545 114.865 158.715 ;
        RECT 115.155 158.545 115.325 158.715 ;
        RECT 61.335 155.825 61.505 155.995 ;
        RECT 61.795 155.825 61.965 155.995 ;
        RECT 62.255 155.825 62.425 155.995 ;
        RECT 62.715 155.825 62.885 155.995 ;
        RECT 63.175 155.825 63.345 155.995 ;
        RECT 63.635 155.825 63.805 155.995 ;
        RECT 64.095 155.825 64.265 155.995 ;
        RECT 64.555 155.825 64.725 155.995 ;
        RECT 65.015 155.825 65.185 155.995 ;
        RECT 65.475 155.825 65.645 155.995 ;
        RECT 65.935 155.825 66.105 155.995 ;
        RECT 66.395 155.825 66.565 155.995 ;
        RECT 66.855 155.825 67.025 155.995 ;
        RECT 67.315 155.825 67.485 155.995 ;
        RECT 67.775 155.825 67.945 155.995 ;
        RECT 68.235 155.825 68.405 155.995 ;
        RECT 68.695 155.825 68.865 155.995 ;
        RECT 69.155 155.825 69.325 155.995 ;
        RECT 69.615 155.825 69.785 155.995 ;
        RECT 70.075 155.825 70.245 155.995 ;
        RECT 70.535 155.825 70.705 155.995 ;
        RECT 70.995 155.825 71.165 155.995 ;
        RECT 71.455 155.825 71.625 155.995 ;
        RECT 71.915 155.825 72.085 155.995 ;
        RECT 72.375 155.825 72.545 155.995 ;
        RECT 72.835 155.825 73.005 155.995 ;
        RECT 73.295 155.825 73.465 155.995 ;
        RECT 73.755 155.825 73.925 155.995 ;
        RECT 74.215 155.825 74.385 155.995 ;
        RECT 74.675 155.825 74.845 155.995 ;
        RECT 75.135 155.825 75.305 155.995 ;
        RECT 75.595 155.825 75.765 155.995 ;
        RECT 76.055 155.825 76.225 155.995 ;
        RECT 76.515 155.825 76.685 155.995 ;
        RECT 76.975 155.825 77.145 155.995 ;
        RECT 77.435 155.825 77.605 155.995 ;
        RECT 77.895 155.825 78.065 155.995 ;
        RECT 78.355 155.825 78.525 155.995 ;
        RECT 78.815 155.825 78.985 155.995 ;
        RECT 79.275 155.825 79.445 155.995 ;
        RECT 79.735 155.825 79.905 155.995 ;
        RECT 80.195 155.825 80.365 155.995 ;
        RECT 80.655 155.825 80.825 155.995 ;
        RECT 81.115 155.825 81.285 155.995 ;
        RECT 81.575 155.825 81.745 155.995 ;
        RECT 82.035 155.825 82.205 155.995 ;
        RECT 82.495 155.825 82.665 155.995 ;
        RECT 82.955 155.825 83.125 155.995 ;
        RECT 83.415 155.825 83.585 155.995 ;
        RECT 83.875 155.825 84.045 155.995 ;
        RECT 84.335 155.825 84.505 155.995 ;
        RECT 84.795 155.825 84.965 155.995 ;
        RECT 85.255 155.825 85.425 155.995 ;
        RECT 85.715 155.825 85.885 155.995 ;
        RECT 86.175 155.825 86.345 155.995 ;
        RECT 86.635 155.825 86.805 155.995 ;
        RECT 87.095 155.825 87.265 155.995 ;
        RECT 87.555 155.825 87.725 155.995 ;
        RECT 88.015 155.825 88.185 155.995 ;
        RECT 88.475 155.825 88.645 155.995 ;
        RECT 88.935 155.825 89.105 155.995 ;
        RECT 89.395 155.825 89.565 155.995 ;
        RECT 89.855 155.825 90.025 155.995 ;
        RECT 90.315 155.825 90.485 155.995 ;
        RECT 90.775 155.825 90.945 155.995 ;
        RECT 91.235 155.825 91.405 155.995 ;
        RECT 91.695 155.825 91.865 155.995 ;
        RECT 92.155 155.825 92.325 155.995 ;
        RECT 92.615 155.825 92.785 155.995 ;
        RECT 93.075 155.825 93.245 155.995 ;
        RECT 93.535 155.825 93.705 155.995 ;
        RECT 93.995 155.825 94.165 155.995 ;
        RECT 94.455 155.825 94.625 155.995 ;
        RECT 94.915 155.825 95.085 155.995 ;
        RECT 95.375 155.825 95.545 155.995 ;
        RECT 95.835 155.825 96.005 155.995 ;
        RECT 96.295 155.825 96.465 155.995 ;
        RECT 96.755 155.825 96.925 155.995 ;
        RECT 97.215 155.825 97.385 155.995 ;
        RECT 97.675 155.825 97.845 155.995 ;
        RECT 98.135 155.825 98.305 155.995 ;
        RECT 98.595 155.825 98.765 155.995 ;
        RECT 99.055 155.825 99.225 155.995 ;
        RECT 99.515 155.825 99.685 155.995 ;
        RECT 99.975 155.825 100.145 155.995 ;
        RECT 100.435 155.825 100.605 155.995 ;
        RECT 100.895 155.825 101.065 155.995 ;
        RECT 101.355 155.825 101.525 155.995 ;
        RECT 101.815 155.825 101.985 155.995 ;
        RECT 102.275 155.825 102.445 155.995 ;
        RECT 102.735 155.825 102.905 155.995 ;
        RECT 103.195 155.825 103.365 155.995 ;
        RECT 103.655 155.825 103.825 155.995 ;
        RECT 104.115 155.825 104.285 155.995 ;
        RECT 104.575 155.825 104.745 155.995 ;
        RECT 105.035 155.825 105.205 155.995 ;
        RECT 105.495 155.825 105.665 155.995 ;
        RECT 105.955 155.825 106.125 155.995 ;
        RECT 106.415 155.825 106.585 155.995 ;
        RECT 106.875 155.825 107.045 155.995 ;
        RECT 107.335 155.825 107.505 155.995 ;
        RECT 107.795 155.825 107.965 155.995 ;
        RECT 108.255 155.825 108.425 155.995 ;
        RECT 108.715 155.825 108.885 155.995 ;
        RECT 109.175 155.825 109.345 155.995 ;
        RECT 109.635 155.825 109.805 155.995 ;
        RECT 110.095 155.825 110.265 155.995 ;
        RECT 110.555 155.825 110.725 155.995 ;
        RECT 111.015 155.825 111.185 155.995 ;
        RECT 111.475 155.825 111.645 155.995 ;
        RECT 111.935 155.825 112.105 155.995 ;
        RECT 112.395 155.825 112.565 155.995 ;
        RECT 112.855 155.825 113.025 155.995 ;
        RECT 113.315 155.825 113.485 155.995 ;
        RECT 113.775 155.825 113.945 155.995 ;
        RECT 114.235 155.825 114.405 155.995 ;
        RECT 114.695 155.825 114.865 155.995 ;
        RECT 115.155 155.825 115.325 155.995 ;
        RECT 61.335 153.105 61.505 153.275 ;
        RECT 61.795 153.105 61.965 153.275 ;
        RECT 62.255 153.105 62.425 153.275 ;
        RECT 62.715 153.105 62.885 153.275 ;
        RECT 63.175 153.105 63.345 153.275 ;
        RECT 63.635 153.105 63.805 153.275 ;
        RECT 64.095 153.105 64.265 153.275 ;
        RECT 64.555 153.105 64.725 153.275 ;
        RECT 65.015 153.105 65.185 153.275 ;
        RECT 65.475 153.105 65.645 153.275 ;
        RECT 65.935 153.105 66.105 153.275 ;
        RECT 66.395 153.105 66.565 153.275 ;
        RECT 66.855 153.105 67.025 153.275 ;
        RECT 67.315 153.105 67.485 153.275 ;
        RECT 67.775 153.105 67.945 153.275 ;
        RECT 68.235 153.105 68.405 153.275 ;
        RECT 68.695 153.105 68.865 153.275 ;
        RECT 69.155 153.105 69.325 153.275 ;
        RECT 69.615 153.105 69.785 153.275 ;
        RECT 70.075 153.105 70.245 153.275 ;
        RECT 70.535 153.105 70.705 153.275 ;
        RECT 70.995 153.105 71.165 153.275 ;
        RECT 71.455 153.105 71.625 153.275 ;
        RECT 71.915 153.105 72.085 153.275 ;
        RECT 72.375 153.105 72.545 153.275 ;
        RECT 72.835 153.105 73.005 153.275 ;
        RECT 73.295 153.105 73.465 153.275 ;
        RECT 73.755 153.105 73.925 153.275 ;
        RECT 74.215 153.105 74.385 153.275 ;
        RECT 74.675 153.105 74.845 153.275 ;
        RECT 75.135 153.105 75.305 153.275 ;
        RECT 75.595 153.105 75.765 153.275 ;
        RECT 76.055 153.105 76.225 153.275 ;
        RECT 76.515 153.105 76.685 153.275 ;
        RECT 76.975 153.105 77.145 153.275 ;
        RECT 77.435 153.105 77.605 153.275 ;
        RECT 77.895 153.105 78.065 153.275 ;
        RECT 78.355 153.105 78.525 153.275 ;
        RECT 78.815 153.105 78.985 153.275 ;
        RECT 79.275 153.105 79.445 153.275 ;
        RECT 79.735 153.105 79.905 153.275 ;
        RECT 80.195 153.105 80.365 153.275 ;
        RECT 80.655 153.105 80.825 153.275 ;
        RECT 81.115 153.105 81.285 153.275 ;
        RECT 81.575 153.105 81.745 153.275 ;
        RECT 82.035 153.105 82.205 153.275 ;
        RECT 82.495 153.105 82.665 153.275 ;
        RECT 82.955 153.105 83.125 153.275 ;
        RECT 83.415 153.105 83.585 153.275 ;
        RECT 83.875 153.105 84.045 153.275 ;
        RECT 84.335 153.105 84.505 153.275 ;
        RECT 84.795 153.105 84.965 153.275 ;
        RECT 85.255 153.105 85.425 153.275 ;
        RECT 85.715 153.105 85.885 153.275 ;
        RECT 86.175 153.105 86.345 153.275 ;
        RECT 86.635 153.105 86.805 153.275 ;
        RECT 87.095 153.105 87.265 153.275 ;
        RECT 87.555 153.105 87.725 153.275 ;
        RECT 88.015 153.105 88.185 153.275 ;
        RECT 88.475 153.105 88.645 153.275 ;
        RECT 88.935 153.105 89.105 153.275 ;
        RECT 89.395 153.105 89.565 153.275 ;
        RECT 89.855 153.105 90.025 153.275 ;
        RECT 90.315 153.105 90.485 153.275 ;
        RECT 90.775 153.105 90.945 153.275 ;
        RECT 91.235 153.105 91.405 153.275 ;
        RECT 91.695 153.105 91.865 153.275 ;
        RECT 92.155 153.105 92.325 153.275 ;
        RECT 92.615 153.105 92.785 153.275 ;
        RECT 93.075 153.105 93.245 153.275 ;
        RECT 93.535 153.105 93.705 153.275 ;
        RECT 93.995 153.105 94.165 153.275 ;
        RECT 94.455 153.105 94.625 153.275 ;
        RECT 94.915 153.105 95.085 153.275 ;
        RECT 95.375 153.105 95.545 153.275 ;
        RECT 95.835 153.105 96.005 153.275 ;
        RECT 96.295 153.105 96.465 153.275 ;
        RECT 96.755 153.105 96.925 153.275 ;
        RECT 97.215 153.105 97.385 153.275 ;
        RECT 97.675 153.105 97.845 153.275 ;
        RECT 98.135 153.105 98.305 153.275 ;
        RECT 98.595 153.105 98.765 153.275 ;
        RECT 99.055 153.105 99.225 153.275 ;
        RECT 99.515 153.105 99.685 153.275 ;
        RECT 99.975 153.105 100.145 153.275 ;
        RECT 100.435 153.105 100.605 153.275 ;
        RECT 100.895 153.105 101.065 153.275 ;
        RECT 101.355 153.105 101.525 153.275 ;
        RECT 101.815 153.105 101.985 153.275 ;
        RECT 102.275 153.105 102.445 153.275 ;
        RECT 102.735 153.105 102.905 153.275 ;
        RECT 103.195 153.105 103.365 153.275 ;
        RECT 103.655 153.105 103.825 153.275 ;
        RECT 104.115 153.105 104.285 153.275 ;
        RECT 104.575 153.105 104.745 153.275 ;
        RECT 105.035 153.105 105.205 153.275 ;
        RECT 105.495 153.105 105.665 153.275 ;
        RECT 105.955 153.105 106.125 153.275 ;
        RECT 106.415 153.105 106.585 153.275 ;
        RECT 106.875 153.105 107.045 153.275 ;
        RECT 107.335 153.105 107.505 153.275 ;
        RECT 107.795 153.105 107.965 153.275 ;
        RECT 108.255 153.105 108.425 153.275 ;
        RECT 108.715 153.105 108.885 153.275 ;
        RECT 109.175 153.105 109.345 153.275 ;
        RECT 109.635 153.105 109.805 153.275 ;
        RECT 110.095 153.105 110.265 153.275 ;
        RECT 110.555 153.105 110.725 153.275 ;
        RECT 111.015 153.105 111.185 153.275 ;
        RECT 111.475 153.105 111.645 153.275 ;
        RECT 111.935 153.105 112.105 153.275 ;
        RECT 112.395 153.105 112.565 153.275 ;
        RECT 112.855 153.105 113.025 153.275 ;
        RECT 113.315 153.105 113.485 153.275 ;
        RECT 113.775 153.105 113.945 153.275 ;
        RECT 114.235 153.105 114.405 153.275 ;
        RECT 114.695 153.105 114.865 153.275 ;
        RECT 115.155 153.105 115.325 153.275 ;
        RECT 106.000 84.080 108.290 86.070 ;
        RECT 115.480 48.920 117.465 49.110 ;
        RECT 140.635 48.920 142.620 49.110 ;
        RECT 115.800 38.735 115.990 40.720 ;
        RECT 115.800 16.580 115.990 18.565 ;
        RECT 119.850 38.935 120.040 40.920 ;
        RECT 119.850 16.780 120.040 18.765 ;
        RECT 125.690 38.110 126.540 41.810 ;
        RECT 126.940 34.810 127.190 41.960 ;
        RECT 127.750 39.985 127.940 41.970 ;
        RECT 127.750 34.930 127.940 36.915 ;
        RECT 126.390 23.560 126.640 32.910 ;
        RECT 127.400 32.270 128.280 32.440 ;
        RECT 126.980 30.290 127.150 32.130 ;
        RECT 128.530 30.290 128.700 32.130 ;
        RECT 127.400 29.980 128.280 30.150 ;
        RECT 126.980 28.000 127.150 29.840 ;
        RECT 128.530 28.000 128.700 29.840 ;
        RECT 127.400 27.690 128.280 27.860 ;
        RECT 126.980 25.710 127.150 27.550 ;
        RECT 128.530 25.710 128.700 27.550 ;
        RECT 127.400 25.400 128.280 25.570 ;
        RECT 126.980 23.420 127.150 25.260 ;
        RECT 128.530 23.420 128.700 25.260 ;
        RECT 130.940 31.210 131.240 43.110 ;
        RECT 132.045 42.900 132.925 43.070 ;
        RECT 131.580 40.920 131.750 42.760 ;
        RECT 133.220 40.920 133.390 42.760 ;
        RECT 132.045 40.610 132.925 40.780 ;
        RECT 131.580 38.630 131.750 40.470 ;
        RECT 133.220 38.630 133.390 40.470 ;
        RECT 132.045 38.320 132.925 38.490 ;
        RECT 131.580 36.340 131.750 38.180 ;
        RECT 133.220 36.340 133.390 38.180 ;
        RECT 132.045 36.030 132.925 36.200 ;
        RECT 131.580 34.050 131.750 35.890 ;
        RECT 133.220 34.050 133.390 35.890 ;
        RECT 132.045 33.740 132.925 33.910 ;
        RECT 131.580 31.760 131.750 33.600 ;
        RECT 133.220 31.760 133.390 33.600 ;
        RECT 132.045 31.450 132.925 31.620 ;
        RECT 131.580 29.470 131.750 31.310 ;
        RECT 133.220 29.470 133.390 31.310 ;
        RECT 132.045 29.160 132.925 29.330 ;
        RECT 138.395 42.900 139.275 43.070 ;
        RECT 137.930 40.920 138.100 42.760 ;
        RECT 139.570 40.920 139.740 42.760 ;
        RECT 138.395 40.610 139.275 40.780 ;
        RECT 137.930 38.630 138.100 40.470 ;
        RECT 139.570 38.630 139.740 40.470 ;
        RECT 138.395 38.320 139.275 38.490 ;
        RECT 137.930 36.340 138.100 38.180 ;
        RECT 139.570 36.340 139.740 38.180 ;
        RECT 138.395 36.030 139.275 36.200 ;
        RECT 137.930 34.050 138.100 35.890 ;
        RECT 139.570 34.050 139.740 35.890 ;
        RECT 138.395 33.740 139.275 33.910 ;
        RECT 137.930 31.760 138.100 33.600 ;
        RECT 139.570 31.760 139.740 33.600 ;
        RECT 138.395 31.450 139.275 31.620 ;
        RECT 137.930 29.470 138.100 31.310 ;
        RECT 139.570 29.470 139.740 31.310 ;
        RECT 140.090 31.210 140.390 43.110 ;
        RECT 138.395 29.160 139.275 29.330 ;
        RECT 132.150 27.100 134.530 27.270 ;
        RECT 131.730 26.620 131.900 26.960 ;
        RECT 134.780 26.620 134.950 26.960 ;
        RECT 132.150 26.310 134.530 26.480 ;
        RECT 141.990 27.810 142.190 43.360 ;
        RECT 142.995 43.160 143.875 43.330 ;
        RECT 142.530 42.680 142.700 43.020 ;
        RECT 144.170 42.680 144.340 43.020 ;
        RECT 142.995 42.370 143.875 42.540 ;
        RECT 142.530 41.890 142.700 42.230 ;
        RECT 144.170 41.890 144.340 42.230 ;
        RECT 142.995 41.580 143.875 41.750 ;
        RECT 142.530 41.100 142.700 41.440 ;
        RECT 144.170 41.100 144.340 41.440 ;
        RECT 142.995 40.790 143.875 40.960 ;
        RECT 142.530 40.310 142.700 40.650 ;
        RECT 144.170 40.310 144.340 40.650 ;
        RECT 142.995 40.000 143.875 40.170 ;
        RECT 142.530 39.520 142.700 39.860 ;
        RECT 144.170 39.520 144.340 39.860 ;
        RECT 142.995 39.210 143.875 39.380 ;
        RECT 142.530 38.730 142.700 39.070 ;
        RECT 144.170 38.730 144.340 39.070 ;
        RECT 142.995 38.420 143.875 38.590 ;
        RECT 142.530 37.940 142.700 38.280 ;
        RECT 144.170 37.940 144.340 38.280 ;
        RECT 142.995 37.630 143.875 37.800 ;
        RECT 142.530 37.150 142.700 37.490 ;
        RECT 144.170 37.150 144.340 37.490 ;
        RECT 142.995 36.840 143.875 37.010 ;
        RECT 142.530 36.360 142.700 36.700 ;
        RECT 144.170 36.360 144.340 36.700 ;
        RECT 142.995 36.050 143.875 36.220 ;
        RECT 142.530 35.570 142.700 35.910 ;
        RECT 144.170 35.570 144.340 35.910 ;
        RECT 142.995 35.260 143.875 35.430 ;
        RECT 142.530 34.780 142.700 35.120 ;
        RECT 144.170 34.780 144.340 35.120 ;
        RECT 142.995 34.470 143.875 34.640 ;
        RECT 142.530 33.990 142.700 34.330 ;
        RECT 144.170 33.990 144.340 34.330 ;
        RECT 142.995 33.680 143.875 33.850 ;
        RECT 142.530 33.200 142.700 33.540 ;
        RECT 144.170 33.200 144.340 33.540 ;
        RECT 142.995 32.890 143.875 33.060 ;
        RECT 142.530 32.410 142.700 32.750 ;
        RECT 144.170 32.410 144.340 32.750 ;
        RECT 142.995 32.100 143.875 32.270 ;
        RECT 142.530 31.620 142.700 31.960 ;
        RECT 144.170 31.620 144.340 31.960 ;
        RECT 142.995 31.310 143.875 31.480 ;
        RECT 142.530 30.830 142.700 31.170 ;
        RECT 144.170 30.830 144.340 31.170 ;
        RECT 142.995 30.520 143.875 30.690 ;
        RECT 142.530 30.040 142.700 30.380 ;
        RECT 144.170 30.040 144.340 30.380 ;
        RECT 142.995 29.730 143.875 29.900 ;
        RECT 142.530 29.250 142.700 29.590 ;
        RECT 144.170 29.250 144.340 29.590 ;
        RECT 142.995 28.940 143.875 29.110 ;
        RECT 142.530 28.460 142.700 28.800 ;
        RECT 144.170 28.460 144.340 28.800 ;
        RECT 142.995 28.150 143.875 28.320 ;
        RECT 136.750 27.100 139.130 27.270 ;
        RECT 136.330 26.620 136.500 26.960 ;
        RECT 139.380 26.620 139.550 26.960 ;
        RECT 136.750 26.310 139.130 26.480 ;
        RECT 142.530 27.670 142.700 28.010 ;
        RECT 144.170 27.670 144.340 28.010 ;
        RECT 142.995 27.360 143.875 27.530 ;
        RECT 146.950 39.190 147.830 39.360 ;
        RECT 146.530 37.210 146.700 39.050 ;
        RECT 148.080 37.210 148.250 39.050 ;
        RECT 146.950 36.900 147.830 37.070 ;
        RECT 146.530 34.920 146.700 36.760 ;
        RECT 148.080 34.920 148.250 36.760 ;
        RECT 146.950 34.610 147.830 34.780 ;
        RECT 146.530 32.630 146.700 34.470 ;
        RECT 148.080 32.630 148.250 34.470 ;
        RECT 146.950 32.320 147.830 32.490 ;
        RECT 146.530 30.340 146.700 32.180 ;
        RECT 148.080 30.340 148.250 32.180 ;
        RECT 146.950 30.030 147.830 30.200 ;
        RECT 146.530 28.050 146.700 29.890 ;
        RECT 148.080 28.050 148.250 29.890 ;
        RECT 146.950 27.740 147.830 27.910 ;
        RECT 146.530 25.760 146.700 27.600 ;
        RECT 148.080 25.760 148.250 27.600 ;
        RECT 146.950 25.450 147.830 25.620 ;
        RECT 127.400 23.110 128.280 23.280 ;
        RECT 131.400 24.650 133.240 24.820 ;
        RECT 133.690 24.650 135.530 24.820 ;
        RECT 135.980 24.650 137.820 24.820 ;
        RECT 138.270 24.650 140.110 24.820 ;
        RECT 131.090 23.520 131.260 24.400 ;
        RECT 133.380 23.520 133.550 24.400 ;
        RECT 135.670 23.520 135.840 24.400 ;
        RECT 137.960 23.520 138.130 24.400 ;
        RECT 140.250 23.520 140.420 24.400 ;
        RECT 131.400 23.100 133.240 23.270 ;
        RECT 133.690 23.100 135.530 23.270 ;
        RECT 135.980 23.100 137.820 23.270 ;
        RECT 138.270 23.100 140.110 23.270 ;
        RECT 145.940 23.060 146.190 24.210 ;
        RECT 146.530 23.470 146.700 25.310 ;
        RECT 148.080 23.470 148.250 25.310 ;
        RECT 146.950 23.160 147.830 23.330 ;
        RECT 148.590 23.060 148.840 24.210 ;
        RECT 126.890 22.460 128.790 22.760 ;
        RECT 130.990 22.510 140.540 22.760 ;
        RECT 146.290 22.560 148.490 22.760 ;
        RECT 128.490 20.810 147.440 21.360 ;
      LAYER met1 ;
        RECT 78.280 208.850 78.600 208.910 ;
        RECT 97.600 208.850 97.920 208.910 ;
        RECT 106.340 208.850 106.660 208.910 ;
        RECT 78.280 208.710 106.660 208.850 ;
        RECT 78.280 208.650 78.600 208.710 ;
        RECT 97.600 208.650 97.920 208.710 ;
        RECT 106.340 208.650 106.660 208.710 ;
        RECT 91.620 208.510 91.940 208.570 ;
        RECT 98.520 208.510 98.840 208.570 ;
        RECT 91.620 208.370 98.840 208.510 ;
        RECT 91.620 208.310 91.940 208.370 ;
        RECT 98.520 208.310 98.840 208.370 ;
        RECT 99.900 208.510 100.220 208.570 ;
        RECT 100.820 208.510 101.140 208.570 ;
        RECT 99.900 208.370 101.140 208.510 ;
        RECT 99.900 208.310 100.220 208.370 ;
        RECT 100.820 208.310 101.140 208.370 ;
        RECT 72.760 208.170 73.080 208.230 ;
        RECT 75.060 208.170 75.380 208.230 ;
        RECT 72.760 208.030 75.380 208.170 ;
        RECT 72.760 207.970 73.080 208.030 ;
        RECT 75.060 207.970 75.380 208.030 ;
        RECT 87.940 208.170 88.260 208.230 ;
        RECT 89.320 208.170 89.640 208.230 ;
        RECT 87.940 208.030 89.640 208.170 ;
        RECT 87.940 207.970 88.260 208.030 ;
        RECT 89.320 207.970 89.640 208.030 ;
        RECT 94.380 208.170 94.700 208.230 ;
        RECT 105.880 208.170 106.200 208.230 ;
        RECT 94.380 208.030 106.200 208.170 ;
        RECT 94.380 207.970 94.700 208.030 ;
        RECT 105.880 207.970 106.200 208.030 ;
        RECT 61.190 207.350 116.270 207.830 ;
        RECT 78.755 207.150 79.045 207.195 ;
        RECT 81.500 207.150 81.820 207.210 ;
        RECT 78.755 207.010 81.820 207.150 ;
        RECT 78.755 206.965 79.045 207.010 ;
        RECT 81.500 206.950 81.820 207.010 ;
        RECT 88.875 207.150 89.165 207.195 ;
        RECT 89.320 207.150 89.640 207.210 ;
        RECT 88.875 207.010 89.640 207.150 ;
        RECT 88.875 206.965 89.165 207.010 ;
        RECT 89.320 206.950 89.640 207.010 ;
        RECT 90.715 207.150 91.005 207.195 ;
        RECT 99.900 207.150 100.220 207.210 ;
        RECT 90.715 207.010 100.220 207.150 ;
        RECT 90.715 206.965 91.005 207.010 ;
        RECT 99.900 206.950 100.220 207.010 ;
        RECT 71.840 206.610 72.160 206.870 ;
        RECT 78.280 206.810 78.600 206.870 ;
        RECT 73.310 206.670 78.600 206.810 ;
        RECT 70.015 206.470 70.305 206.515 ;
        RECT 73.310 206.470 73.450 206.670 ;
        RECT 78.280 206.610 78.600 206.670 ;
        RECT 92.095 206.625 92.385 206.855 ;
        RECT 93.175 206.810 93.465 206.855 ;
        RECT 96.680 206.810 97.000 206.870 ;
        RECT 113.700 206.810 114.020 206.870 ;
        RECT 93.175 206.670 97.000 206.810 ;
        RECT 93.175 206.625 93.465 206.670 ;
        RECT 70.015 206.330 73.450 206.470 ;
        RECT 73.680 206.470 74.000 206.530 ;
        RECT 75.995 206.470 76.285 206.515 ;
        RECT 77.835 206.470 78.125 206.515 ;
        RECT 79.675 206.470 79.965 206.515 ;
        RECT 73.680 206.330 76.285 206.470 ;
        RECT 70.015 206.285 70.305 206.330 ;
        RECT 73.680 206.270 74.000 206.330 ;
        RECT 75.995 206.285 76.285 206.330 ;
        RECT 76.530 206.330 79.965 206.470 ;
        RECT 76.530 206.190 76.670 206.330 ;
        RECT 77.835 206.285 78.125 206.330 ;
        RECT 79.675 206.285 79.965 206.330 ;
        RECT 84.260 206.270 84.580 206.530 ;
        RECT 89.795 206.285 90.085 206.515 ;
        RECT 75.535 205.945 75.825 206.175 ;
        RECT 74.615 205.790 74.905 205.835 ;
        RECT 71.930 205.650 74.905 205.790 ;
        RECT 75.610 205.790 75.750 205.945 ;
        RECT 76.440 205.930 76.760 206.190 ;
        RECT 76.915 206.130 77.205 206.175 ;
        RECT 77.360 206.130 77.680 206.190 ;
        RECT 76.915 205.990 77.680 206.130 ;
        RECT 76.915 205.945 77.205 205.990 ;
        RECT 77.360 205.930 77.680 205.990 ;
        RECT 82.895 206.130 83.185 206.175 ;
        RECT 85.655 206.130 85.945 206.175 ;
        RECT 82.895 205.990 85.945 206.130 ;
        RECT 89.870 206.130 90.010 206.285 ;
        RECT 91.620 206.270 91.940 206.530 ;
        RECT 92.170 206.470 92.310 206.625 ;
        RECT 96.680 206.610 97.000 206.670 ;
        RECT 100.450 206.670 114.020 206.810 ;
        RECT 93.920 206.470 94.240 206.530 ;
        RECT 95.775 206.470 96.065 206.515 ;
        RECT 92.170 206.330 93.690 206.470 ;
        RECT 93.550 206.190 93.690 206.330 ;
        RECT 93.920 206.330 96.065 206.470 ;
        RECT 93.920 206.270 94.240 206.330 ;
        RECT 95.775 206.285 96.065 206.330 ;
        RECT 96.220 206.270 96.540 206.530 ;
        RECT 97.155 206.470 97.445 206.515 ;
        RECT 97.600 206.470 97.920 206.530 ;
        RECT 97.155 206.330 97.920 206.470 ;
        RECT 97.155 206.285 97.445 206.330 ;
        RECT 97.600 206.270 97.920 206.330 ;
        RECT 98.520 206.270 98.840 206.530 ;
        RECT 100.450 206.515 100.590 206.670 ;
        RECT 113.700 206.610 114.020 206.670 ;
        RECT 100.375 206.285 100.665 206.515 ;
        RECT 101.710 206.470 102.000 206.515 ;
        RECT 103.120 206.470 103.440 206.530 ;
        RECT 101.710 206.330 103.440 206.470 ;
        RECT 101.710 206.285 102.000 206.330 ;
        RECT 103.120 206.270 103.440 206.330 ;
        RECT 93.000 206.130 93.320 206.190 ;
        RECT 89.870 205.990 93.320 206.130 ;
        RECT 82.895 205.945 83.185 205.990 ;
        RECT 85.655 205.945 85.945 205.990 ;
        RECT 93.000 205.930 93.320 205.990 ;
        RECT 93.460 205.930 93.780 206.190 ;
        RECT 94.380 205.930 94.700 206.190 ;
        RECT 95.315 206.130 95.605 206.175 ;
        RECT 98.980 206.130 99.300 206.190 ;
        RECT 95.315 205.990 99.300 206.130 ;
        RECT 95.315 205.945 95.605 205.990 ;
        RECT 98.980 205.930 99.300 205.990 ;
        RECT 99.455 205.945 99.745 206.175 ;
        RECT 101.255 206.130 101.545 206.175 ;
        RECT 102.445 206.130 102.735 206.175 ;
        RECT 104.965 206.130 105.255 206.175 ;
        RECT 110.495 206.130 110.785 206.175 ;
        RECT 101.255 205.990 105.255 206.130 ;
        RECT 101.255 205.945 101.545 205.990 ;
        RECT 102.445 205.945 102.735 205.990 ;
        RECT 104.965 205.945 105.255 205.990 ;
        RECT 107.350 205.990 110.785 206.130 ;
        RECT 85.195 205.790 85.485 205.835 ;
        RECT 75.610 205.650 85.485 205.790 ;
        RECT 71.930 205.495 72.070 205.650 ;
        RECT 74.615 205.605 74.905 205.650 ;
        RECT 76.990 205.510 77.130 205.650 ;
        RECT 85.195 205.605 85.485 205.650 ;
        RECT 86.100 205.790 86.420 205.850 ;
        RECT 93.935 205.790 94.225 205.835 ;
        RECT 94.840 205.790 95.160 205.850 ;
        RECT 86.100 205.650 95.160 205.790 ;
        RECT 86.100 205.590 86.420 205.650 ;
        RECT 93.935 205.605 94.225 205.650 ;
        RECT 94.840 205.590 95.160 205.650 ;
        RECT 95.775 205.790 96.065 205.835 ;
        RECT 96.680 205.790 97.000 205.850 ;
        RECT 95.775 205.650 97.000 205.790 ;
        RECT 95.775 205.605 96.065 205.650 ;
        RECT 96.680 205.590 97.000 205.650 ;
        RECT 98.060 205.790 98.380 205.850 ;
        RECT 99.530 205.790 99.670 205.945 ;
        RECT 98.060 205.650 99.670 205.790 ;
        RECT 98.060 205.590 98.380 205.650 ;
        RECT 71.855 205.265 72.145 205.495 ;
        RECT 72.775 205.450 73.065 205.495 ;
        RECT 73.220 205.450 73.540 205.510 ;
        RECT 72.775 205.310 73.540 205.450 ;
        RECT 72.775 205.265 73.065 205.310 ;
        RECT 73.220 205.250 73.540 205.310 ;
        RECT 76.900 205.250 77.220 205.510 ;
        RECT 83.340 205.250 83.660 205.510 ;
        RECT 92.080 205.450 92.400 205.510 ;
        RECT 93.015 205.450 93.305 205.495 ;
        RECT 92.080 205.310 93.305 205.450 ;
        RECT 92.080 205.250 92.400 205.310 ;
        RECT 93.015 205.265 93.305 205.310 ;
        RECT 96.220 205.250 96.540 205.510 ;
        RECT 97.140 205.450 97.460 205.510 ;
        RECT 97.615 205.450 97.905 205.495 ;
        RECT 97.140 205.310 97.905 205.450 ;
        RECT 99.530 205.450 99.670 205.650 ;
        RECT 100.860 205.790 101.150 205.835 ;
        RECT 102.960 205.790 103.250 205.835 ;
        RECT 104.530 205.790 104.820 205.835 ;
        RECT 100.860 205.650 104.820 205.790 ;
        RECT 100.860 205.605 101.150 205.650 ;
        RECT 102.960 205.605 103.250 205.650 ;
        RECT 104.530 205.605 104.820 205.650 ;
        RECT 107.350 205.495 107.490 205.990 ;
        RECT 110.495 205.945 110.785 205.990 ;
        RECT 112.320 205.930 112.640 206.190 ;
        RECT 107.275 205.450 107.565 205.495 ;
        RECT 99.530 205.310 107.565 205.450 ;
        RECT 97.140 205.250 97.460 205.310 ;
        RECT 97.615 205.265 97.905 205.310 ;
        RECT 107.275 205.265 107.565 205.310 ;
        RECT 107.735 205.450 108.025 205.495 ;
        RECT 109.560 205.450 109.880 205.510 ;
        RECT 107.735 205.310 109.880 205.450 ;
        RECT 107.735 205.265 108.025 205.310 ;
        RECT 109.560 205.250 109.880 205.310 ;
        RECT 61.190 204.630 115.470 205.110 ;
        RECT 62.180 204.430 62.500 204.490 ;
        RECT 64.955 204.430 65.245 204.475 ;
        RECT 62.180 204.290 65.245 204.430 ;
        RECT 62.180 204.230 62.500 204.290 ;
        RECT 64.955 204.245 65.245 204.290 ;
        RECT 66.795 204.430 67.085 204.475 ;
        RECT 69.080 204.430 69.400 204.490 ;
        RECT 66.795 204.290 69.400 204.430 ;
        RECT 66.795 204.245 67.085 204.290 ;
        RECT 69.080 204.230 69.400 204.290 ;
        RECT 72.760 204.230 73.080 204.490 ;
        RECT 73.680 204.430 74.000 204.490 ;
        RECT 92.080 204.430 92.400 204.490 ;
        RECT 99.900 204.430 100.220 204.490 ;
        RECT 73.680 204.290 78.970 204.430 ;
        RECT 73.680 204.230 74.000 204.290 ;
        RECT 78.830 204.150 78.970 204.290 ;
        RECT 92.080 204.290 100.220 204.430 ;
        RECT 92.080 204.230 92.400 204.290 ;
        RECT 63.560 204.090 63.880 204.150 ;
        RECT 75.995 204.090 76.285 204.135 ;
        RECT 63.560 203.950 76.285 204.090 ;
        RECT 63.560 203.890 63.880 203.950 ;
        RECT 75.995 203.905 76.285 203.950 ;
        RECT 77.360 203.890 77.680 204.150 ;
        RECT 78.740 203.890 79.060 204.150 ;
        RECT 85.220 204.090 85.510 204.135 ;
        RECT 87.320 204.090 87.610 204.135 ;
        RECT 88.890 204.090 89.180 204.135 ;
        RECT 85.220 203.950 89.180 204.090 ;
        RECT 85.220 203.905 85.510 203.950 ;
        RECT 87.320 203.905 87.610 203.950 ;
        RECT 88.890 203.905 89.180 203.950 ;
        RECT 91.635 204.090 91.925 204.135 ;
        RECT 93.000 204.090 93.320 204.150 ;
        RECT 91.635 203.950 95.530 204.090 ;
        RECT 91.635 203.905 91.925 203.950 ;
        RECT 93.000 203.890 93.320 203.950 ;
        RECT 68.175 203.750 68.465 203.795 ;
        RECT 77.450 203.750 77.590 203.890 ;
        RECT 65.950 203.610 68.465 203.750 ;
        RECT 64.940 203.410 65.260 203.470 ;
        RECT 65.950 203.455 66.090 203.610 ;
        RECT 68.175 203.565 68.465 203.610 ;
        RECT 71.930 203.610 77.590 203.750 ;
        RECT 77.835 203.750 78.125 203.795 ;
        RECT 78.830 203.750 78.970 203.890 ;
        RECT 82.435 203.750 82.725 203.795 ;
        RECT 85.615 203.750 85.905 203.795 ;
        RECT 86.805 203.750 87.095 203.795 ;
        RECT 89.325 203.750 89.615 203.795 ;
        RECT 77.835 203.610 82.725 203.750 ;
        RECT 65.875 203.410 66.165 203.455 ;
        RECT 64.940 203.270 66.165 203.410 ;
        RECT 64.940 203.210 65.260 203.270 ;
        RECT 65.875 203.225 66.165 203.270 ;
        RECT 66.780 203.410 67.100 203.470 ;
        RECT 67.715 203.410 68.005 203.455 ;
        RECT 71.930 203.410 72.070 203.610 ;
        RECT 77.835 203.565 78.125 203.610 ;
        RECT 82.435 203.565 82.725 203.610 ;
        RECT 84.350 203.610 85.410 203.750 ;
        RECT 66.780 203.270 72.070 203.410 ;
        RECT 66.780 203.210 67.100 203.270 ;
        RECT 67.715 203.225 68.005 203.270 ;
        RECT 73.680 203.210 74.000 203.470 ;
        RECT 74.600 203.210 74.920 203.470 ;
        RECT 75.075 203.410 75.365 203.455 ;
        RECT 76.440 203.410 76.760 203.470 ;
        RECT 75.075 203.270 76.760 203.410 ;
        RECT 75.075 203.225 75.365 203.270 ;
        RECT 76.440 203.210 76.760 203.270 ;
        RECT 76.900 203.410 77.220 203.470 ;
        RECT 77.375 203.410 77.665 203.455 ;
        RECT 76.900 203.270 77.665 203.410 ;
        RECT 76.900 203.210 77.220 203.270 ;
        RECT 77.375 203.225 77.665 203.270 ;
        RECT 78.280 203.210 78.600 203.470 ;
        RECT 78.755 203.410 79.045 203.455 ;
        RECT 79.200 203.410 79.520 203.470 ;
        RECT 84.350 203.455 84.490 203.610 ;
        RECT 78.755 203.270 79.520 203.410 ;
        RECT 78.755 203.225 79.045 203.270 ;
        RECT 79.200 203.210 79.520 203.270 ;
        RECT 84.275 203.225 84.565 203.455 ;
        RECT 84.735 203.225 85.025 203.455 ;
        RECT 85.270 203.410 85.410 203.610 ;
        RECT 85.615 203.610 89.615 203.750 ;
        RECT 85.615 203.565 85.905 203.610 ;
        RECT 86.805 203.565 87.095 203.610 ;
        RECT 89.325 203.565 89.615 203.610 ;
        RECT 95.390 203.455 95.530 203.950 ;
        RECT 97.690 203.795 97.830 204.290 ;
        RECT 99.900 204.230 100.220 204.290 ;
        RECT 99.440 203.890 99.760 204.150 ;
        RECT 107.835 204.090 108.125 204.135 ;
        RECT 110.955 204.090 111.245 204.135 ;
        RECT 112.845 204.090 113.135 204.135 ;
        RECT 107.835 203.950 113.135 204.090 ;
        RECT 107.835 203.905 108.125 203.950 ;
        RECT 110.955 203.905 111.245 203.950 ;
        RECT 112.845 203.905 113.135 203.950 ;
        RECT 97.615 203.565 97.905 203.795 ;
        RECT 98.520 203.750 98.840 203.810 ;
        RECT 103.135 203.750 103.425 203.795 ;
        RECT 98.520 203.610 103.425 203.750 ;
        RECT 95.315 203.410 95.605 203.455 ;
        RECT 95.760 203.410 96.080 203.470 ;
        RECT 85.270 203.270 87.250 203.410 ;
        RECT 64.480 203.070 64.800 203.130 ;
        RECT 75.995 203.070 76.285 203.115 ;
        RECT 79.675 203.070 79.965 203.115 ;
        RECT 64.480 202.930 75.750 203.070 ;
        RECT 64.480 202.870 64.800 202.930 ;
        RECT 71.380 202.530 71.700 202.790 ;
        RECT 75.610 202.730 75.750 202.930 ;
        RECT 75.995 202.930 79.965 203.070 ;
        RECT 75.995 202.885 76.285 202.930 ;
        RECT 79.675 202.885 79.965 202.930 ;
        RECT 82.420 203.070 82.740 203.130 ;
        RECT 84.810 203.070 84.950 203.225 ;
        RECT 87.110 203.130 87.250 203.270 ;
        RECT 95.315 203.270 96.080 203.410 ;
        RECT 95.315 203.225 95.605 203.270 ;
        RECT 95.760 203.210 96.080 203.270 ;
        RECT 96.695 203.410 96.985 203.455 ;
        RECT 97.140 203.410 97.460 203.470 ;
        RECT 96.695 203.270 97.460 203.410 ;
        RECT 97.690 203.410 97.830 203.565 ;
        RECT 98.520 203.550 98.840 203.610 ;
        RECT 103.135 203.565 103.425 203.610 ;
        RECT 112.320 203.550 112.640 203.810 ;
        RECT 98.075 203.410 98.365 203.455 ;
        RECT 97.690 203.270 98.365 203.410 ;
        RECT 96.695 203.225 96.985 203.270 ;
        RECT 97.140 203.210 97.460 203.270 ;
        RECT 98.075 203.225 98.365 203.270 ;
        RECT 98.610 203.270 101.050 203.410 ;
        RECT 82.420 202.930 84.950 203.070 ;
        RECT 85.180 203.070 85.500 203.130 ;
        RECT 85.960 203.070 86.250 203.115 ;
        RECT 85.180 202.930 86.250 203.070 ;
        RECT 82.420 202.870 82.740 202.930 ;
        RECT 85.180 202.870 85.500 202.930 ;
        RECT 85.960 202.885 86.250 202.930 ;
        RECT 87.020 202.870 87.340 203.130 ;
        RECT 98.610 203.070 98.750 203.270 ;
        RECT 91.250 202.930 98.750 203.070 ;
        RECT 99.455 203.070 99.745 203.115 ;
        RECT 100.375 203.070 100.665 203.115 ;
        RECT 99.455 202.930 100.665 203.070 ;
        RECT 100.910 203.070 101.050 203.270 ;
        RECT 106.755 203.115 107.045 203.430 ;
        RECT 107.835 203.410 108.125 203.455 ;
        RECT 111.415 203.410 111.705 203.455 ;
        RECT 113.250 203.410 113.540 203.455 ;
        RECT 107.835 203.270 113.540 203.410 ;
        RECT 107.835 203.225 108.125 203.270 ;
        RECT 111.415 203.225 111.705 203.270 ;
        RECT 113.250 203.225 113.540 203.270 ;
        RECT 113.700 203.210 114.020 203.470 ;
        RECT 106.455 203.070 107.045 203.115 ;
        RECT 109.695 203.070 110.345 203.115 ;
        RECT 100.910 202.930 110.345 203.070 ;
        RECT 76.455 202.730 76.745 202.775 ;
        RECT 75.610 202.590 76.745 202.730 ;
        RECT 76.455 202.545 76.745 202.590 ;
        RECT 83.815 202.730 84.105 202.775 ;
        RECT 91.250 202.730 91.390 202.930 ;
        RECT 99.455 202.885 99.745 202.930 ;
        RECT 100.375 202.885 100.665 202.930 ;
        RECT 106.455 202.885 106.745 202.930 ;
        RECT 109.695 202.885 110.345 202.930 ;
        RECT 83.815 202.590 91.390 202.730 ;
        RECT 83.815 202.545 84.105 202.590 ;
        RECT 92.080 202.530 92.400 202.790 ;
        RECT 93.920 202.730 94.240 202.790 ;
        RECT 95.775 202.730 96.065 202.775 ;
        RECT 93.920 202.590 96.065 202.730 ;
        RECT 93.920 202.530 94.240 202.590 ;
        RECT 95.775 202.545 96.065 202.590 ;
        RECT 98.060 202.730 98.380 202.790 ;
        RECT 98.535 202.730 98.825 202.775 ;
        RECT 98.060 202.590 98.825 202.730 ;
        RECT 98.060 202.530 98.380 202.590 ;
        RECT 98.535 202.545 98.825 202.590 ;
        RECT 104.960 202.530 105.280 202.790 ;
        RECT 61.190 201.910 116.270 202.390 ;
        RECT 71.840 201.710 72.160 201.770 ;
        RECT 74.615 201.710 74.905 201.755 ;
        RECT 75.980 201.710 76.300 201.770 ;
        RECT 76.900 201.710 77.220 201.770 ;
        RECT 84.275 201.710 84.565 201.755 ;
        RECT 85.180 201.710 85.500 201.770 ;
        RECT 96.220 201.710 96.540 201.770 ;
        RECT 65.950 201.570 74.905 201.710 ;
        RECT 64.020 201.370 64.340 201.430 ;
        RECT 65.415 201.370 65.705 201.415 ;
        RECT 64.020 201.230 65.705 201.370 ;
        RECT 64.020 201.170 64.340 201.230 ;
        RECT 65.415 201.185 65.705 201.230 ;
        RECT 63.560 200.830 63.880 201.090 ;
        RECT 64.480 200.830 64.800 201.090 ;
        RECT 64.955 201.030 65.245 201.075 ;
        RECT 65.950 201.030 66.090 201.570 ;
        RECT 71.840 201.510 72.160 201.570 ;
        RECT 74.615 201.525 74.905 201.570 ;
        RECT 75.610 201.570 84.030 201.710 ;
        RECT 72.760 201.370 73.080 201.430 ;
        RECT 72.760 201.230 74.370 201.370 ;
        RECT 72.760 201.170 73.080 201.230 ;
        RECT 64.955 200.890 66.090 201.030 ;
        RECT 66.335 201.030 66.625 201.075 ;
        RECT 70.460 201.030 70.780 201.090 ;
        RECT 66.335 200.890 70.780 201.030 ;
        RECT 64.955 200.845 65.245 200.890 ;
        RECT 66.335 200.845 66.625 200.890 ;
        RECT 70.460 200.830 70.780 200.890 ;
        RECT 72.300 201.075 72.620 201.090 ;
        RECT 74.230 201.075 74.370 201.230 ;
        RECT 75.610 201.090 75.750 201.570 ;
        RECT 75.980 201.510 76.300 201.570 ;
        RECT 76.900 201.510 77.220 201.570 ;
        RECT 81.210 201.370 81.500 201.415 ;
        RECT 83.340 201.370 83.660 201.430 ;
        RECT 81.210 201.230 83.660 201.370 ;
        RECT 81.210 201.185 81.500 201.230 ;
        RECT 83.340 201.170 83.660 201.230 ;
        RECT 72.300 200.845 72.650 201.075 ;
        RECT 74.155 200.845 74.445 201.075 ;
        RECT 75.075 201.030 75.365 201.075 ;
        RECT 75.520 201.030 75.840 201.090 ;
        RECT 75.075 200.890 75.840 201.030 ;
        RECT 75.075 200.845 75.365 200.890 ;
        RECT 72.300 200.830 72.620 200.845 ;
        RECT 75.520 200.830 75.840 200.890 ;
        RECT 79.200 201.030 79.520 201.090 ;
        RECT 83.890 201.075 84.030 201.570 ;
        RECT 84.275 201.570 85.500 201.710 ;
        RECT 84.275 201.525 84.565 201.570 ;
        RECT 85.180 201.510 85.500 201.570 ;
        RECT 92.630 201.570 96.540 201.710 ;
        RECT 92.080 201.370 92.400 201.430 ;
        RECT 86.650 201.230 92.400 201.370 ;
        RECT 82.895 201.030 83.185 201.075 ;
        RECT 79.200 200.890 83.185 201.030 ;
        RECT 79.200 200.830 79.520 200.890 ;
        RECT 82.895 200.845 83.185 200.890 ;
        RECT 83.815 200.845 84.105 201.075 ;
        RECT 85.195 200.845 85.485 201.075 ;
        RECT 69.105 200.690 69.395 200.735 ;
        RECT 71.625 200.690 71.915 200.735 ;
        RECT 72.815 200.690 73.105 200.735 ;
        RECT 69.105 200.550 73.105 200.690 ;
        RECT 69.105 200.505 69.395 200.550 ;
        RECT 71.625 200.505 71.915 200.550 ;
        RECT 72.815 200.505 73.105 200.550 ;
        RECT 73.680 200.490 74.000 200.750 ;
        RECT 77.845 200.690 78.135 200.735 ;
        RECT 80.365 200.690 80.655 200.735 ;
        RECT 81.555 200.690 81.845 200.735 ;
        RECT 77.845 200.550 81.845 200.690 ;
        RECT 77.845 200.505 78.135 200.550 ;
        RECT 80.365 200.505 80.655 200.550 ;
        RECT 81.555 200.505 81.845 200.550 ;
        RECT 82.420 200.490 82.740 200.750 ;
        RECT 83.355 200.690 83.645 200.735 ;
        RECT 85.270 200.690 85.410 200.845 ;
        RECT 86.100 200.830 86.420 201.090 ;
        RECT 86.650 201.075 86.790 201.230 ;
        RECT 92.080 201.170 92.400 201.230 ;
        RECT 86.575 200.845 86.865 201.075 ;
        RECT 88.415 201.030 88.705 201.075 ;
        RECT 92.630 201.030 92.770 201.570 ;
        RECT 96.220 201.510 96.540 201.570 ;
        RECT 98.980 201.710 99.300 201.770 ;
        RECT 101.295 201.710 101.585 201.755 ;
        RECT 98.980 201.570 101.585 201.710 ;
        RECT 98.980 201.510 99.300 201.570 ;
        RECT 101.295 201.525 101.585 201.570 ;
        RECT 105.880 201.510 106.200 201.770 ;
        RECT 106.340 201.710 106.660 201.770 ;
        RECT 106.340 201.570 112.550 201.710 ;
        RECT 106.340 201.510 106.660 201.570 ;
        RECT 106.800 201.370 107.120 201.430 ;
        RECT 94.010 201.230 107.120 201.370 ;
        RECT 88.415 200.890 92.770 201.030 ;
        RECT 88.415 200.845 88.705 200.890 ;
        RECT 93.460 200.830 93.780 201.090 ;
        RECT 94.010 201.075 94.150 201.230 ;
        RECT 106.800 201.170 107.120 201.230 ;
        RECT 93.935 200.845 94.225 201.075 ;
        RECT 95.270 201.030 95.560 201.075 ;
        RECT 96.680 201.030 97.000 201.090 ;
        RECT 95.270 200.890 97.000 201.030 ;
        RECT 95.270 200.845 95.560 200.890 ;
        RECT 96.680 200.830 97.000 200.890 ;
        RECT 97.600 201.030 97.920 201.090 ;
        RECT 99.440 201.030 99.760 201.090 ;
        RECT 112.410 201.075 112.550 201.570 ;
        RECT 104.055 201.030 104.345 201.075 ;
        RECT 97.600 200.890 99.210 201.030 ;
        RECT 97.600 200.830 97.920 200.890 ;
        RECT 83.355 200.550 85.410 200.690 ;
        RECT 89.795 200.690 90.085 200.735 ;
        RECT 90.255 200.690 90.545 200.735 ;
        RECT 89.795 200.550 90.545 200.690 ;
        RECT 83.355 200.505 83.645 200.550 ;
        RECT 89.795 200.505 90.085 200.550 ;
        RECT 90.255 200.505 90.545 200.550 ;
        RECT 94.815 200.690 95.105 200.735 ;
        RECT 96.005 200.690 96.295 200.735 ;
        RECT 98.525 200.690 98.815 200.735 ;
        RECT 94.815 200.550 98.815 200.690 ;
        RECT 99.070 200.690 99.210 200.890 ;
        RECT 99.440 200.890 104.345 201.030 ;
        RECT 99.440 200.830 99.760 200.890 ;
        RECT 104.055 200.845 104.345 200.890 ;
        RECT 104.975 200.845 105.265 201.075 ;
        RECT 111.415 201.030 111.705 201.075 ;
        RECT 109.650 200.890 111.705 201.030 ;
        RECT 105.050 200.690 105.190 200.845 ;
        RECT 109.650 200.735 109.790 200.890 ;
        RECT 111.415 200.845 111.705 200.890 ;
        RECT 112.335 200.845 112.625 201.075 ;
        RECT 99.070 200.550 105.190 200.690 ;
        RECT 94.815 200.505 95.105 200.550 ;
        RECT 96.005 200.505 96.295 200.550 ;
        RECT 98.525 200.505 98.815 200.550 ;
        RECT 109.575 200.505 109.865 200.735 ;
        RECT 66.780 200.150 67.100 200.410 ;
        RECT 69.540 200.350 69.830 200.395 ;
        RECT 71.110 200.350 71.400 200.395 ;
        RECT 73.210 200.350 73.500 200.395 ;
        RECT 69.540 200.210 73.500 200.350 ;
        RECT 69.540 200.165 69.830 200.210 ;
        RECT 71.110 200.165 71.400 200.210 ;
        RECT 73.210 200.165 73.500 200.210 ;
        RECT 78.280 200.350 78.570 200.395 ;
        RECT 79.850 200.350 80.140 200.395 ;
        RECT 81.950 200.350 82.240 200.395 ;
        RECT 78.280 200.210 82.240 200.350 ;
        RECT 78.280 200.165 78.570 200.210 ;
        RECT 79.850 200.165 80.140 200.210 ;
        RECT 81.950 200.165 82.240 200.210 ;
        RECT 89.335 200.350 89.625 200.395 ;
        RECT 93.920 200.350 94.240 200.410 ;
        RECT 89.335 200.210 94.240 200.350 ;
        RECT 89.335 200.165 89.625 200.210 ;
        RECT 93.920 200.150 94.240 200.210 ;
        RECT 94.420 200.350 94.710 200.395 ;
        RECT 96.520 200.350 96.810 200.395 ;
        RECT 98.090 200.350 98.380 200.395 ;
        RECT 94.420 200.210 98.380 200.350 ;
        RECT 94.420 200.165 94.710 200.210 ;
        RECT 96.520 200.165 96.810 200.210 ;
        RECT 98.090 200.165 98.380 200.210 ;
        RECT 99.900 200.350 100.220 200.410 ;
        RECT 109.650 200.350 109.790 200.505 ;
        RECT 110.940 200.490 111.260 200.750 ;
        RECT 99.900 200.210 109.790 200.350 ;
        RECT 99.900 200.150 100.220 200.210 ;
        RECT 64.480 199.810 64.800 200.070 ;
        RECT 66.320 199.810 66.640 200.070 ;
        RECT 75.535 200.010 75.825 200.055 ;
        RECT 76.440 200.010 76.760 200.070 ;
        RECT 77.820 200.010 78.140 200.070 ;
        RECT 75.535 199.870 78.140 200.010 ;
        RECT 75.535 199.825 75.825 199.870 ;
        RECT 76.440 199.810 76.760 199.870 ;
        RECT 77.820 199.810 78.140 199.870 ;
        RECT 87.480 199.810 87.800 200.070 ;
        RECT 93.460 200.010 93.780 200.070 ;
        RECT 97.140 200.010 97.460 200.070 ;
        RECT 93.460 199.870 97.460 200.010 ;
        RECT 93.460 199.810 93.780 199.870 ;
        RECT 97.140 199.810 97.460 199.870 ;
        RECT 98.520 200.010 98.840 200.070 ;
        RECT 100.835 200.010 101.125 200.055 ;
        RECT 98.520 199.870 101.125 200.010 ;
        RECT 98.520 199.810 98.840 199.870 ;
        RECT 100.835 199.825 101.125 199.870 ;
        RECT 107.260 200.010 107.580 200.070 ;
        RECT 111.415 200.010 111.705 200.055 ;
        RECT 107.260 199.870 111.705 200.010 ;
        RECT 107.260 199.810 107.580 199.870 ;
        RECT 111.415 199.825 111.705 199.870 ;
        RECT 61.190 199.190 115.470 199.670 ;
        RECT 64.940 198.790 65.260 199.050 ;
        RECT 84.735 198.990 85.025 199.035 ;
        RECT 73.310 198.850 80.350 198.990 ;
        RECT 64.020 198.450 64.340 198.710 ;
        RECT 67.700 198.650 67.990 198.695 ;
        RECT 69.270 198.650 69.560 198.695 ;
        RECT 71.370 198.650 71.660 198.695 ;
        RECT 67.700 198.510 71.660 198.650 ;
        RECT 67.700 198.465 67.990 198.510 ;
        RECT 69.270 198.465 69.560 198.510 ;
        RECT 71.370 198.465 71.660 198.510 ;
        RECT 72.775 198.650 73.065 198.695 ;
        RECT 73.310 198.650 73.450 198.850 ;
        RECT 72.775 198.510 73.450 198.650 ;
        RECT 72.775 198.465 73.065 198.510 ;
        RECT 73.680 198.450 74.000 198.710 ;
        RECT 76.020 198.650 76.310 198.695 ;
        RECT 78.120 198.650 78.410 198.695 ;
        RECT 79.690 198.650 79.980 198.695 ;
        RECT 76.020 198.510 79.980 198.650 ;
        RECT 80.210 198.650 80.350 198.850 ;
        RECT 84.735 198.850 91.390 198.990 ;
        RECT 84.735 198.805 85.025 198.850 ;
        RECT 82.880 198.650 83.200 198.710 ;
        RECT 80.210 198.510 83.200 198.650 ;
        RECT 76.020 198.465 76.310 198.510 ;
        RECT 78.120 198.465 78.410 198.510 ;
        RECT 79.690 198.465 79.980 198.510 ;
        RECT 82.880 198.450 83.200 198.510 ;
        RECT 83.355 198.650 83.645 198.695 ;
        RECT 85.640 198.650 85.960 198.710 ;
        RECT 83.355 198.510 85.960 198.650 ;
        RECT 83.355 198.465 83.645 198.510 ;
        RECT 85.640 198.450 85.960 198.510 ;
        RECT 87.060 198.650 87.350 198.695 ;
        RECT 89.160 198.650 89.450 198.695 ;
        RECT 90.730 198.650 91.020 198.695 ;
        RECT 87.060 198.510 91.020 198.650 ;
        RECT 91.250 198.650 91.390 198.850 ;
        RECT 93.460 198.790 93.780 199.050 ;
        RECT 98.075 198.990 98.365 199.035 ;
        RECT 99.440 198.990 99.760 199.050 ;
        RECT 98.075 198.850 99.760 198.990 ;
        RECT 98.075 198.805 98.365 198.850 ;
        RECT 99.440 198.790 99.760 198.850 ;
        RECT 102.675 198.990 102.965 199.035 ;
        RECT 103.120 198.990 103.440 199.050 ;
        RECT 102.675 198.850 103.440 198.990 ;
        RECT 102.675 198.805 102.965 198.850 ;
        RECT 103.120 198.790 103.440 198.850 ;
        RECT 94.840 198.650 95.160 198.710 ;
        RECT 91.250 198.510 95.160 198.650 ;
        RECT 87.060 198.465 87.350 198.510 ;
        RECT 89.160 198.465 89.450 198.510 ;
        RECT 90.730 198.465 91.020 198.510 ;
        RECT 94.840 198.450 95.160 198.510 ;
        RECT 96.695 198.650 96.985 198.695 ;
        RECT 99.900 198.650 100.220 198.710 ;
        RECT 100.835 198.650 101.125 198.695 ;
        RECT 96.695 198.510 97.370 198.650 ;
        RECT 96.695 198.465 96.985 198.510 ;
        RECT 67.265 198.310 67.555 198.355 ;
        RECT 69.785 198.310 70.075 198.355 ;
        RECT 70.975 198.310 71.265 198.355 ;
        RECT 67.265 198.170 71.265 198.310 ;
        RECT 67.265 198.125 67.555 198.170 ;
        RECT 69.785 198.125 70.075 198.170 ;
        RECT 70.975 198.125 71.265 198.170 ;
        RECT 71.855 198.310 72.145 198.355 ;
        RECT 73.770 198.310 73.910 198.450 ;
        RECT 97.230 198.370 97.370 198.510 ;
        RECT 97.690 198.510 101.125 198.650 ;
        RECT 76.415 198.310 76.705 198.355 ;
        RECT 77.605 198.310 77.895 198.355 ;
        RECT 80.125 198.310 80.415 198.355 ;
        RECT 82.420 198.310 82.740 198.370 ;
        RECT 86.575 198.310 86.865 198.355 ;
        RECT 71.855 198.170 75.750 198.310 ;
        RECT 71.855 198.125 72.145 198.170 ;
        RECT 64.495 197.785 64.785 198.015 ;
        RECT 66.320 197.970 66.640 198.030 ;
        RECT 70.520 197.970 70.810 198.015 ;
        RECT 66.320 197.830 70.810 197.970 ;
        RECT 64.570 197.290 64.710 197.785 ;
        RECT 66.320 197.770 66.640 197.830 ;
        RECT 70.520 197.785 70.810 197.830 ;
        RECT 73.680 197.770 74.000 198.030 ;
        RECT 75.610 198.015 75.750 198.170 ;
        RECT 76.415 198.170 80.415 198.310 ;
        RECT 76.415 198.125 76.705 198.170 ;
        RECT 77.605 198.125 77.895 198.170 ;
        RECT 80.125 198.125 80.415 198.170 ;
        RECT 80.670 198.170 86.865 198.310 ;
        RECT 75.535 197.970 75.825 198.015 ;
        RECT 75.980 197.970 76.300 198.030 ;
        RECT 80.670 197.970 80.810 198.170 ;
        RECT 82.420 198.110 82.740 198.170 ;
        RECT 86.575 198.125 86.865 198.170 ;
        RECT 87.455 198.310 87.745 198.355 ;
        RECT 88.645 198.310 88.935 198.355 ;
        RECT 91.165 198.310 91.455 198.355 ;
        RECT 87.455 198.170 91.455 198.310 ;
        RECT 87.455 198.125 87.745 198.170 ;
        RECT 88.645 198.125 88.935 198.170 ;
        RECT 91.165 198.125 91.455 198.170 ;
        RECT 97.140 198.110 97.460 198.370 ;
        RECT 75.535 197.830 80.810 197.970 ;
        RECT 84.275 197.970 84.565 198.015 ;
        RECT 85.640 197.970 85.960 198.030 ;
        RECT 84.275 197.830 85.960 197.970 ;
        RECT 75.535 197.785 75.825 197.830 ;
        RECT 75.980 197.770 76.300 197.830 ;
        RECT 84.275 197.785 84.565 197.830 ;
        RECT 85.640 197.770 85.960 197.830 ;
        RECT 86.115 197.970 86.405 198.015 ;
        RECT 95.315 197.970 95.605 198.015 ;
        RECT 96.310 197.970 96.910 197.980 ;
        RECT 97.690 197.970 97.830 198.510 ;
        RECT 99.900 198.450 100.220 198.510 ;
        RECT 100.835 198.465 101.125 198.510 ;
        RECT 103.620 198.650 103.910 198.695 ;
        RECT 105.720 198.650 106.010 198.695 ;
        RECT 107.290 198.650 107.580 198.695 ;
        RECT 103.620 198.510 107.580 198.650 ;
        RECT 103.620 198.465 103.910 198.510 ;
        RECT 105.720 198.465 106.010 198.510 ;
        RECT 107.290 198.465 107.580 198.510 ;
        RECT 110.035 198.650 110.325 198.695 ;
        RECT 111.400 198.650 111.720 198.710 ;
        RECT 110.035 198.510 113.470 198.650 ;
        RECT 110.035 198.465 110.325 198.510 ;
        RECT 111.400 198.450 111.720 198.510 ;
        RECT 113.330 198.355 113.470 198.510 ;
        RECT 104.015 198.310 104.305 198.355 ;
        RECT 105.205 198.310 105.495 198.355 ;
        RECT 107.725 198.310 108.015 198.355 ;
        RECT 104.015 198.170 108.015 198.310 ;
        RECT 104.015 198.125 104.305 198.170 ;
        RECT 105.205 198.125 105.495 198.170 ;
        RECT 107.725 198.125 108.015 198.170 ;
        RECT 113.255 198.125 113.545 198.355 ;
        RECT 100.375 197.970 100.665 198.015 ;
        RECT 86.115 197.840 97.830 197.970 ;
        RECT 86.115 197.830 96.450 197.840 ;
        RECT 96.770 197.830 97.830 197.840 ;
        RECT 98.610 197.830 100.665 197.970 ;
        RECT 86.115 197.785 86.405 197.830 ;
        RECT 95.315 197.785 95.605 197.830 ;
        RECT 75.060 197.630 75.380 197.690 ;
        RECT 76.760 197.630 77.050 197.675 ;
        RECT 75.060 197.490 77.050 197.630 ;
        RECT 75.060 197.430 75.380 197.490 ;
        RECT 76.760 197.445 77.050 197.490 ;
        RECT 82.880 197.630 83.200 197.690 ;
        RECT 84.720 197.630 85.040 197.690 ;
        RECT 87.940 197.675 88.260 197.690 ;
        RECT 82.880 197.490 85.040 197.630 ;
        RECT 82.880 197.430 83.200 197.490 ;
        RECT 84.720 197.430 85.040 197.490 ;
        RECT 87.910 197.445 88.260 197.675 ;
        RECT 95.775 197.630 96.065 197.675 ;
        RECT 96.220 197.630 96.540 197.690 ;
        RECT 98.610 197.630 98.750 197.830 ;
        RECT 100.375 197.785 100.665 197.830 ;
        RECT 87.940 197.430 88.260 197.445 ;
        RECT 93.550 197.490 95.530 197.630 ;
        RECT 71.380 197.290 71.700 197.350 ;
        RECT 64.570 197.150 71.700 197.290 ;
        RECT 71.380 197.090 71.700 197.150 ;
        RECT 78.740 197.290 79.060 197.350 ;
        RECT 82.435 197.290 82.725 197.335 ;
        RECT 78.740 197.150 82.725 197.290 ;
        RECT 78.740 197.090 79.060 197.150 ;
        RECT 82.435 197.105 82.725 197.150 ;
        RECT 85.655 197.290 85.945 197.335 ;
        RECT 93.550 197.290 93.690 197.490 ;
        RECT 85.655 197.150 93.690 197.290 ;
        RECT 85.655 197.105 85.945 197.150 ;
        RECT 93.920 197.090 94.240 197.350 ;
        RECT 94.840 197.090 95.160 197.350 ;
        RECT 95.390 197.290 95.530 197.490 ;
        RECT 95.775 197.490 96.540 197.630 ;
        RECT 95.775 197.445 96.065 197.490 ;
        RECT 96.220 197.430 96.540 197.490 ;
        RECT 96.770 197.490 98.750 197.630 ;
        RECT 96.770 197.290 96.910 197.490 ;
        RECT 98.980 197.430 99.300 197.690 ;
        RECT 95.390 197.150 96.910 197.290 ;
        RECT 97.140 197.090 97.460 197.350 ;
        RECT 97.995 197.290 98.285 197.335 ;
        RECT 98.520 197.290 98.840 197.350 ;
        RECT 97.995 197.150 98.840 197.290 ;
        RECT 100.450 197.290 100.590 197.785 ;
        RECT 101.740 197.770 102.060 198.030 ;
        RECT 103.135 197.970 103.425 198.015 ;
        RECT 106.800 197.970 107.120 198.030 ;
        RECT 110.020 197.970 110.340 198.030 ;
        RECT 103.135 197.830 110.340 197.970 ;
        RECT 103.135 197.785 103.425 197.830 ;
        RECT 106.800 197.770 107.120 197.830 ;
        RECT 110.020 197.770 110.340 197.830 ;
        RECT 103.580 197.630 103.900 197.690 ;
        RECT 104.360 197.630 104.650 197.675 ;
        RECT 103.580 197.490 104.650 197.630 ;
        RECT 103.580 197.430 103.900 197.490 ;
        RECT 104.360 197.445 104.650 197.490 ;
        RECT 109.560 197.290 109.880 197.350 ;
        RECT 100.450 197.150 109.880 197.290 ;
        RECT 97.995 197.105 98.285 197.150 ;
        RECT 98.520 197.090 98.840 197.150 ;
        RECT 109.560 197.090 109.880 197.150 ;
        RECT 110.480 197.090 110.800 197.350 ;
        RECT 61.190 196.470 116.270 196.950 ;
        RECT 70.460 196.070 70.780 196.330 ;
        RECT 72.760 196.270 73.080 196.330 ;
        RECT 74.615 196.270 74.905 196.315 ;
        RECT 72.160 196.130 74.905 196.270 ;
        RECT 71.395 195.590 71.685 195.635 ;
        RECT 72.160 195.590 72.300 196.130 ;
        RECT 72.760 196.070 73.080 196.130 ;
        RECT 74.615 196.085 74.905 196.130 ;
        RECT 75.455 196.270 75.745 196.315 ;
        RECT 77.360 196.270 77.680 196.330 ;
        RECT 75.455 196.130 77.680 196.270 ;
        RECT 75.455 196.085 75.745 196.130 ;
        RECT 77.360 196.070 77.680 196.130 ;
        RECT 87.020 196.270 87.340 196.330 ;
        RECT 87.495 196.270 87.785 196.315 ;
        RECT 87.020 196.130 87.785 196.270 ;
        RECT 87.020 196.070 87.340 196.130 ;
        RECT 87.495 196.085 87.785 196.130 ;
        RECT 91.175 196.085 91.465 196.315 ;
        RECT 98.535 196.270 98.825 196.315 ;
        RECT 103.580 196.270 103.900 196.330 ;
        RECT 98.535 196.130 103.900 196.270 ;
        RECT 98.535 196.085 98.825 196.130 ;
        RECT 76.455 195.930 76.745 195.975 ;
        RECT 78.280 195.930 78.600 195.990 ;
        RECT 76.455 195.790 78.600 195.930 ;
        RECT 76.455 195.745 76.745 195.790 ;
        RECT 78.280 195.730 78.600 195.790 ;
        RECT 85.655 195.930 85.945 195.975 ;
        RECT 91.250 195.930 91.390 196.085 ;
        RECT 103.580 196.070 103.900 196.130 ;
        RECT 101.295 195.930 101.585 195.975 ;
        RECT 85.655 195.790 101.585 195.930 ;
        RECT 85.655 195.745 85.945 195.790 ;
        RECT 101.295 195.745 101.585 195.790 ;
        RECT 110.020 195.930 110.340 195.990 ;
        RECT 113.700 195.930 114.020 195.990 ;
        RECT 110.020 195.790 114.020 195.930 ;
        RECT 110.020 195.730 110.340 195.790 ;
        RECT 113.700 195.730 114.020 195.790 ;
        RECT 71.395 195.450 72.300 195.590 ;
        RECT 72.775 195.590 73.065 195.635 ;
        RECT 79.200 195.590 79.520 195.650 ;
        RECT 72.775 195.450 79.520 195.590 ;
        RECT 71.395 195.405 71.685 195.450 ;
        RECT 72.775 195.405 73.065 195.450 ;
        RECT 79.200 195.390 79.520 195.450 ;
        RECT 88.415 195.590 88.705 195.635 ;
        RECT 90.240 195.590 90.560 195.650 ;
        RECT 88.415 195.450 90.560 195.590 ;
        RECT 88.415 195.405 88.705 195.450 ;
        RECT 90.240 195.390 90.560 195.450 ;
        RECT 97.600 195.390 97.920 195.650 ;
        RECT 99.455 195.405 99.745 195.635 ;
        RECT 100.835 195.590 101.125 195.635 ;
        RECT 110.480 195.590 110.800 195.650 ;
        RECT 100.835 195.450 110.800 195.590 ;
        RECT 100.835 195.405 101.125 195.450 ;
        RECT 71.855 195.250 72.145 195.295 ;
        RECT 71.010 195.110 72.145 195.250 ;
        RECT 71.010 194.570 71.150 195.110 ;
        RECT 71.855 195.065 72.145 195.110 ;
        RECT 72.315 195.065 72.605 195.295 ;
        RECT 71.380 194.910 71.700 194.970 ;
        RECT 72.390 194.910 72.530 195.065 ;
        RECT 76.900 195.050 77.220 195.310 ;
        RECT 85.640 195.250 85.960 195.310 ;
        RECT 98.060 195.250 98.380 195.310 ;
        RECT 85.640 195.110 98.380 195.250 ;
        RECT 99.530 195.250 99.670 195.405 ;
        RECT 110.480 195.390 110.800 195.450 ;
        RECT 111.415 195.405 111.705 195.635 ;
        RECT 107.260 195.250 107.580 195.310 ;
        RECT 99.530 195.110 107.580 195.250 ;
        RECT 85.640 195.050 85.960 195.110 ;
        RECT 98.060 195.050 98.380 195.110 ;
        RECT 107.260 195.050 107.580 195.110 ;
        RECT 109.560 195.250 109.880 195.310 ;
        RECT 111.490 195.250 111.630 195.405 ;
        RECT 109.560 195.110 111.630 195.250 ;
        RECT 109.560 195.050 109.880 195.110 ;
        RECT 112.320 195.050 112.640 195.310 ;
        RECT 71.380 194.770 72.530 194.910 ;
        RECT 71.380 194.710 71.700 194.770 ;
        RECT 75.060 194.570 75.380 194.630 ;
        RECT 71.010 194.430 75.380 194.570 ;
        RECT 75.060 194.370 75.380 194.430 ;
        RECT 75.535 194.570 75.825 194.615 ;
        RECT 78.740 194.570 79.060 194.630 ;
        RECT 75.535 194.430 79.060 194.570 ;
        RECT 75.535 194.385 75.825 194.430 ;
        RECT 78.740 194.370 79.060 194.430 ;
        RECT 96.680 194.570 97.000 194.630 ;
        RECT 98.980 194.570 99.300 194.630 ;
        RECT 96.680 194.430 99.300 194.570 ;
        RECT 96.680 194.370 97.000 194.430 ;
        RECT 98.980 194.370 99.300 194.430 ;
        RECT 99.900 194.570 100.220 194.630 ;
        RECT 100.375 194.570 100.665 194.615 ;
        RECT 99.900 194.430 100.665 194.570 ;
        RECT 99.900 194.370 100.220 194.430 ;
        RECT 100.375 194.385 100.665 194.430 ;
        RECT 110.480 194.370 110.800 194.630 ;
        RECT 61.190 193.750 115.470 194.230 ;
        RECT 72.300 193.550 72.620 193.610 ;
        RECT 72.775 193.550 73.065 193.595 ;
        RECT 79.675 193.550 79.965 193.595 ;
        RECT 72.300 193.410 73.065 193.550 ;
        RECT 72.300 193.350 72.620 193.410 ;
        RECT 72.775 193.365 73.065 193.410 ;
        RECT 75.150 193.410 79.965 193.550 ;
        RECT 73.220 192.530 73.540 192.590 ;
        RECT 73.695 192.530 73.985 192.575 ;
        RECT 73.220 192.390 73.985 192.530 ;
        RECT 73.220 192.330 73.540 192.390 ;
        RECT 73.695 192.345 73.985 192.390 ;
        RECT 74.615 192.530 74.905 192.575 ;
        RECT 75.150 192.530 75.290 193.410 ;
        RECT 79.675 193.365 79.965 193.410 ;
        RECT 93.460 193.550 93.780 193.610 ;
        RECT 95.775 193.550 96.065 193.595 ;
        RECT 93.460 193.410 96.065 193.550 ;
        RECT 93.460 193.350 93.780 193.410 ;
        RECT 95.775 193.365 96.065 193.410 ;
        RECT 97.140 193.550 97.460 193.610 ;
        RECT 102.215 193.550 102.505 193.595 ;
        RECT 97.140 193.410 102.505 193.550 ;
        RECT 75.535 193.210 75.825 193.255 ;
        RECT 75.980 193.210 76.300 193.270 ;
        RECT 78.740 193.210 79.060 193.270 ;
        RECT 75.535 193.070 76.300 193.210 ;
        RECT 75.535 193.025 75.825 193.070 ;
        RECT 75.980 193.010 76.300 193.070 ;
        RECT 76.990 193.070 79.060 193.210 ;
        RECT 76.990 192.870 77.130 193.070 ;
        RECT 78.740 193.010 79.060 193.070 ;
        RECT 79.215 193.210 79.505 193.255 ;
        RECT 84.260 193.210 84.580 193.270 ;
        RECT 90.255 193.210 90.545 193.255 ;
        RECT 95.850 193.210 95.990 193.365 ;
        RECT 97.140 193.350 97.460 193.410 ;
        RECT 102.215 193.365 102.505 193.410 ;
        RECT 98.995 193.210 99.285 193.255 ;
        RECT 79.215 193.070 84.580 193.210 ;
        RECT 79.215 193.025 79.505 193.070 ;
        RECT 84.260 193.010 84.580 193.070 ;
        RECT 87.110 193.070 95.070 193.210 ;
        RECT 95.850 193.070 99.285 193.210 ;
        RECT 81.960 192.870 82.280 192.930 ;
        RECT 86.575 192.870 86.865 192.915 ;
        RECT 76.070 192.730 77.130 192.870 ;
        RECT 77.450 192.730 82.280 192.870 ;
        RECT 76.070 192.575 76.210 192.730 ;
        RECT 74.615 192.390 75.290 192.530 ;
        RECT 75.535 192.530 75.825 192.575 ;
        RECT 75.995 192.530 76.285 192.575 ;
        RECT 75.535 192.390 76.285 192.530 ;
        RECT 74.615 192.345 74.905 192.390 ;
        RECT 75.535 192.345 75.825 192.390 ;
        RECT 75.995 192.345 76.285 192.390 ;
        RECT 76.440 192.530 76.760 192.590 ;
        RECT 77.450 192.575 77.590 192.730 ;
        RECT 81.960 192.670 82.280 192.730 ;
        RECT 82.510 192.730 86.865 192.870 ;
        RECT 76.915 192.530 77.205 192.575 ;
        RECT 76.440 192.390 77.205 192.530 ;
        RECT 73.220 191.850 73.540 191.910 ;
        RECT 74.690 191.850 74.830 192.345 ;
        RECT 76.440 192.330 76.760 192.390 ;
        RECT 76.915 192.345 77.205 192.390 ;
        RECT 77.375 192.345 77.665 192.575 ;
        RECT 77.835 192.345 78.125 192.575 ;
        RECT 75.060 192.190 75.380 192.250 ;
        RECT 77.910 192.190 78.050 192.345 ;
        RECT 78.280 192.330 78.600 192.590 ;
        RECT 82.510 192.530 82.650 192.730 ;
        RECT 86.575 192.685 86.865 192.730 ;
        RECT 87.110 192.590 87.250 193.070 ;
        RECT 90.255 193.025 90.545 193.070 ;
        RECT 93.920 192.870 94.240 192.930 ;
        RECT 87.570 192.730 94.240 192.870 ;
        RECT 78.830 192.390 82.650 192.530 ;
        RECT 78.830 192.190 78.970 192.390 ;
        RECT 82.895 192.345 83.185 192.575 ;
        RECT 86.115 192.530 86.405 192.575 ;
        RECT 87.020 192.530 87.340 192.590 ;
        RECT 87.570 192.575 87.710 192.730 ;
        RECT 93.920 192.670 94.240 192.730 ;
        RECT 86.115 192.390 87.340 192.530 ;
        RECT 86.115 192.345 86.405 192.390 ;
        RECT 75.060 192.050 78.970 192.190 ;
        RECT 79.200 192.190 79.520 192.250 ;
        RECT 82.420 192.190 82.740 192.250 ;
        RECT 79.200 192.050 82.740 192.190 ;
        RECT 82.970 192.190 83.110 192.345 ;
        RECT 87.020 192.330 87.340 192.390 ;
        RECT 87.495 192.345 87.785 192.575 ;
        RECT 89.335 192.530 89.625 192.575 ;
        RECT 89.780 192.530 90.100 192.590 ;
        RECT 89.335 192.390 90.100 192.530 ;
        RECT 89.335 192.345 89.625 192.390 ;
        RECT 89.780 192.330 90.100 192.390 ;
        RECT 90.700 192.330 91.020 192.590 ;
        RECT 92.095 192.345 92.385 192.575 ;
        RECT 83.340 192.190 83.660 192.250 ;
        RECT 82.970 192.050 83.660 192.190 ;
        RECT 75.060 191.990 75.380 192.050 ;
        RECT 79.200 191.990 79.520 192.050 ;
        RECT 82.420 191.990 82.740 192.050 ;
        RECT 83.340 191.990 83.660 192.050 ;
        RECT 83.800 192.190 84.120 192.250 ;
        RECT 85.195 192.190 85.485 192.235 ;
        RECT 83.800 192.050 85.485 192.190 ;
        RECT 83.800 191.990 84.120 192.050 ;
        RECT 85.195 192.005 85.485 192.050 ;
        RECT 91.175 192.190 91.465 192.235 ;
        RECT 91.620 192.190 91.940 192.250 ;
        RECT 91.175 192.050 91.940 192.190 ;
        RECT 92.170 192.190 92.310 192.345 ;
        RECT 92.540 192.330 92.860 192.590 ;
        RECT 93.000 192.330 93.320 192.590 ;
        RECT 94.380 192.330 94.700 192.590 ;
        RECT 94.930 192.575 95.070 193.070 ;
        RECT 98.995 193.025 99.285 193.070 ;
        RECT 103.620 193.210 103.910 193.255 ;
        RECT 105.720 193.210 106.010 193.255 ;
        RECT 107.290 193.210 107.580 193.255 ;
        RECT 103.620 193.070 107.580 193.210 ;
        RECT 103.620 193.025 103.910 193.070 ;
        RECT 105.720 193.025 106.010 193.070 ;
        RECT 107.290 193.025 107.580 193.070 ;
        RECT 104.015 192.870 104.305 192.915 ;
        RECT 105.205 192.870 105.495 192.915 ;
        RECT 107.725 192.870 108.015 192.915 ;
        RECT 104.015 192.730 108.015 192.870 ;
        RECT 104.015 192.685 104.305 192.730 ;
        RECT 105.205 192.685 105.495 192.730 ;
        RECT 107.725 192.685 108.015 192.730 ;
        RECT 94.855 192.530 95.145 192.575 ;
        RECT 95.760 192.530 96.080 192.590 ;
        RECT 94.855 192.390 96.080 192.530 ;
        RECT 94.855 192.345 95.145 192.390 ;
        RECT 95.760 192.330 96.080 192.390 ;
        RECT 97.140 192.330 97.460 192.590 ;
        RECT 98.060 192.330 98.380 192.590 ;
        RECT 99.440 192.330 99.760 192.590 ;
        RECT 101.295 192.345 101.585 192.575 ;
        RECT 97.230 192.190 97.370 192.330 ;
        RECT 92.170 192.050 97.370 192.190 ;
        RECT 91.175 192.005 91.465 192.050 ;
        RECT 91.620 191.990 91.940 192.050 ;
        RECT 100.360 191.990 100.680 192.250 ;
        RECT 73.220 191.710 74.830 191.850 ;
        RECT 73.220 191.650 73.540 191.710 ;
        RECT 77.360 191.650 77.680 191.910 ;
        RECT 84.260 191.650 84.580 191.910 ;
        RECT 84.720 191.650 85.040 191.910 ;
        RECT 88.415 191.850 88.705 191.895 ;
        RECT 89.320 191.850 89.640 191.910 ;
        RECT 88.415 191.710 89.640 191.850 ;
        RECT 88.415 191.665 88.705 191.710 ;
        RECT 89.320 191.650 89.640 191.710 ;
        RECT 92.540 191.850 92.860 191.910 ;
        RECT 97.155 191.850 97.445 191.895 ;
        RECT 92.540 191.710 97.445 191.850 ;
        RECT 101.370 191.850 101.510 192.345 ;
        RECT 102.660 192.330 102.980 192.590 ;
        RECT 103.135 192.530 103.425 192.575 ;
        RECT 106.800 192.530 107.120 192.590 ;
        RECT 110.020 192.530 110.340 192.590 ;
        RECT 103.135 192.390 110.340 192.530 ;
        RECT 103.135 192.345 103.425 192.390 ;
        RECT 106.800 192.330 107.120 192.390 ;
        RECT 110.020 192.330 110.340 192.390 ;
        RECT 113.240 192.330 113.560 192.590 ;
        RECT 103.580 192.190 103.900 192.250 ;
        RECT 104.360 192.190 104.650 192.235 ;
        RECT 103.580 192.050 104.650 192.190 ;
        RECT 103.580 191.990 103.900 192.050 ;
        RECT 104.360 192.005 104.650 192.050 ;
        RECT 105.880 192.190 106.200 192.250 ;
        RECT 110.495 192.190 110.785 192.235 ;
        RECT 105.880 192.050 110.785 192.190 ;
        RECT 105.880 191.990 106.200 192.050 ;
        RECT 110.495 192.005 110.785 192.050 ;
        RECT 104.960 191.850 105.280 191.910 ;
        RECT 101.370 191.710 105.280 191.850 ;
        RECT 92.540 191.650 92.860 191.710 ;
        RECT 97.155 191.665 97.445 191.710 ;
        RECT 104.960 191.650 105.280 191.710 ;
        RECT 110.035 191.850 110.325 191.895 ;
        RECT 113.240 191.850 113.560 191.910 ;
        RECT 110.035 191.710 113.560 191.850 ;
        RECT 110.035 191.665 110.325 191.710 ;
        RECT 113.240 191.650 113.560 191.710 ;
        RECT 61.190 191.030 116.270 191.510 ;
        RECT 81.960 190.830 82.280 190.890 ;
        RECT 82.435 190.830 82.725 190.875 ;
        RECT 81.960 190.690 82.725 190.830 ;
        RECT 81.960 190.630 82.280 190.690 ;
        RECT 82.435 190.645 82.725 190.690 ;
        RECT 90.700 190.830 91.020 190.890 ;
        RECT 92.095 190.830 92.385 190.875 ;
        RECT 90.700 190.690 92.385 190.830 ;
        RECT 90.700 190.630 91.020 190.690 ;
        RECT 92.095 190.645 92.385 190.690 ;
        RECT 93.000 190.830 93.320 190.890 ;
        RECT 95.775 190.830 96.065 190.875 ;
        RECT 93.000 190.690 96.065 190.830 ;
        RECT 93.000 190.630 93.320 190.690 ;
        RECT 95.775 190.645 96.065 190.690 ;
        RECT 96.220 190.830 96.540 190.890 ;
        RECT 98.980 190.830 99.300 190.890 ;
        RECT 100.375 190.830 100.665 190.875 ;
        RECT 96.220 190.690 100.665 190.830 ;
        RECT 96.220 190.630 96.540 190.690 ;
        RECT 98.980 190.630 99.300 190.690 ;
        RECT 100.375 190.645 100.665 190.690 ;
        RECT 103.120 190.630 103.440 190.890 ;
        RECT 109.575 190.830 109.865 190.875 ;
        RECT 110.940 190.830 111.260 190.890 ;
        RECT 109.575 190.690 111.260 190.830 ;
        RECT 109.575 190.645 109.865 190.690 ;
        RECT 110.940 190.630 111.260 190.690 ;
        RECT 111.400 190.630 111.720 190.890 ;
        RECT 76.900 190.490 77.220 190.550 ;
        RECT 74.230 190.350 77.220 190.490 ;
        RECT 72.300 189.950 72.620 190.210 ;
        RECT 73.220 190.150 73.540 190.210 ;
        RECT 74.230 190.195 74.370 190.350 ;
        RECT 76.900 190.290 77.220 190.350 ;
        RECT 96.680 190.490 97.000 190.550 ;
        RECT 98.520 190.490 98.840 190.550 ;
        RECT 100.835 190.490 101.125 190.535 ;
        RECT 96.680 190.350 101.125 190.490 ;
        RECT 96.680 190.290 97.000 190.350 ;
        RECT 98.520 190.290 98.840 190.350 ;
        RECT 100.835 190.305 101.125 190.350 ;
        RECT 103.210 190.350 108.870 190.490 ;
        RECT 103.210 190.210 103.350 190.350 ;
        RECT 75.520 190.195 75.840 190.210 ;
        RECT 73.695 190.150 73.985 190.195 ;
        RECT 73.220 190.010 73.985 190.150 ;
        RECT 73.220 189.950 73.540 190.010 ;
        RECT 73.695 189.965 73.985 190.010 ;
        RECT 74.155 189.965 74.445 190.195 ;
        RECT 75.490 190.150 75.840 190.195 ;
        RECT 75.325 190.010 75.840 190.150 ;
        RECT 75.490 189.965 75.840 190.010 ;
        RECT 75.520 189.950 75.840 189.965 ;
        RECT 84.720 190.150 85.040 190.210 ;
        RECT 90.255 190.150 90.545 190.195 ;
        RECT 84.720 190.010 90.545 190.150 ;
        RECT 84.720 189.950 85.040 190.010 ;
        RECT 90.255 189.965 90.545 190.010 ;
        RECT 96.220 190.150 96.540 190.210 ;
        RECT 97.155 190.150 97.445 190.195 ;
        RECT 96.220 190.010 97.445 190.150 ;
        RECT 96.220 189.950 96.540 190.010 ;
        RECT 97.155 189.965 97.445 190.010 ;
        RECT 97.615 190.150 97.905 190.195 ;
        RECT 98.995 190.150 99.285 190.195 ;
        RECT 97.615 190.010 99.285 190.150 ;
        RECT 97.615 189.965 97.905 190.010 ;
        RECT 98.995 189.965 99.285 190.010 ;
        RECT 99.915 189.965 100.205 190.195 ;
        RECT 75.035 189.810 75.325 189.855 ;
        RECT 76.225 189.810 76.515 189.855 ;
        RECT 78.745 189.810 79.035 189.855 ;
        RECT 75.035 189.670 79.035 189.810 ;
        RECT 75.035 189.625 75.325 189.670 ;
        RECT 76.225 189.625 76.515 189.670 ;
        RECT 78.745 189.625 79.035 189.670 ;
        RECT 85.640 189.610 85.960 189.870 ;
        RECT 94.380 189.810 94.700 189.870 ;
        RECT 95.315 189.810 95.605 189.855 ;
        RECT 94.380 189.670 95.605 189.810 ;
        RECT 94.380 189.610 94.700 189.670 ;
        RECT 95.315 189.625 95.605 189.670 ;
        RECT 95.760 189.810 96.080 189.870 ;
        RECT 96.695 189.810 96.985 189.855 ;
        RECT 97.690 189.810 97.830 189.965 ;
        RECT 95.760 189.670 96.985 189.810 ;
        RECT 74.640 189.470 74.930 189.515 ;
        RECT 76.740 189.470 77.030 189.515 ;
        RECT 78.310 189.470 78.600 189.515 ;
        RECT 74.640 189.330 78.600 189.470 ;
        RECT 95.390 189.470 95.530 189.625 ;
        RECT 95.760 189.610 96.080 189.670 ;
        RECT 96.695 189.625 96.985 189.670 ;
        RECT 97.230 189.670 97.830 189.810 ;
        RECT 98.075 189.810 98.365 189.855 ;
        RECT 99.440 189.810 99.760 189.870 ;
        RECT 98.075 189.670 99.760 189.810 ;
        RECT 99.990 189.810 100.130 189.965 ;
        RECT 103.120 189.950 103.440 190.210 ;
        RECT 105.420 190.150 105.740 190.210 ;
        RECT 108.730 190.195 108.870 190.350 ;
        RECT 110.480 190.290 110.800 190.550 ;
        RECT 107.735 190.150 108.025 190.195 ;
        RECT 105.420 190.010 108.025 190.150 ;
        RECT 105.420 189.950 105.740 190.010 ;
        RECT 107.735 189.965 108.025 190.010 ;
        RECT 108.655 190.150 108.945 190.195 ;
        RECT 110.955 190.150 111.245 190.195 ;
        RECT 108.655 190.010 111.245 190.150 ;
        RECT 108.655 189.965 108.945 190.010 ;
        RECT 110.955 189.965 111.245 190.010 ;
        RECT 104.040 189.810 104.360 189.870 ;
        RECT 105.895 189.810 106.185 189.855 ;
        RECT 99.990 189.670 106.185 189.810 ;
        RECT 97.230 189.530 97.370 189.670 ;
        RECT 98.075 189.625 98.365 189.670 ;
        RECT 99.440 189.610 99.760 189.670 ;
        RECT 104.040 189.610 104.360 189.670 ;
        RECT 105.895 189.625 106.185 189.670 ;
        RECT 107.260 189.810 107.580 189.870 ;
        RECT 109.115 189.810 109.405 189.855 ;
        RECT 114.160 189.810 114.480 189.870 ;
        RECT 107.260 189.670 109.405 189.810 ;
        RECT 107.260 189.610 107.580 189.670 ;
        RECT 109.115 189.625 109.405 189.670 ;
        RECT 109.650 189.670 114.480 189.810 ;
        RECT 97.140 189.470 97.460 189.530 ;
        RECT 109.650 189.470 109.790 189.670 ;
        RECT 114.160 189.610 114.480 189.670 ;
        RECT 95.390 189.330 97.460 189.470 ;
        RECT 74.640 189.285 74.930 189.330 ;
        RECT 76.740 189.285 77.030 189.330 ;
        RECT 78.310 189.285 78.600 189.330 ;
        RECT 97.140 189.270 97.460 189.330 ;
        RECT 98.150 189.330 109.790 189.470 ;
        RECT 112.335 189.470 112.625 189.515 ;
        RECT 113.240 189.470 113.560 189.530 ;
        RECT 112.335 189.330 113.560 189.470 ;
        RECT 71.380 188.930 71.700 189.190 ;
        RECT 73.220 188.930 73.540 189.190 ;
        RECT 75.060 189.130 75.380 189.190 ;
        RECT 81.055 189.130 81.345 189.175 ;
        RECT 83.340 189.130 83.660 189.190 ;
        RECT 85.180 189.130 85.500 189.190 ;
        RECT 75.060 188.990 85.500 189.130 ;
        RECT 75.060 188.930 75.380 188.990 ;
        RECT 81.055 188.945 81.345 188.990 ;
        RECT 83.340 188.930 83.660 188.990 ;
        RECT 85.180 188.930 85.500 188.990 ;
        RECT 86.100 189.130 86.420 189.190 ;
        RECT 87.495 189.130 87.785 189.175 ;
        RECT 86.100 188.990 87.785 189.130 ;
        RECT 86.100 188.930 86.420 188.990 ;
        RECT 87.495 188.945 87.785 188.990 ;
        RECT 90.240 189.130 90.560 189.190 ;
        RECT 98.150 189.130 98.290 189.330 ;
        RECT 112.335 189.285 112.625 189.330 ;
        RECT 113.240 189.270 113.560 189.330 ;
        RECT 90.240 188.990 98.290 189.130 ;
        RECT 101.755 189.130 102.045 189.175 ;
        RECT 104.500 189.130 104.820 189.190 ;
        RECT 101.755 188.990 104.820 189.130 ;
        RECT 90.240 188.930 90.560 188.990 ;
        RECT 101.755 188.945 102.045 188.990 ;
        RECT 104.500 188.930 104.820 188.990 ;
        RECT 106.340 189.130 106.660 189.190 ;
        RECT 106.815 189.130 107.105 189.175 ;
        RECT 106.340 188.990 107.105 189.130 ;
        RECT 106.340 188.930 106.660 188.990 ;
        RECT 106.815 188.945 107.105 188.990 ;
        RECT 61.190 188.310 115.470 188.790 ;
        RECT 70.475 188.110 70.765 188.155 ;
        RECT 73.220 188.110 73.540 188.170 ;
        RECT 70.475 187.970 73.540 188.110 ;
        RECT 70.475 187.925 70.765 187.970 ;
        RECT 73.220 187.910 73.540 187.970 ;
        RECT 75.535 188.110 75.825 188.155 ;
        RECT 75.980 188.110 76.300 188.170 ;
        RECT 84.260 188.110 84.580 188.170 ;
        RECT 75.535 187.970 84.580 188.110 ;
        RECT 75.535 187.925 75.825 187.970 ;
        RECT 67.255 187.430 67.545 187.475 ;
        RECT 71.380 187.430 71.700 187.490 ;
        RECT 67.255 187.290 71.700 187.430 ;
        RECT 67.255 187.245 67.545 187.290 ;
        RECT 71.380 187.230 71.700 187.290 ;
        RECT 73.695 187.430 73.985 187.475 ;
        RECT 75.610 187.430 75.750 187.925 ;
        RECT 75.980 187.910 76.300 187.970 ;
        RECT 84.260 187.910 84.580 187.970 ;
        RECT 85.640 187.910 85.960 188.170 ;
        RECT 93.475 188.110 93.765 188.155 ;
        RECT 93.920 188.110 94.240 188.170 ;
        RECT 93.475 187.970 94.240 188.110 ;
        RECT 93.475 187.925 93.765 187.970 ;
        RECT 93.920 187.910 94.240 187.970 ;
        RECT 95.315 188.110 95.605 188.155 ;
        RECT 98.060 188.110 98.380 188.170 ;
        RECT 95.315 187.970 98.380 188.110 ;
        RECT 95.315 187.925 95.605 187.970 ;
        RECT 98.060 187.910 98.380 187.970 ;
        RECT 99.440 187.910 99.760 188.170 ;
        RECT 104.960 187.910 105.280 188.170 ;
        RECT 77.400 187.770 77.690 187.815 ;
        RECT 79.500 187.770 79.790 187.815 ;
        RECT 81.070 187.770 81.360 187.815 ;
        RECT 77.400 187.630 81.360 187.770 ;
        RECT 77.400 187.585 77.690 187.630 ;
        RECT 79.500 187.585 79.790 187.630 ;
        RECT 81.070 187.585 81.360 187.630 ;
        RECT 87.060 187.770 87.350 187.815 ;
        RECT 89.160 187.770 89.450 187.815 ;
        RECT 90.730 187.770 91.020 187.815 ;
        RECT 87.060 187.630 91.020 187.770 ;
        RECT 87.060 187.585 87.350 187.630 ;
        RECT 89.160 187.585 89.450 187.630 ;
        RECT 90.730 187.585 91.020 187.630 ;
        RECT 73.695 187.290 75.750 187.430 ;
        RECT 77.795 187.430 78.085 187.475 ;
        RECT 78.985 187.430 79.275 187.475 ;
        RECT 81.505 187.430 81.795 187.475 ;
        RECT 77.795 187.290 81.795 187.430 ;
        RECT 73.695 187.245 73.985 187.290 ;
        RECT 77.795 187.245 78.085 187.290 ;
        RECT 78.985 187.245 79.275 187.290 ;
        RECT 81.505 187.245 81.795 187.290 ;
        RECT 87.455 187.430 87.745 187.475 ;
        RECT 88.645 187.430 88.935 187.475 ;
        RECT 91.165 187.430 91.455 187.475 ;
        RECT 87.455 187.290 91.455 187.430 ;
        RECT 87.455 187.245 87.745 187.290 ;
        RECT 88.645 187.245 88.935 187.290 ;
        RECT 91.165 187.245 91.455 187.290 ;
        RECT 104.500 187.230 104.820 187.490 ;
        RECT 109.575 187.430 109.865 187.475 ;
        RECT 112.320 187.430 112.640 187.490 ;
        RECT 109.575 187.290 112.640 187.430 ;
        RECT 109.575 187.245 109.865 187.290 ;
        RECT 112.320 187.230 112.640 187.290 ;
        RECT 76.900 186.890 77.220 187.150 ;
        RECT 77.360 187.090 77.680 187.150 ;
        RECT 78.195 187.090 78.485 187.135 ;
        RECT 77.360 186.950 78.485 187.090 ;
        RECT 77.360 186.890 77.680 186.950 ;
        RECT 78.195 186.905 78.485 186.950 ;
        RECT 84.260 186.890 84.580 187.150 ;
        RECT 84.720 186.890 85.040 187.150 ;
        RECT 85.655 187.090 85.945 187.135 ;
        RECT 86.100 187.090 86.420 187.150 ;
        RECT 85.655 186.950 86.420 187.090 ;
        RECT 85.655 186.905 85.945 186.950 ;
        RECT 86.100 186.890 86.420 186.950 ;
        RECT 86.560 186.890 86.880 187.150 ;
        RECT 87.910 187.090 88.200 187.135 ;
        RECT 89.320 187.090 89.640 187.150 ;
        RECT 87.910 186.950 89.640 187.090 ;
        RECT 87.910 186.905 88.200 186.950 ;
        RECT 89.320 186.890 89.640 186.950 ;
        RECT 93.920 186.890 94.240 187.150 ;
        RECT 96.695 187.090 96.985 187.135 ;
        RECT 97.140 187.090 97.460 187.150 ;
        RECT 96.695 186.950 97.460 187.090 ;
        RECT 96.695 186.905 96.985 186.950 ;
        RECT 97.140 186.890 97.460 186.950 ;
        RECT 103.120 187.090 103.440 187.150 ;
        RECT 104.975 187.090 105.265 187.135 ;
        RECT 103.120 186.950 105.265 187.090 ;
        RECT 103.120 186.890 103.440 186.950 ;
        RECT 104.975 186.905 105.265 186.950 ;
        RECT 105.895 186.905 106.185 187.135 ;
        RECT 110.495 187.090 110.785 187.135 ;
        RECT 110.940 187.090 111.260 187.150 ;
        RECT 110.495 186.950 111.260 187.090 ;
        RECT 110.495 186.905 110.785 186.950 ;
        RECT 70.015 186.750 70.305 186.795 ;
        RECT 70.920 186.750 71.240 186.810 ;
        RECT 70.015 186.610 71.240 186.750 ;
        RECT 70.015 186.565 70.305 186.610 ;
        RECT 70.920 186.550 71.240 186.610 ;
        RECT 73.220 186.750 73.540 186.810 ;
        RECT 74.615 186.750 74.905 186.795 ;
        RECT 75.060 186.750 75.380 186.810 ;
        RECT 73.220 186.610 75.380 186.750 ;
        RECT 73.220 186.550 73.540 186.610 ;
        RECT 74.615 186.565 74.905 186.610 ;
        RECT 75.060 186.550 75.380 186.610 ;
        RECT 75.695 186.750 75.985 186.795 ;
        RECT 84.810 186.750 84.950 186.890 ;
        RECT 75.695 186.610 84.950 186.750 ;
        RECT 92.080 186.750 92.400 186.810 ;
        RECT 95.315 186.750 95.605 186.795 ;
        RECT 98.060 186.750 98.380 186.810 ;
        RECT 92.080 186.610 98.380 186.750 ;
        RECT 75.695 186.565 75.985 186.610 ;
        RECT 76.440 186.210 76.760 186.470 ;
        RECT 83.890 186.455 84.030 186.610 ;
        RECT 92.080 186.550 92.400 186.610 ;
        RECT 95.315 186.565 95.605 186.610 ;
        RECT 98.060 186.550 98.380 186.610 ;
        RECT 99.440 186.750 99.760 186.810 ;
        RECT 105.970 186.750 106.110 186.905 ;
        RECT 110.940 186.890 111.260 186.950 ;
        RECT 99.440 186.610 106.110 186.750 ;
        RECT 99.440 186.550 99.760 186.610 ;
        RECT 83.815 186.225 84.105 186.455 ;
        RECT 84.735 186.410 85.025 186.455 ;
        RECT 85.180 186.410 85.500 186.470 ;
        RECT 84.735 186.270 85.500 186.410 ;
        RECT 84.735 186.225 85.025 186.270 ;
        RECT 85.180 186.210 85.500 186.270 ;
        RECT 94.395 186.410 94.685 186.455 ;
        RECT 98.980 186.410 99.300 186.470 ;
        RECT 94.395 186.270 99.300 186.410 ;
        RECT 94.395 186.225 94.685 186.270 ;
        RECT 98.980 186.210 99.300 186.270 ;
        RECT 104.500 186.410 104.820 186.470 ;
        RECT 106.355 186.410 106.645 186.455 ;
        RECT 107.260 186.410 107.580 186.470 ;
        RECT 104.500 186.270 107.580 186.410 ;
        RECT 104.500 186.210 104.820 186.270 ;
        RECT 106.355 186.225 106.645 186.270 ;
        RECT 107.260 186.210 107.580 186.270 ;
        RECT 111.860 186.410 112.180 186.470 ;
        RECT 113.255 186.410 113.545 186.455 ;
        RECT 111.860 186.270 113.545 186.410 ;
        RECT 111.860 186.210 112.180 186.270 ;
        RECT 113.255 186.225 113.545 186.270 ;
        RECT 61.190 185.590 116.270 186.070 ;
        RECT 75.980 185.390 76.300 185.450 ;
        RECT 76.455 185.390 76.745 185.435 ;
        RECT 75.980 185.250 76.745 185.390 ;
        RECT 75.980 185.190 76.300 185.250 ;
        RECT 76.455 185.205 76.745 185.250 ;
        RECT 104.040 185.390 104.360 185.450 ;
        RECT 104.515 185.390 104.805 185.435 ;
        RECT 104.040 185.250 104.805 185.390 ;
        RECT 104.040 185.190 104.360 185.250 ;
        RECT 104.515 185.205 104.805 185.250 ;
        RECT 111.875 185.390 112.165 185.435 ;
        RECT 112.320 185.390 112.640 185.450 ;
        RECT 111.875 185.250 112.640 185.390 ;
        RECT 111.875 185.205 112.165 185.250 ;
        RECT 112.320 185.190 112.640 185.250 ;
        RECT 86.560 185.050 86.880 185.110 ;
        RECT 93.920 185.050 94.240 185.110 ;
        RECT 69.630 184.910 86.880 185.050 ;
        RECT 69.630 184.755 69.770 184.910 ;
        RECT 70.920 184.755 71.240 184.770 ;
        RECT 69.555 184.525 69.845 184.755 ;
        RECT 70.890 184.710 71.240 184.755 ;
        RECT 77.910 184.710 78.050 184.910 ;
        RECT 86.560 184.850 86.880 184.910 ;
        RECT 90.790 184.910 94.240 185.050 ;
        RECT 78.280 184.755 78.600 184.770 ;
        RECT 70.890 184.570 71.390 184.710 ;
        RECT 77.450 184.570 78.050 184.710 ;
        RECT 70.890 184.525 71.240 184.570 ;
        RECT 70.920 184.510 71.240 184.525 ;
        RECT 70.435 184.370 70.725 184.415 ;
        RECT 71.625 184.370 71.915 184.415 ;
        RECT 74.145 184.370 74.435 184.415 ;
        RECT 70.435 184.230 74.435 184.370 ;
        RECT 70.435 184.185 70.725 184.230 ;
        RECT 71.625 184.185 71.915 184.230 ;
        RECT 74.145 184.185 74.435 184.230 ;
        RECT 76.900 184.370 77.220 184.430 ;
        RECT 77.450 184.370 77.590 184.570 ;
        RECT 78.250 184.525 78.600 184.755 ;
        RECT 78.280 184.510 78.600 184.525 ;
        RECT 79.660 184.710 79.980 184.770 ;
        RECT 84.275 184.710 84.565 184.755 ;
        RECT 79.660 184.570 84.565 184.710 ;
        RECT 79.660 184.510 79.980 184.570 ;
        RECT 84.275 184.525 84.565 184.570 ;
        RECT 85.195 184.710 85.485 184.755 ;
        RECT 87.020 184.710 87.340 184.770 ;
        RECT 85.195 184.570 87.340 184.710 ;
        RECT 85.195 184.525 85.485 184.570 ;
        RECT 76.900 184.230 77.590 184.370 ;
        RECT 77.795 184.370 78.085 184.415 ;
        RECT 78.985 184.370 79.275 184.415 ;
        RECT 81.505 184.370 81.795 184.415 ;
        RECT 77.795 184.230 81.795 184.370 ;
        RECT 84.350 184.370 84.490 184.525 ;
        RECT 87.020 184.510 87.340 184.570 ;
        RECT 88.860 184.510 89.180 184.770 ;
        RECT 89.795 184.710 90.085 184.755 ;
        RECT 90.790 184.710 90.930 184.910 ;
        RECT 93.920 184.850 94.240 184.910 ;
        RECT 91.620 184.755 91.940 184.770 ;
        RECT 91.590 184.710 91.940 184.755 ;
        RECT 89.795 184.570 90.930 184.710 ;
        RECT 91.425 184.570 91.940 184.710 ;
        RECT 89.795 184.525 90.085 184.570 ;
        RECT 91.590 184.525 91.940 184.570 ;
        RECT 98.950 184.710 99.240 184.755 ;
        RECT 100.360 184.710 100.680 184.770 ;
        RECT 106.340 184.755 106.660 184.770 ;
        RECT 106.310 184.710 106.660 184.755 ;
        RECT 98.950 184.570 100.680 184.710 ;
        RECT 106.145 184.570 106.660 184.710 ;
        RECT 98.950 184.525 99.240 184.570 ;
        RECT 91.620 184.510 91.940 184.525 ;
        RECT 100.360 184.510 100.680 184.570 ;
        RECT 106.310 184.525 106.660 184.570 ;
        RECT 106.340 184.510 106.660 184.525 ;
        RECT 88.905 184.370 89.045 184.510 ;
        RECT 84.350 184.230 89.045 184.370 ;
        RECT 76.900 184.170 77.220 184.230 ;
        RECT 77.795 184.185 78.085 184.230 ;
        RECT 78.985 184.185 79.275 184.230 ;
        RECT 81.505 184.185 81.795 184.230 ;
        RECT 90.255 184.185 90.545 184.415 ;
        RECT 91.135 184.370 91.425 184.415 ;
        RECT 92.325 184.370 92.615 184.415 ;
        RECT 94.845 184.370 95.135 184.415 ;
        RECT 91.135 184.230 95.135 184.370 ;
        RECT 91.135 184.185 91.425 184.230 ;
        RECT 92.325 184.185 92.615 184.230 ;
        RECT 94.845 184.185 95.135 184.230 ;
        RECT 97.615 184.185 97.905 184.415 ;
        RECT 98.495 184.370 98.785 184.415 ;
        RECT 99.685 184.370 99.975 184.415 ;
        RECT 102.205 184.370 102.495 184.415 ;
        RECT 98.495 184.230 102.495 184.370 ;
        RECT 98.495 184.185 98.785 184.230 ;
        RECT 99.685 184.185 99.975 184.230 ;
        RECT 102.205 184.185 102.495 184.230 ;
        RECT 104.975 184.185 105.265 184.415 ;
        RECT 105.855 184.370 106.145 184.415 ;
        RECT 107.045 184.370 107.335 184.415 ;
        RECT 109.565 184.370 109.855 184.415 ;
        RECT 105.855 184.230 109.855 184.370 ;
        RECT 105.855 184.185 106.145 184.230 ;
        RECT 107.045 184.185 107.335 184.230 ;
        RECT 109.565 184.185 109.855 184.230 ;
        RECT 70.040 184.030 70.330 184.075 ;
        RECT 72.140 184.030 72.430 184.075 ;
        RECT 73.710 184.030 74.000 184.075 ;
        RECT 70.040 183.890 74.000 184.030 ;
        RECT 70.040 183.845 70.330 183.890 ;
        RECT 72.140 183.845 72.430 183.890 ;
        RECT 73.710 183.845 74.000 183.890 ;
        RECT 77.400 184.030 77.690 184.075 ;
        RECT 79.500 184.030 79.790 184.075 ;
        RECT 81.070 184.030 81.360 184.075 ;
        RECT 77.400 183.890 81.360 184.030 ;
        RECT 77.400 183.845 77.690 183.890 ;
        RECT 79.500 183.845 79.790 183.890 ;
        RECT 81.070 183.845 81.360 183.890 ;
        RECT 83.800 183.830 84.120 184.090 ;
        RECT 89.780 183.830 90.100 184.090 ;
        RECT 85.180 183.490 85.500 183.750 ;
        RECT 90.330 183.690 90.470 184.185 ;
        RECT 90.740 184.030 91.030 184.075 ;
        RECT 92.840 184.030 93.130 184.075 ;
        RECT 94.410 184.030 94.700 184.075 ;
        RECT 97.690 184.030 97.830 184.185 ;
        RECT 90.740 183.890 94.700 184.030 ;
        RECT 90.740 183.845 91.030 183.890 ;
        RECT 92.840 183.845 93.130 183.890 ;
        RECT 94.410 183.845 94.700 183.890 ;
        RECT 94.930 183.890 97.830 184.030 ;
        RECT 94.930 183.690 95.070 183.890 ;
        RECT 90.330 183.550 95.070 183.690 ;
        RECT 97.140 183.490 97.460 183.750 ;
        RECT 97.690 183.690 97.830 183.890 ;
        RECT 98.100 184.030 98.390 184.075 ;
        RECT 100.200 184.030 100.490 184.075 ;
        RECT 101.770 184.030 102.060 184.075 ;
        RECT 105.050 184.030 105.190 184.185 ;
        RECT 98.100 183.890 102.060 184.030 ;
        RECT 98.100 183.845 98.390 183.890 ;
        RECT 100.200 183.845 100.490 183.890 ;
        RECT 101.770 183.845 102.060 183.890 ;
        RECT 102.290 183.890 105.190 184.030 ;
        RECT 102.290 183.690 102.430 183.890 ;
        RECT 97.690 183.550 102.430 183.690 ;
        RECT 105.050 183.690 105.190 183.890 ;
        RECT 105.460 184.030 105.750 184.075 ;
        RECT 107.560 184.030 107.850 184.075 ;
        RECT 109.130 184.030 109.420 184.075 ;
        RECT 105.460 183.890 109.420 184.030 ;
        RECT 105.460 183.845 105.750 183.890 ;
        RECT 107.560 183.845 107.850 183.890 ;
        RECT 109.130 183.845 109.420 183.890 ;
        RECT 106.800 183.690 107.120 183.750 ;
        RECT 105.050 183.550 107.120 183.690 ;
        RECT 106.800 183.490 107.120 183.550 ;
        RECT 61.190 182.870 115.470 183.350 ;
        RECT 72.300 182.670 72.620 182.730 ;
        RECT 76.915 182.670 77.205 182.715 ;
        RECT 72.300 182.530 77.205 182.670 ;
        RECT 72.300 182.470 72.620 182.530 ;
        RECT 76.915 182.485 77.205 182.530 ;
        RECT 78.280 182.670 78.600 182.730 ;
        RECT 79.215 182.670 79.505 182.715 ;
        RECT 78.280 182.530 79.505 182.670 ;
        RECT 78.280 182.470 78.600 182.530 ;
        RECT 79.215 182.485 79.505 182.530 ;
        RECT 88.860 182.670 89.180 182.730 ;
        RECT 88.860 182.530 95.070 182.670 ;
        RECT 88.860 182.470 89.180 182.530 ;
        RECT 76.440 182.330 76.760 182.390 ;
        RECT 81.055 182.330 81.345 182.375 ;
        RECT 76.440 182.190 81.345 182.330 ;
        RECT 76.440 182.130 76.760 182.190 ;
        RECT 81.055 182.145 81.345 182.190 ;
        RECT 87.980 182.330 88.270 182.375 ;
        RECT 90.080 182.330 90.370 182.375 ;
        RECT 91.650 182.330 91.940 182.375 ;
        RECT 87.980 182.190 91.940 182.330 ;
        RECT 87.980 182.145 88.270 182.190 ;
        RECT 90.080 182.145 90.370 182.190 ;
        RECT 91.650 182.145 91.940 182.190 ;
        RECT 94.395 182.145 94.685 182.375 ;
        RECT 94.930 182.330 95.070 182.530 ;
        RECT 98.980 182.470 99.300 182.730 ;
        RECT 103.135 182.670 103.425 182.715 ;
        RECT 103.580 182.670 103.900 182.730 ;
        RECT 103.135 182.530 103.900 182.670 ;
        RECT 103.135 182.485 103.425 182.530 ;
        RECT 103.580 182.470 103.900 182.530 ;
        RECT 105.895 182.670 106.185 182.715 ;
        RECT 107.720 182.670 108.040 182.730 ;
        RECT 109.560 182.670 109.880 182.730 ;
        RECT 105.895 182.530 109.880 182.670 ;
        RECT 105.895 182.485 106.185 182.530 ;
        RECT 107.720 182.470 108.040 182.530 ;
        RECT 109.560 182.470 109.880 182.530 ;
        RECT 99.440 182.330 99.760 182.390 ;
        RECT 100.360 182.330 100.680 182.390 ;
        RECT 101.755 182.330 102.045 182.375 ;
        RECT 94.930 182.190 102.045 182.330 ;
        RECT 85.180 181.990 85.500 182.050 ;
        RECT 80.210 181.850 85.500 181.990 ;
        RECT 75.980 181.650 76.300 181.710 ;
        RECT 80.210 181.695 80.350 181.850 ;
        RECT 85.180 181.790 85.500 181.850 ;
        RECT 86.560 181.990 86.880 182.050 ;
        RECT 87.495 181.990 87.785 182.035 ;
        RECT 86.560 181.850 87.785 181.990 ;
        RECT 86.560 181.790 86.880 181.850 ;
        RECT 87.495 181.805 87.785 181.850 ;
        RECT 88.375 181.990 88.665 182.035 ;
        RECT 89.565 181.990 89.855 182.035 ;
        RECT 92.085 181.990 92.375 182.035 ;
        RECT 88.375 181.850 92.375 181.990 ;
        RECT 94.470 181.990 94.610 182.145 ;
        RECT 99.440 182.130 99.760 182.190 ;
        RECT 100.360 182.130 100.680 182.190 ;
        RECT 101.755 182.145 102.045 182.190 ;
        RECT 108.640 182.330 108.930 182.375 ;
        RECT 110.210 182.330 110.500 182.375 ;
        RECT 112.310 182.330 112.600 182.375 ;
        RECT 108.640 182.190 112.600 182.330 ;
        RECT 108.640 182.145 108.930 182.190 ;
        RECT 110.210 182.145 110.500 182.190 ;
        RECT 112.310 182.145 112.600 182.190 ;
        RECT 96.220 181.990 96.540 182.050 ;
        RECT 94.470 181.850 96.540 181.990 ;
        RECT 88.375 181.805 88.665 181.850 ;
        RECT 89.565 181.805 89.855 181.850 ;
        RECT 92.085 181.805 92.375 181.850 ;
        RECT 96.220 181.790 96.540 181.850 ;
        RECT 105.435 181.990 105.725 182.035 ;
        RECT 105.880 181.990 106.200 182.050 ;
        RECT 105.435 181.850 106.200 181.990 ;
        RECT 105.435 181.805 105.725 181.850 ;
        RECT 105.880 181.790 106.200 181.850 ;
        RECT 108.205 181.990 108.495 182.035 ;
        RECT 110.725 181.990 111.015 182.035 ;
        RECT 111.915 181.990 112.205 182.035 ;
        RECT 108.205 181.850 112.205 181.990 ;
        RECT 108.205 181.805 108.495 181.850 ;
        RECT 110.725 181.805 111.015 181.850 ;
        RECT 111.915 181.805 112.205 181.850 ;
        RECT 78.295 181.650 78.585 181.695 ;
        RECT 75.980 181.510 78.585 181.650 ;
        RECT 75.980 181.450 76.300 181.510 ;
        RECT 78.295 181.465 78.585 181.510 ;
        RECT 80.135 181.465 80.425 181.695 ;
        RECT 81.515 181.650 81.805 181.695 ;
        RECT 82.895 181.650 83.185 181.695 ;
        RECT 81.515 181.510 83.185 181.650 ;
        RECT 81.515 181.465 81.805 181.510 ;
        RECT 82.895 181.465 83.185 181.510 ;
        RECT 83.800 181.650 84.120 181.710 ;
        RECT 85.655 181.650 85.945 181.695 ;
        RECT 83.800 181.510 85.945 181.650 ;
        RECT 83.800 181.450 84.120 181.510 ;
        RECT 85.655 181.465 85.945 181.510 ;
        RECT 88.830 181.650 89.120 181.695 ;
        RECT 92.540 181.650 92.860 181.710 ;
        RECT 88.830 181.510 92.860 181.650 ;
        RECT 88.830 181.465 89.120 181.510 ;
        RECT 92.540 181.450 92.860 181.510 ;
        RECT 102.660 181.450 102.980 181.710 ;
        RECT 104.040 181.450 104.360 181.710 ;
        RECT 104.975 181.465 105.265 181.695 ;
        RECT 106.800 181.650 107.120 181.710 ;
        RECT 112.795 181.650 113.085 181.695 ;
        RECT 106.800 181.510 113.085 181.650 ;
        RECT 76.915 181.310 77.205 181.355 ;
        RECT 79.200 181.310 79.520 181.370 ;
        RECT 76.915 181.170 79.520 181.310 ;
        RECT 105.050 181.310 105.190 181.465 ;
        RECT 106.800 181.450 107.120 181.510 ;
        RECT 112.795 181.465 113.085 181.510 ;
        RECT 110.020 181.310 110.340 181.370 ;
        RECT 105.050 181.170 110.340 181.310 ;
        RECT 76.915 181.125 77.205 181.170 ;
        RECT 79.200 181.110 79.520 181.170 ;
        RECT 110.020 181.110 110.340 181.170 ;
        RECT 111.570 181.310 111.860 181.355 ;
        RECT 112.320 181.310 112.640 181.370 ;
        RECT 111.570 181.170 112.640 181.310 ;
        RECT 111.570 181.125 111.860 181.170 ;
        RECT 112.320 181.110 112.640 181.170 ;
        RECT 73.220 180.970 73.540 181.030 ;
        RECT 77.835 180.970 78.125 181.015 ;
        RECT 73.220 180.830 78.125 180.970 ;
        RECT 73.220 180.770 73.540 180.830 ;
        RECT 77.835 180.785 78.125 180.830 ;
        RECT 98.060 180.970 98.380 181.030 ;
        RECT 105.880 180.970 106.200 181.030 ;
        RECT 98.060 180.830 106.200 180.970 ;
        RECT 98.060 180.770 98.380 180.830 ;
        RECT 105.880 180.770 106.200 180.830 ;
        RECT 61.190 180.150 116.270 180.630 ;
        RECT 96.680 179.750 97.000 180.010 ;
        RECT 102.215 179.950 102.505 179.995 ;
        RECT 104.040 179.950 104.360 180.010 ;
        RECT 102.215 179.810 104.360 179.950 ;
        RECT 102.215 179.765 102.505 179.810 ;
        RECT 104.040 179.750 104.360 179.810 ;
        RECT 104.500 179.750 104.820 180.010 ;
        RECT 111.875 179.950 112.165 179.995 ;
        RECT 112.780 179.950 113.100 180.010 ;
        RECT 111.875 179.810 113.100 179.950 ;
        RECT 111.875 179.765 112.165 179.810 ;
        RECT 112.780 179.750 113.100 179.810 ;
        RECT 96.220 179.610 96.540 179.670 ;
        RECT 95.390 179.470 96.540 179.610 ;
        RECT 95.390 179.315 95.530 179.470 ;
        RECT 96.220 179.410 96.540 179.470 ;
        RECT 99.900 179.610 100.220 179.670 ;
        RECT 109.560 179.610 109.880 179.670 ;
        RECT 99.900 179.470 109.880 179.610 ;
        RECT 99.900 179.410 100.220 179.470 ;
        RECT 95.315 179.085 95.605 179.315 ;
        RECT 95.775 179.270 96.065 179.315 ;
        RECT 97.140 179.270 97.460 179.330 ;
        RECT 95.775 179.130 97.460 179.270 ;
        RECT 95.775 179.085 96.065 179.130 ;
        RECT 97.140 179.070 97.460 179.130 ;
        RECT 100.360 179.270 100.680 179.330 ;
        RECT 102.750 179.315 102.890 179.470 ;
        RECT 109.560 179.410 109.880 179.470 ;
        RECT 101.755 179.270 102.045 179.315 ;
        RECT 100.360 179.130 102.045 179.270 ;
        RECT 100.360 179.070 100.680 179.130 ;
        RECT 101.755 179.085 102.045 179.130 ;
        RECT 102.675 179.085 102.965 179.315 ;
        RECT 103.120 179.270 103.440 179.330 ;
        RECT 104.055 179.270 104.345 179.315 ;
        RECT 103.120 179.130 104.345 179.270 ;
        RECT 103.120 179.070 103.440 179.130 ;
        RECT 104.055 179.085 104.345 179.130 ;
        RECT 105.435 179.270 105.725 179.315 ;
        RECT 105.880 179.270 106.200 179.330 ;
        RECT 105.435 179.130 106.200 179.270 ;
        RECT 105.435 179.085 105.725 179.130 ;
        RECT 104.130 178.930 104.270 179.085 ;
        RECT 105.880 179.070 106.200 179.130 ;
        RECT 107.720 179.070 108.040 179.330 ;
        RECT 110.495 179.270 110.785 179.315 ;
        RECT 110.955 179.270 111.245 179.315 ;
        RECT 110.495 179.130 111.245 179.270 ;
        RECT 110.495 179.085 110.785 179.130 ;
        RECT 110.955 179.085 111.245 179.130 ;
        RECT 112.335 179.085 112.625 179.315 ;
        RECT 111.400 178.930 111.720 178.990 ;
        RECT 112.410 178.930 112.550 179.085 ;
        RECT 104.130 178.790 112.550 178.930 ;
        RECT 111.400 178.730 111.720 178.790 ;
        RECT 105.420 178.390 105.740 178.650 ;
        RECT 110.940 178.390 111.260 178.650 ;
        RECT 61.190 177.430 115.470 177.910 ;
        RECT 110.020 177.030 110.340 177.290 ;
        RECT 111.400 177.030 111.720 177.290 ;
        RECT 109.560 176.890 109.880 176.950 ;
        RECT 110.495 176.890 110.785 176.935 ;
        RECT 109.560 176.750 110.785 176.890 ;
        RECT 109.560 176.690 109.880 176.750 ;
        RECT 110.495 176.705 110.785 176.750 ;
        RECT 108.195 176.550 108.485 176.595 ;
        RECT 111.490 176.550 111.630 177.030 ;
        RECT 108.195 176.410 111.630 176.550 ;
        RECT 108.195 176.365 108.485 176.410 ;
        RECT 109.115 176.210 109.405 176.255 ;
        RECT 110.480 176.210 110.800 176.270 ;
        RECT 109.115 176.070 110.800 176.210 ;
        RECT 109.115 176.025 109.405 176.070 ;
        RECT 110.480 176.010 110.800 176.070 ;
        RECT 110.570 175.870 110.710 176.010 ;
        RECT 111.255 175.870 111.545 175.915 ;
        RECT 110.570 175.730 111.545 175.870 ;
        RECT 111.255 175.685 111.545 175.730 ;
        RECT 112.335 175.870 112.625 175.915 ;
        RECT 113.240 175.870 113.560 175.930 ;
        RECT 112.335 175.730 113.560 175.870 ;
        RECT 112.335 175.685 112.625 175.730 ;
        RECT 113.240 175.670 113.560 175.730 ;
        RECT 61.190 174.710 116.270 175.190 ;
        RECT 112.320 174.310 112.640 174.570 ;
        RECT 110.020 174.170 110.340 174.230 ;
        RECT 110.020 174.030 112.550 174.170 ;
        RECT 110.020 173.970 110.340 174.030 ;
        RECT 105.880 173.830 106.200 173.890 ;
        RECT 110.955 173.830 111.245 173.875 ;
        RECT 105.880 173.690 111.245 173.830 ;
        RECT 105.880 173.630 106.200 173.690 ;
        RECT 110.955 173.645 111.245 173.690 ;
        RECT 111.860 173.630 112.180 173.890 ;
        RECT 112.410 173.875 112.550 174.030 ;
        RECT 112.335 173.645 112.625 173.875 ;
        RECT 61.190 171.990 115.470 172.470 ;
        RECT 61.190 169.270 116.270 169.750 ;
        RECT 61.190 166.550 115.470 167.030 ;
        RECT 61.190 163.830 116.270 164.310 ;
        RECT 61.190 161.110 115.470 161.590 ;
        RECT 61.190 158.390 116.270 158.870 ;
        RECT 61.190 155.670 115.470 156.150 ;
        RECT 61.190 152.950 116.270 153.430 ;
        RECT 131.490 98.910 133.920 98.960 ;
        RECT 129.770 98.230 133.920 98.910 ;
        RECT 104.440 92.920 106.710 93.690 ;
        RECT 102.780 92.780 106.710 92.920 ;
        RECT 129.770 92.810 130.450 98.230 ;
        RECT 131.490 98.210 133.920 98.230 ;
        RECT 139.405 95.040 144.820 95.775 ;
        RECT 144.085 92.815 144.820 95.040 ;
        RECT 147.310 94.310 149.580 94.370 ;
        RECT 147.310 93.015 153.090 94.310 ;
        RECT 147.130 92.815 153.090 93.015 ;
        RECT 102.780 92.040 115.580 92.780 ;
        RECT 125.530 92.130 130.550 92.810 ;
        RECT 102.780 91.895 106.710 92.040 ;
        RECT 102.780 91.370 103.805 91.895 ;
        RECT 102.750 90.345 103.835 91.370 ;
        RECT 104.440 91.180 106.710 91.895 ;
        RECT 110.160 86.890 110.900 92.040 ;
        RECT 125.530 89.380 126.210 92.130 ;
        RECT 144.070 92.055 153.090 92.815 ;
        RECT 147.170 92.010 153.090 92.055 ;
        RECT 147.170 91.910 150.090 92.010 ;
        RECT 147.170 91.860 149.580 91.910 ;
        RECT 120.800 88.700 127.820 89.380 ;
        RECT 147.170 86.960 148.115 91.860 ;
        RECT 105.850 83.410 108.490 86.470 ;
        RECT 110.160 86.150 118.220 86.890 ;
        RECT 93.750 83.250 95.250 83.280 ;
        RECT 104.980 83.260 108.490 83.410 ;
        RECT 99.690 83.250 108.490 83.260 ;
        RECT 93.750 81.760 108.490 83.250 ;
        RECT 93.750 81.750 99.710 81.760 ;
        RECT 93.750 81.720 95.250 81.750 ;
        RECT 104.980 81.000 108.490 81.760 ;
        RECT 104.980 80.900 107.250 81.000 ;
        RECT 105.470 69.245 106.660 80.900 ;
        RECT 105.470 68.055 112.985 69.245 ;
        RECT 105.470 49.420 106.660 68.055 ;
        RECT 107.200 68.050 110.280 68.055 ;
        RECT 117.490 67.730 118.210 86.150 ;
        RECT 147.090 83.120 148.190 86.960 ;
        RECT 147.060 82.020 148.220 83.120 ;
        RECT 112.460 67.010 118.210 67.730 ;
        RECT 144.780 49.500 145.700 49.530 ;
        RECT 105.470 48.665 117.695 49.420 ;
        RECT 143.530 49.380 145.700 49.500 ;
        RECT 105.470 40.655 106.660 48.665 ;
        RECT 140.380 48.600 145.700 49.380 ;
        RECT 143.530 48.580 145.700 48.600 ;
        RECT 144.780 48.550 145.700 48.580 ;
        RECT 111.440 45.260 112.940 45.290 ;
        RECT 125.090 45.260 149.340 45.910 ;
        RECT 111.440 43.760 149.340 45.260 ;
        RECT 111.440 43.730 112.940 43.760 ;
        RECT 115.770 40.655 116.020 40.780 ;
        RECT 105.470 39.465 116.285 40.655 ;
        RECT 105.470 21.605 106.660 39.465 ;
        RECT 115.770 38.675 116.020 39.465 ;
        RECT 119.540 38.710 120.240 43.760 ;
        RECT 125.090 43.560 149.340 43.760 ;
        RECT 125.090 34.660 127.290 42.410 ;
        RECT 127.440 39.660 128.390 43.560 ;
        RECT 127.720 36.960 127.970 36.975 ;
        RECT 125.090 22.810 126.740 34.660 ;
        RECT 127.590 34.460 129.440 36.960 ;
        RECT 127.340 32.210 128.340 32.560 ;
        RECT 126.950 31.760 127.180 32.190 ;
        RECT 128.490 31.760 129.440 34.460 ;
        RECT 126.940 30.610 129.440 31.760 ;
        RECT 129.590 31.060 131.340 43.560 ;
        RECT 131.940 42.860 137.290 43.210 ;
        RECT 138.290 42.860 139.390 43.160 ;
        RECT 131.550 42.460 131.780 42.820 ;
        RECT 133.140 42.810 137.290 42.860 ;
        RECT 133.140 42.460 137.640 42.810 ;
        RECT 137.900 42.460 138.130 42.820 ;
        RECT 139.540 42.460 139.770 42.820 ;
        RECT 131.540 41.660 139.770 42.460 ;
        RECT 131.540 41.260 135.140 41.660 ;
        RECT 131.550 40.860 131.780 41.260 ;
        RECT 133.140 41.210 135.140 41.260 ;
        RECT 133.190 40.860 135.140 41.210 ;
        RECT 131.990 40.810 132.990 40.860 ;
        RECT 131.985 40.580 132.990 40.810 ;
        RECT 131.990 40.560 132.990 40.580 ;
        RECT 133.240 40.530 135.140 40.860 ;
        RECT 131.550 40.110 131.780 40.530 ;
        RECT 133.190 40.110 135.140 40.530 ;
        RECT 131.540 38.860 135.140 40.110 ;
        RECT 131.550 38.570 131.780 38.860 ;
        RECT 133.140 38.560 135.140 38.860 ;
        RECT 131.940 38.260 135.140 38.560 ;
        RECT 131.550 37.960 131.780 38.240 ;
        RECT 133.140 37.960 135.140 38.260 ;
        RECT 131.540 36.760 135.140 37.960 ;
        RECT 131.550 36.280 131.780 36.760 ;
        RECT 131.990 36.230 132.990 36.260 ;
        RECT 131.985 36.000 132.990 36.230 ;
        RECT 131.990 35.960 132.990 36.000 ;
        RECT 131.550 35.660 131.780 35.950 ;
        RECT 133.140 35.660 135.140 36.760 ;
        RECT 131.540 34.460 135.140 35.660 ;
        RECT 131.550 33.990 131.780 34.460 ;
        RECT 133.140 33.960 135.140 34.460 ;
        RECT 131.940 33.710 135.140 33.960 ;
        RECT 131.550 33.260 131.780 33.660 ;
        RECT 133.140 33.260 135.140 33.710 ;
        RECT 131.540 32.060 135.140 33.260 ;
        RECT 131.550 31.700 131.780 32.060 ;
        RECT 131.990 31.650 132.990 31.710 ;
        RECT 131.985 31.420 132.990 31.650 ;
        RECT 131.990 31.410 132.990 31.420 ;
        RECT 131.550 31.010 131.780 31.370 ;
        RECT 133.140 31.010 135.140 32.060 ;
        RECT 126.950 30.230 127.180 30.610 ;
        RECT 128.490 30.210 129.440 30.610 ;
        RECT 127.340 29.910 129.440 30.210 ;
        RECT 126.950 29.510 127.180 29.900 ;
        RECT 128.490 29.510 129.440 29.910 ;
        RECT 131.540 29.810 135.140 31.010 ;
        RECT 126.940 28.360 129.440 29.510 ;
        RECT 131.550 29.410 131.780 29.810 ;
        RECT 133.140 29.360 135.140 29.810 ;
        RECT 131.940 29.160 135.140 29.360 ;
        RECT 136.140 41.260 139.770 41.660 ;
        RECT 136.140 40.060 137.640 41.260 ;
        RECT 137.900 40.860 138.130 41.260 ;
        RECT 139.540 40.860 139.770 41.260 ;
        RECT 138.340 40.810 139.390 40.860 ;
        RECT 138.335 40.580 139.390 40.810 ;
        RECT 138.340 40.560 139.390 40.580 ;
        RECT 137.900 40.060 138.130 40.530 ;
        RECT 139.540 40.060 139.770 40.530 ;
        RECT 136.140 38.860 139.770 40.060 ;
        RECT 136.140 37.960 137.640 38.860 ;
        RECT 137.900 38.570 138.130 38.860 ;
        RECT 139.540 38.570 139.770 38.860 ;
        RECT 138.290 38.260 139.390 38.560 ;
        RECT 137.900 37.960 138.130 38.240 ;
        RECT 139.540 37.960 139.770 38.240 ;
        RECT 136.140 36.760 139.770 37.960 ;
        RECT 136.140 35.660 137.640 36.760 ;
        RECT 137.900 36.280 138.130 36.760 ;
        RECT 139.540 36.280 139.770 36.760 ;
        RECT 138.340 36.230 139.390 36.260 ;
        RECT 138.335 36.000 139.390 36.230 ;
        RECT 138.340 35.960 139.390 36.000 ;
        RECT 137.900 35.660 138.130 35.950 ;
        RECT 139.540 35.660 139.770 35.950 ;
        RECT 136.140 34.460 139.770 35.660 ;
        RECT 136.140 33.260 137.640 34.460 ;
        RECT 137.900 33.990 138.130 34.460 ;
        RECT 139.540 33.990 139.770 34.460 ;
        RECT 138.290 33.660 139.390 33.960 ;
        RECT 137.900 33.260 138.130 33.660 ;
        RECT 139.540 33.260 139.770 33.660 ;
        RECT 136.140 32.060 139.770 33.260 ;
        RECT 136.140 31.010 137.640 32.060 ;
        RECT 137.900 31.700 138.130 32.060 ;
        RECT 138.340 31.650 139.390 31.710 ;
        RECT 139.540 31.700 139.770 32.060 ;
        RECT 138.335 31.420 139.390 31.650 ;
        RECT 138.340 31.410 139.390 31.420 ;
        RECT 137.900 31.010 138.130 31.370 ;
        RECT 139.540 31.010 139.770 31.370 ;
        RECT 139.940 31.060 142.240 43.560 ;
        RECT 142.890 43.110 143.940 43.410 ;
        RECT 136.140 29.810 139.770 31.010 ;
        RECT 136.140 29.160 137.640 29.810 ;
        RECT 137.900 29.410 138.130 29.810 ;
        RECT 139.540 29.410 139.770 29.810 ;
        RECT 138.615 29.360 139.165 29.390 ;
        RECT 131.940 29.110 137.640 29.160 ;
        RECT 126.950 27.940 127.180 28.360 ;
        RECT 127.340 27.610 128.340 27.960 ;
        RECT 126.950 27.210 127.180 27.610 ;
        RECT 128.490 27.210 129.440 28.360 ;
        RECT 133.140 28.210 137.640 29.110 ;
        RECT 138.290 29.060 139.390 29.360 ;
        RECT 138.390 28.810 139.340 29.060 ;
        RECT 138.615 28.780 139.165 28.810 ;
        RECT 133.140 27.410 135.490 28.210 ;
        RECT 138.340 27.710 139.340 28.110 ;
        RECT 132.240 27.300 135.490 27.410 ;
        RECT 136.790 27.460 139.340 27.710 ;
        RECT 136.790 27.300 139.190 27.460 ;
        RECT 140.390 27.410 142.240 31.060 ;
        RECT 142.390 30.310 142.740 43.110 ;
        RECT 144.140 42.620 144.370 43.080 ;
        RECT 142.940 42.570 143.990 42.610 ;
        RECT 142.935 42.340 143.990 42.570 ;
        RECT 142.940 42.310 143.990 42.340 ;
        RECT 144.740 42.510 149.340 42.660 ;
        RECT 150.790 42.510 153.090 92.010 ;
        RECT 144.740 42.500 153.350 42.510 ;
        RECT 144.140 41.830 144.370 42.290 ;
        RECT 142.890 41.510 143.940 41.810 ;
        RECT 144.740 41.700 155.700 42.500 ;
        RECT 144.140 41.040 144.370 41.500 ;
        RECT 142.940 40.990 143.990 41.010 ;
        RECT 142.935 40.760 143.990 40.990 ;
        RECT 142.940 40.710 143.990 40.760 ;
        RECT 144.740 40.800 157.310 41.700 ;
        RECT 142.890 39.960 143.940 40.260 ;
        RECT 144.140 40.250 144.370 40.710 ;
        RECT 144.740 40.210 155.700 40.800 ;
        RECT 156.410 40.600 157.310 40.800 ;
        RECT 144.140 39.460 144.370 39.920 ;
        RECT 144.740 39.460 149.340 40.210 ;
        RECT 152.660 40.200 155.700 40.210 ;
        RECT 156.380 39.700 157.340 40.600 ;
        RECT 142.940 39.410 143.990 39.460 ;
        RECT 142.935 39.180 143.990 39.410 ;
        RECT 142.940 39.160 143.990 39.180 ;
        RECT 144.740 39.410 148.090 39.460 ;
        RECT 144.140 38.670 144.370 39.130 ;
        RECT 142.890 38.360 143.940 38.660 ;
        RECT 144.140 37.880 144.370 38.340 ;
        RECT 142.940 37.830 143.990 37.860 ;
        RECT 142.935 37.600 143.990 37.830 ;
        RECT 142.940 37.560 143.990 37.600 ;
        RECT 144.140 37.090 144.370 37.550 ;
        RECT 142.890 36.760 143.940 37.060 ;
        RECT 144.140 36.300 144.370 36.760 ;
        RECT 142.940 36.250 143.990 36.260 ;
        RECT 142.935 36.020 143.990 36.250 ;
        RECT 142.940 35.960 143.990 36.020 ;
        RECT 144.140 35.510 144.370 35.970 ;
        RECT 142.890 35.210 143.940 35.510 ;
        RECT 144.140 34.720 144.370 35.180 ;
        RECT 142.940 34.670 143.990 34.710 ;
        RECT 142.935 34.440 143.990 34.670 ;
        RECT 142.940 34.410 143.990 34.440 ;
        RECT 144.140 33.930 144.370 34.390 ;
        RECT 142.890 33.610 143.940 33.910 ;
        RECT 142.940 33.090 143.990 33.160 ;
        RECT 144.140 33.140 144.370 33.600 ;
        RECT 142.935 32.860 143.990 33.090 ;
        RECT 142.890 32.060 143.940 32.360 ;
        RECT 144.140 32.350 144.370 32.810 ;
        RECT 144.140 31.560 144.370 32.020 ;
        RECT 142.940 31.510 143.990 31.560 ;
        RECT 142.935 31.280 143.990 31.510 ;
        RECT 142.940 31.260 143.990 31.280 ;
        RECT 144.140 30.770 144.370 31.230 ;
        RECT 142.890 30.460 143.940 30.760 ;
        RECT 142.390 29.410 142.790 30.310 ;
        RECT 144.140 29.980 144.370 30.440 ;
        RECT 142.940 29.930 143.990 29.960 ;
        RECT 142.935 29.700 143.990 29.930 ;
        RECT 142.940 29.660 143.990 29.700 ;
        RECT 142.390 27.560 142.740 29.410 ;
        RECT 144.140 29.190 144.370 29.650 ;
        RECT 142.890 28.860 143.940 29.160 ;
        RECT 142.940 28.350 143.990 28.410 ;
        RECT 144.140 28.400 144.370 28.860 ;
        RECT 142.935 28.120 143.990 28.350 ;
        RECT 142.940 28.110 143.990 28.120 ;
        RECT 144.140 27.610 144.370 28.070 ;
        RECT 142.890 27.310 143.940 27.610 ;
        RECT 126.940 26.060 129.440 27.210 ;
        RECT 130.240 26.870 131.240 27.260 ;
        RECT 132.090 27.160 135.490 27.300 ;
        RECT 132.090 27.070 134.590 27.160 ;
        RECT 136.690 27.070 139.190 27.300 ;
        RECT 132.240 27.060 134.540 27.070 ;
        RECT 131.700 26.960 131.930 27.020 ;
        RECT 134.750 26.960 134.980 27.020 ;
        RECT 136.300 26.960 136.530 27.020 ;
        RECT 139.350 26.960 139.580 27.020 ;
        RECT 131.590 26.870 131.990 26.960 ;
        RECT 134.690 26.870 135.090 26.960 ;
        RECT 130.240 26.655 135.090 26.870 ;
        RECT 130.240 26.260 131.240 26.655 ;
        RECT 131.590 26.610 131.990 26.655 ;
        RECT 134.690 26.610 135.090 26.655 ;
        RECT 136.190 26.885 136.590 26.960 ;
        RECT 139.290 26.885 139.690 26.960 ;
        RECT 140.090 26.885 141.090 27.260 ;
        RECT 136.190 26.660 141.090 26.885 ;
        RECT 136.190 26.610 136.590 26.660 ;
        RECT 139.290 26.640 141.090 26.660 ;
        RECT 139.290 26.610 139.690 26.640 ;
        RECT 131.700 26.560 131.930 26.610 ;
        RECT 134.750 26.560 134.980 26.610 ;
        RECT 136.300 26.560 136.530 26.610 ;
        RECT 139.350 26.560 139.580 26.610 ;
        RECT 132.090 26.410 134.590 26.510 ;
        RECT 136.690 26.410 139.190 26.510 ;
        RECT 132.090 26.280 139.190 26.410 ;
        RECT 132.290 26.060 138.940 26.280 ;
        RECT 140.090 26.260 141.090 26.640 ;
        RECT 144.740 26.610 146.040 39.410 ;
        RECT 146.840 39.260 147.890 39.410 ;
        RECT 146.890 39.160 147.890 39.260 ;
        RECT 146.500 38.760 146.730 39.110 ;
        RECT 146.390 38.560 146.740 38.760 ;
        RECT 148.050 38.560 148.280 39.110 ;
        RECT 146.390 37.610 148.280 38.560 ;
        RECT 146.390 36.310 146.740 37.610 ;
        RECT 146.890 36.860 147.890 37.160 ;
        RECT 148.050 37.150 148.280 37.610 ;
        RECT 148.050 36.310 148.280 36.820 ;
        RECT 146.390 35.360 148.280 36.310 ;
        RECT 146.390 33.960 146.740 35.360 ;
        RECT 148.050 34.860 148.280 35.360 ;
        RECT 146.890 34.560 147.890 34.860 ;
        RECT 148.050 33.960 148.280 34.530 ;
        RECT 146.390 33.010 148.280 33.960 ;
        RECT 146.390 31.810 146.740 33.010 ;
        RECT 148.050 32.570 148.280 33.010 ;
        RECT 146.890 32.260 147.890 32.560 ;
        RECT 148.050 31.810 148.280 32.240 ;
        RECT 146.390 30.860 148.280 31.810 ;
        RECT 146.390 29.510 146.740 30.860 ;
        RECT 146.890 29.960 147.890 30.310 ;
        RECT 148.050 30.280 148.280 30.860 ;
        RECT 148.050 29.510 148.280 29.950 ;
        RECT 146.390 28.560 148.280 29.510 ;
        RECT 146.390 27.260 146.740 28.560 ;
        RECT 146.890 27.660 147.890 28.010 ;
        RECT 148.050 27.990 148.280 28.560 ;
        RECT 148.050 27.260 148.280 27.660 ;
        RECT 146.390 26.310 148.280 27.260 ;
        RECT 126.950 25.650 127.180 26.060 ;
        RECT 128.490 25.810 129.440 26.060 ;
        RECT 128.490 25.660 129.820 25.810 ;
        RECT 131.140 25.660 132.140 25.960 ;
        RECT 127.340 25.360 129.820 25.660 ;
        RECT 126.950 24.960 127.180 25.320 ;
        RECT 128.490 25.160 129.820 25.360 ;
        RECT 128.490 24.960 129.440 25.160 ;
        RECT 133.140 25.110 138.390 26.060 ;
        RECT 139.290 25.660 140.290 25.960 ;
        RECT 144.245 25.930 145.135 25.960 ;
        RECT 146.390 25.930 146.740 26.310 ;
        RECT 144.245 25.040 146.740 25.930 ;
        RECT 148.050 25.700 148.280 26.310 ;
        RECT 146.990 25.650 147.890 25.660 ;
        RECT 146.890 25.420 147.890 25.650 ;
        RECT 146.990 25.360 147.890 25.420 ;
        RECT 144.245 25.010 145.135 25.040 ;
        RECT 126.940 23.810 129.440 24.960 ;
        RECT 146.390 24.910 146.740 25.040 ;
        RECT 148.050 24.910 148.280 25.370 ;
        RECT 131.340 24.620 133.300 24.850 ;
        RECT 133.630 24.620 135.590 24.850 ;
        RECT 135.920 24.620 137.880 24.850 ;
        RECT 138.210 24.620 140.170 24.850 ;
        RECT 131.060 24.410 131.290 24.460 ;
        RECT 126.950 23.360 127.180 23.810 ;
        RECT 128.490 23.360 129.440 23.810 ;
        RECT 130.940 23.510 131.340 24.410 ;
        RECT 131.060 23.460 131.290 23.510 ;
        RECT 128.540 23.310 129.440 23.360 ;
        RECT 131.790 23.310 132.690 24.620 ;
        RECT 133.350 24.310 133.580 24.460 ;
        RECT 133.240 23.610 133.690 24.310 ;
        RECT 133.350 23.460 133.580 23.610 ;
        RECT 134.190 23.310 135.090 24.620 ;
        RECT 135.640 24.310 135.870 24.460 ;
        RECT 135.540 23.610 135.990 24.310 ;
        RECT 135.640 23.460 135.870 23.610 ;
        RECT 136.490 23.310 137.390 24.620 ;
        RECT 137.930 24.310 138.160 24.460 ;
        RECT 137.840 23.610 138.290 24.310 ;
        RECT 137.930 23.460 138.160 23.610 ;
        RECT 138.740 23.310 139.640 24.620 ;
        RECT 140.220 24.410 140.450 24.460 ;
        RECT 140.140 23.510 140.540 24.410 ;
        RECT 140.220 23.460 140.450 23.510 ;
        RECT 127.340 22.960 128.340 23.310 ;
        RECT 128.540 23.300 140.140 23.310 ;
        RECT 128.540 23.070 140.170 23.300 ;
        RECT 128.540 23.010 140.140 23.070 ;
        RECT 140.740 22.810 142.090 24.860 ;
        RECT 144.540 22.810 146.240 24.310 ;
        RECT 146.390 23.960 148.340 24.910 ;
        RECT 148.590 24.310 149.340 37.260 ;
        RECT 146.390 23.460 146.740 23.960 ;
        RECT 146.500 23.410 146.730 23.460 ;
        RECT 148.050 23.410 148.280 23.960 ;
        RECT 146.890 23.060 147.890 23.410 ;
        RECT 148.490 22.810 149.340 24.310 ;
        RECT 125.140 21.605 149.340 22.810 ;
        RECT 105.470 20.460 149.340 21.605 ;
        RECT 105.470 20.415 118.640 20.460 ;
        RECT 122.640 20.415 130.285 20.460 ;
        RECT 115.540 20.410 116.290 20.415 ;
        RECT 115.770 18.310 116.020 18.625 ;
        RECT 119.820 18.310 120.070 18.825 ;
        RECT 115.540 17.110 120.340 18.310 ;
        RECT 115.770 16.520 116.020 17.110 ;
        RECT 117.340 14.860 118.540 17.110 ;
        RECT 119.820 16.720 120.070 17.110 ;
        RECT 150.940 14.860 152.140 14.890 ;
        RECT 117.340 13.660 152.140 14.860 ;
        RECT 150.940 13.630 152.140 13.660 ;
      LAYER via ;
        RECT 78.310 208.650 78.570 208.910 ;
        RECT 97.630 208.650 97.890 208.910 ;
        RECT 106.370 208.650 106.630 208.910 ;
        RECT 91.650 208.310 91.910 208.570 ;
        RECT 98.550 208.310 98.810 208.570 ;
        RECT 99.930 208.310 100.190 208.570 ;
        RECT 100.850 208.310 101.110 208.570 ;
        RECT 72.790 207.970 73.050 208.230 ;
        RECT 75.090 207.970 75.350 208.230 ;
        RECT 87.970 207.970 88.230 208.230 ;
        RECT 89.350 207.970 89.610 208.230 ;
        RECT 94.410 207.970 94.670 208.230 ;
        RECT 105.910 207.970 106.170 208.230 ;
        RECT 73.990 207.460 74.250 207.720 ;
        RECT 74.310 207.460 74.570 207.720 ;
        RECT 74.630 207.460 74.890 207.720 ;
        RECT 74.950 207.460 75.210 207.720 ;
        RECT 75.270 207.460 75.530 207.720 ;
        RECT 87.560 207.460 87.820 207.720 ;
        RECT 87.880 207.460 88.140 207.720 ;
        RECT 88.200 207.460 88.460 207.720 ;
        RECT 88.520 207.460 88.780 207.720 ;
        RECT 88.840 207.460 89.100 207.720 ;
        RECT 101.130 207.460 101.390 207.720 ;
        RECT 101.450 207.460 101.710 207.720 ;
        RECT 101.770 207.460 102.030 207.720 ;
        RECT 102.090 207.460 102.350 207.720 ;
        RECT 102.410 207.460 102.670 207.720 ;
        RECT 114.700 207.460 114.960 207.720 ;
        RECT 115.020 207.460 115.280 207.720 ;
        RECT 115.340 207.460 115.600 207.720 ;
        RECT 115.660 207.460 115.920 207.720 ;
        RECT 115.980 207.460 116.240 207.720 ;
        RECT 81.530 206.950 81.790 207.210 ;
        RECT 89.350 206.950 89.610 207.210 ;
        RECT 99.930 206.950 100.190 207.210 ;
        RECT 71.870 206.610 72.130 206.870 ;
        RECT 78.310 206.610 78.570 206.870 ;
        RECT 73.710 206.270 73.970 206.530 ;
        RECT 84.290 206.270 84.550 206.530 ;
        RECT 76.470 205.930 76.730 206.190 ;
        RECT 77.390 205.930 77.650 206.190 ;
        RECT 91.650 206.270 91.910 206.530 ;
        RECT 96.710 206.610 96.970 206.870 ;
        RECT 93.950 206.270 94.210 206.530 ;
        RECT 96.250 206.270 96.510 206.530 ;
        RECT 97.630 206.270 97.890 206.530 ;
        RECT 98.550 206.270 98.810 206.530 ;
        RECT 113.730 206.610 113.990 206.870 ;
        RECT 103.150 206.270 103.410 206.530 ;
        RECT 93.030 205.930 93.290 206.190 ;
        RECT 93.490 205.930 93.750 206.190 ;
        RECT 94.410 205.930 94.670 206.190 ;
        RECT 99.010 205.930 99.270 206.190 ;
        RECT 86.130 205.590 86.390 205.850 ;
        RECT 94.870 205.590 95.130 205.850 ;
        RECT 96.710 205.590 96.970 205.850 ;
        RECT 98.090 205.590 98.350 205.850 ;
        RECT 73.250 205.250 73.510 205.510 ;
        RECT 76.930 205.250 77.190 205.510 ;
        RECT 83.370 205.250 83.630 205.510 ;
        RECT 92.110 205.250 92.370 205.510 ;
        RECT 96.250 205.250 96.510 205.510 ;
        RECT 97.170 205.250 97.430 205.510 ;
        RECT 112.350 205.930 112.610 206.190 ;
        RECT 109.590 205.250 109.850 205.510 ;
        RECT 67.205 204.740 67.465 205.000 ;
        RECT 67.525 204.740 67.785 205.000 ;
        RECT 67.845 204.740 68.105 205.000 ;
        RECT 68.165 204.740 68.425 205.000 ;
        RECT 68.485 204.740 68.745 205.000 ;
        RECT 80.775 204.740 81.035 205.000 ;
        RECT 81.095 204.740 81.355 205.000 ;
        RECT 81.415 204.740 81.675 205.000 ;
        RECT 81.735 204.740 81.995 205.000 ;
        RECT 82.055 204.740 82.315 205.000 ;
        RECT 94.345 204.740 94.605 205.000 ;
        RECT 94.665 204.740 94.925 205.000 ;
        RECT 94.985 204.740 95.245 205.000 ;
        RECT 95.305 204.740 95.565 205.000 ;
        RECT 95.625 204.740 95.885 205.000 ;
        RECT 107.915 204.740 108.175 205.000 ;
        RECT 108.235 204.740 108.495 205.000 ;
        RECT 108.555 204.740 108.815 205.000 ;
        RECT 108.875 204.740 109.135 205.000 ;
        RECT 109.195 204.740 109.455 205.000 ;
        RECT 62.210 204.230 62.470 204.490 ;
        RECT 69.110 204.230 69.370 204.490 ;
        RECT 72.790 204.230 73.050 204.490 ;
        RECT 73.710 204.230 73.970 204.490 ;
        RECT 92.110 204.230 92.370 204.490 ;
        RECT 63.590 203.890 63.850 204.150 ;
        RECT 77.390 203.890 77.650 204.150 ;
        RECT 78.770 203.890 79.030 204.150 ;
        RECT 93.030 203.890 93.290 204.150 ;
        RECT 64.970 203.210 65.230 203.470 ;
        RECT 66.810 203.210 67.070 203.470 ;
        RECT 73.710 203.210 73.970 203.470 ;
        RECT 74.630 203.210 74.890 203.470 ;
        RECT 76.470 203.210 76.730 203.470 ;
        RECT 76.930 203.210 77.190 203.470 ;
        RECT 78.310 203.210 78.570 203.470 ;
        RECT 79.230 203.210 79.490 203.470 ;
        RECT 99.930 204.230 100.190 204.490 ;
        RECT 99.470 203.890 99.730 204.150 ;
        RECT 64.510 202.870 64.770 203.130 ;
        RECT 71.410 202.530 71.670 202.790 ;
        RECT 82.450 202.870 82.710 203.130 ;
        RECT 95.790 203.210 96.050 203.470 ;
        RECT 97.170 203.210 97.430 203.470 ;
        RECT 98.550 203.550 98.810 203.810 ;
        RECT 112.350 203.550 112.610 203.810 ;
        RECT 85.210 202.870 85.470 203.130 ;
        RECT 87.050 202.870 87.310 203.130 ;
        RECT 113.730 203.210 113.990 203.470 ;
        RECT 92.110 202.530 92.370 202.790 ;
        RECT 93.950 202.530 94.210 202.790 ;
        RECT 98.090 202.530 98.350 202.790 ;
        RECT 104.990 202.530 105.250 202.790 ;
        RECT 73.990 202.020 74.250 202.280 ;
        RECT 74.310 202.020 74.570 202.280 ;
        RECT 74.630 202.020 74.890 202.280 ;
        RECT 74.950 202.020 75.210 202.280 ;
        RECT 75.270 202.020 75.530 202.280 ;
        RECT 87.560 202.020 87.820 202.280 ;
        RECT 87.880 202.020 88.140 202.280 ;
        RECT 88.200 202.020 88.460 202.280 ;
        RECT 88.520 202.020 88.780 202.280 ;
        RECT 88.840 202.020 89.100 202.280 ;
        RECT 101.130 202.020 101.390 202.280 ;
        RECT 101.450 202.020 101.710 202.280 ;
        RECT 101.770 202.020 102.030 202.280 ;
        RECT 102.090 202.020 102.350 202.280 ;
        RECT 102.410 202.020 102.670 202.280 ;
        RECT 114.700 202.020 114.960 202.280 ;
        RECT 115.020 202.020 115.280 202.280 ;
        RECT 115.340 202.020 115.600 202.280 ;
        RECT 115.660 202.020 115.920 202.280 ;
        RECT 115.980 202.020 116.240 202.280 ;
        RECT 64.050 201.170 64.310 201.430 ;
        RECT 63.590 200.830 63.850 201.090 ;
        RECT 64.510 200.830 64.770 201.090 ;
        RECT 71.870 201.510 72.130 201.770 ;
        RECT 72.790 201.170 73.050 201.430 ;
        RECT 70.490 200.830 70.750 201.090 ;
        RECT 72.330 200.830 72.590 201.090 ;
        RECT 76.010 201.510 76.270 201.770 ;
        RECT 76.930 201.510 77.190 201.770 ;
        RECT 83.370 201.170 83.630 201.430 ;
        RECT 75.550 200.830 75.810 201.090 ;
        RECT 79.230 200.830 79.490 201.090 ;
        RECT 85.210 201.510 85.470 201.770 ;
        RECT 73.710 200.490 73.970 200.750 ;
        RECT 82.450 200.490 82.710 200.750 ;
        RECT 86.130 200.830 86.390 201.090 ;
        RECT 92.110 201.170 92.370 201.430 ;
        RECT 96.250 201.510 96.510 201.770 ;
        RECT 99.010 201.510 99.270 201.770 ;
        RECT 105.910 201.510 106.170 201.770 ;
        RECT 106.370 201.510 106.630 201.770 ;
        RECT 93.490 200.830 93.750 201.090 ;
        RECT 106.830 201.170 107.090 201.430 ;
        RECT 96.710 200.830 96.970 201.090 ;
        RECT 97.630 200.830 97.890 201.090 ;
        RECT 99.470 200.830 99.730 201.090 ;
        RECT 66.810 200.150 67.070 200.410 ;
        RECT 93.950 200.150 94.210 200.410 ;
        RECT 99.930 200.150 100.190 200.410 ;
        RECT 110.970 200.490 111.230 200.750 ;
        RECT 64.510 199.810 64.770 200.070 ;
        RECT 66.350 199.810 66.610 200.070 ;
        RECT 76.470 199.810 76.730 200.070 ;
        RECT 77.850 199.810 78.110 200.070 ;
        RECT 87.510 199.810 87.770 200.070 ;
        RECT 93.490 199.810 93.750 200.070 ;
        RECT 97.170 199.810 97.430 200.070 ;
        RECT 98.550 199.810 98.810 200.070 ;
        RECT 107.290 199.810 107.550 200.070 ;
        RECT 67.205 199.300 67.465 199.560 ;
        RECT 67.525 199.300 67.785 199.560 ;
        RECT 67.845 199.300 68.105 199.560 ;
        RECT 68.165 199.300 68.425 199.560 ;
        RECT 68.485 199.300 68.745 199.560 ;
        RECT 80.775 199.300 81.035 199.560 ;
        RECT 81.095 199.300 81.355 199.560 ;
        RECT 81.415 199.300 81.675 199.560 ;
        RECT 81.735 199.300 81.995 199.560 ;
        RECT 82.055 199.300 82.315 199.560 ;
        RECT 94.345 199.300 94.605 199.560 ;
        RECT 94.665 199.300 94.925 199.560 ;
        RECT 94.985 199.300 95.245 199.560 ;
        RECT 95.305 199.300 95.565 199.560 ;
        RECT 95.625 199.300 95.885 199.560 ;
        RECT 107.915 199.300 108.175 199.560 ;
        RECT 108.235 199.300 108.495 199.560 ;
        RECT 108.555 199.300 108.815 199.560 ;
        RECT 108.875 199.300 109.135 199.560 ;
        RECT 109.195 199.300 109.455 199.560 ;
        RECT 64.970 198.790 65.230 199.050 ;
        RECT 64.050 198.450 64.310 198.710 ;
        RECT 73.710 198.450 73.970 198.710 ;
        RECT 82.910 198.450 83.170 198.710 ;
        RECT 85.670 198.450 85.930 198.710 ;
        RECT 93.490 198.790 93.750 199.050 ;
        RECT 99.470 198.790 99.730 199.050 ;
        RECT 103.150 198.790 103.410 199.050 ;
        RECT 94.870 198.450 95.130 198.710 ;
        RECT 66.350 197.770 66.610 198.030 ;
        RECT 73.710 197.770 73.970 198.030 ;
        RECT 76.010 197.770 76.270 198.030 ;
        RECT 82.450 198.110 82.710 198.370 ;
        RECT 97.170 198.110 97.430 198.370 ;
        RECT 85.670 197.770 85.930 198.030 ;
        RECT 99.930 198.450 100.190 198.710 ;
        RECT 111.430 198.450 111.690 198.710 ;
        RECT 75.090 197.430 75.350 197.690 ;
        RECT 82.910 197.430 83.170 197.690 ;
        RECT 84.750 197.430 85.010 197.690 ;
        RECT 87.970 197.430 88.230 197.690 ;
        RECT 71.410 197.090 71.670 197.350 ;
        RECT 78.770 197.090 79.030 197.350 ;
        RECT 93.950 197.090 94.210 197.350 ;
        RECT 94.870 197.090 95.130 197.350 ;
        RECT 96.250 197.430 96.510 197.690 ;
        RECT 99.010 197.430 99.270 197.690 ;
        RECT 97.170 197.090 97.430 197.350 ;
        RECT 98.550 197.090 98.810 197.350 ;
        RECT 101.770 197.770 102.030 198.030 ;
        RECT 106.830 197.770 107.090 198.030 ;
        RECT 110.050 197.770 110.310 198.030 ;
        RECT 103.610 197.430 103.870 197.690 ;
        RECT 109.590 197.090 109.850 197.350 ;
        RECT 110.510 197.090 110.770 197.350 ;
        RECT 73.990 196.580 74.250 196.840 ;
        RECT 74.310 196.580 74.570 196.840 ;
        RECT 74.630 196.580 74.890 196.840 ;
        RECT 74.950 196.580 75.210 196.840 ;
        RECT 75.270 196.580 75.530 196.840 ;
        RECT 87.560 196.580 87.820 196.840 ;
        RECT 87.880 196.580 88.140 196.840 ;
        RECT 88.200 196.580 88.460 196.840 ;
        RECT 88.520 196.580 88.780 196.840 ;
        RECT 88.840 196.580 89.100 196.840 ;
        RECT 101.130 196.580 101.390 196.840 ;
        RECT 101.450 196.580 101.710 196.840 ;
        RECT 101.770 196.580 102.030 196.840 ;
        RECT 102.090 196.580 102.350 196.840 ;
        RECT 102.410 196.580 102.670 196.840 ;
        RECT 114.700 196.580 114.960 196.840 ;
        RECT 115.020 196.580 115.280 196.840 ;
        RECT 115.340 196.580 115.600 196.840 ;
        RECT 115.660 196.580 115.920 196.840 ;
        RECT 115.980 196.580 116.240 196.840 ;
        RECT 70.490 196.070 70.750 196.330 ;
        RECT 72.790 196.070 73.050 196.330 ;
        RECT 77.390 196.070 77.650 196.330 ;
        RECT 87.050 196.070 87.310 196.330 ;
        RECT 78.310 195.730 78.570 195.990 ;
        RECT 103.610 196.070 103.870 196.330 ;
        RECT 110.050 195.730 110.310 195.990 ;
        RECT 113.730 195.730 113.990 195.990 ;
        RECT 79.230 195.390 79.490 195.650 ;
        RECT 90.270 195.390 90.530 195.650 ;
        RECT 97.630 195.390 97.890 195.650 ;
        RECT 71.410 194.710 71.670 194.970 ;
        RECT 76.930 195.050 77.190 195.310 ;
        RECT 85.670 195.050 85.930 195.310 ;
        RECT 98.090 195.050 98.350 195.310 ;
        RECT 110.510 195.390 110.770 195.650 ;
        RECT 107.290 195.050 107.550 195.310 ;
        RECT 109.590 195.050 109.850 195.310 ;
        RECT 112.350 195.050 112.610 195.310 ;
        RECT 75.090 194.370 75.350 194.630 ;
        RECT 78.770 194.370 79.030 194.630 ;
        RECT 96.710 194.370 96.970 194.630 ;
        RECT 99.010 194.370 99.270 194.630 ;
        RECT 99.930 194.370 100.190 194.630 ;
        RECT 110.510 194.370 110.770 194.630 ;
        RECT 67.205 193.860 67.465 194.120 ;
        RECT 67.525 193.860 67.785 194.120 ;
        RECT 67.845 193.860 68.105 194.120 ;
        RECT 68.165 193.860 68.425 194.120 ;
        RECT 68.485 193.860 68.745 194.120 ;
        RECT 80.775 193.860 81.035 194.120 ;
        RECT 81.095 193.860 81.355 194.120 ;
        RECT 81.415 193.860 81.675 194.120 ;
        RECT 81.735 193.860 81.995 194.120 ;
        RECT 82.055 193.860 82.315 194.120 ;
        RECT 94.345 193.860 94.605 194.120 ;
        RECT 94.665 193.860 94.925 194.120 ;
        RECT 94.985 193.860 95.245 194.120 ;
        RECT 95.305 193.860 95.565 194.120 ;
        RECT 95.625 193.860 95.885 194.120 ;
        RECT 107.915 193.860 108.175 194.120 ;
        RECT 108.235 193.860 108.495 194.120 ;
        RECT 108.555 193.860 108.815 194.120 ;
        RECT 108.875 193.860 109.135 194.120 ;
        RECT 109.195 193.860 109.455 194.120 ;
        RECT 72.330 193.350 72.590 193.610 ;
        RECT 73.250 192.330 73.510 192.590 ;
        RECT 93.490 193.350 93.750 193.610 ;
        RECT 76.010 193.010 76.270 193.270 ;
        RECT 78.770 193.010 79.030 193.270 ;
        RECT 84.290 193.010 84.550 193.270 ;
        RECT 97.170 193.350 97.430 193.610 ;
        RECT 73.250 191.650 73.510 191.910 ;
        RECT 76.470 192.330 76.730 192.590 ;
        RECT 81.990 192.670 82.250 192.930 ;
        RECT 75.090 191.990 75.350 192.250 ;
        RECT 78.310 192.330 78.570 192.590 ;
        RECT 79.230 191.990 79.490 192.250 ;
        RECT 82.450 191.990 82.710 192.250 ;
        RECT 87.050 192.330 87.310 192.590 ;
        RECT 93.950 192.670 94.210 192.930 ;
        RECT 89.810 192.330 90.070 192.590 ;
        RECT 90.730 192.330 90.990 192.590 ;
        RECT 83.370 191.990 83.630 192.250 ;
        RECT 83.830 191.990 84.090 192.250 ;
        RECT 91.650 191.990 91.910 192.250 ;
        RECT 92.570 192.330 92.830 192.590 ;
        RECT 93.030 192.330 93.290 192.590 ;
        RECT 94.410 192.330 94.670 192.590 ;
        RECT 95.790 192.330 96.050 192.590 ;
        RECT 97.170 192.330 97.430 192.590 ;
        RECT 98.090 192.330 98.350 192.590 ;
        RECT 99.470 192.330 99.730 192.590 ;
        RECT 100.390 191.990 100.650 192.250 ;
        RECT 77.390 191.650 77.650 191.910 ;
        RECT 84.290 191.650 84.550 191.910 ;
        RECT 84.750 191.650 85.010 191.910 ;
        RECT 89.350 191.650 89.610 191.910 ;
        RECT 92.570 191.650 92.830 191.910 ;
        RECT 102.690 192.330 102.950 192.590 ;
        RECT 106.830 192.330 107.090 192.590 ;
        RECT 110.050 192.330 110.310 192.590 ;
        RECT 113.270 192.330 113.530 192.590 ;
        RECT 103.610 191.990 103.870 192.250 ;
        RECT 105.910 191.990 106.170 192.250 ;
        RECT 104.990 191.650 105.250 191.910 ;
        RECT 113.270 191.650 113.530 191.910 ;
        RECT 73.990 191.140 74.250 191.400 ;
        RECT 74.310 191.140 74.570 191.400 ;
        RECT 74.630 191.140 74.890 191.400 ;
        RECT 74.950 191.140 75.210 191.400 ;
        RECT 75.270 191.140 75.530 191.400 ;
        RECT 87.560 191.140 87.820 191.400 ;
        RECT 87.880 191.140 88.140 191.400 ;
        RECT 88.200 191.140 88.460 191.400 ;
        RECT 88.520 191.140 88.780 191.400 ;
        RECT 88.840 191.140 89.100 191.400 ;
        RECT 101.130 191.140 101.390 191.400 ;
        RECT 101.450 191.140 101.710 191.400 ;
        RECT 101.770 191.140 102.030 191.400 ;
        RECT 102.090 191.140 102.350 191.400 ;
        RECT 102.410 191.140 102.670 191.400 ;
        RECT 114.700 191.140 114.960 191.400 ;
        RECT 115.020 191.140 115.280 191.400 ;
        RECT 115.340 191.140 115.600 191.400 ;
        RECT 115.660 191.140 115.920 191.400 ;
        RECT 115.980 191.140 116.240 191.400 ;
        RECT 81.990 190.630 82.250 190.890 ;
        RECT 90.730 190.630 90.990 190.890 ;
        RECT 93.030 190.630 93.290 190.890 ;
        RECT 96.250 190.630 96.510 190.890 ;
        RECT 99.010 190.630 99.270 190.890 ;
        RECT 103.150 190.630 103.410 190.890 ;
        RECT 110.970 190.630 111.230 190.890 ;
        RECT 111.430 190.630 111.690 190.890 ;
        RECT 72.330 189.950 72.590 190.210 ;
        RECT 73.250 189.950 73.510 190.210 ;
        RECT 76.930 190.290 77.190 190.550 ;
        RECT 96.710 190.290 96.970 190.550 ;
        RECT 98.550 190.290 98.810 190.550 ;
        RECT 75.550 189.950 75.810 190.210 ;
        RECT 84.750 189.950 85.010 190.210 ;
        RECT 96.250 189.950 96.510 190.210 ;
        RECT 85.670 189.610 85.930 189.870 ;
        RECT 94.410 189.610 94.670 189.870 ;
        RECT 95.790 189.610 96.050 189.870 ;
        RECT 99.470 189.610 99.730 189.870 ;
        RECT 103.150 189.950 103.410 190.210 ;
        RECT 105.450 189.950 105.710 190.210 ;
        RECT 110.510 190.290 110.770 190.550 ;
        RECT 104.070 189.610 104.330 189.870 ;
        RECT 107.290 189.610 107.550 189.870 ;
        RECT 97.170 189.270 97.430 189.530 ;
        RECT 114.190 189.610 114.450 189.870 ;
        RECT 71.410 188.930 71.670 189.190 ;
        RECT 73.250 188.930 73.510 189.190 ;
        RECT 75.090 188.930 75.350 189.190 ;
        RECT 83.370 188.930 83.630 189.190 ;
        RECT 85.210 188.930 85.470 189.190 ;
        RECT 86.130 188.930 86.390 189.190 ;
        RECT 90.270 188.930 90.530 189.190 ;
        RECT 113.270 189.270 113.530 189.530 ;
        RECT 104.530 188.930 104.790 189.190 ;
        RECT 106.370 188.930 106.630 189.190 ;
        RECT 67.205 188.420 67.465 188.680 ;
        RECT 67.525 188.420 67.785 188.680 ;
        RECT 67.845 188.420 68.105 188.680 ;
        RECT 68.165 188.420 68.425 188.680 ;
        RECT 68.485 188.420 68.745 188.680 ;
        RECT 80.775 188.420 81.035 188.680 ;
        RECT 81.095 188.420 81.355 188.680 ;
        RECT 81.415 188.420 81.675 188.680 ;
        RECT 81.735 188.420 81.995 188.680 ;
        RECT 82.055 188.420 82.315 188.680 ;
        RECT 94.345 188.420 94.605 188.680 ;
        RECT 94.665 188.420 94.925 188.680 ;
        RECT 94.985 188.420 95.245 188.680 ;
        RECT 95.305 188.420 95.565 188.680 ;
        RECT 95.625 188.420 95.885 188.680 ;
        RECT 107.915 188.420 108.175 188.680 ;
        RECT 108.235 188.420 108.495 188.680 ;
        RECT 108.555 188.420 108.815 188.680 ;
        RECT 108.875 188.420 109.135 188.680 ;
        RECT 109.195 188.420 109.455 188.680 ;
        RECT 73.250 187.910 73.510 188.170 ;
        RECT 71.410 187.230 71.670 187.490 ;
        RECT 76.010 187.910 76.270 188.170 ;
        RECT 84.290 187.910 84.550 188.170 ;
        RECT 85.670 187.910 85.930 188.170 ;
        RECT 93.950 187.910 94.210 188.170 ;
        RECT 98.090 187.910 98.350 188.170 ;
        RECT 99.470 187.910 99.730 188.170 ;
        RECT 104.990 187.910 105.250 188.170 ;
        RECT 104.530 187.230 104.790 187.490 ;
        RECT 112.350 187.230 112.610 187.490 ;
        RECT 76.930 186.890 77.190 187.150 ;
        RECT 77.390 186.890 77.650 187.150 ;
        RECT 84.290 186.890 84.550 187.150 ;
        RECT 84.750 186.890 85.010 187.150 ;
        RECT 86.130 186.890 86.390 187.150 ;
        RECT 86.590 186.890 86.850 187.150 ;
        RECT 89.350 186.890 89.610 187.150 ;
        RECT 93.950 186.890 94.210 187.150 ;
        RECT 97.170 186.890 97.430 187.150 ;
        RECT 103.150 186.890 103.410 187.150 ;
        RECT 70.950 186.550 71.210 186.810 ;
        RECT 73.250 186.550 73.510 186.810 ;
        RECT 75.090 186.550 75.350 186.810 ;
        RECT 76.470 186.210 76.730 186.470 ;
        RECT 92.110 186.550 92.370 186.810 ;
        RECT 98.090 186.550 98.350 186.810 ;
        RECT 99.470 186.550 99.730 186.810 ;
        RECT 110.970 186.890 111.230 187.150 ;
        RECT 85.210 186.210 85.470 186.470 ;
        RECT 99.010 186.210 99.270 186.470 ;
        RECT 104.530 186.210 104.790 186.470 ;
        RECT 107.290 186.210 107.550 186.470 ;
        RECT 111.890 186.210 112.150 186.470 ;
        RECT 73.990 185.700 74.250 185.960 ;
        RECT 74.310 185.700 74.570 185.960 ;
        RECT 74.630 185.700 74.890 185.960 ;
        RECT 74.950 185.700 75.210 185.960 ;
        RECT 75.270 185.700 75.530 185.960 ;
        RECT 87.560 185.700 87.820 185.960 ;
        RECT 87.880 185.700 88.140 185.960 ;
        RECT 88.200 185.700 88.460 185.960 ;
        RECT 88.520 185.700 88.780 185.960 ;
        RECT 88.840 185.700 89.100 185.960 ;
        RECT 101.130 185.700 101.390 185.960 ;
        RECT 101.450 185.700 101.710 185.960 ;
        RECT 101.770 185.700 102.030 185.960 ;
        RECT 102.090 185.700 102.350 185.960 ;
        RECT 102.410 185.700 102.670 185.960 ;
        RECT 114.700 185.700 114.960 185.960 ;
        RECT 115.020 185.700 115.280 185.960 ;
        RECT 115.340 185.700 115.600 185.960 ;
        RECT 115.660 185.700 115.920 185.960 ;
        RECT 115.980 185.700 116.240 185.960 ;
        RECT 76.010 185.190 76.270 185.450 ;
        RECT 104.070 185.190 104.330 185.450 ;
        RECT 112.350 185.190 112.610 185.450 ;
        RECT 70.950 184.510 71.210 184.770 ;
        RECT 86.590 184.850 86.850 185.110 ;
        RECT 76.930 184.170 77.190 184.430 ;
        RECT 78.310 184.510 78.570 184.770 ;
        RECT 79.690 184.510 79.950 184.770 ;
        RECT 87.050 184.510 87.310 184.770 ;
        RECT 88.890 184.510 89.150 184.770 ;
        RECT 93.950 184.850 94.210 185.110 ;
        RECT 91.650 184.510 91.910 184.770 ;
        RECT 100.390 184.510 100.650 184.770 ;
        RECT 106.370 184.510 106.630 184.770 ;
        RECT 83.830 183.830 84.090 184.090 ;
        RECT 89.810 183.830 90.070 184.090 ;
        RECT 85.210 183.490 85.470 183.750 ;
        RECT 97.170 183.490 97.430 183.750 ;
        RECT 106.830 183.490 107.090 183.750 ;
        RECT 67.205 182.980 67.465 183.240 ;
        RECT 67.525 182.980 67.785 183.240 ;
        RECT 67.845 182.980 68.105 183.240 ;
        RECT 68.165 182.980 68.425 183.240 ;
        RECT 68.485 182.980 68.745 183.240 ;
        RECT 80.775 182.980 81.035 183.240 ;
        RECT 81.095 182.980 81.355 183.240 ;
        RECT 81.415 182.980 81.675 183.240 ;
        RECT 81.735 182.980 81.995 183.240 ;
        RECT 82.055 182.980 82.315 183.240 ;
        RECT 94.345 182.980 94.605 183.240 ;
        RECT 94.665 182.980 94.925 183.240 ;
        RECT 94.985 182.980 95.245 183.240 ;
        RECT 95.305 182.980 95.565 183.240 ;
        RECT 95.625 182.980 95.885 183.240 ;
        RECT 107.915 182.980 108.175 183.240 ;
        RECT 108.235 182.980 108.495 183.240 ;
        RECT 108.555 182.980 108.815 183.240 ;
        RECT 108.875 182.980 109.135 183.240 ;
        RECT 109.195 182.980 109.455 183.240 ;
        RECT 72.330 182.470 72.590 182.730 ;
        RECT 78.310 182.470 78.570 182.730 ;
        RECT 88.890 182.470 89.150 182.730 ;
        RECT 76.470 182.130 76.730 182.390 ;
        RECT 99.010 182.470 99.270 182.730 ;
        RECT 103.610 182.470 103.870 182.730 ;
        RECT 107.750 182.470 108.010 182.730 ;
        RECT 109.590 182.470 109.850 182.730 ;
        RECT 76.010 181.450 76.270 181.710 ;
        RECT 85.210 181.790 85.470 182.050 ;
        RECT 86.590 181.790 86.850 182.050 ;
        RECT 99.470 182.130 99.730 182.390 ;
        RECT 100.390 182.130 100.650 182.390 ;
        RECT 96.250 181.790 96.510 182.050 ;
        RECT 105.910 181.790 106.170 182.050 ;
        RECT 83.830 181.450 84.090 181.710 ;
        RECT 92.570 181.450 92.830 181.710 ;
        RECT 102.690 181.450 102.950 181.710 ;
        RECT 104.070 181.450 104.330 181.710 ;
        RECT 79.230 181.110 79.490 181.370 ;
        RECT 106.830 181.450 107.090 181.710 ;
        RECT 110.050 181.110 110.310 181.370 ;
        RECT 112.350 181.110 112.610 181.370 ;
        RECT 73.250 180.770 73.510 181.030 ;
        RECT 98.090 180.770 98.350 181.030 ;
        RECT 105.910 180.770 106.170 181.030 ;
        RECT 73.990 180.260 74.250 180.520 ;
        RECT 74.310 180.260 74.570 180.520 ;
        RECT 74.630 180.260 74.890 180.520 ;
        RECT 74.950 180.260 75.210 180.520 ;
        RECT 75.270 180.260 75.530 180.520 ;
        RECT 87.560 180.260 87.820 180.520 ;
        RECT 87.880 180.260 88.140 180.520 ;
        RECT 88.200 180.260 88.460 180.520 ;
        RECT 88.520 180.260 88.780 180.520 ;
        RECT 88.840 180.260 89.100 180.520 ;
        RECT 101.130 180.260 101.390 180.520 ;
        RECT 101.450 180.260 101.710 180.520 ;
        RECT 101.770 180.260 102.030 180.520 ;
        RECT 102.090 180.260 102.350 180.520 ;
        RECT 102.410 180.260 102.670 180.520 ;
        RECT 114.700 180.260 114.960 180.520 ;
        RECT 115.020 180.260 115.280 180.520 ;
        RECT 115.340 180.260 115.600 180.520 ;
        RECT 115.660 180.260 115.920 180.520 ;
        RECT 115.980 180.260 116.240 180.520 ;
        RECT 96.710 179.750 96.970 180.010 ;
        RECT 104.070 179.750 104.330 180.010 ;
        RECT 104.530 179.750 104.790 180.010 ;
        RECT 112.810 179.750 113.070 180.010 ;
        RECT 96.250 179.410 96.510 179.670 ;
        RECT 99.930 179.410 100.190 179.670 ;
        RECT 97.170 179.070 97.430 179.330 ;
        RECT 100.390 179.070 100.650 179.330 ;
        RECT 109.590 179.410 109.850 179.670 ;
        RECT 103.150 179.070 103.410 179.330 ;
        RECT 105.910 179.070 106.170 179.330 ;
        RECT 107.750 179.070 108.010 179.330 ;
        RECT 111.430 178.730 111.690 178.990 ;
        RECT 105.450 178.390 105.710 178.650 ;
        RECT 110.970 178.390 111.230 178.650 ;
        RECT 67.205 177.540 67.465 177.800 ;
        RECT 67.525 177.540 67.785 177.800 ;
        RECT 67.845 177.540 68.105 177.800 ;
        RECT 68.165 177.540 68.425 177.800 ;
        RECT 68.485 177.540 68.745 177.800 ;
        RECT 80.775 177.540 81.035 177.800 ;
        RECT 81.095 177.540 81.355 177.800 ;
        RECT 81.415 177.540 81.675 177.800 ;
        RECT 81.735 177.540 81.995 177.800 ;
        RECT 82.055 177.540 82.315 177.800 ;
        RECT 94.345 177.540 94.605 177.800 ;
        RECT 94.665 177.540 94.925 177.800 ;
        RECT 94.985 177.540 95.245 177.800 ;
        RECT 95.305 177.540 95.565 177.800 ;
        RECT 95.625 177.540 95.885 177.800 ;
        RECT 107.915 177.540 108.175 177.800 ;
        RECT 108.235 177.540 108.495 177.800 ;
        RECT 108.555 177.540 108.815 177.800 ;
        RECT 108.875 177.540 109.135 177.800 ;
        RECT 109.195 177.540 109.455 177.800 ;
        RECT 110.050 177.030 110.310 177.290 ;
        RECT 111.430 177.030 111.690 177.290 ;
        RECT 109.590 176.690 109.850 176.950 ;
        RECT 110.510 176.010 110.770 176.270 ;
        RECT 113.270 175.670 113.530 175.930 ;
        RECT 73.990 174.820 74.250 175.080 ;
        RECT 74.310 174.820 74.570 175.080 ;
        RECT 74.630 174.820 74.890 175.080 ;
        RECT 74.950 174.820 75.210 175.080 ;
        RECT 75.270 174.820 75.530 175.080 ;
        RECT 87.560 174.820 87.820 175.080 ;
        RECT 87.880 174.820 88.140 175.080 ;
        RECT 88.200 174.820 88.460 175.080 ;
        RECT 88.520 174.820 88.780 175.080 ;
        RECT 88.840 174.820 89.100 175.080 ;
        RECT 101.130 174.820 101.390 175.080 ;
        RECT 101.450 174.820 101.710 175.080 ;
        RECT 101.770 174.820 102.030 175.080 ;
        RECT 102.090 174.820 102.350 175.080 ;
        RECT 102.410 174.820 102.670 175.080 ;
        RECT 114.700 174.820 114.960 175.080 ;
        RECT 115.020 174.820 115.280 175.080 ;
        RECT 115.340 174.820 115.600 175.080 ;
        RECT 115.660 174.820 115.920 175.080 ;
        RECT 115.980 174.820 116.240 175.080 ;
        RECT 112.350 174.310 112.610 174.570 ;
        RECT 110.050 173.970 110.310 174.230 ;
        RECT 105.910 173.630 106.170 173.890 ;
        RECT 111.890 173.630 112.150 173.890 ;
        RECT 67.205 172.100 67.465 172.360 ;
        RECT 67.525 172.100 67.785 172.360 ;
        RECT 67.845 172.100 68.105 172.360 ;
        RECT 68.165 172.100 68.425 172.360 ;
        RECT 68.485 172.100 68.745 172.360 ;
        RECT 80.775 172.100 81.035 172.360 ;
        RECT 81.095 172.100 81.355 172.360 ;
        RECT 81.415 172.100 81.675 172.360 ;
        RECT 81.735 172.100 81.995 172.360 ;
        RECT 82.055 172.100 82.315 172.360 ;
        RECT 94.345 172.100 94.605 172.360 ;
        RECT 94.665 172.100 94.925 172.360 ;
        RECT 94.985 172.100 95.245 172.360 ;
        RECT 95.305 172.100 95.565 172.360 ;
        RECT 95.625 172.100 95.885 172.360 ;
        RECT 107.915 172.100 108.175 172.360 ;
        RECT 108.235 172.100 108.495 172.360 ;
        RECT 108.555 172.100 108.815 172.360 ;
        RECT 108.875 172.100 109.135 172.360 ;
        RECT 109.195 172.100 109.455 172.360 ;
        RECT 73.990 169.380 74.250 169.640 ;
        RECT 74.310 169.380 74.570 169.640 ;
        RECT 74.630 169.380 74.890 169.640 ;
        RECT 74.950 169.380 75.210 169.640 ;
        RECT 75.270 169.380 75.530 169.640 ;
        RECT 87.560 169.380 87.820 169.640 ;
        RECT 87.880 169.380 88.140 169.640 ;
        RECT 88.200 169.380 88.460 169.640 ;
        RECT 88.520 169.380 88.780 169.640 ;
        RECT 88.840 169.380 89.100 169.640 ;
        RECT 101.130 169.380 101.390 169.640 ;
        RECT 101.450 169.380 101.710 169.640 ;
        RECT 101.770 169.380 102.030 169.640 ;
        RECT 102.090 169.380 102.350 169.640 ;
        RECT 102.410 169.380 102.670 169.640 ;
        RECT 114.700 169.380 114.960 169.640 ;
        RECT 115.020 169.380 115.280 169.640 ;
        RECT 115.340 169.380 115.600 169.640 ;
        RECT 115.660 169.380 115.920 169.640 ;
        RECT 115.980 169.380 116.240 169.640 ;
        RECT 67.205 166.660 67.465 166.920 ;
        RECT 67.525 166.660 67.785 166.920 ;
        RECT 67.845 166.660 68.105 166.920 ;
        RECT 68.165 166.660 68.425 166.920 ;
        RECT 68.485 166.660 68.745 166.920 ;
        RECT 80.775 166.660 81.035 166.920 ;
        RECT 81.095 166.660 81.355 166.920 ;
        RECT 81.415 166.660 81.675 166.920 ;
        RECT 81.735 166.660 81.995 166.920 ;
        RECT 82.055 166.660 82.315 166.920 ;
        RECT 94.345 166.660 94.605 166.920 ;
        RECT 94.665 166.660 94.925 166.920 ;
        RECT 94.985 166.660 95.245 166.920 ;
        RECT 95.305 166.660 95.565 166.920 ;
        RECT 95.625 166.660 95.885 166.920 ;
        RECT 107.915 166.660 108.175 166.920 ;
        RECT 108.235 166.660 108.495 166.920 ;
        RECT 108.555 166.660 108.815 166.920 ;
        RECT 108.875 166.660 109.135 166.920 ;
        RECT 109.195 166.660 109.455 166.920 ;
        RECT 73.990 163.940 74.250 164.200 ;
        RECT 74.310 163.940 74.570 164.200 ;
        RECT 74.630 163.940 74.890 164.200 ;
        RECT 74.950 163.940 75.210 164.200 ;
        RECT 75.270 163.940 75.530 164.200 ;
        RECT 87.560 163.940 87.820 164.200 ;
        RECT 87.880 163.940 88.140 164.200 ;
        RECT 88.200 163.940 88.460 164.200 ;
        RECT 88.520 163.940 88.780 164.200 ;
        RECT 88.840 163.940 89.100 164.200 ;
        RECT 101.130 163.940 101.390 164.200 ;
        RECT 101.450 163.940 101.710 164.200 ;
        RECT 101.770 163.940 102.030 164.200 ;
        RECT 102.090 163.940 102.350 164.200 ;
        RECT 102.410 163.940 102.670 164.200 ;
        RECT 114.700 163.940 114.960 164.200 ;
        RECT 115.020 163.940 115.280 164.200 ;
        RECT 115.340 163.940 115.600 164.200 ;
        RECT 115.660 163.940 115.920 164.200 ;
        RECT 115.980 163.940 116.240 164.200 ;
        RECT 67.205 161.220 67.465 161.480 ;
        RECT 67.525 161.220 67.785 161.480 ;
        RECT 67.845 161.220 68.105 161.480 ;
        RECT 68.165 161.220 68.425 161.480 ;
        RECT 68.485 161.220 68.745 161.480 ;
        RECT 80.775 161.220 81.035 161.480 ;
        RECT 81.095 161.220 81.355 161.480 ;
        RECT 81.415 161.220 81.675 161.480 ;
        RECT 81.735 161.220 81.995 161.480 ;
        RECT 82.055 161.220 82.315 161.480 ;
        RECT 94.345 161.220 94.605 161.480 ;
        RECT 94.665 161.220 94.925 161.480 ;
        RECT 94.985 161.220 95.245 161.480 ;
        RECT 95.305 161.220 95.565 161.480 ;
        RECT 95.625 161.220 95.885 161.480 ;
        RECT 107.915 161.220 108.175 161.480 ;
        RECT 108.235 161.220 108.495 161.480 ;
        RECT 108.555 161.220 108.815 161.480 ;
        RECT 108.875 161.220 109.135 161.480 ;
        RECT 109.195 161.220 109.455 161.480 ;
        RECT 73.990 158.500 74.250 158.760 ;
        RECT 74.310 158.500 74.570 158.760 ;
        RECT 74.630 158.500 74.890 158.760 ;
        RECT 74.950 158.500 75.210 158.760 ;
        RECT 75.270 158.500 75.530 158.760 ;
        RECT 87.560 158.500 87.820 158.760 ;
        RECT 87.880 158.500 88.140 158.760 ;
        RECT 88.200 158.500 88.460 158.760 ;
        RECT 88.520 158.500 88.780 158.760 ;
        RECT 88.840 158.500 89.100 158.760 ;
        RECT 101.130 158.500 101.390 158.760 ;
        RECT 101.450 158.500 101.710 158.760 ;
        RECT 101.770 158.500 102.030 158.760 ;
        RECT 102.090 158.500 102.350 158.760 ;
        RECT 102.410 158.500 102.670 158.760 ;
        RECT 114.700 158.500 114.960 158.760 ;
        RECT 115.020 158.500 115.280 158.760 ;
        RECT 115.340 158.500 115.600 158.760 ;
        RECT 115.660 158.500 115.920 158.760 ;
        RECT 115.980 158.500 116.240 158.760 ;
        RECT 67.205 155.780 67.465 156.040 ;
        RECT 67.525 155.780 67.785 156.040 ;
        RECT 67.845 155.780 68.105 156.040 ;
        RECT 68.165 155.780 68.425 156.040 ;
        RECT 68.485 155.780 68.745 156.040 ;
        RECT 80.775 155.780 81.035 156.040 ;
        RECT 81.095 155.780 81.355 156.040 ;
        RECT 81.415 155.780 81.675 156.040 ;
        RECT 81.735 155.780 81.995 156.040 ;
        RECT 82.055 155.780 82.315 156.040 ;
        RECT 94.345 155.780 94.605 156.040 ;
        RECT 94.665 155.780 94.925 156.040 ;
        RECT 94.985 155.780 95.245 156.040 ;
        RECT 95.305 155.780 95.565 156.040 ;
        RECT 95.625 155.780 95.885 156.040 ;
        RECT 107.915 155.780 108.175 156.040 ;
        RECT 108.235 155.780 108.495 156.040 ;
        RECT 108.555 155.780 108.815 156.040 ;
        RECT 108.875 155.780 109.135 156.040 ;
        RECT 109.195 155.780 109.455 156.040 ;
        RECT 73.990 153.060 74.250 153.320 ;
        RECT 74.310 153.060 74.570 153.320 ;
        RECT 74.630 153.060 74.890 153.320 ;
        RECT 74.950 153.060 75.210 153.320 ;
        RECT 75.270 153.060 75.530 153.320 ;
        RECT 87.560 153.060 87.820 153.320 ;
        RECT 87.880 153.060 88.140 153.320 ;
        RECT 88.200 153.060 88.460 153.320 ;
        RECT 88.520 153.060 88.780 153.320 ;
        RECT 88.840 153.060 89.100 153.320 ;
        RECT 101.130 153.060 101.390 153.320 ;
        RECT 101.450 153.060 101.710 153.320 ;
        RECT 101.770 153.060 102.030 153.320 ;
        RECT 102.090 153.060 102.350 153.320 ;
        RECT 102.410 153.060 102.670 153.320 ;
        RECT 114.700 153.060 114.960 153.320 ;
        RECT 115.020 153.060 115.280 153.320 ;
        RECT 115.340 153.060 115.600 153.320 ;
        RECT 115.660 153.060 115.920 153.320 ;
        RECT 115.980 153.060 116.240 153.320 ;
        RECT 102.780 90.345 103.805 91.370 ;
        RECT 127.110 88.700 127.790 89.380 ;
        RECT 111.765 68.055 112.955 69.245 ;
        RECT 147.090 82.020 148.190 83.120 ;
        RECT 112.490 67.010 113.210 67.730 ;
        RECT 144.780 48.580 145.700 49.500 ;
        RECT 138.340 42.860 139.340 43.160 ;
        RECT 129.890 40.860 130.740 41.210 ;
        RECT 129.790 40.560 130.740 40.860 ;
        RECT 125.290 22.910 126.090 32.710 ;
        RECT 127.390 32.210 128.290 32.560 ;
        RECT 129.890 36.260 130.740 40.560 ;
        RECT 129.790 35.960 130.740 36.260 ;
        RECT 129.890 31.710 130.740 35.960 ;
        RECT 129.790 31.410 130.740 31.710 ;
        RECT 129.890 31.260 130.740 31.410 ;
        RECT 132.040 40.560 132.940 40.860 ;
        RECT 132.040 35.960 132.940 36.260 ;
        RECT 132.040 31.410 132.940 31.710 ;
        RECT 138.440 40.560 139.340 40.860 ;
        RECT 138.340 38.260 139.340 38.560 ;
        RECT 138.440 35.960 139.340 36.260 ;
        RECT 138.340 33.660 139.340 33.960 ;
        RECT 138.440 31.410 139.340 31.710 ;
        RECT 140.640 33.960 141.490 43.610 ;
        RECT 142.940 43.110 143.890 43.410 ;
        RECT 140.640 33.560 141.540 33.960 ;
        RECT 140.640 32.410 141.490 33.560 ;
        RECT 140.640 32.010 141.540 32.410 ;
        RECT 127.390 27.610 128.290 27.960 ;
        RECT 138.340 29.060 139.340 29.360 ;
        RECT 138.615 28.810 139.165 29.060 ;
        RECT 138.390 27.460 139.240 28.110 ;
        RECT 140.640 30.810 141.490 32.010 ;
        RECT 140.640 27.810 141.540 30.810 ;
        RECT 140.640 27.460 141.890 27.810 ;
        RECT 140.740 27.410 141.890 27.460 ;
        RECT 142.990 42.310 143.940 42.610 ;
        RECT 142.940 41.510 143.890 41.810 ;
        RECT 142.990 40.710 143.940 41.010 ;
        RECT 142.940 39.960 143.890 40.260 ;
        RECT 142.990 39.160 143.940 39.460 ;
        RECT 142.940 38.360 143.890 38.660 ;
        RECT 142.990 37.560 143.940 37.860 ;
        RECT 142.940 36.760 143.890 37.060 ;
        RECT 142.990 35.960 143.940 36.260 ;
        RECT 142.940 35.210 143.890 35.510 ;
        RECT 142.990 34.410 143.940 34.710 ;
        RECT 142.940 33.610 143.890 33.910 ;
        RECT 142.990 32.860 143.940 33.160 ;
        RECT 142.940 32.060 143.890 32.360 ;
        RECT 142.990 31.260 143.940 31.560 ;
        RECT 142.940 30.460 143.890 30.760 ;
        RECT 142.440 29.610 142.740 30.010 ;
        RECT 142.990 29.660 143.940 29.960 ;
        RECT 142.940 28.860 143.890 29.160 ;
        RECT 142.990 28.110 143.940 28.410 ;
        RECT 142.940 27.310 143.890 27.610 ;
        RECT 130.340 27.040 131.040 27.060 ;
        RECT 130.315 26.485 131.040 27.040 ;
        RECT 130.340 26.460 131.040 26.485 ;
        RECT 131.640 26.610 131.940 26.960 ;
        RECT 134.740 26.610 135.040 26.960 ;
        RECT 136.240 26.610 136.540 26.960 ;
        RECT 139.340 26.610 139.640 26.960 ;
        RECT 140.365 26.490 140.915 27.040 ;
        RECT 145.090 26.610 145.690 42.460 ;
        RECT 148.790 39.760 149.190 42.460 ;
        RECT 156.410 39.700 157.310 40.600 ;
        RECT 146.890 39.260 147.840 39.560 ;
        RECT 147.040 39.160 147.790 39.260 ;
        RECT 146.940 36.860 147.840 37.160 ;
        RECT 146.940 34.560 147.840 34.860 ;
        RECT 146.940 32.260 147.840 32.560 ;
        RECT 146.940 29.960 147.840 30.310 ;
        RECT 146.940 27.660 147.840 28.010 ;
        RECT 129.140 25.160 129.790 25.810 ;
        RECT 131.190 25.660 132.090 25.960 ;
        RECT 133.290 25.410 133.690 26.110 ;
        RECT 137.840 25.410 138.240 26.110 ;
        RECT 139.340 25.660 140.240 25.960 ;
        RECT 147.040 25.360 147.840 25.660 ;
        RECT 130.990 23.510 131.290 24.410 ;
        RECT 133.290 23.610 133.640 24.310 ;
        RECT 135.590 23.610 135.940 24.310 ;
        RECT 137.890 23.610 138.240 24.310 ;
        RECT 140.190 23.510 140.490 24.410 ;
        RECT 127.390 22.960 128.290 23.310 ;
        RECT 148.740 24.610 149.140 37.110 ;
        RECT 146.940 23.060 147.840 23.410 ;
        RECT 130.840 22.260 131.340 22.360 ;
        RECT 135.590 22.260 135.940 22.360 ;
        RECT 139.990 22.260 140.490 22.360 ;
        RECT 130.840 21.910 140.490 22.260 ;
        RECT 130.840 21.610 140.440 21.910 ;
        RECT 150.940 13.660 152.140 14.860 ;
      LAYER met2 ;
        RECT 94.380 218.550 94.680 218.560 ;
        RECT 94.345 218.270 94.715 218.550 ;
        RECT 87.950 217.340 88.250 217.350 ;
        RECT 87.915 217.060 88.285 217.340 ;
        RECT 81.540 216.070 81.840 216.080 ;
        RECT 81.505 215.790 81.875 216.070 ;
        RECT 75.080 214.480 75.380 214.490 ;
        RECT 75.045 214.200 75.415 214.480 ;
        RECT 68.620 213.130 68.920 213.140 ;
        RECT 62.070 213.020 62.370 213.030 ;
        RECT 62.035 212.740 62.405 213.020 ;
        RECT 68.585 212.850 68.955 213.130 ;
        RECT 62.070 210.470 62.370 212.740 ;
        RECT 62.070 209.470 62.480 210.470 ;
        RECT 68.620 209.710 68.920 212.850 ;
        RECT 62.200 208.470 62.480 209.470 ;
        RECT 68.640 208.470 68.920 209.710 ;
        RECT 75.080 209.450 75.380 214.200 ;
        RECT 81.540 210.470 81.840 215.790 ;
        RECT 81.520 209.530 81.840 210.470 ;
        RECT 87.950 209.550 88.250 217.060 ;
        RECT 94.380 209.740 94.680 218.270 ;
        RECT 107.330 215.800 107.630 215.810 ;
        RECT 107.295 215.520 107.665 215.800 ;
        RECT 100.840 214.190 101.140 214.200 ;
        RECT 100.805 213.910 101.175 214.190 ;
        RECT 75.080 208.470 75.360 209.450 ;
        RECT 78.310 208.620 78.570 208.940 ;
        RECT 62.270 204.520 62.410 208.470 ;
        RECT 68.710 205.960 68.850 208.470 ;
        RECT 75.150 208.260 75.290 208.470 ;
        RECT 72.790 207.940 73.050 208.260 ;
        RECT 75.090 207.940 75.350 208.260 ;
        RECT 71.870 206.580 72.130 206.900 ;
        RECT 68.710 205.820 69.310 205.960 ;
        RECT 67.205 204.685 68.745 205.055 ;
        RECT 69.170 204.520 69.310 205.820 ;
        RECT 62.210 204.200 62.470 204.520 ;
        RECT 69.110 204.200 69.370 204.520 ;
        RECT 63.590 203.860 63.850 204.180 ;
        RECT 63.650 201.120 63.790 203.860 ;
        RECT 64.970 203.180 65.230 203.500 ;
        RECT 66.810 203.180 67.070 203.500 ;
        RECT 64.510 202.840 64.770 203.160 ;
        RECT 64.050 201.140 64.310 201.460 ;
        RECT 63.590 200.800 63.850 201.120 ;
        RECT 64.110 198.740 64.250 201.140 ;
        RECT 64.570 201.120 64.710 202.840 ;
        RECT 64.510 200.800 64.770 201.120 ;
        RECT 64.510 199.780 64.770 200.100 ;
        RECT 64.050 198.420 64.310 198.740 ;
        RECT 64.570 198.595 64.710 199.780 ;
        RECT 65.030 199.080 65.170 203.180 ;
        RECT 66.870 200.440 67.010 203.180 ;
        RECT 71.410 202.500 71.670 202.820 ;
        RECT 70.490 200.800 70.750 201.120 ;
        RECT 66.810 200.120 67.070 200.440 ;
        RECT 66.350 199.780 66.610 200.100 ;
        RECT 64.970 198.760 65.230 199.080 ;
        RECT 64.500 198.225 64.780 198.595 ;
        RECT 66.410 198.060 66.550 199.780 ;
        RECT 67.205 199.245 68.745 199.615 ;
        RECT 66.350 197.740 66.610 198.060 ;
        RECT 70.550 196.360 70.690 200.800 ;
        RECT 71.470 197.380 71.610 202.500 ;
        RECT 71.930 201.800 72.070 206.580 ;
        RECT 72.850 204.520 72.990 207.940 ;
        RECT 73.990 207.405 75.530 207.775 ;
        RECT 78.370 206.900 78.510 208.620 ;
        RECT 81.520 208.470 81.800 209.530 ;
        RECT 87.960 208.470 88.240 209.550 ;
        RECT 81.590 207.240 81.730 208.470 ;
        RECT 88.030 208.260 88.170 208.470 ;
        RECT 91.650 208.280 91.910 208.600 ;
        RECT 94.400 208.470 94.680 209.740 ;
        RECT 100.840 209.660 101.140 213.910 ;
        RECT 107.330 210.470 107.630 215.520 ;
        RECT 113.700 211.310 114.000 211.320 ;
        RECT 113.665 211.030 114.035 211.310 ;
        RECT 113.700 210.860 114.000 211.030 ;
        RECT 107.280 209.790 107.630 210.470 ;
        RECT 97.630 208.620 97.890 208.940 ;
        RECT 87.970 207.940 88.230 208.260 ;
        RECT 89.350 207.940 89.610 208.260 ;
        RECT 87.560 207.405 89.100 207.775 ;
        RECT 89.410 207.240 89.550 207.940 ;
        RECT 81.530 206.920 81.790 207.240 ;
        RECT 89.350 206.920 89.610 207.240 ;
        RECT 78.310 206.580 78.570 206.900 ;
        RECT 73.710 206.240 73.970 206.560 ;
        RECT 73.250 205.220 73.510 205.540 ;
        RECT 72.790 204.200 73.050 204.520 ;
        RECT 71.870 201.480 72.130 201.800 ;
        RECT 72.790 201.140 73.050 201.460 ;
        RECT 72.330 200.800 72.590 201.120 ;
        RECT 71.410 197.060 71.670 197.380 ;
        RECT 70.490 196.040 70.750 196.360 ;
        RECT 71.470 195.000 71.610 197.060 ;
        RECT 71.410 194.680 71.670 195.000 ;
        RECT 67.205 193.805 68.745 194.175 ;
        RECT 72.390 193.640 72.530 200.800 ;
        RECT 72.850 196.360 72.990 201.140 ;
        RECT 72.790 196.040 73.050 196.360 ;
        RECT 72.330 193.320 72.590 193.640 ;
        RECT 73.310 192.620 73.450 205.220 ;
        RECT 73.770 204.520 73.910 206.240 ;
        RECT 76.470 205.900 76.730 206.220 ;
        RECT 77.390 205.900 77.650 206.220 ;
        RECT 73.710 204.200 73.970 204.520 ;
        RECT 73.770 203.500 73.910 204.200 ;
        RECT 76.530 203.500 76.670 205.900 ;
        RECT 76.930 205.220 77.190 205.540 ;
        RECT 76.990 203.500 77.130 205.220 ;
        RECT 77.450 204.180 77.590 205.900 ;
        RECT 78.370 204.600 78.510 206.580 ;
        RECT 91.710 206.560 91.850 208.280 ;
        RECT 94.470 208.260 94.610 208.470 ;
        RECT 94.410 207.940 94.670 208.260 ;
        RECT 93.550 207.180 94.610 207.320 ;
        RECT 93.550 206.640 93.690 207.180 ;
        RECT 84.290 206.240 84.550 206.560 ;
        RECT 91.650 206.240 91.910 206.560 ;
        RECT 92.630 206.500 93.690 206.640 ;
        RECT 83.370 205.220 83.630 205.540 ;
        RECT 80.775 204.685 82.315 205.055 ;
        RECT 78.370 204.460 79.430 204.600 ;
        RECT 77.390 203.860 77.650 204.180 ;
        RECT 78.770 203.860 79.030 204.180 ;
        RECT 73.710 203.180 73.970 203.500 ;
        RECT 74.630 203.180 74.890 203.500 ;
        RECT 76.470 203.180 76.730 203.500 ;
        RECT 76.930 203.180 77.190 203.500 ;
        RECT 74.690 202.730 74.830 203.180 ;
        RECT 74.690 202.590 76.210 202.730 ;
        RECT 73.990 201.965 75.530 202.335 ;
        RECT 76.070 201.800 76.210 202.590 ;
        RECT 76.010 201.480 76.270 201.800 ;
        RECT 75.550 200.800 75.810 201.120 ;
        RECT 73.710 200.460 73.970 200.780 ;
        RECT 73.770 198.740 73.910 200.460 ;
        RECT 73.710 198.420 73.970 198.740 ;
        RECT 75.080 198.225 75.360 198.595 ;
        RECT 73.710 197.915 73.970 198.060 ;
        RECT 73.700 197.545 73.980 197.915 ;
        RECT 75.150 197.720 75.290 198.225 ;
        RECT 75.090 197.400 75.350 197.720 ;
        RECT 75.610 197.630 75.750 200.800 ;
        RECT 76.530 200.100 76.670 203.180 ;
        RECT 76.990 201.800 77.130 203.180 ;
        RECT 76.930 201.480 77.190 201.800 ;
        RECT 76.470 199.780 76.730 200.100 ;
        RECT 76.010 197.800 76.270 198.060 ;
        RECT 76.010 197.740 77.130 197.800 ;
        RECT 76.070 197.660 77.130 197.740 ;
        RECT 75.610 197.490 75.910 197.630 ;
        RECT 75.770 197.290 75.910 197.490 ;
        RECT 75.770 197.150 76.210 197.290 ;
        RECT 73.990 196.525 75.530 196.895 ;
        RECT 75.090 194.570 75.350 194.660 ;
        RECT 76.070 194.570 76.210 197.150 ;
        RECT 76.990 195.340 77.130 197.660 ;
        RECT 77.450 196.360 77.590 203.860 ;
        RECT 78.310 203.180 78.570 203.500 ;
        RECT 77.850 199.840 78.110 200.100 ;
        RECT 78.370 199.840 78.510 203.180 ;
        RECT 77.850 199.780 78.510 199.840 ;
        RECT 77.910 199.700 78.510 199.780 ;
        RECT 77.390 196.040 77.650 196.360 ;
        RECT 78.370 196.020 78.510 199.700 ;
        RECT 78.830 197.380 78.970 203.860 ;
        RECT 79.290 203.500 79.430 204.460 ;
        RECT 79.230 203.180 79.490 203.500 ;
        RECT 79.290 201.120 79.430 203.180 ;
        RECT 82.450 202.840 82.710 203.160 ;
        RECT 79.230 200.800 79.490 201.120 ;
        RECT 78.770 197.060 79.030 197.380 ;
        RECT 78.310 195.700 78.570 196.020 ;
        RECT 76.930 195.020 77.190 195.340 ;
        RECT 75.090 194.430 76.210 194.570 ;
        RECT 75.090 194.340 75.350 194.430 ;
        RECT 73.250 192.300 73.510 192.620 ;
        RECT 75.150 192.280 75.290 194.340 ;
        RECT 76.010 192.980 76.270 193.300 ;
        RECT 75.090 191.960 75.350 192.280 ;
        RECT 73.250 191.620 73.510 191.940 ;
        RECT 73.310 190.240 73.450 191.620 ;
        RECT 73.990 191.085 75.530 191.455 ;
        RECT 76.070 190.320 76.210 192.980 ;
        RECT 76.470 192.300 76.730 192.620 ;
        RECT 75.610 190.240 76.210 190.320 ;
        RECT 72.330 189.920 72.590 190.240 ;
        RECT 73.250 189.920 73.510 190.240 ;
        RECT 75.550 190.180 76.210 190.240 ;
        RECT 75.550 189.920 75.810 190.180 ;
        RECT 71.410 188.900 71.670 189.220 ;
        RECT 67.205 188.365 68.745 188.735 ;
        RECT 71.470 187.520 71.610 188.900 ;
        RECT 71.410 187.200 71.670 187.520 ;
        RECT 70.950 186.520 71.210 186.840 ;
        RECT 71.010 184.800 71.150 186.520 ;
        RECT 70.950 184.480 71.210 184.800 ;
        RECT 67.205 182.925 68.745 183.295 ;
        RECT 72.390 182.760 72.530 189.920 ;
        RECT 73.250 188.900 73.510 189.220 ;
        RECT 75.090 188.900 75.350 189.220 ;
        RECT 73.310 188.200 73.450 188.900 ;
        RECT 73.250 187.880 73.510 188.200 ;
        RECT 75.150 186.840 75.290 188.900 ;
        RECT 76.010 187.880 76.270 188.200 ;
        RECT 73.250 186.520 73.510 186.840 ;
        RECT 75.090 186.520 75.350 186.840 ;
        RECT 72.330 182.440 72.590 182.760 ;
        RECT 73.310 181.060 73.450 186.520 ;
        RECT 73.990 185.645 75.530 186.015 ;
        RECT 76.070 185.480 76.210 187.880 ;
        RECT 76.530 186.500 76.670 192.300 ;
        RECT 76.990 190.580 77.130 195.020 ;
        RECT 78.370 192.620 78.510 195.700 ;
        RECT 78.830 194.660 78.970 197.060 ;
        RECT 79.290 195.680 79.430 200.800 ;
        RECT 82.510 200.780 82.650 202.840 ;
        RECT 83.430 201.460 83.570 205.220 ;
        RECT 83.370 201.140 83.630 201.460 ;
        RECT 82.450 200.460 82.710 200.780 ;
        RECT 80.775 199.245 82.315 199.615 ;
        RECT 82.510 198.400 82.650 200.460 ;
        RECT 82.910 198.420 83.170 198.740 ;
        RECT 82.450 198.080 82.710 198.400 ;
        RECT 82.970 197.720 83.110 198.420 ;
        RECT 82.910 197.400 83.170 197.720 ;
        RECT 79.230 195.590 79.490 195.680 ;
        RECT 79.230 195.450 79.890 195.590 ;
        RECT 79.230 195.360 79.490 195.450 ;
        RECT 78.770 194.340 79.030 194.660 ;
        RECT 78.770 193.210 79.030 193.300 ;
        RECT 78.770 193.070 79.430 193.210 ;
        RECT 78.770 192.980 79.030 193.070 ;
        RECT 78.310 192.300 78.570 192.620 ;
        RECT 79.290 192.280 79.430 193.070 ;
        RECT 79.230 191.960 79.490 192.280 ;
        RECT 77.390 191.620 77.650 191.940 ;
        RECT 76.930 190.260 77.190 190.580 ;
        RECT 76.990 187.180 77.130 190.260 ;
        RECT 77.450 187.180 77.590 191.620 ;
        RECT 76.930 186.860 77.190 187.180 ;
        RECT 77.390 186.860 77.650 187.180 ;
        RECT 76.470 186.180 76.730 186.500 ;
        RECT 76.010 185.160 76.270 185.480 ;
        RECT 76.070 181.740 76.210 185.160 ;
        RECT 76.530 182.420 76.670 186.180 ;
        RECT 76.990 184.460 77.130 186.860 ;
        RECT 78.310 184.480 78.570 184.800 ;
        RECT 76.930 184.140 77.190 184.460 ;
        RECT 78.370 182.760 78.510 184.480 ;
        RECT 78.310 182.440 78.570 182.760 ;
        RECT 76.470 182.100 76.730 182.420 ;
        RECT 76.010 181.420 76.270 181.740 ;
        RECT 79.290 181.400 79.430 191.960 ;
        RECT 79.750 184.800 79.890 195.450 ;
        RECT 80.775 193.805 82.315 194.175 ;
        RECT 81.990 192.640 82.250 192.960 ;
        RECT 82.050 190.920 82.190 192.640 ;
        RECT 82.450 192.190 82.710 192.280 ;
        RECT 82.970 192.190 83.110 197.400 ;
        RECT 84.350 193.300 84.490 206.240 ;
        RECT 86.130 205.560 86.390 205.880 ;
        RECT 85.210 202.840 85.470 203.160 ;
        RECT 85.270 201.800 85.410 202.840 ;
        RECT 85.210 201.480 85.470 201.800 ;
        RECT 86.190 201.120 86.330 205.560 ;
        RECT 92.110 205.220 92.370 205.540 ;
        RECT 92.170 204.520 92.310 205.220 ;
        RECT 92.110 204.200 92.370 204.520 ;
        RECT 92.630 203.240 92.770 206.500 ;
        RECT 93.950 206.240 94.210 206.560 ;
        RECT 93.030 205.900 93.290 206.220 ;
        RECT 93.490 205.900 93.750 206.220 ;
        RECT 93.090 204.180 93.230 205.900 ;
        RECT 93.030 203.860 93.290 204.180 ;
        RECT 87.050 202.840 87.310 203.160 ;
        RECT 92.630 203.100 93.230 203.240 ;
        RECT 86.130 200.800 86.390 201.120 ;
        RECT 85.660 200.265 85.940 200.635 ;
        RECT 85.730 198.740 85.870 200.265 ;
        RECT 85.670 198.420 85.930 198.740 ;
        RECT 84.740 197.545 85.020 197.915 ;
        RECT 85.670 197.740 85.930 198.060 ;
        RECT 84.750 197.400 85.010 197.545 ;
        RECT 85.730 195.340 85.870 197.740 ;
        RECT 87.110 196.360 87.250 202.840 ;
        RECT 92.110 202.500 92.370 202.820 ;
        RECT 87.560 201.965 89.100 202.335 ;
        RECT 92.170 201.460 92.310 202.500 ;
        RECT 92.110 201.140 92.370 201.460 ;
        RECT 87.510 199.780 87.770 200.100 ;
        RECT 87.570 198.840 87.710 199.780 ;
        RECT 93.090 198.840 93.230 203.100 ;
        RECT 93.550 201.120 93.690 205.900 ;
        RECT 94.010 202.820 94.150 206.240 ;
        RECT 94.470 206.220 94.610 207.180 ;
        RECT 96.710 206.810 96.970 206.900 ;
        RECT 96.710 206.670 97.370 206.810 ;
        RECT 96.710 206.580 96.970 206.670 ;
        RECT 96.250 206.240 96.510 206.560 ;
        RECT 94.410 205.900 94.670 206.220 ;
        RECT 96.310 205.960 96.450 206.240 ;
        RECT 94.930 205.880 96.450 205.960 ;
        RECT 94.870 205.820 96.450 205.880 ;
        RECT 94.870 205.560 95.130 205.820 ;
        RECT 96.710 205.560 96.970 205.880 ;
        RECT 96.250 205.220 96.510 205.540 ;
        RECT 94.345 204.685 95.885 205.055 ;
        RECT 95.790 203.180 96.050 203.500 ;
        RECT 93.950 202.500 94.210 202.820 ;
        RECT 93.490 200.800 93.750 201.120 ;
        RECT 93.550 200.100 93.690 200.800 ;
        RECT 94.010 200.440 94.150 202.500 ;
        RECT 95.850 201.200 95.990 203.180 ;
        RECT 96.310 201.800 96.450 205.220 ;
        RECT 96.250 201.480 96.510 201.800 ;
        RECT 95.850 201.060 96.450 201.200 ;
        RECT 96.770 201.120 96.910 205.560 ;
        RECT 97.230 205.540 97.370 206.670 ;
        RECT 97.690 206.560 97.830 208.620 ;
        RECT 98.550 208.280 98.810 208.600 ;
        RECT 99.930 208.280 100.190 208.600 ;
        RECT 100.840 208.470 101.120 209.660 ;
        RECT 106.370 208.620 106.630 208.940 ;
        RECT 100.850 208.280 101.110 208.470 ;
        RECT 98.610 206.560 98.750 208.280 ;
        RECT 99.990 207.240 100.130 208.280 ;
        RECT 105.910 207.940 106.170 208.260 ;
        RECT 101.130 207.405 102.670 207.775 ;
        RECT 99.930 206.920 100.190 207.240 ;
        RECT 97.630 206.240 97.890 206.560 ;
        RECT 98.550 206.240 98.810 206.560 ;
        RECT 103.150 206.240 103.410 206.560 ;
        RECT 98.090 205.560 98.350 205.880 ;
        RECT 97.170 205.220 97.430 205.540 ;
        RECT 97.230 203.500 97.370 205.220 ;
        RECT 97.170 203.180 97.430 203.500 ;
        RECT 93.950 200.120 94.210 200.440 ;
        RECT 93.490 199.780 93.750 200.100 ;
        RECT 93.550 199.080 93.690 199.780 ;
        RECT 94.345 199.245 95.885 199.615 ;
        RECT 87.570 198.700 88.170 198.840 ;
        RECT 88.030 197.720 88.170 198.700 ;
        RECT 92.630 198.700 93.230 198.840 ;
        RECT 93.490 198.760 93.750 199.080 ;
        RECT 92.630 197.915 92.770 198.700 ;
        RECT 94.870 198.420 95.130 198.740 ;
        RECT 94.930 197.915 95.070 198.420 ;
        RECT 87.970 197.400 88.230 197.720 ;
        RECT 92.560 197.545 92.840 197.915 ;
        RECT 94.860 197.545 95.140 197.915 ;
        RECT 96.310 197.720 96.450 201.060 ;
        RECT 96.710 200.800 96.970 201.120 ;
        RECT 97.230 200.520 97.370 203.180 ;
        RECT 98.150 202.820 98.290 205.560 ;
        RECT 98.610 203.840 98.750 206.240 ;
        RECT 99.010 205.900 99.270 206.220 ;
        RECT 98.550 203.520 98.810 203.840 ;
        RECT 98.090 202.500 98.350 202.820 ;
        RECT 97.630 200.800 97.890 201.120 ;
        RECT 96.770 200.380 97.370 200.520 ;
        RECT 87.560 196.525 89.100 196.895 ;
        RECT 87.050 196.040 87.310 196.360 ;
        RECT 90.270 195.360 90.530 195.680 ;
        RECT 85.670 195.020 85.930 195.340 ;
        RECT 84.290 192.980 84.550 193.300 ;
        RECT 87.050 192.300 87.310 192.620 ;
        RECT 89.810 192.300 90.070 192.620 ;
        RECT 82.450 192.050 83.110 192.190 ;
        RECT 82.450 191.960 82.710 192.050 ;
        RECT 83.370 191.960 83.630 192.280 ;
        RECT 83.830 191.960 84.090 192.280 ;
        RECT 81.990 190.600 82.250 190.920 ;
        RECT 83.430 189.220 83.570 191.960 ;
        RECT 83.370 188.900 83.630 189.220 ;
        RECT 80.775 188.365 82.315 188.735 ;
        RECT 79.690 184.480 79.950 184.800 ;
        RECT 83.890 184.120 84.030 191.960 ;
        RECT 84.290 191.620 84.550 191.940 ;
        RECT 84.750 191.620 85.010 191.940 ;
        RECT 84.350 188.200 84.490 191.620 ;
        RECT 84.810 190.240 84.950 191.620 ;
        RECT 84.750 189.920 85.010 190.240 ;
        RECT 84.290 187.880 84.550 188.200 ;
        RECT 84.350 187.180 84.490 187.880 ;
        RECT 84.810 187.180 84.950 189.920 ;
        RECT 85.670 189.580 85.930 189.900 ;
        RECT 85.210 188.900 85.470 189.220 ;
        RECT 84.290 186.860 84.550 187.180 ;
        RECT 84.750 186.860 85.010 187.180 ;
        RECT 85.270 186.500 85.410 188.900 ;
        RECT 85.730 188.200 85.870 189.580 ;
        RECT 86.130 188.900 86.390 189.220 ;
        RECT 85.670 187.880 85.930 188.200 ;
        RECT 86.190 187.180 86.330 188.900 ;
        RECT 86.130 186.860 86.390 187.180 ;
        RECT 86.590 186.860 86.850 187.180 ;
        RECT 85.210 186.180 85.470 186.500 ;
        RECT 86.650 185.140 86.790 186.860 ;
        RECT 86.590 184.820 86.850 185.140 ;
        RECT 83.830 183.800 84.090 184.120 ;
        RECT 80.775 182.925 82.315 183.295 ;
        RECT 83.890 181.740 84.030 183.800 ;
        RECT 85.210 183.460 85.470 183.780 ;
        RECT 85.270 182.080 85.410 183.460 ;
        RECT 86.650 182.080 86.790 184.820 ;
        RECT 87.110 184.800 87.250 192.300 ;
        RECT 89.350 191.620 89.610 191.940 ;
        RECT 87.560 191.085 89.100 191.455 ;
        RECT 89.410 187.180 89.550 191.620 ;
        RECT 89.350 186.860 89.610 187.180 ;
        RECT 87.560 185.645 89.100 186.015 ;
        RECT 87.050 184.480 87.310 184.800 ;
        RECT 88.890 184.480 89.150 184.800 ;
        RECT 88.950 182.760 89.090 184.480 ;
        RECT 89.870 184.120 90.010 192.300 ;
        RECT 90.330 189.220 90.470 195.360 ;
        RECT 92.630 192.620 92.770 197.545 ;
        RECT 96.250 197.400 96.510 197.720 ;
        RECT 93.950 197.060 94.210 197.380 ;
        RECT 94.870 197.120 95.130 197.380 ;
        RECT 96.770 197.120 96.910 200.380 ;
        RECT 97.170 199.840 97.430 200.100 ;
        RECT 97.690 199.840 97.830 200.800 ;
        RECT 97.170 199.780 97.830 199.840 ;
        RECT 97.230 199.700 97.830 199.780 ;
        RECT 97.230 198.400 97.370 199.700 ;
        RECT 97.170 198.080 97.430 198.400 ;
        RECT 94.870 197.060 96.910 197.120 ;
        RECT 97.170 197.060 97.430 197.380 ;
        RECT 93.490 193.320 93.750 193.640 ;
        RECT 90.730 192.300 90.990 192.620 ;
        RECT 92.570 192.530 92.830 192.620 ;
        RECT 92.170 192.390 92.830 192.530 ;
        RECT 90.790 190.920 90.930 192.300 ;
        RECT 91.650 191.960 91.910 192.280 ;
        RECT 90.730 190.600 90.990 190.920 ;
        RECT 90.270 188.900 90.530 189.220 ;
        RECT 91.710 184.800 91.850 191.960 ;
        RECT 92.170 186.840 92.310 192.390 ;
        RECT 92.570 192.300 92.830 192.390 ;
        RECT 93.030 192.300 93.290 192.620 ;
        RECT 92.570 191.620 92.830 191.940 ;
        RECT 92.110 186.520 92.370 186.840 ;
        RECT 91.650 184.480 91.910 184.800 ;
        RECT 89.810 183.800 90.070 184.120 ;
        RECT 88.890 182.440 89.150 182.760 ;
        RECT 85.210 181.760 85.470 182.080 ;
        RECT 86.590 181.760 86.850 182.080 ;
        RECT 92.630 181.740 92.770 191.620 ;
        RECT 93.090 190.920 93.230 192.300 ;
        RECT 93.030 190.600 93.290 190.920 ;
        RECT 93.550 187.600 93.690 193.320 ;
        RECT 94.010 192.960 94.150 197.060 ;
        RECT 94.930 196.980 96.910 197.060 ;
        RECT 96.710 194.340 96.970 194.660 ;
        RECT 94.345 193.805 95.885 194.175 ;
        RECT 93.950 192.640 94.210 192.960 ;
        RECT 94.410 192.300 94.670 192.620 ;
        RECT 95.790 192.300 96.050 192.620 ;
        RECT 94.470 189.900 94.610 192.300 ;
        RECT 95.850 191.000 95.990 192.300 ;
        RECT 96.770 191.000 96.910 194.340 ;
        RECT 97.230 193.640 97.370 197.060 ;
        RECT 97.630 195.360 97.890 195.680 ;
        RECT 97.170 193.320 97.430 193.640 ;
        RECT 97.230 192.620 97.370 193.320 ;
        RECT 97.170 192.300 97.430 192.620 ;
        RECT 95.850 190.920 96.450 191.000 ;
        RECT 95.850 190.860 96.510 190.920 ;
        RECT 96.770 190.860 97.370 191.000 ;
        RECT 95.850 189.900 95.990 190.860 ;
        RECT 96.250 190.600 96.510 190.860 ;
        RECT 96.710 190.260 96.970 190.580 ;
        RECT 96.250 189.920 96.510 190.240 ;
        RECT 94.410 189.580 94.670 189.900 ;
        RECT 95.790 189.580 96.050 189.900 ;
        RECT 94.470 189.130 94.610 189.580 ;
        RECT 94.010 188.990 94.610 189.130 ;
        RECT 94.010 188.200 94.150 188.990 ;
        RECT 94.345 188.365 95.885 188.735 ;
        RECT 93.950 187.880 94.210 188.200 ;
        RECT 93.550 187.460 94.150 187.600 ;
        RECT 94.010 187.180 94.150 187.460 ;
        RECT 93.950 186.860 94.210 187.180 ;
        RECT 94.010 185.140 94.150 186.860 ;
        RECT 93.950 184.820 94.210 185.140 ;
        RECT 94.345 182.925 95.885 183.295 ;
        RECT 96.310 182.080 96.450 189.920 ;
        RECT 96.250 181.760 96.510 182.080 ;
        RECT 83.830 181.420 84.090 181.740 ;
        RECT 92.570 181.420 92.830 181.740 ;
        RECT 79.230 181.080 79.490 181.400 ;
        RECT 73.250 180.740 73.510 181.060 ;
        RECT 73.990 180.205 75.530 180.575 ;
        RECT 87.560 180.205 89.100 180.575 ;
        RECT 96.310 179.700 96.450 181.760 ;
        RECT 96.770 180.040 96.910 190.260 ;
        RECT 97.230 189.560 97.370 190.860 ;
        RECT 97.170 189.240 97.430 189.560 ;
        RECT 97.170 186.860 97.430 187.180 ;
        RECT 97.230 183.780 97.370 186.860 ;
        RECT 97.170 183.460 97.430 183.780 ;
        RECT 96.710 179.720 96.970 180.040 ;
        RECT 96.250 179.380 96.510 179.700 ;
        RECT 97.230 179.360 97.370 183.460 ;
        RECT 97.690 179.555 97.830 195.360 ;
        RECT 98.150 195.340 98.290 202.500 ;
        RECT 98.610 200.100 98.750 203.520 ;
        RECT 99.070 201.800 99.210 205.900 ;
        RECT 99.930 204.200 100.190 204.520 ;
        RECT 99.470 203.860 99.730 204.180 ;
        RECT 99.010 201.480 99.270 201.800 ;
        RECT 99.530 201.120 99.670 203.860 ;
        RECT 99.470 200.800 99.730 201.120 ;
        RECT 99.990 200.440 100.130 204.200 ;
        RECT 101.130 201.965 102.670 202.335 ;
        RECT 99.930 200.120 100.190 200.440 ;
        RECT 98.550 199.780 98.810 200.100 ;
        RECT 99.470 198.760 99.730 199.080 ;
        RECT 99.010 197.400 99.270 197.720 ;
        RECT 98.550 197.060 98.810 197.380 ;
        RECT 98.090 195.020 98.350 195.340 ;
        RECT 98.090 192.300 98.350 192.620 ;
        RECT 98.150 188.200 98.290 192.300 ;
        RECT 98.610 190.580 98.750 197.060 ;
        RECT 99.070 194.660 99.210 197.400 ;
        RECT 99.010 194.340 99.270 194.660 ;
        RECT 99.530 193.720 99.670 198.760 ;
        RECT 99.990 198.740 100.130 200.120 ;
        RECT 103.210 199.080 103.350 206.240 ;
        RECT 104.990 202.500 105.250 202.820 ;
        RECT 103.150 198.760 103.410 199.080 ;
        RECT 99.930 198.420 100.190 198.740 ;
        RECT 105.050 198.595 105.190 202.500 ;
        RECT 105.970 201.800 106.110 207.940 ;
        RECT 106.430 201.800 106.570 208.620 ;
        RECT 107.280 208.470 107.560 209.790 ;
        RECT 113.720 208.470 114.000 210.860 ;
        RECT 105.910 201.480 106.170 201.800 ;
        RECT 106.370 201.480 106.630 201.800 ;
        RECT 106.830 201.140 107.090 201.460 ;
        RECT 104.980 198.225 105.260 198.595 ;
        RECT 106.890 198.060 107.030 201.140 ;
        RECT 107.350 200.635 107.490 208.470 ;
        RECT 113.790 207.320 113.930 208.470 ;
        RECT 114.700 207.405 116.240 207.775 ;
        RECT 113.790 207.180 114.390 207.320 ;
        RECT 113.730 206.580 113.990 206.900 ;
        RECT 112.350 205.900 112.610 206.220 ;
        RECT 109.590 205.220 109.850 205.540 ;
        RECT 107.915 204.685 109.455 205.055 ;
        RECT 107.280 200.265 107.560 200.635 ;
        RECT 107.290 199.780 107.550 200.100 ;
        RECT 101.770 197.915 102.030 198.060 ;
        RECT 101.760 197.545 102.040 197.915 ;
        RECT 106.830 197.740 107.090 198.060 ;
        RECT 103.610 197.400 103.870 197.720 ;
        RECT 101.130 196.525 102.670 196.895 ;
        RECT 103.670 196.360 103.810 197.400 ;
        RECT 103.610 196.040 103.870 196.360 ;
        RECT 107.350 195.340 107.490 199.780 ;
        RECT 107.915 199.245 109.455 199.615 ;
        RECT 109.650 197.380 109.790 205.220 ;
        RECT 112.410 203.840 112.550 205.900 ;
        RECT 112.350 203.520 112.610 203.840 ;
        RECT 113.790 203.500 113.930 206.580 ;
        RECT 113.730 203.180 113.990 203.500 ;
        RECT 110.970 200.460 111.230 200.780 ;
        RECT 110.050 197.740 110.310 198.060 ;
        RECT 109.590 197.060 109.850 197.380 ;
        RECT 110.110 196.020 110.250 197.740 ;
        RECT 110.510 197.060 110.770 197.380 ;
        RECT 110.050 195.700 110.310 196.020 ;
        RECT 107.290 195.020 107.550 195.340 ;
        RECT 109.590 195.020 109.850 195.340 ;
        RECT 99.930 194.340 100.190 194.660 ;
        RECT 99.070 193.580 99.670 193.720 ;
        RECT 99.070 190.920 99.210 193.580 ;
        RECT 99.470 192.300 99.730 192.620 ;
        RECT 99.010 190.600 99.270 190.920 ;
        RECT 98.550 190.260 98.810 190.580 ;
        RECT 99.530 190.320 99.670 192.300 ;
        RECT 99.070 190.180 99.670 190.320 ;
        RECT 98.090 187.880 98.350 188.200 ;
        RECT 98.090 186.520 98.350 186.840 ;
        RECT 98.150 181.060 98.290 186.520 ;
        RECT 99.070 186.500 99.210 190.180 ;
        RECT 99.470 189.580 99.730 189.900 ;
        RECT 99.530 188.200 99.670 189.580 ;
        RECT 99.470 187.880 99.730 188.200 ;
        RECT 99.470 186.520 99.730 186.840 ;
        RECT 99.010 186.180 99.270 186.500 ;
        RECT 99.070 182.760 99.210 186.180 ;
        RECT 99.010 182.440 99.270 182.760 ;
        RECT 99.530 182.420 99.670 186.520 ;
        RECT 99.470 182.100 99.730 182.420 ;
        RECT 98.090 180.740 98.350 181.060 ;
        RECT 99.990 179.700 100.130 194.340 ;
        RECT 107.915 193.805 109.455 194.175 ;
        RECT 102.690 192.360 102.950 192.620 ;
        RECT 102.690 192.300 103.350 192.360 ;
        RECT 106.830 192.300 107.090 192.620 ;
        RECT 100.390 191.960 100.650 192.280 ;
        RECT 102.750 192.220 103.350 192.300 ;
        RECT 100.450 184.800 100.590 191.960 ;
        RECT 101.130 191.085 102.670 191.455 ;
        RECT 103.210 190.920 103.350 192.220 ;
        RECT 103.610 191.960 103.870 192.280 ;
        RECT 105.910 191.960 106.170 192.280 ;
        RECT 103.150 190.600 103.410 190.920 ;
        RECT 103.150 189.920 103.410 190.240 ;
        RECT 103.210 187.180 103.350 189.920 ;
        RECT 103.150 186.860 103.410 187.180 ;
        RECT 101.130 185.645 102.670 186.015 ;
        RECT 100.390 184.480 100.650 184.800 ;
        RECT 100.390 182.100 100.650 182.420 ;
        RECT 97.170 179.040 97.430 179.360 ;
        RECT 97.620 179.185 97.900 179.555 ;
        RECT 99.930 179.380 100.190 179.700 ;
        RECT 100.450 179.360 100.590 182.100 ;
        RECT 102.680 181.905 102.960 182.275 ;
        RECT 102.750 181.740 102.890 181.905 ;
        RECT 102.690 181.420 102.950 181.740 ;
        RECT 101.130 180.205 102.670 180.575 ;
        RECT 103.210 179.360 103.350 186.860 ;
        RECT 103.670 182.760 103.810 191.960 ;
        RECT 104.990 191.620 105.250 191.940 ;
        RECT 104.070 189.580 104.330 189.900 ;
        RECT 104.130 185.480 104.270 189.580 ;
        RECT 104.530 188.900 104.790 189.220 ;
        RECT 104.590 187.520 104.730 188.900 ;
        RECT 105.050 188.200 105.190 191.620 ;
        RECT 105.450 189.920 105.710 190.240 ;
        RECT 104.990 187.880 105.250 188.200 ;
        RECT 104.530 187.200 104.790 187.520 ;
        RECT 104.530 186.180 104.790 186.500 ;
        RECT 104.070 185.160 104.330 185.480 ;
        RECT 103.610 182.440 103.870 182.760 ;
        RECT 104.070 181.420 104.330 181.740 ;
        RECT 104.130 180.040 104.270 181.420 ;
        RECT 104.590 180.040 104.730 186.180 ;
        RECT 104.070 179.720 104.330 180.040 ;
        RECT 104.530 179.720 104.790 180.040 ;
        RECT 100.390 179.040 100.650 179.360 ;
        RECT 103.150 179.040 103.410 179.360 ;
        RECT 105.510 178.680 105.650 189.920 ;
        RECT 105.970 182.080 106.110 191.960 ;
        RECT 106.370 188.900 106.630 189.220 ;
        RECT 106.430 184.800 106.570 188.900 ;
        RECT 106.370 184.480 106.630 184.800 ;
        RECT 106.890 183.780 107.030 192.300 ;
        RECT 107.290 189.580 107.550 189.900 ;
        RECT 107.350 186.500 107.490 189.580 ;
        RECT 107.915 188.365 109.455 188.735 ;
        RECT 107.290 186.180 107.550 186.500 ;
        RECT 106.830 183.460 107.090 183.780 ;
        RECT 105.910 181.760 106.170 182.080 ;
        RECT 106.890 181.740 107.030 183.460 ;
        RECT 107.915 182.925 109.455 183.295 ;
        RECT 109.650 182.760 109.790 195.020 ;
        RECT 110.110 192.620 110.250 195.700 ;
        RECT 110.570 195.680 110.710 197.060 ;
        RECT 110.510 195.360 110.770 195.680 ;
        RECT 110.510 194.340 110.770 194.660 ;
        RECT 110.050 192.300 110.310 192.620 ;
        RECT 110.570 190.580 110.710 194.340 ;
        RECT 111.030 190.920 111.170 200.460 ;
        RECT 111.430 198.420 111.690 198.740 ;
        RECT 111.490 190.920 111.630 198.420 ;
        RECT 113.790 196.020 113.930 203.180 ;
        RECT 113.730 195.700 113.990 196.020 ;
        RECT 112.350 195.020 112.610 195.340 ;
        RECT 110.970 190.600 111.230 190.920 ;
        RECT 111.430 190.600 111.690 190.920 ;
        RECT 110.510 190.260 110.770 190.580 ;
        RECT 107.750 182.440 108.010 182.760 ;
        RECT 109.590 182.440 109.850 182.760 ;
        RECT 106.830 181.420 107.090 181.740 ;
        RECT 105.910 180.740 106.170 181.060 ;
        RECT 105.970 179.360 106.110 180.740 ;
        RECT 107.810 179.360 107.950 182.440 ;
        RECT 110.050 181.080 110.310 181.400 ;
        RECT 109.590 179.380 109.850 179.700 ;
        RECT 105.910 179.040 106.170 179.360 ;
        RECT 107.750 179.040 108.010 179.360 ;
        RECT 105.450 178.360 105.710 178.680 ;
        RECT 67.205 177.485 68.745 177.855 ;
        RECT 80.775 177.485 82.315 177.855 ;
        RECT 94.345 177.485 95.885 177.855 ;
        RECT 73.990 174.765 75.530 175.135 ;
        RECT 87.560 174.765 89.100 175.135 ;
        RECT 101.130 174.765 102.670 175.135 ;
        RECT 105.970 173.920 106.110 179.040 ;
        RECT 107.915 177.485 109.455 177.855 ;
        RECT 109.650 176.980 109.790 179.380 ;
        RECT 110.110 177.320 110.250 181.080 ;
        RECT 110.050 177.000 110.310 177.320 ;
        RECT 109.590 176.660 109.850 176.980 ;
        RECT 110.110 174.260 110.250 177.000 ;
        RECT 110.570 176.300 110.710 190.260 ;
        RECT 112.410 187.520 112.550 195.020 ;
        RECT 113.270 192.300 113.530 192.620 ;
        RECT 113.330 191.940 113.470 192.300 ;
        RECT 113.270 191.620 113.530 191.940 ;
        RECT 113.330 189.560 113.470 191.620 ;
        RECT 114.250 189.900 114.390 207.180 ;
        RECT 114.700 201.965 116.240 202.335 ;
        RECT 114.700 196.525 116.240 196.895 ;
        RECT 114.700 191.085 116.240 191.455 ;
        RECT 114.190 189.580 114.450 189.900 ;
        RECT 113.270 189.240 113.530 189.560 ;
        RECT 112.350 187.200 112.610 187.520 ;
        RECT 110.970 186.860 111.230 187.180 ;
        RECT 111.030 178.680 111.170 186.860 ;
        RECT 111.890 186.180 112.150 186.500 ;
        RECT 111.430 178.700 111.690 179.020 ;
        RECT 110.970 178.360 111.230 178.680 ;
        RECT 111.490 177.320 111.630 178.700 ;
        RECT 111.430 177.000 111.690 177.320 ;
        RECT 110.510 175.980 110.770 176.300 ;
        RECT 110.050 173.940 110.310 174.260 ;
        RECT 111.950 173.920 112.090 186.180 ;
        RECT 112.410 185.480 112.550 187.200 ;
        RECT 112.350 185.160 112.610 185.480 ;
        RECT 112.410 182.160 112.550 185.160 ;
        RECT 112.410 182.020 113.010 182.160 ;
        RECT 112.350 181.080 112.610 181.400 ;
        RECT 112.410 174.600 112.550 181.080 ;
        RECT 112.870 180.040 113.010 182.020 ;
        RECT 112.810 179.720 113.070 180.040 ;
        RECT 113.330 175.960 113.470 189.240 ;
        RECT 114.700 185.645 116.240 186.015 ;
        RECT 114.700 180.205 116.240 180.575 ;
        RECT 113.270 175.640 113.530 175.960 ;
        RECT 114.700 174.765 116.240 175.135 ;
        RECT 112.350 174.280 112.610 174.600 ;
        RECT 105.910 173.600 106.170 173.920 ;
        RECT 111.890 173.600 112.150 173.920 ;
        RECT 67.205 172.045 68.745 172.415 ;
        RECT 80.775 172.045 82.315 172.415 ;
        RECT 94.345 172.045 95.885 172.415 ;
        RECT 107.915 172.045 109.455 172.415 ;
        RECT 73.990 169.325 75.530 169.695 ;
        RECT 87.560 169.325 89.100 169.695 ;
        RECT 101.130 169.325 102.670 169.695 ;
        RECT 114.700 169.325 116.240 169.695 ;
        RECT 67.205 166.605 68.745 166.975 ;
        RECT 80.775 166.605 82.315 166.975 ;
        RECT 94.345 166.605 95.885 166.975 ;
        RECT 107.915 166.605 109.455 166.975 ;
        RECT 73.990 163.885 75.530 164.255 ;
        RECT 87.560 163.885 89.100 164.255 ;
        RECT 101.130 163.885 102.670 164.255 ;
        RECT 114.700 163.885 116.240 164.255 ;
        RECT 67.205 161.165 68.745 161.535 ;
        RECT 80.775 161.165 82.315 161.535 ;
        RECT 94.345 161.165 95.885 161.535 ;
        RECT 107.915 161.165 109.455 161.535 ;
        RECT 73.990 158.445 75.530 158.815 ;
        RECT 87.560 158.445 89.100 158.815 ;
        RECT 101.130 158.445 102.670 158.815 ;
        RECT 114.700 158.445 116.240 158.815 ;
        RECT 67.205 155.725 68.745 156.095 ;
        RECT 80.775 155.725 82.315 156.095 ;
        RECT 94.345 155.725 95.885 156.095 ;
        RECT 107.915 155.725 109.455 156.095 ;
        RECT 73.990 153.005 75.530 153.375 ;
        RECT 87.560 153.005 89.100 153.375 ;
        RECT 101.130 153.005 102.670 153.375 ;
        RECT 114.700 153.005 116.240 153.375 ;
        RECT 102.780 89.445 103.805 91.400 ;
        RECT 102.760 88.470 103.825 89.445 ;
        RECT 102.780 88.445 103.805 88.470 ;
        RECT 127.110 87.575 127.790 89.410 ;
        RECT 90.275 83.250 91.725 83.270 ;
        RECT 90.250 81.750 95.280 83.250 ;
        RECT 90.275 81.730 91.725 81.750 ;
        RECT 147.090 79.605 148.190 83.150 ;
        RECT 147.070 78.555 148.210 79.605 ;
        RECT 147.090 78.530 148.190 78.555 ;
        RECT 111.765 69.245 112.955 69.275 ;
        RECT 111.765 68.055 114.840 69.245 ;
        RECT 111.765 68.025 112.955 68.055 ;
        RECT 107.760 67.730 108.480 67.775 ;
        RECT 112.490 67.730 113.210 67.760 ;
        RECT 107.760 67.010 113.210 67.730 ;
        RECT 107.760 66.965 108.480 67.010 ;
        RECT 112.490 66.980 113.210 67.010 ;
        RECT 144.750 49.475 146.470 49.500 ;
        RECT 144.750 48.605 146.490 49.475 ;
        RECT 144.750 48.580 146.470 48.605 ;
        RECT 66.775 45.250 68.225 45.270 ;
        RECT 98.970 45.250 112.970 45.260 ;
        RECT 66.750 43.760 112.970 45.250 ;
        RECT 66.750 43.750 99.710 43.760 ;
        RECT 66.775 43.730 68.225 43.750 ;
        RECT 140.640 43.460 141.490 43.660 ;
        RECT 134.750 43.410 136.530 43.450 ;
        RECT 134.740 43.160 139.390 43.410 ;
        RECT 134.750 42.860 139.390 43.160 ;
        RECT 140.640 43.060 143.940 43.460 ;
        RECT 134.750 42.820 139.340 42.860 ;
        RECT 129.890 40.910 130.740 41.260 ;
        RECT 129.790 40.860 130.740 40.910 ;
        RECT 132.040 40.860 132.940 40.910 ;
        RECT 129.740 40.560 133.190 40.860 ;
        RECT 129.790 40.510 130.740 40.560 ;
        RECT 132.040 40.510 132.940 40.560 ;
        RECT 129.890 36.310 130.740 40.510 ;
        RECT 134.750 38.600 136.530 42.820 ;
        RECT 138.340 42.810 139.340 42.820 ;
        RECT 140.640 41.860 141.490 43.060 ;
        RECT 142.940 42.260 149.340 42.660 ;
        RECT 140.640 41.460 143.940 41.860 ;
        RECT 140.640 40.910 141.490 41.460 ;
        RECT 144.740 41.010 149.340 42.260 ;
        RECT 138.440 40.560 141.490 40.910 ;
        RECT 142.940 40.710 149.340 41.010 ;
        RECT 138.440 40.510 139.340 40.560 ;
        RECT 140.640 40.310 141.490 40.560 ;
        RECT 140.640 39.910 143.940 40.310 ;
        RECT 140.640 38.710 141.490 39.910 ;
        RECT 144.790 39.460 149.340 40.710 ;
        RECT 142.940 39.160 148.040 39.460 ;
        RECT 144.740 39.010 148.040 39.160 ;
        RECT 138.340 38.600 139.340 38.610 ;
        RECT 134.750 38.220 139.390 38.600 ;
        RECT 140.640 38.310 143.940 38.710 ;
        RECT 129.790 36.260 130.740 36.310 ;
        RECT 132.040 36.260 132.940 36.310 ;
        RECT 129.740 35.960 133.190 36.260 ;
        RECT 129.790 35.910 130.740 35.960 ;
        RECT 132.040 35.910 132.940 35.960 ;
        RECT 125.290 32.710 126.090 32.760 ;
        RECT 125.290 32.060 128.440 32.710 ;
        RECT 125.290 28.160 126.090 32.060 ;
        RECT 129.890 31.760 130.740 35.910 ;
        RECT 134.750 34.000 136.530 38.220 ;
        RECT 138.340 38.210 139.340 38.220 ;
        RECT 140.640 37.110 141.490 38.310 ;
        RECT 144.740 37.860 146.040 39.010 ;
        RECT 142.940 37.560 146.040 37.860 ;
        RECT 140.640 36.710 143.890 37.110 ;
        RECT 140.640 36.360 141.490 36.710 ;
        RECT 138.440 35.960 141.490 36.360 ;
        RECT 144.740 36.310 146.040 37.560 ;
        RECT 146.890 36.710 149.340 37.260 ;
        RECT 142.940 35.960 146.040 36.310 ;
        RECT 138.440 35.910 139.340 35.960 ;
        RECT 140.640 35.560 141.490 35.960 ;
        RECT 140.640 35.160 143.890 35.560 ;
        RECT 138.340 34.000 139.340 34.010 ;
        RECT 134.750 33.620 139.340 34.000 ;
        RECT 129.790 31.710 130.740 31.760 ;
        RECT 132.040 31.710 132.940 31.760 ;
        RECT 129.740 31.410 133.190 31.710 ;
        RECT 129.790 31.360 130.740 31.410 ;
        RECT 132.040 31.360 132.940 31.410 ;
        RECT 129.890 31.210 130.740 31.360 ;
        RECT 134.750 30.120 136.530 33.620 ;
        RECT 138.340 33.610 139.340 33.620 ;
        RECT 140.640 33.960 141.490 35.160 ;
        RECT 144.740 34.960 146.040 35.960 ;
        RECT 144.740 34.710 148.040 34.960 ;
        RECT 142.940 34.410 148.040 34.710 ;
        RECT 142.940 34.360 146.040 34.410 ;
        RECT 140.640 33.560 143.940 33.960 ;
        RECT 140.640 32.410 141.490 33.560 ;
        RECT 144.740 33.160 146.040 34.360 ;
        RECT 142.940 32.810 146.040 33.160 ;
        RECT 140.640 32.010 143.940 32.410 ;
        RECT 140.640 31.760 141.490 32.010 ;
        RECT 138.440 31.410 141.490 31.760 ;
        RECT 144.740 31.560 146.040 32.810 ;
        RECT 148.590 32.710 149.340 36.710 ;
        RECT 156.410 34.925 157.310 40.630 ;
        RECT 156.390 34.075 157.330 34.925 ;
        RECT 156.410 34.050 157.310 34.075 ;
        RECT 146.890 32.160 149.340 32.710 ;
        RECT 138.440 31.360 139.340 31.410 ;
        RECT 140.640 30.810 141.490 31.410 ;
        RECT 142.940 31.210 146.040 31.560 ;
        RECT 140.640 30.410 143.940 30.810 ;
        RECT 134.760 28.880 136.520 30.120 ;
        RECT 138.615 29.410 139.165 29.980 ;
        RECT 125.290 27.510 128.440 28.160 ;
        RECT 138.340 27.860 139.340 29.410 ;
        RECT 140.640 29.210 141.540 30.410 ;
        RECT 144.740 30.360 146.040 31.210 ;
        RECT 141.740 29.560 142.740 30.060 ;
        RECT 144.740 30.010 148.040 30.360 ;
        RECT 142.940 29.810 148.040 30.010 ;
        RECT 142.940 29.610 146.040 29.810 ;
        RECT 141.740 29.510 142.440 29.560 ;
        RECT 140.640 28.810 143.890 29.210 ;
        RECT 140.640 27.860 141.540 28.810 ;
        RECT 144.740 28.460 146.040 29.610 ;
        RECT 142.940 28.060 146.040 28.460 ;
        RECT 148.590 28.110 149.340 32.160 ;
        RECT 125.290 23.560 126.090 27.510 ;
        RECT 129.940 27.040 131.140 27.760 ;
        RECT 138.390 27.410 139.240 27.860 ;
        RECT 140.640 27.710 141.890 27.860 ;
        RECT 140.640 27.410 143.890 27.710 ;
        RECT 141.790 27.260 143.890 27.410 ;
        RECT 140.290 27.040 141.590 27.260 ;
        RECT 129.940 27.010 135.015 27.040 ;
        RECT 136.265 27.010 141.590 27.040 ;
        RECT 129.940 26.560 135.040 27.010 ;
        RECT 136.240 26.560 141.590 27.010 ;
        RECT 144.740 27.210 146.040 28.060 ;
        RECT 146.890 27.560 149.340 28.110 ;
        RECT 144.740 26.610 147.840 27.210 ;
        RECT 129.940 26.485 135.015 26.560 ;
        RECT 136.265 26.490 141.590 26.560 ;
        RECT 129.940 26.310 131.140 26.485 ;
        RECT 140.290 26.260 141.590 26.490 ;
        RECT 129.140 25.810 129.790 25.840 ;
        RECT 129.140 25.160 130.510 25.810 ;
        RECT 130.790 25.560 132.140 26.010 ;
        RECT 129.140 25.130 129.790 25.160 ;
        RECT 125.290 22.910 128.440 23.560 ;
        RECT 125.290 22.860 126.090 22.910 ;
        RECT 130.790 22.360 131.440 25.560 ;
        RECT 133.190 23.460 133.790 26.210 ;
        RECT 135.490 22.360 136.040 24.460 ;
        RECT 137.740 23.460 138.340 26.210 ;
        RECT 139.240 25.560 140.590 26.010 ;
        RECT 143.225 25.930 144.065 26.105 ;
        RECT 139.940 22.360 140.590 25.560 ;
        RECT 143.200 25.040 145.165 25.930 ;
        RECT 147.040 25.310 147.840 26.610 ;
        RECT 143.225 24.865 144.065 25.040 ;
        RECT 148.590 23.560 149.340 27.560 ;
        RECT 146.890 23.010 149.340 23.560 ;
        RECT 130.790 21.460 140.590 22.360 ;
        RECT 150.940 14.860 152.140 22.155 ;
        RECT 150.910 13.660 152.170 14.860 ;
      LAYER via2 ;
        RECT 94.390 218.270 94.670 218.550 ;
        RECT 87.960 217.060 88.240 217.340 ;
        RECT 81.550 215.790 81.830 216.070 ;
        RECT 75.090 214.200 75.370 214.480 ;
        RECT 62.080 212.740 62.360 213.020 ;
        RECT 68.630 212.850 68.910 213.130 ;
        RECT 107.340 215.520 107.620 215.800 ;
        RECT 100.850 213.910 101.130 214.190 ;
        RECT 67.235 204.730 67.515 205.010 ;
        RECT 67.635 204.730 67.915 205.010 ;
        RECT 68.035 204.730 68.315 205.010 ;
        RECT 68.435 204.730 68.715 205.010 ;
        RECT 64.500 198.270 64.780 198.550 ;
        RECT 67.235 199.290 67.515 199.570 ;
        RECT 67.635 199.290 67.915 199.570 ;
        RECT 68.035 199.290 68.315 199.570 ;
        RECT 68.435 199.290 68.715 199.570 ;
        RECT 74.020 207.450 74.300 207.730 ;
        RECT 74.420 207.450 74.700 207.730 ;
        RECT 74.820 207.450 75.100 207.730 ;
        RECT 75.220 207.450 75.500 207.730 ;
        RECT 113.710 211.030 113.990 211.310 ;
        RECT 87.590 207.450 87.870 207.730 ;
        RECT 87.990 207.450 88.270 207.730 ;
        RECT 88.390 207.450 88.670 207.730 ;
        RECT 88.790 207.450 89.070 207.730 ;
        RECT 67.235 193.850 67.515 194.130 ;
        RECT 67.635 193.850 67.915 194.130 ;
        RECT 68.035 193.850 68.315 194.130 ;
        RECT 68.435 193.850 68.715 194.130 ;
        RECT 80.805 204.730 81.085 205.010 ;
        RECT 81.205 204.730 81.485 205.010 ;
        RECT 81.605 204.730 81.885 205.010 ;
        RECT 82.005 204.730 82.285 205.010 ;
        RECT 74.020 202.010 74.300 202.290 ;
        RECT 74.420 202.010 74.700 202.290 ;
        RECT 74.820 202.010 75.100 202.290 ;
        RECT 75.220 202.010 75.500 202.290 ;
        RECT 75.080 198.270 75.360 198.550 ;
        RECT 73.700 197.590 73.980 197.870 ;
        RECT 74.020 196.570 74.300 196.850 ;
        RECT 74.420 196.570 74.700 196.850 ;
        RECT 74.820 196.570 75.100 196.850 ;
        RECT 75.220 196.570 75.500 196.850 ;
        RECT 74.020 191.130 74.300 191.410 ;
        RECT 74.420 191.130 74.700 191.410 ;
        RECT 74.820 191.130 75.100 191.410 ;
        RECT 75.220 191.130 75.500 191.410 ;
        RECT 67.235 188.410 67.515 188.690 ;
        RECT 67.635 188.410 67.915 188.690 ;
        RECT 68.035 188.410 68.315 188.690 ;
        RECT 68.435 188.410 68.715 188.690 ;
        RECT 67.235 182.970 67.515 183.250 ;
        RECT 67.635 182.970 67.915 183.250 ;
        RECT 68.035 182.970 68.315 183.250 ;
        RECT 68.435 182.970 68.715 183.250 ;
        RECT 74.020 185.690 74.300 185.970 ;
        RECT 74.420 185.690 74.700 185.970 ;
        RECT 74.820 185.690 75.100 185.970 ;
        RECT 75.220 185.690 75.500 185.970 ;
        RECT 80.805 199.290 81.085 199.570 ;
        RECT 81.205 199.290 81.485 199.570 ;
        RECT 81.605 199.290 81.885 199.570 ;
        RECT 82.005 199.290 82.285 199.570 ;
        RECT 80.805 193.850 81.085 194.130 ;
        RECT 81.205 193.850 81.485 194.130 ;
        RECT 81.605 193.850 81.885 194.130 ;
        RECT 82.005 193.850 82.285 194.130 ;
        RECT 85.660 200.310 85.940 200.590 ;
        RECT 84.740 197.590 85.020 197.870 ;
        RECT 87.590 202.010 87.870 202.290 ;
        RECT 87.990 202.010 88.270 202.290 ;
        RECT 88.390 202.010 88.670 202.290 ;
        RECT 88.790 202.010 89.070 202.290 ;
        RECT 94.375 204.730 94.655 205.010 ;
        RECT 94.775 204.730 95.055 205.010 ;
        RECT 95.175 204.730 95.455 205.010 ;
        RECT 95.575 204.730 95.855 205.010 ;
        RECT 101.160 207.450 101.440 207.730 ;
        RECT 101.560 207.450 101.840 207.730 ;
        RECT 101.960 207.450 102.240 207.730 ;
        RECT 102.360 207.450 102.640 207.730 ;
        RECT 94.375 199.290 94.655 199.570 ;
        RECT 94.775 199.290 95.055 199.570 ;
        RECT 95.175 199.290 95.455 199.570 ;
        RECT 95.575 199.290 95.855 199.570 ;
        RECT 92.560 197.590 92.840 197.870 ;
        RECT 94.860 197.590 95.140 197.870 ;
        RECT 87.590 196.570 87.870 196.850 ;
        RECT 87.990 196.570 88.270 196.850 ;
        RECT 88.390 196.570 88.670 196.850 ;
        RECT 88.790 196.570 89.070 196.850 ;
        RECT 80.805 188.410 81.085 188.690 ;
        RECT 81.205 188.410 81.485 188.690 ;
        RECT 81.605 188.410 81.885 188.690 ;
        RECT 82.005 188.410 82.285 188.690 ;
        RECT 80.805 182.970 81.085 183.250 ;
        RECT 81.205 182.970 81.485 183.250 ;
        RECT 81.605 182.970 81.885 183.250 ;
        RECT 82.005 182.970 82.285 183.250 ;
        RECT 87.590 191.130 87.870 191.410 ;
        RECT 87.990 191.130 88.270 191.410 ;
        RECT 88.390 191.130 88.670 191.410 ;
        RECT 88.790 191.130 89.070 191.410 ;
        RECT 87.590 185.690 87.870 185.970 ;
        RECT 87.990 185.690 88.270 185.970 ;
        RECT 88.390 185.690 88.670 185.970 ;
        RECT 88.790 185.690 89.070 185.970 ;
        RECT 94.375 193.850 94.655 194.130 ;
        RECT 94.775 193.850 95.055 194.130 ;
        RECT 95.175 193.850 95.455 194.130 ;
        RECT 95.575 193.850 95.855 194.130 ;
        RECT 94.375 188.410 94.655 188.690 ;
        RECT 94.775 188.410 95.055 188.690 ;
        RECT 95.175 188.410 95.455 188.690 ;
        RECT 95.575 188.410 95.855 188.690 ;
        RECT 94.375 182.970 94.655 183.250 ;
        RECT 94.775 182.970 95.055 183.250 ;
        RECT 95.175 182.970 95.455 183.250 ;
        RECT 95.575 182.970 95.855 183.250 ;
        RECT 74.020 180.250 74.300 180.530 ;
        RECT 74.420 180.250 74.700 180.530 ;
        RECT 74.820 180.250 75.100 180.530 ;
        RECT 75.220 180.250 75.500 180.530 ;
        RECT 87.590 180.250 87.870 180.530 ;
        RECT 87.990 180.250 88.270 180.530 ;
        RECT 88.390 180.250 88.670 180.530 ;
        RECT 88.790 180.250 89.070 180.530 ;
        RECT 101.160 202.010 101.440 202.290 ;
        RECT 101.560 202.010 101.840 202.290 ;
        RECT 101.960 202.010 102.240 202.290 ;
        RECT 102.360 202.010 102.640 202.290 ;
        RECT 104.980 198.270 105.260 198.550 ;
        RECT 114.730 207.450 115.010 207.730 ;
        RECT 115.130 207.450 115.410 207.730 ;
        RECT 115.530 207.450 115.810 207.730 ;
        RECT 115.930 207.450 116.210 207.730 ;
        RECT 107.945 204.730 108.225 205.010 ;
        RECT 108.345 204.730 108.625 205.010 ;
        RECT 108.745 204.730 109.025 205.010 ;
        RECT 109.145 204.730 109.425 205.010 ;
        RECT 107.280 200.310 107.560 200.590 ;
        RECT 101.760 197.590 102.040 197.870 ;
        RECT 101.160 196.570 101.440 196.850 ;
        RECT 101.560 196.570 101.840 196.850 ;
        RECT 101.960 196.570 102.240 196.850 ;
        RECT 102.360 196.570 102.640 196.850 ;
        RECT 107.945 199.290 108.225 199.570 ;
        RECT 108.345 199.290 108.625 199.570 ;
        RECT 108.745 199.290 109.025 199.570 ;
        RECT 109.145 199.290 109.425 199.570 ;
        RECT 107.945 193.850 108.225 194.130 ;
        RECT 108.345 193.850 108.625 194.130 ;
        RECT 108.745 193.850 109.025 194.130 ;
        RECT 109.145 193.850 109.425 194.130 ;
        RECT 101.160 191.130 101.440 191.410 ;
        RECT 101.560 191.130 101.840 191.410 ;
        RECT 101.960 191.130 102.240 191.410 ;
        RECT 102.360 191.130 102.640 191.410 ;
        RECT 101.160 185.690 101.440 185.970 ;
        RECT 101.560 185.690 101.840 185.970 ;
        RECT 101.960 185.690 102.240 185.970 ;
        RECT 102.360 185.690 102.640 185.970 ;
        RECT 97.620 179.230 97.900 179.510 ;
        RECT 102.680 181.950 102.960 182.230 ;
        RECT 101.160 180.250 101.440 180.530 ;
        RECT 101.560 180.250 101.840 180.530 ;
        RECT 101.960 180.250 102.240 180.530 ;
        RECT 102.360 180.250 102.640 180.530 ;
        RECT 107.945 188.410 108.225 188.690 ;
        RECT 108.345 188.410 108.625 188.690 ;
        RECT 108.745 188.410 109.025 188.690 ;
        RECT 109.145 188.410 109.425 188.690 ;
        RECT 107.945 182.970 108.225 183.250 ;
        RECT 108.345 182.970 108.625 183.250 ;
        RECT 108.745 182.970 109.025 183.250 ;
        RECT 109.145 182.970 109.425 183.250 ;
        RECT 67.235 177.530 67.515 177.810 ;
        RECT 67.635 177.530 67.915 177.810 ;
        RECT 68.035 177.530 68.315 177.810 ;
        RECT 68.435 177.530 68.715 177.810 ;
        RECT 80.805 177.530 81.085 177.810 ;
        RECT 81.205 177.530 81.485 177.810 ;
        RECT 81.605 177.530 81.885 177.810 ;
        RECT 82.005 177.530 82.285 177.810 ;
        RECT 94.375 177.530 94.655 177.810 ;
        RECT 94.775 177.530 95.055 177.810 ;
        RECT 95.175 177.530 95.455 177.810 ;
        RECT 95.575 177.530 95.855 177.810 ;
        RECT 74.020 174.810 74.300 175.090 ;
        RECT 74.420 174.810 74.700 175.090 ;
        RECT 74.820 174.810 75.100 175.090 ;
        RECT 75.220 174.810 75.500 175.090 ;
        RECT 87.590 174.810 87.870 175.090 ;
        RECT 87.990 174.810 88.270 175.090 ;
        RECT 88.390 174.810 88.670 175.090 ;
        RECT 88.790 174.810 89.070 175.090 ;
        RECT 101.160 174.810 101.440 175.090 ;
        RECT 101.560 174.810 101.840 175.090 ;
        RECT 101.960 174.810 102.240 175.090 ;
        RECT 102.360 174.810 102.640 175.090 ;
        RECT 107.945 177.530 108.225 177.810 ;
        RECT 108.345 177.530 108.625 177.810 ;
        RECT 108.745 177.530 109.025 177.810 ;
        RECT 109.145 177.530 109.425 177.810 ;
        RECT 114.730 202.010 115.010 202.290 ;
        RECT 115.130 202.010 115.410 202.290 ;
        RECT 115.530 202.010 115.810 202.290 ;
        RECT 115.930 202.010 116.210 202.290 ;
        RECT 114.730 196.570 115.010 196.850 ;
        RECT 115.130 196.570 115.410 196.850 ;
        RECT 115.530 196.570 115.810 196.850 ;
        RECT 115.930 196.570 116.210 196.850 ;
        RECT 114.730 191.130 115.010 191.410 ;
        RECT 115.130 191.130 115.410 191.410 ;
        RECT 115.530 191.130 115.810 191.410 ;
        RECT 115.930 191.130 116.210 191.410 ;
        RECT 114.730 185.690 115.010 185.970 ;
        RECT 115.130 185.690 115.410 185.970 ;
        RECT 115.530 185.690 115.810 185.970 ;
        RECT 115.930 185.690 116.210 185.970 ;
        RECT 114.730 180.250 115.010 180.530 ;
        RECT 115.130 180.250 115.410 180.530 ;
        RECT 115.530 180.250 115.810 180.530 ;
        RECT 115.930 180.250 116.210 180.530 ;
        RECT 114.730 174.810 115.010 175.090 ;
        RECT 115.130 174.810 115.410 175.090 ;
        RECT 115.530 174.810 115.810 175.090 ;
        RECT 115.930 174.810 116.210 175.090 ;
        RECT 67.235 172.090 67.515 172.370 ;
        RECT 67.635 172.090 67.915 172.370 ;
        RECT 68.035 172.090 68.315 172.370 ;
        RECT 68.435 172.090 68.715 172.370 ;
        RECT 80.805 172.090 81.085 172.370 ;
        RECT 81.205 172.090 81.485 172.370 ;
        RECT 81.605 172.090 81.885 172.370 ;
        RECT 82.005 172.090 82.285 172.370 ;
        RECT 94.375 172.090 94.655 172.370 ;
        RECT 94.775 172.090 95.055 172.370 ;
        RECT 95.175 172.090 95.455 172.370 ;
        RECT 95.575 172.090 95.855 172.370 ;
        RECT 107.945 172.090 108.225 172.370 ;
        RECT 108.345 172.090 108.625 172.370 ;
        RECT 108.745 172.090 109.025 172.370 ;
        RECT 109.145 172.090 109.425 172.370 ;
        RECT 74.020 169.370 74.300 169.650 ;
        RECT 74.420 169.370 74.700 169.650 ;
        RECT 74.820 169.370 75.100 169.650 ;
        RECT 75.220 169.370 75.500 169.650 ;
        RECT 87.590 169.370 87.870 169.650 ;
        RECT 87.990 169.370 88.270 169.650 ;
        RECT 88.390 169.370 88.670 169.650 ;
        RECT 88.790 169.370 89.070 169.650 ;
        RECT 101.160 169.370 101.440 169.650 ;
        RECT 101.560 169.370 101.840 169.650 ;
        RECT 101.960 169.370 102.240 169.650 ;
        RECT 102.360 169.370 102.640 169.650 ;
        RECT 114.730 169.370 115.010 169.650 ;
        RECT 115.130 169.370 115.410 169.650 ;
        RECT 115.530 169.370 115.810 169.650 ;
        RECT 115.930 169.370 116.210 169.650 ;
        RECT 67.235 166.650 67.515 166.930 ;
        RECT 67.635 166.650 67.915 166.930 ;
        RECT 68.035 166.650 68.315 166.930 ;
        RECT 68.435 166.650 68.715 166.930 ;
        RECT 80.805 166.650 81.085 166.930 ;
        RECT 81.205 166.650 81.485 166.930 ;
        RECT 81.605 166.650 81.885 166.930 ;
        RECT 82.005 166.650 82.285 166.930 ;
        RECT 94.375 166.650 94.655 166.930 ;
        RECT 94.775 166.650 95.055 166.930 ;
        RECT 95.175 166.650 95.455 166.930 ;
        RECT 95.575 166.650 95.855 166.930 ;
        RECT 107.945 166.650 108.225 166.930 ;
        RECT 108.345 166.650 108.625 166.930 ;
        RECT 108.745 166.650 109.025 166.930 ;
        RECT 109.145 166.650 109.425 166.930 ;
        RECT 74.020 163.930 74.300 164.210 ;
        RECT 74.420 163.930 74.700 164.210 ;
        RECT 74.820 163.930 75.100 164.210 ;
        RECT 75.220 163.930 75.500 164.210 ;
        RECT 87.590 163.930 87.870 164.210 ;
        RECT 87.990 163.930 88.270 164.210 ;
        RECT 88.390 163.930 88.670 164.210 ;
        RECT 88.790 163.930 89.070 164.210 ;
        RECT 101.160 163.930 101.440 164.210 ;
        RECT 101.560 163.930 101.840 164.210 ;
        RECT 101.960 163.930 102.240 164.210 ;
        RECT 102.360 163.930 102.640 164.210 ;
        RECT 114.730 163.930 115.010 164.210 ;
        RECT 115.130 163.930 115.410 164.210 ;
        RECT 115.530 163.930 115.810 164.210 ;
        RECT 115.930 163.930 116.210 164.210 ;
        RECT 67.235 161.210 67.515 161.490 ;
        RECT 67.635 161.210 67.915 161.490 ;
        RECT 68.035 161.210 68.315 161.490 ;
        RECT 68.435 161.210 68.715 161.490 ;
        RECT 80.805 161.210 81.085 161.490 ;
        RECT 81.205 161.210 81.485 161.490 ;
        RECT 81.605 161.210 81.885 161.490 ;
        RECT 82.005 161.210 82.285 161.490 ;
        RECT 94.375 161.210 94.655 161.490 ;
        RECT 94.775 161.210 95.055 161.490 ;
        RECT 95.175 161.210 95.455 161.490 ;
        RECT 95.575 161.210 95.855 161.490 ;
        RECT 107.945 161.210 108.225 161.490 ;
        RECT 108.345 161.210 108.625 161.490 ;
        RECT 108.745 161.210 109.025 161.490 ;
        RECT 109.145 161.210 109.425 161.490 ;
        RECT 74.020 158.490 74.300 158.770 ;
        RECT 74.420 158.490 74.700 158.770 ;
        RECT 74.820 158.490 75.100 158.770 ;
        RECT 75.220 158.490 75.500 158.770 ;
        RECT 87.590 158.490 87.870 158.770 ;
        RECT 87.990 158.490 88.270 158.770 ;
        RECT 88.390 158.490 88.670 158.770 ;
        RECT 88.790 158.490 89.070 158.770 ;
        RECT 101.160 158.490 101.440 158.770 ;
        RECT 101.560 158.490 101.840 158.770 ;
        RECT 101.960 158.490 102.240 158.770 ;
        RECT 102.360 158.490 102.640 158.770 ;
        RECT 114.730 158.490 115.010 158.770 ;
        RECT 115.130 158.490 115.410 158.770 ;
        RECT 115.530 158.490 115.810 158.770 ;
        RECT 115.930 158.490 116.210 158.770 ;
        RECT 67.235 155.770 67.515 156.050 ;
        RECT 67.635 155.770 67.915 156.050 ;
        RECT 68.035 155.770 68.315 156.050 ;
        RECT 68.435 155.770 68.715 156.050 ;
        RECT 80.805 155.770 81.085 156.050 ;
        RECT 81.205 155.770 81.485 156.050 ;
        RECT 81.605 155.770 81.885 156.050 ;
        RECT 82.005 155.770 82.285 156.050 ;
        RECT 94.375 155.770 94.655 156.050 ;
        RECT 94.775 155.770 95.055 156.050 ;
        RECT 95.175 155.770 95.455 156.050 ;
        RECT 95.575 155.770 95.855 156.050 ;
        RECT 107.945 155.770 108.225 156.050 ;
        RECT 108.345 155.770 108.625 156.050 ;
        RECT 108.745 155.770 109.025 156.050 ;
        RECT 109.145 155.770 109.425 156.050 ;
        RECT 74.020 153.050 74.300 153.330 ;
        RECT 74.420 153.050 74.700 153.330 ;
        RECT 74.820 153.050 75.100 153.330 ;
        RECT 75.220 153.050 75.500 153.330 ;
        RECT 87.590 153.050 87.870 153.330 ;
        RECT 87.990 153.050 88.270 153.330 ;
        RECT 88.390 153.050 88.670 153.330 ;
        RECT 88.790 153.050 89.070 153.330 ;
        RECT 101.160 153.050 101.440 153.330 ;
        RECT 101.560 153.050 101.840 153.330 ;
        RECT 101.960 153.050 102.240 153.330 ;
        RECT 102.360 153.050 102.640 153.330 ;
        RECT 114.730 153.050 115.010 153.330 ;
        RECT 115.130 153.050 115.410 153.330 ;
        RECT 115.530 153.050 115.810 153.330 ;
        RECT 115.930 153.050 116.210 153.330 ;
        RECT 102.805 88.470 103.780 89.445 ;
        RECT 127.110 87.620 127.790 88.300 ;
        RECT 90.275 81.775 91.725 83.225 ;
        RECT 147.115 78.555 148.165 79.605 ;
        RECT 113.605 68.055 114.795 69.245 ;
        RECT 145.575 48.605 146.445 49.475 ;
        RECT 66.775 43.775 68.225 45.225 ;
        RECT 156.435 34.075 157.285 34.925 ;
        RECT 134.990 29.360 136.440 30.160 ;
        RECT 138.615 29.385 139.165 29.935 ;
        RECT 130.040 27.110 130.640 27.660 ;
        RECT 140.890 26.460 141.490 27.160 ;
        RECT 129.815 25.160 130.465 25.810 ;
        RECT 143.225 24.910 144.065 26.060 ;
        RECT 150.940 20.910 152.140 22.110 ;
      LAYER met3 ;
        RECT 107.290 220.690 107.670 221.010 ;
        RECT 100.800 219.420 101.180 219.740 ;
        RECT 81.260 218.560 81.580 218.600 ;
        RECT 94.365 218.560 94.695 218.575 ;
        RECT 81.260 218.260 94.695 218.560 ;
        RECT 81.260 218.220 81.580 218.260 ;
        RECT 94.365 218.245 94.695 218.260 ;
        RECT 77.580 217.350 77.900 217.390 ;
        RECT 87.935 217.350 88.265 217.365 ;
        RECT 77.580 217.050 88.265 217.350 ;
        RECT 77.580 217.010 77.900 217.050 ;
        RECT 87.935 217.035 88.265 217.050 ;
        RECT 73.900 216.080 74.220 216.120 ;
        RECT 81.525 216.080 81.855 216.095 ;
        RECT 73.900 215.780 81.855 216.080 ;
        RECT 73.900 215.740 74.220 215.780 ;
        RECT 81.525 215.765 81.855 215.780 ;
        RECT 70.220 214.490 70.540 214.530 ;
        RECT 75.065 214.490 75.395 214.505 ;
        RECT 70.220 214.190 75.395 214.490 ;
        RECT 100.840 214.215 101.140 219.420 ;
        RECT 107.330 215.825 107.630 220.690 ;
        RECT 107.315 215.495 107.645 215.825 ;
        RECT 70.220 214.150 70.540 214.190 ;
        RECT 75.065 214.175 75.395 214.190 ;
        RECT 100.825 213.885 101.155 214.215 ;
        RECT 66.540 213.140 66.860 213.180 ;
        RECT 68.605 213.140 68.935 213.155 ;
        RECT 62.055 213.030 62.385 213.045 ;
        RECT 62.830 213.030 63.210 213.040 ;
        RECT 62.055 212.730 63.210 213.030 ;
        RECT 66.540 212.840 68.935 213.140 ;
        RECT 66.540 212.800 66.860 212.840 ;
        RECT 68.605 212.825 68.935 212.840 ;
        RECT 62.055 212.715 62.385 212.730 ;
        RECT 62.830 212.720 63.210 212.730 ;
        RECT 113.660 212.020 114.040 212.340 ;
        RECT 113.700 211.335 114.000 212.020 ;
        RECT 113.685 211.005 114.015 211.335 ;
        RECT 73.970 207.425 75.550 207.755 ;
        RECT 87.540 207.425 89.120 207.755 ;
        RECT 101.110 207.425 102.690 207.755 ;
        RECT 114.680 207.425 116.260 207.755 ;
        RECT 67.185 204.705 68.765 205.035 ;
        RECT 80.755 204.705 82.335 205.035 ;
        RECT 94.325 204.705 95.905 205.035 ;
        RECT 107.895 204.705 109.475 205.035 ;
        RECT 73.970 201.985 75.550 202.315 ;
        RECT 87.540 201.985 89.120 202.315 ;
        RECT 101.110 201.985 102.690 202.315 ;
        RECT 114.680 201.985 116.260 202.315 ;
        RECT 85.635 200.600 85.965 200.615 ;
        RECT 107.255 200.600 107.585 200.615 ;
        RECT 85.635 200.300 107.585 200.600 ;
        RECT 85.635 200.285 85.965 200.300 ;
        RECT 107.255 200.285 107.585 200.300 ;
        RECT 67.185 199.265 68.765 199.595 ;
        RECT 80.755 199.265 82.335 199.595 ;
        RECT 94.325 199.265 95.905 199.595 ;
        RECT 107.895 199.265 109.475 199.595 ;
        RECT 64.475 198.560 64.805 198.575 ;
        RECT 75.055 198.560 75.385 198.575 ;
        RECT 103.780 198.560 104.160 198.570 ;
        RECT 104.955 198.560 105.285 198.575 ;
        RECT 64.475 198.260 75.385 198.560 ;
        RECT 64.475 198.245 64.805 198.260 ;
        RECT 75.055 198.245 75.385 198.260 ;
        RECT 83.580 198.260 105.285 198.560 ;
        RECT 73.675 197.880 74.005 197.895 ;
        RECT 83.580 197.880 83.880 198.260 ;
        RECT 103.780 198.250 104.160 198.260 ;
        RECT 104.955 198.245 105.285 198.260 ;
        RECT 73.675 197.580 83.880 197.880 ;
        RECT 84.715 197.880 85.045 197.895 ;
        RECT 92.535 197.880 92.865 197.895 ;
        RECT 84.715 197.580 92.865 197.880 ;
        RECT 73.675 197.565 74.005 197.580 ;
        RECT 84.715 197.565 85.045 197.580 ;
        RECT 92.535 197.565 92.865 197.580 ;
        RECT 94.835 197.880 95.165 197.895 ;
        RECT 101.735 197.880 102.065 197.895 ;
        RECT 94.835 197.580 102.065 197.880 ;
        RECT 94.835 197.565 95.165 197.580 ;
        RECT 101.735 197.565 102.065 197.580 ;
        RECT 73.970 196.545 75.550 196.875 ;
        RECT 87.540 196.545 89.120 196.875 ;
        RECT 101.110 196.545 102.690 196.875 ;
        RECT 114.680 196.545 116.260 196.875 ;
        RECT 67.185 193.825 68.765 194.155 ;
        RECT 80.755 193.825 82.335 194.155 ;
        RECT 94.325 193.825 95.905 194.155 ;
        RECT 107.895 193.825 109.475 194.155 ;
        RECT 73.970 191.105 75.550 191.435 ;
        RECT 87.540 191.105 89.120 191.435 ;
        RECT 101.110 191.105 102.690 191.435 ;
        RECT 114.680 191.105 116.260 191.435 ;
        RECT 67.185 188.385 68.765 188.715 ;
        RECT 80.755 188.385 82.335 188.715 ;
        RECT 94.325 188.385 95.905 188.715 ;
        RECT 107.895 188.385 109.475 188.715 ;
        RECT 73.970 185.665 75.550 185.995 ;
        RECT 87.540 185.665 89.120 185.995 ;
        RECT 101.110 185.665 102.690 185.995 ;
        RECT 114.680 185.665 116.260 185.995 ;
        RECT 67.185 182.945 68.765 183.275 ;
        RECT 80.755 182.945 82.335 183.275 ;
        RECT 94.325 182.945 95.905 183.275 ;
        RECT 107.895 182.945 109.475 183.275 ;
        RECT 102.655 182.240 102.985 182.255 ;
        RECT 103.780 182.240 104.160 182.250 ;
        RECT 102.655 181.940 104.160 182.240 ;
        RECT 102.655 181.925 102.985 181.940 ;
        RECT 103.780 181.930 104.160 181.940 ;
        RECT 73.970 180.225 75.550 180.555 ;
        RECT 87.540 180.225 89.120 180.555 ;
        RECT 101.110 180.225 102.690 180.555 ;
        RECT 114.680 180.225 116.260 180.555 ;
        RECT 116.430 179.630 118.430 179.670 ;
        RECT 97.595 179.520 97.925 179.535 ;
        RECT 116.430 179.520 158.870 179.630 ;
        RECT 97.595 179.220 158.870 179.520 ;
        RECT 97.595 179.205 97.925 179.220 ;
        RECT 116.430 179.070 158.870 179.220 ;
        RECT 117.270 178.730 158.870 179.070 ;
        RECT 67.185 177.505 68.765 177.835 ;
        RECT 80.755 177.505 82.335 177.835 ;
        RECT 94.325 177.505 95.905 177.835 ;
        RECT 107.895 177.505 109.475 177.835 ;
        RECT 73.970 174.785 75.550 175.115 ;
        RECT 87.540 174.785 89.120 175.115 ;
        RECT 101.110 174.785 102.690 175.115 ;
        RECT 114.680 174.785 116.260 175.115 ;
        RECT 67.185 172.065 68.765 172.395 ;
        RECT 80.755 172.065 82.335 172.395 ;
        RECT 94.325 172.065 95.905 172.395 ;
        RECT 107.895 172.065 109.475 172.395 ;
        RECT 73.970 169.345 75.550 169.675 ;
        RECT 87.540 169.345 89.120 169.675 ;
        RECT 101.110 169.345 102.690 169.675 ;
        RECT 114.680 169.345 116.260 169.675 ;
        RECT 67.185 166.625 68.765 166.955 ;
        RECT 80.755 166.625 82.335 166.955 ;
        RECT 94.325 166.625 95.905 166.955 ;
        RECT 107.895 166.625 109.475 166.955 ;
        RECT 73.970 163.905 75.550 164.235 ;
        RECT 87.540 163.905 89.120 164.235 ;
        RECT 101.110 163.905 102.690 164.235 ;
        RECT 114.680 163.905 116.260 164.235 ;
        RECT 67.185 161.185 68.765 161.515 ;
        RECT 80.755 161.185 82.335 161.515 ;
        RECT 94.325 161.185 95.905 161.515 ;
        RECT 107.895 161.185 109.475 161.515 ;
        RECT 73.970 158.465 75.550 158.795 ;
        RECT 87.540 158.465 89.120 158.795 ;
        RECT 101.110 158.465 102.690 158.795 ;
        RECT 114.680 158.465 116.260 158.795 ;
        RECT 67.185 155.745 68.765 156.075 ;
        RECT 80.755 155.745 82.335 156.075 ;
        RECT 94.325 155.745 95.905 156.075 ;
        RECT 107.895 155.745 109.475 156.075 ;
        RECT 73.970 153.025 75.550 153.355 ;
        RECT 87.540 153.025 89.120 153.355 ;
        RECT 101.110 153.025 102.690 153.355 ;
        RECT 114.680 153.025 116.260 153.355 ;
        RECT 24.565 142.560 26.055 142.585 ;
        RECT 24.560 141.060 68.650 142.560 ;
        RECT 24.565 141.035 26.055 141.060 ;
        RECT 87.255 83.250 88.745 83.275 ;
        RECT 87.250 81.750 91.750 83.250 ;
        RECT 87.255 81.725 88.745 81.750 ;
        RECT 28.255 45.250 29.745 45.275 ;
        RECT 28.250 43.750 68.250 45.250 ;
        RECT 28.255 43.725 29.745 43.750 ;
        RECT 102.780 27.510 103.805 89.470 ;
        RECT 127.085 87.595 127.815 88.325 ;
        RECT 127.110 86.800 127.790 87.595 ;
        RECT 110.070 70.460 126.930 85.860 ;
        RECT 128.770 69.750 145.630 85.150 ;
        RECT 113.580 69.245 114.820 69.270 ;
        RECT 113.580 68.055 116.365 69.245 ;
        RECT 113.580 68.030 114.820 68.055 ;
        RECT 147.090 67.995 148.190 79.630 ;
        RECT 107.735 66.985 108.505 67.755 ;
        RECT 107.760 63.150 108.480 66.985 ;
        RECT 109.980 51.340 126.840 66.740 ;
        RECT 128.940 51.540 145.800 66.940 ;
        RECT 147.065 66.905 148.215 67.995 ;
        RECT 147.090 66.900 148.190 66.905 ;
        RECT 145.550 50.065 146.470 50.070 ;
        RECT 145.525 49.155 146.495 50.065 ;
        RECT 145.550 48.580 146.470 49.155 ;
        RECT 156.410 32.940 157.310 34.950 ;
        RECT 157.970 32.940 158.870 178.730 ;
        RECT 156.410 32.040 158.870 32.940 ;
        RECT 134.890 30.175 141.840 30.210 ;
        RECT 134.890 29.985 142.405 30.175 ;
        RECT 134.890 29.535 142.440 29.985 ;
        RECT 134.890 29.350 142.405 29.535 ;
        RECT 134.890 29.260 141.840 29.350 ;
        RECT 137.190 28.760 140.040 29.260 ;
        RECT 123.990 27.510 130.840 27.860 ;
        RECT 102.780 26.960 130.840 27.510 ;
        RECT 140.840 27.310 150.690 27.410 ;
        RECT 102.780 26.510 124.640 26.960 ;
        RECT 140.840 26.610 152.140 27.310 ;
        RECT 102.780 26.500 103.805 26.510 ;
        RECT 140.840 26.410 141.640 26.610 ;
        RECT 149.840 26.110 152.140 26.610 ;
        RECT 129.540 24.885 144.090 26.085 ;
        RECT 150.940 22.135 152.140 26.110 ;
        RECT 150.915 20.885 152.165 22.135 ;
        RECT 156.410 8.645 157.310 32.040 ;
        RECT 156.385 7.755 157.335 8.645 ;
        RECT 156.410 7.750 157.310 7.755 ;
      LAYER via3 ;
        RECT 107.320 220.690 107.640 221.010 ;
        RECT 100.830 219.420 101.150 219.740 ;
        RECT 81.260 218.250 81.580 218.570 ;
        RECT 77.580 217.040 77.900 217.360 ;
        RECT 73.900 215.770 74.220 216.090 ;
        RECT 70.220 214.180 70.540 214.500 ;
        RECT 62.860 212.720 63.180 213.040 ;
        RECT 66.540 212.830 66.860 213.150 ;
        RECT 113.690 212.020 114.010 212.340 ;
        RECT 74.000 207.430 74.320 207.750 ;
        RECT 74.400 207.430 74.720 207.750 ;
        RECT 74.800 207.430 75.120 207.750 ;
        RECT 75.200 207.430 75.520 207.750 ;
        RECT 87.570 207.430 87.890 207.750 ;
        RECT 87.970 207.430 88.290 207.750 ;
        RECT 88.370 207.430 88.690 207.750 ;
        RECT 88.770 207.430 89.090 207.750 ;
        RECT 101.140 207.430 101.460 207.750 ;
        RECT 101.540 207.430 101.860 207.750 ;
        RECT 101.940 207.430 102.260 207.750 ;
        RECT 102.340 207.430 102.660 207.750 ;
        RECT 114.710 207.430 115.030 207.750 ;
        RECT 115.110 207.430 115.430 207.750 ;
        RECT 115.510 207.430 115.830 207.750 ;
        RECT 115.910 207.430 116.230 207.750 ;
        RECT 67.215 204.710 67.535 205.030 ;
        RECT 67.615 204.710 67.935 205.030 ;
        RECT 68.015 204.710 68.335 205.030 ;
        RECT 68.415 204.710 68.735 205.030 ;
        RECT 80.785 204.710 81.105 205.030 ;
        RECT 81.185 204.710 81.505 205.030 ;
        RECT 81.585 204.710 81.905 205.030 ;
        RECT 81.985 204.710 82.305 205.030 ;
        RECT 94.355 204.710 94.675 205.030 ;
        RECT 94.755 204.710 95.075 205.030 ;
        RECT 95.155 204.710 95.475 205.030 ;
        RECT 95.555 204.710 95.875 205.030 ;
        RECT 107.925 204.710 108.245 205.030 ;
        RECT 108.325 204.710 108.645 205.030 ;
        RECT 108.725 204.710 109.045 205.030 ;
        RECT 109.125 204.710 109.445 205.030 ;
        RECT 74.000 201.990 74.320 202.310 ;
        RECT 74.400 201.990 74.720 202.310 ;
        RECT 74.800 201.990 75.120 202.310 ;
        RECT 75.200 201.990 75.520 202.310 ;
        RECT 87.570 201.990 87.890 202.310 ;
        RECT 87.970 201.990 88.290 202.310 ;
        RECT 88.370 201.990 88.690 202.310 ;
        RECT 88.770 201.990 89.090 202.310 ;
        RECT 101.140 201.990 101.460 202.310 ;
        RECT 101.540 201.990 101.860 202.310 ;
        RECT 101.940 201.990 102.260 202.310 ;
        RECT 102.340 201.990 102.660 202.310 ;
        RECT 114.710 201.990 115.030 202.310 ;
        RECT 115.110 201.990 115.430 202.310 ;
        RECT 115.510 201.990 115.830 202.310 ;
        RECT 115.910 201.990 116.230 202.310 ;
        RECT 67.215 199.270 67.535 199.590 ;
        RECT 67.615 199.270 67.935 199.590 ;
        RECT 68.015 199.270 68.335 199.590 ;
        RECT 68.415 199.270 68.735 199.590 ;
        RECT 80.785 199.270 81.105 199.590 ;
        RECT 81.185 199.270 81.505 199.590 ;
        RECT 81.585 199.270 81.905 199.590 ;
        RECT 81.985 199.270 82.305 199.590 ;
        RECT 94.355 199.270 94.675 199.590 ;
        RECT 94.755 199.270 95.075 199.590 ;
        RECT 95.155 199.270 95.475 199.590 ;
        RECT 95.555 199.270 95.875 199.590 ;
        RECT 107.925 199.270 108.245 199.590 ;
        RECT 108.325 199.270 108.645 199.590 ;
        RECT 108.725 199.270 109.045 199.590 ;
        RECT 109.125 199.270 109.445 199.590 ;
        RECT 103.810 198.250 104.130 198.570 ;
        RECT 74.000 196.550 74.320 196.870 ;
        RECT 74.400 196.550 74.720 196.870 ;
        RECT 74.800 196.550 75.120 196.870 ;
        RECT 75.200 196.550 75.520 196.870 ;
        RECT 87.570 196.550 87.890 196.870 ;
        RECT 87.970 196.550 88.290 196.870 ;
        RECT 88.370 196.550 88.690 196.870 ;
        RECT 88.770 196.550 89.090 196.870 ;
        RECT 101.140 196.550 101.460 196.870 ;
        RECT 101.540 196.550 101.860 196.870 ;
        RECT 101.940 196.550 102.260 196.870 ;
        RECT 102.340 196.550 102.660 196.870 ;
        RECT 114.710 196.550 115.030 196.870 ;
        RECT 115.110 196.550 115.430 196.870 ;
        RECT 115.510 196.550 115.830 196.870 ;
        RECT 115.910 196.550 116.230 196.870 ;
        RECT 67.215 193.830 67.535 194.150 ;
        RECT 67.615 193.830 67.935 194.150 ;
        RECT 68.015 193.830 68.335 194.150 ;
        RECT 68.415 193.830 68.735 194.150 ;
        RECT 80.785 193.830 81.105 194.150 ;
        RECT 81.185 193.830 81.505 194.150 ;
        RECT 81.585 193.830 81.905 194.150 ;
        RECT 81.985 193.830 82.305 194.150 ;
        RECT 94.355 193.830 94.675 194.150 ;
        RECT 94.755 193.830 95.075 194.150 ;
        RECT 95.155 193.830 95.475 194.150 ;
        RECT 95.555 193.830 95.875 194.150 ;
        RECT 107.925 193.830 108.245 194.150 ;
        RECT 108.325 193.830 108.645 194.150 ;
        RECT 108.725 193.830 109.045 194.150 ;
        RECT 109.125 193.830 109.445 194.150 ;
        RECT 74.000 191.110 74.320 191.430 ;
        RECT 74.400 191.110 74.720 191.430 ;
        RECT 74.800 191.110 75.120 191.430 ;
        RECT 75.200 191.110 75.520 191.430 ;
        RECT 87.570 191.110 87.890 191.430 ;
        RECT 87.970 191.110 88.290 191.430 ;
        RECT 88.370 191.110 88.690 191.430 ;
        RECT 88.770 191.110 89.090 191.430 ;
        RECT 101.140 191.110 101.460 191.430 ;
        RECT 101.540 191.110 101.860 191.430 ;
        RECT 101.940 191.110 102.260 191.430 ;
        RECT 102.340 191.110 102.660 191.430 ;
        RECT 114.710 191.110 115.030 191.430 ;
        RECT 115.110 191.110 115.430 191.430 ;
        RECT 115.510 191.110 115.830 191.430 ;
        RECT 115.910 191.110 116.230 191.430 ;
        RECT 67.215 188.390 67.535 188.710 ;
        RECT 67.615 188.390 67.935 188.710 ;
        RECT 68.015 188.390 68.335 188.710 ;
        RECT 68.415 188.390 68.735 188.710 ;
        RECT 80.785 188.390 81.105 188.710 ;
        RECT 81.185 188.390 81.505 188.710 ;
        RECT 81.585 188.390 81.905 188.710 ;
        RECT 81.985 188.390 82.305 188.710 ;
        RECT 94.355 188.390 94.675 188.710 ;
        RECT 94.755 188.390 95.075 188.710 ;
        RECT 95.155 188.390 95.475 188.710 ;
        RECT 95.555 188.390 95.875 188.710 ;
        RECT 107.925 188.390 108.245 188.710 ;
        RECT 108.325 188.390 108.645 188.710 ;
        RECT 108.725 188.390 109.045 188.710 ;
        RECT 109.125 188.390 109.445 188.710 ;
        RECT 74.000 185.670 74.320 185.990 ;
        RECT 74.400 185.670 74.720 185.990 ;
        RECT 74.800 185.670 75.120 185.990 ;
        RECT 75.200 185.670 75.520 185.990 ;
        RECT 87.570 185.670 87.890 185.990 ;
        RECT 87.970 185.670 88.290 185.990 ;
        RECT 88.370 185.670 88.690 185.990 ;
        RECT 88.770 185.670 89.090 185.990 ;
        RECT 101.140 185.670 101.460 185.990 ;
        RECT 101.540 185.670 101.860 185.990 ;
        RECT 101.940 185.670 102.260 185.990 ;
        RECT 102.340 185.670 102.660 185.990 ;
        RECT 114.710 185.670 115.030 185.990 ;
        RECT 115.110 185.670 115.430 185.990 ;
        RECT 115.510 185.670 115.830 185.990 ;
        RECT 115.910 185.670 116.230 185.990 ;
        RECT 67.215 182.950 67.535 183.270 ;
        RECT 67.615 182.950 67.935 183.270 ;
        RECT 68.015 182.950 68.335 183.270 ;
        RECT 68.415 182.950 68.735 183.270 ;
        RECT 80.785 182.950 81.105 183.270 ;
        RECT 81.185 182.950 81.505 183.270 ;
        RECT 81.585 182.950 81.905 183.270 ;
        RECT 81.985 182.950 82.305 183.270 ;
        RECT 94.355 182.950 94.675 183.270 ;
        RECT 94.755 182.950 95.075 183.270 ;
        RECT 95.155 182.950 95.475 183.270 ;
        RECT 95.555 182.950 95.875 183.270 ;
        RECT 107.925 182.950 108.245 183.270 ;
        RECT 108.325 182.950 108.645 183.270 ;
        RECT 108.725 182.950 109.045 183.270 ;
        RECT 109.125 182.950 109.445 183.270 ;
        RECT 103.810 181.930 104.130 182.250 ;
        RECT 74.000 180.230 74.320 180.550 ;
        RECT 74.400 180.230 74.720 180.550 ;
        RECT 74.800 180.230 75.120 180.550 ;
        RECT 75.200 180.230 75.520 180.550 ;
        RECT 87.570 180.230 87.890 180.550 ;
        RECT 87.970 180.230 88.290 180.550 ;
        RECT 88.370 180.230 88.690 180.550 ;
        RECT 88.770 180.230 89.090 180.550 ;
        RECT 101.140 180.230 101.460 180.550 ;
        RECT 101.540 180.230 101.860 180.550 ;
        RECT 101.940 180.230 102.260 180.550 ;
        RECT 102.340 180.230 102.660 180.550 ;
        RECT 114.710 180.230 115.030 180.550 ;
        RECT 115.110 180.230 115.430 180.550 ;
        RECT 115.510 180.230 115.830 180.550 ;
        RECT 115.910 180.230 116.230 180.550 ;
        RECT 67.215 177.510 67.535 177.830 ;
        RECT 67.615 177.510 67.935 177.830 ;
        RECT 68.015 177.510 68.335 177.830 ;
        RECT 68.415 177.510 68.735 177.830 ;
        RECT 80.785 177.510 81.105 177.830 ;
        RECT 81.185 177.510 81.505 177.830 ;
        RECT 81.585 177.510 81.905 177.830 ;
        RECT 81.985 177.510 82.305 177.830 ;
        RECT 94.355 177.510 94.675 177.830 ;
        RECT 94.755 177.510 95.075 177.830 ;
        RECT 95.155 177.510 95.475 177.830 ;
        RECT 95.555 177.510 95.875 177.830 ;
        RECT 107.925 177.510 108.245 177.830 ;
        RECT 108.325 177.510 108.645 177.830 ;
        RECT 108.725 177.510 109.045 177.830 ;
        RECT 109.125 177.510 109.445 177.830 ;
        RECT 74.000 174.790 74.320 175.110 ;
        RECT 74.400 174.790 74.720 175.110 ;
        RECT 74.800 174.790 75.120 175.110 ;
        RECT 75.200 174.790 75.520 175.110 ;
        RECT 87.570 174.790 87.890 175.110 ;
        RECT 87.970 174.790 88.290 175.110 ;
        RECT 88.370 174.790 88.690 175.110 ;
        RECT 88.770 174.790 89.090 175.110 ;
        RECT 101.140 174.790 101.460 175.110 ;
        RECT 101.540 174.790 101.860 175.110 ;
        RECT 101.940 174.790 102.260 175.110 ;
        RECT 102.340 174.790 102.660 175.110 ;
        RECT 114.710 174.790 115.030 175.110 ;
        RECT 115.110 174.790 115.430 175.110 ;
        RECT 115.510 174.790 115.830 175.110 ;
        RECT 115.910 174.790 116.230 175.110 ;
        RECT 67.215 172.070 67.535 172.390 ;
        RECT 67.615 172.070 67.935 172.390 ;
        RECT 68.015 172.070 68.335 172.390 ;
        RECT 68.415 172.070 68.735 172.390 ;
        RECT 80.785 172.070 81.105 172.390 ;
        RECT 81.185 172.070 81.505 172.390 ;
        RECT 81.585 172.070 81.905 172.390 ;
        RECT 81.985 172.070 82.305 172.390 ;
        RECT 94.355 172.070 94.675 172.390 ;
        RECT 94.755 172.070 95.075 172.390 ;
        RECT 95.155 172.070 95.475 172.390 ;
        RECT 95.555 172.070 95.875 172.390 ;
        RECT 107.925 172.070 108.245 172.390 ;
        RECT 108.325 172.070 108.645 172.390 ;
        RECT 108.725 172.070 109.045 172.390 ;
        RECT 109.125 172.070 109.445 172.390 ;
        RECT 74.000 169.350 74.320 169.670 ;
        RECT 74.400 169.350 74.720 169.670 ;
        RECT 74.800 169.350 75.120 169.670 ;
        RECT 75.200 169.350 75.520 169.670 ;
        RECT 87.570 169.350 87.890 169.670 ;
        RECT 87.970 169.350 88.290 169.670 ;
        RECT 88.370 169.350 88.690 169.670 ;
        RECT 88.770 169.350 89.090 169.670 ;
        RECT 101.140 169.350 101.460 169.670 ;
        RECT 101.540 169.350 101.860 169.670 ;
        RECT 101.940 169.350 102.260 169.670 ;
        RECT 102.340 169.350 102.660 169.670 ;
        RECT 114.710 169.350 115.030 169.670 ;
        RECT 115.110 169.350 115.430 169.670 ;
        RECT 115.510 169.350 115.830 169.670 ;
        RECT 115.910 169.350 116.230 169.670 ;
        RECT 67.215 166.630 67.535 166.950 ;
        RECT 67.615 166.630 67.935 166.950 ;
        RECT 68.015 166.630 68.335 166.950 ;
        RECT 68.415 166.630 68.735 166.950 ;
        RECT 80.785 166.630 81.105 166.950 ;
        RECT 81.185 166.630 81.505 166.950 ;
        RECT 81.585 166.630 81.905 166.950 ;
        RECT 81.985 166.630 82.305 166.950 ;
        RECT 94.355 166.630 94.675 166.950 ;
        RECT 94.755 166.630 95.075 166.950 ;
        RECT 95.155 166.630 95.475 166.950 ;
        RECT 95.555 166.630 95.875 166.950 ;
        RECT 107.925 166.630 108.245 166.950 ;
        RECT 108.325 166.630 108.645 166.950 ;
        RECT 108.725 166.630 109.045 166.950 ;
        RECT 109.125 166.630 109.445 166.950 ;
        RECT 74.000 163.910 74.320 164.230 ;
        RECT 74.400 163.910 74.720 164.230 ;
        RECT 74.800 163.910 75.120 164.230 ;
        RECT 75.200 163.910 75.520 164.230 ;
        RECT 87.570 163.910 87.890 164.230 ;
        RECT 87.970 163.910 88.290 164.230 ;
        RECT 88.370 163.910 88.690 164.230 ;
        RECT 88.770 163.910 89.090 164.230 ;
        RECT 101.140 163.910 101.460 164.230 ;
        RECT 101.540 163.910 101.860 164.230 ;
        RECT 101.940 163.910 102.260 164.230 ;
        RECT 102.340 163.910 102.660 164.230 ;
        RECT 114.710 163.910 115.030 164.230 ;
        RECT 115.110 163.910 115.430 164.230 ;
        RECT 115.510 163.910 115.830 164.230 ;
        RECT 115.910 163.910 116.230 164.230 ;
        RECT 67.215 161.190 67.535 161.510 ;
        RECT 67.615 161.190 67.935 161.510 ;
        RECT 68.015 161.190 68.335 161.510 ;
        RECT 68.415 161.190 68.735 161.510 ;
        RECT 80.785 161.190 81.105 161.510 ;
        RECT 81.185 161.190 81.505 161.510 ;
        RECT 81.585 161.190 81.905 161.510 ;
        RECT 81.985 161.190 82.305 161.510 ;
        RECT 94.355 161.190 94.675 161.510 ;
        RECT 94.755 161.190 95.075 161.510 ;
        RECT 95.155 161.190 95.475 161.510 ;
        RECT 95.555 161.190 95.875 161.510 ;
        RECT 107.925 161.190 108.245 161.510 ;
        RECT 108.325 161.190 108.645 161.510 ;
        RECT 108.725 161.190 109.045 161.510 ;
        RECT 109.125 161.190 109.445 161.510 ;
        RECT 74.000 158.470 74.320 158.790 ;
        RECT 74.400 158.470 74.720 158.790 ;
        RECT 74.800 158.470 75.120 158.790 ;
        RECT 75.200 158.470 75.520 158.790 ;
        RECT 87.570 158.470 87.890 158.790 ;
        RECT 87.970 158.470 88.290 158.790 ;
        RECT 88.370 158.470 88.690 158.790 ;
        RECT 88.770 158.470 89.090 158.790 ;
        RECT 101.140 158.470 101.460 158.790 ;
        RECT 101.540 158.470 101.860 158.790 ;
        RECT 101.940 158.470 102.260 158.790 ;
        RECT 102.340 158.470 102.660 158.790 ;
        RECT 114.710 158.470 115.030 158.790 ;
        RECT 115.110 158.470 115.430 158.790 ;
        RECT 115.510 158.470 115.830 158.790 ;
        RECT 115.910 158.470 116.230 158.790 ;
        RECT 67.215 155.750 67.535 156.070 ;
        RECT 67.615 155.750 67.935 156.070 ;
        RECT 68.015 155.750 68.335 156.070 ;
        RECT 68.415 155.750 68.735 156.070 ;
        RECT 80.785 155.750 81.105 156.070 ;
        RECT 81.185 155.750 81.505 156.070 ;
        RECT 81.585 155.750 81.905 156.070 ;
        RECT 81.985 155.750 82.305 156.070 ;
        RECT 94.355 155.750 94.675 156.070 ;
        RECT 94.755 155.750 95.075 156.070 ;
        RECT 95.155 155.750 95.475 156.070 ;
        RECT 95.555 155.750 95.875 156.070 ;
        RECT 107.925 155.750 108.245 156.070 ;
        RECT 108.325 155.750 108.645 156.070 ;
        RECT 108.725 155.750 109.045 156.070 ;
        RECT 109.125 155.750 109.445 156.070 ;
        RECT 74.000 153.030 74.320 153.350 ;
        RECT 74.400 153.030 74.720 153.350 ;
        RECT 74.800 153.030 75.120 153.350 ;
        RECT 75.200 153.030 75.520 153.350 ;
        RECT 87.570 153.030 87.890 153.350 ;
        RECT 87.970 153.030 88.290 153.350 ;
        RECT 88.370 153.030 88.690 153.350 ;
        RECT 88.770 153.030 89.090 153.350 ;
        RECT 101.140 153.030 101.460 153.350 ;
        RECT 101.540 153.030 101.860 153.350 ;
        RECT 101.940 153.030 102.260 153.350 ;
        RECT 102.340 153.030 102.660 153.350 ;
        RECT 114.710 153.030 115.030 153.350 ;
        RECT 115.110 153.030 115.430 153.350 ;
        RECT 115.510 153.030 115.830 153.350 ;
        RECT 115.910 153.030 116.230 153.350 ;
        RECT 24.565 141.065 26.055 142.555 ;
        RECT 67.120 141.060 68.620 142.560 ;
        RECT 87.255 81.755 88.745 83.245 ;
        RECT 28.255 43.755 29.745 45.245 ;
        RECT 127.110 86.830 127.790 87.510 ;
        RECT 126.510 70.600 126.830 85.720 ;
        RECT 145.210 69.890 145.530 85.010 ;
        RECT 115.145 68.055 116.335 69.245 ;
        RECT 147.095 66.905 148.185 67.995 ;
        RECT 107.760 63.180 108.480 63.900 ;
        RECT 126.420 51.480 126.740 66.600 ;
        RECT 145.380 51.680 145.700 66.800 ;
        RECT 145.555 49.155 146.465 50.065 ;
        RECT 156.415 7.755 157.305 8.645 ;
      LAYER met4 ;
        RECT 3.990 223.800 4.290 224.760 ;
        RECT 7.670 223.800 7.970 224.760 ;
        RECT 11.350 223.800 11.650 224.760 ;
        RECT 15.030 223.800 15.330 224.760 ;
        RECT 18.710 223.800 19.010 224.760 ;
        RECT 22.390 223.800 22.690 224.760 ;
        RECT 26.070 223.800 26.370 224.760 ;
        RECT 29.750 223.800 30.050 224.760 ;
        RECT 33.430 223.800 33.730 224.760 ;
        RECT 37.110 223.800 37.410 224.760 ;
        RECT 40.790 223.800 41.090 224.760 ;
        RECT 44.470 223.800 44.770 224.760 ;
        RECT 48.150 223.800 48.450 224.760 ;
        RECT 51.830 223.800 52.130 224.760 ;
        RECT 55.510 223.800 55.810 224.760 ;
        RECT 59.190 223.800 59.490 224.760 ;
        RECT 3.200 223.500 59.920 223.800 ;
        RECT 49.000 220.760 50.500 223.500 ;
        RECT 62.870 213.045 63.170 224.760 ;
        RECT 66.550 213.155 66.850 224.760 ;
        RECT 70.230 214.505 70.530 224.760 ;
        RECT 73.910 216.095 74.210 224.760 ;
        RECT 77.590 217.365 77.890 224.760 ;
        RECT 81.270 218.575 81.570 224.760 ;
        RECT 84.950 219.730 85.250 224.760 ;
        RECT 88.630 221.000 88.930 224.760 ;
        RECT 107.315 221.000 107.645 221.015 ;
        RECT 88.630 220.700 107.645 221.000 ;
        RECT 107.315 220.685 107.645 220.700 ;
        RECT 100.825 219.730 101.155 219.745 ;
        RECT 84.950 219.430 101.155 219.730 ;
        RECT 100.825 219.415 101.155 219.430 ;
        RECT 81.255 218.245 81.585 218.575 ;
        RECT 77.575 217.035 77.905 217.365 ;
        RECT 73.895 215.765 74.225 216.095 ;
        RECT 70.215 214.175 70.545 214.505 ;
        RECT 62.855 212.715 63.185 213.045 ;
        RECT 66.535 212.825 66.865 213.155 ;
        RECT 113.685 212.330 114.015 212.345 ;
        RECT 151.190 212.330 151.490 224.760 ;
        RECT 113.685 212.030 151.490 212.330 ;
        RECT 113.685 212.015 114.015 212.030 ;
        RECT 67.175 155.880 68.775 207.830 ;
        RECT 73.960 158.100 75.560 207.830 ;
        RECT 67.120 152.950 68.775 155.880 ;
        RECT 73.930 152.950 75.560 158.100 ;
        RECT 80.745 152.950 82.345 207.830 ;
        RECT 87.530 152.950 89.130 207.830 ;
        RECT 94.315 152.950 95.915 207.830 ;
        RECT 101.100 152.950 102.700 207.830 ;
        RECT 103.805 198.245 104.135 198.575 ;
        RECT 103.820 182.255 104.120 198.245 ;
        RECT 103.805 181.925 104.135 182.255 ;
        RECT 107.885 152.950 109.485 207.830 ;
        RECT 114.670 152.950 116.270 207.830 ;
        RECT 67.120 142.565 68.620 152.950 ;
        RECT 2.500 141.060 26.060 142.560 ;
        RECT 67.115 141.055 68.625 142.565 ;
        RECT 73.930 138.480 75.430 152.950 ;
        RECT 50.500 136.980 75.430 138.480 ;
        RECT 127.105 87.020 127.795 87.515 ;
        RECT 125.990 85.840 145.960 87.020 ;
        RECT 50.500 81.750 88.750 83.250 ;
        RECT 110.465 70.855 125.075 85.465 ;
        RECT 125.990 80.000 127.170 85.840 ;
        RECT 116.860 69.285 117.990 70.855 ;
        RECT 126.430 70.520 126.910 80.000 ;
        RECT 129.165 70.145 143.775 84.755 ;
        RECT 144.780 79.440 145.960 85.840 ;
        RECT 136.855 69.285 137.985 70.145 ;
        RECT 145.130 69.810 145.610 79.440 ;
        RECT 115.140 69.245 116.340 69.250 ;
        RECT 116.860 69.245 137.985 69.285 ;
        RECT 115.140 68.155 137.985 69.245 ;
        RECT 115.140 68.055 117.785 68.155 ;
        RECT 115.140 68.050 116.340 68.055 ;
        RECT 144.950 66.900 148.190 68.000 ;
        RECT 107.755 63.900 108.485 63.905 ;
        RECT 110.375 63.900 124.985 66.345 ;
        RECT 126.340 66.220 126.820 66.680 ;
        RECT 129.335 66.220 143.945 66.545 ;
        RECT 107.755 63.180 124.985 63.900 ;
        RECT 107.755 63.175 108.485 63.180 ;
        RECT 110.375 51.735 124.985 63.180 ;
        RECT 126.100 61.410 143.945 66.220 ;
        RECT 144.950 62.060 146.050 66.900 ;
        RECT 126.340 51.400 126.820 61.410 ;
        RECT 127.380 50.790 128.300 61.410 ;
        RECT 129.335 51.935 143.945 61.410 ;
        RECT 145.300 51.600 145.780 62.060 ;
        RECT 127.380 49.870 146.470 50.790 ;
        RECT 145.550 49.150 146.470 49.870 ;
        RECT 2.500 43.750 29.750 45.250 ;
        RECT 156.410 1.000 157.310 8.650 ;
  END
END tt_um_twin_tee_opamp_osc
END LIBRARY

