MACRO tt_um_brucemack_sb_mixer
  CLASS BLOCK ;
  FOREIGN tt_um_brucemack_sb_mixer ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.435600 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 79.824295 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 110.740 63.630 126.560 65.640 ;
        RECT 136.490 63.630 152.310 65.640 ;
        RECT 110.750 53.990 122.850 57.950 ;
        RECT 99.620 50.650 106.130 53.000 ;
        RECT 130.170 49.150 134.130 61.250 ;
        RECT 110.830 44.150 122.930 48.110 ;
      LAYER nwell ;
        RECT 128.980 39.930 130.585 42.530 ;
      LAYER pwell ;
        RECT 130.875 41.275 131.785 42.100 ;
        RECT 130.875 41.170 131.975 41.275 ;
        RECT 131.805 41.105 131.975 41.170 ;
        RECT 130.915 40.135 131.700 40.565 ;
      LAYER nwell ;
        RECT 134.980 39.930 136.585 42.530 ;
      LAYER pwell ;
        RECT 136.875 41.275 137.785 42.100 ;
        RECT 136.875 41.170 137.975 41.275 ;
        RECT 137.805 41.105 137.975 41.170 ;
        RECT 136.915 40.135 137.700 40.565 ;
        RECT 110.830 35.190 122.930 39.150 ;
        RECT 129.620 37.060 131.660 39.100 ;
        RECT 143.300 35.600 154.130 47.700 ;
        RECT 149.060 35.120 150.630 35.600 ;
        RECT 151.370 35.130 152.940 35.600 ;
        RECT 99.620 31.470 106.130 33.820 ;
        RECT 110.830 26.230 122.930 30.190 ;
        RECT 130.170 22.050 134.130 34.150 ;
        RECT 132.100 20.940 132.880 22.050 ;
        RECT 142.740 21.230 143.450 22.900 ;
        RECT 142.740 20.880 144.210 21.230 ;
        RECT 144.980 20.880 146.630 21.220 ;
        RECT 147.420 20.880 148.730 21.210 ;
        RECT 149.520 20.880 151.230 21.200 ;
        RECT 111.940 17.670 137.760 18.360 ;
        RECT 141.530 17.670 152.360 20.880 ;
        RECT 111.940 17.050 152.360 17.670 ;
        RECT 111.940 16.350 137.760 17.050 ;
        RECT 141.530 13.780 152.360 17.050 ;
      LAYER li1 ;
        RECT 110.920 65.290 126.380 65.460 ;
        RECT 110.920 63.980 111.090 65.290 ;
        RECT 111.570 64.460 113.730 64.810 ;
        RECT 123.570 64.460 125.730 64.810 ;
        RECT 111.410 63.980 112.110 64.080 ;
        RECT 126.210 63.980 126.380 65.290 ;
        RECT 110.920 63.810 126.380 63.980 ;
        RECT 136.670 65.290 152.130 65.460 ;
        RECT 136.670 63.980 136.840 65.290 ;
        RECT 151.960 65.050 152.130 65.290 ;
        RECT 137.320 64.460 139.480 64.810 ;
        RECT 149.320 64.460 151.480 64.810 ;
        RECT 151.860 64.250 152.260 65.050 ;
        RECT 151.960 63.980 152.130 64.250 ;
        RECT 136.670 63.810 152.130 63.980 ;
        RECT 111.410 63.620 112.110 63.810 ;
        RECT 130.350 60.900 133.950 61.070 ;
        RECT 110.930 57.600 122.670 57.770 ;
        RECT 110.930 57.250 111.100 57.600 ;
        RECT 110.790 54.720 111.190 57.250 ;
        RECT 111.780 57.030 121.820 57.200 ;
        RECT 111.440 54.970 111.610 56.970 ;
        RECT 121.990 54.970 122.160 56.970 ;
        RECT 111.780 54.740 121.820 54.910 ;
        RECT 110.930 54.340 111.100 54.720 ;
        RECT 122.500 54.340 122.670 57.600 ;
        RECT 110.930 54.170 122.670 54.340 ;
        RECT 103.720 52.820 104.820 52.910 ;
        RECT 99.800 52.650 105.950 52.820 ;
        RECT 99.800 51.000 99.970 52.650 ;
        RECT 103.720 52.560 104.820 52.650 ;
        RECT 100.450 51.480 102.610 52.170 ;
        RECT 103.140 51.480 105.300 52.170 ;
        RECT 105.780 51.000 105.950 52.650 ;
        RECT 99.800 50.830 105.950 51.000 ;
        RECT 130.350 49.500 130.520 60.900 ;
        RECT 131.150 60.390 133.150 60.560 ;
        RECT 130.920 50.180 131.090 60.220 ;
        RECT 133.210 50.180 133.380 60.220 ;
        RECT 131.150 49.840 133.150 50.010 ;
        RECT 131.100 49.500 133.100 49.560 ;
        RECT 133.780 49.500 133.950 60.900 ;
        RECT 130.350 49.330 133.950 49.500 ;
        RECT 131.100 49.240 133.100 49.330 ;
        RECT 111.010 47.760 122.750 47.930 ;
        RECT 111.010 47.360 111.180 47.760 ;
        RECT 110.890 44.880 111.280 47.360 ;
        RECT 111.860 47.190 121.900 47.360 ;
        RECT 111.520 45.130 111.690 47.130 ;
        RECT 122.070 45.130 122.240 47.130 ;
        RECT 111.860 44.900 121.900 45.070 ;
        RECT 111.010 44.500 111.180 44.880 ;
        RECT 122.580 44.500 122.750 47.760 ;
        RECT 111.010 44.330 122.750 44.500 ;
        RECT 143.480 47.350 153.950 47.520 ;
        RECT 129.085 41.510 129.255 42.340 ;
        RECT 129.425 41.780 131.635 42.010 ;
        RECT 129.425 41.680 130.405 41.780 ;
        RECT 131.005 41.680 131.635 41.780 ;
        RECT 129.085 41.300 130.395 41.510 ;
        RECT 129.085 40.960 129.255 41.300 ;
        RECT 130.575 41.280 130.815 41.610 ;
        RECT 131.805 41.510 131.975 42.340 ;
        RECT 130.985 41.280 131.975 41.510 ;
        RECT 131.805 40.960 131.975 41.280 ;
        RECT 135.085 41.510 135.255 42.340 ;
        RECT 135.425 41.780 137.635 42.010 ;
        RECT 135.425 41.680 136.405 41.780 ;
        RECT 137.005 41.680 137.635 41.780 ;
        RECT 135.085 41.300 136.395 41.510 ;
        RECT 135.085 40.960 135.255 41.300 ;
        RECT 136.575 41.280 136.815 41.610 ;
        RECT 137.805 41.510 137.975 42.340 ;
        RECT 136.985 41.280 137.975 41.510 ;
        RECT 137.805 40.960 137.975 41.280 ;
        RECT 129.085 40.495 129.255 40.580 ;
        RECT 131.805 40.495 131.975 40.580 ;
        RECT 129.085 40.205 130.420 40.495 ;
        RECT 131.080 40.205 131.975 40.495 ;
        RECT 129.085 40.120 129.255 40.205 ;
        RECT 131.805 40.120 131.975 40.205 ;
        RECT 135.085 40.495 135.255 40.580 ;
        RECT 137.805 40.495 137.975 40.580 ;
        RECT 135.085 40.205 136.420 40.495 ;
        RECT 137.080 40.205 137.975 40.495 ;
        RECT 135.085 40.120 135.255 40.205 ;
        RECT 137.805 40.120 137.975 40.205 ;
        RECT 111.010 38.800 122.750 38.970 ;
        RECT 111.010 38.430 111.180 38.800 ;
        RECT 110.900 35.940 111.250 38.430 ;
        RECT 111.860 38.230 121.900 38.400 ;
        RECT 111.520 36.170 111.690 38.170 ;
        RECT 122.070 36.170 122.240 38.170 ;
        RECT 111.860 35.940 121.900 36.110 ;
        RECT 111.010 35.540 111.180 35.940 ;
        RECT 122.580 35.540 122.750 38.800 ;
        RECT 129.800 38.750 131.480 38.920 ;
        RECT 129.800 37.410 129.970 38.750 ;
        RECT 131.310 38.510 131.480 38.750 ;
        RECT 130.370 37.730 130.910 38.430 ;
        RECT 131.250 37.680 131.560 38.510 ;
        RECT 131.310 37.410 131.480 37.680 ;
        RECT 129.800 37.240 131.480 37.410 ;
        RECT 143.480 35.950 143.650 47.350 ;
        RECT 144.280 46.840 146.280 47.010 ;
        RECT 146.570 46.840 148.570 47.010 ;
        RECT 148.860 46.840 150.860 47.010 ;
        RECT 151.150 46.840 153.150 47.010 ;
        RECT 144.050 36.630 144.220 46.670 ;
        RECT 146.340 36.630 146.510 46.670 ;
        RECT 148.630 36.630 148.800 46.670 ;
        RECT 150.920 36.630 151.090 46.670 ;
        RECT 153.210 36.630 153.380 46.670 ;
        RECT 153.780 41.960 153.950 47.350 ;
        RECT 153.660 40.420 154.040 41.960 ;
        RECT 144.280 36.290 146.280 36.460 ;
        RECT 146.570 36.290 148.570 36.460 ;
        RECT 148.860 36.290 150.860 36.460 ;
        RECT 151.150 36.290 153.150 36.460 ;
        RECT 153.780 35.950 153.950 40.420 ;
        RECT 143.480 35.780 153.950 35.950 ;
        RECT 111.010 35.370 122.750 35.540 ;
        RECT 130.940 33.970 133.120 34.090 ;
        RECT 130.350 33.800 133.950 33.970 ;
        RECT 99.800 33.470 105.950 33.640 ;
        RECT 99.800 31.820 99.970 33.470 ;
        RECT 100.450 32.300 102.610 32.990 ;
        RECT 103.140 32.300 105.300 32.990 ;
        RECT 103.910 31.820 105.210 31.940 ;
        RECT 105.780 31.820 105.950 33.470 ;
        RECT 99.800 31.650 105.950 31.820 ;
        RECT 103.910 31.540 105.210 31.650 ;
        RECT 111.010 29.840 122.750 30.010 ;
        RECT 111.010 29.400 111.180 29.840 ;
        RECT 110.950 27.040 111.280 29.400 ;
        RECT 111.860 29.270 121.900 29.440 ;
        RECT 111.520 27.210 111.690 29.210 ;
        RECT 122.070 27.210 122.240 29.210 ;
        RECT 111.010 26.580 111.180 27.040 ;
        RECT 111.860 26.980 121.900 27.150 ;
        RECT 122.580 26.580 122.750 29.840 ;
        RECT 111.010 26.410 122.750 26.580 ;
        RECT 130.350 22.400 130.520 33.800 ;
        RECT 130.940 33.710 133.120 33.800 ;
        RECT 131.150 33.290 133.150 33.460 ;
        RECT 130.920 23.080 131.090 33.120 ;
        RECT 133.210 23.080 133.380 33.120 ;
        RECT 131.150 22.740 133.150 22.910 ;
        RECT 133.780 22.400 133.950 33.800 ;
        RECT 130.350 22.230 133.950 22.400 ;
        RECT 141.710 20.530 152.180 20.700 ;
        RECT 113.630 18.180 114.840 18.310 ;
        RECT 112.120 18.010 137.580 18.180 ;
        RECT 112.120 16.700 112.290 18.010 ;
        RECT 113.630 17.890 114.840 18.010 ;
        RECT 112.770 17.180 114.930 17.530 ;
        RECT 134.770 17.180 136.930 17.530 ;
        RECT 137.410 16.700 137.580 18.010 ;
        RECT 112.120 16.530 137.580 16.700 ;
        RECT 141.710 14.130 141.880 20.530 ;
        RECT 142.510 20.020 144.510 20.190 ;
        RECT 144.800 20.020 146.800 20.190 ;
        RECT 147.090 20.020 149.090 20.190 ;
        RECT 149.380 20.020 151.380 20.190 ;
        RECT 142.280 14.810 142.450 19.850 ;
        RECT 144.570 14.810 144.740 19.850 ;
        RECT 146.860 14.810 147.030 19.850 ;
        RECT 149.150 14.810 149.320 19.850 ;
        RECT 151.440 14.810 151.610 19.850 ;
        RECT 152.010 18.370 152.180 20.530 ;
        RECT 151.940 14.900 152.340 18.370 ;
        RECT 142.510 14.470 144.510 14.640 ;
        RECT 144.800 14.470 146.800 14.640 ;
        RECT 147.090 14.470 149.090 14.640 ;
        RECT 149.380 14.470 151.380 14.640 ;
        RECT 152.010 14.130 152.180 14.900 ;
        RECT 141.710 13.960 152.180 14.130 ;
      LAYER met1 ;
        RECT 109.270 64.900 110.040 65.510 ;
        RECT 109.270 64.330 113.800 64.900 ;
        RECT 123.660 64.760 139.600 65.050 ;
        RECT 149.680 64.980 151.000 65.030 ;
        RECT 123.595 64.510 139.600 64.760 ;
        RECT 109.270 63.740 110.040 64.330 ;
        RECT 123.660 64.300 139.600 64.510 ;
        RECT 149.290 64.310 151.630 64.980 ;
        RECT 111.370 63.130 112.200 64.140 ;
        RECT 111.510 62.710 111.960 63.130 ;
        RECT 112.190 60.585 113.120 60.610 ;
        RECT 131.320 60.590 132.890 64.300 ;
        RECT 149.680 64.260 151.000 64.310 ;
        RECT 151.770 64.170 152.480 65.160 ;
        RECT 108.705 59.655 113.120 60.585 ;
        RECT 131.170 60.360 133.130 60.590 ;
        RECT 130.890 60.070 131.120 60.200 ;
        RECT 104.190 53.520 104.600 53.800 ;
        RECT 103.660 52.500 104.910 53.520 ;
        RECT 98.140 52.330 99.120 52.370 ;
        RECT 98.130 51.360 102.660 52.330 ;
        RECT 108.705 52.310 109.635 59.655 ;
        RECT 112.190 58.260 113.120 59.655 ;
        RECT 110.570 56.530 111.250 57.310 ;
        RECT 111.990 57.230 121.630 58.260 ;
        RECT 111.800 57.000 121.800 57.230 ;
        RECT 109.900 55.190 111.250 56.530 ;
        RECT 110.570 54.640 111.250 55.190 ;
        RECT 111.410 54.990 111.640 56.950 ;
        RECT 111.990 56.890 121.630 57.000 ;
        RECT 121.960 56.740 122.190 56.950 ;
        RECT 121.960 55.130 124.860 56.740 ;
        RECT 111.980 54.940 121.600 55.030 ;
        RECT 121.960 54.990 122.190 55.130 ;
        RECT 111.800 54.710 121.800 54.940 ;
        RECT 111.980 53.660 121.600 54.710 ;
        RECT 123.100 53.915 124.850 55.130 ;
        RECT 107.850 52.300 109.710 52.310 ;
        RECT 98.140 51.290 99.120 51.360 ;
        RECT 103.120 51.280 109.710 52.300 ;
        RECT 107.850 51.270 109.710 51.280 ;
        RECT 108.670 45.740 109.710 51.270 ;
        RECT 120.710 51.740 121.520 53.660 ;
        RECT 123.070 52.165 124.880 53.915 ;
        RECT 129.970 51.740 131.150 60.070 ;
        RECT 120.710 50.330 131.150 51.740 ;
        RECT 120.710 50.280 130.660 50.330 ;
        RECT 120.710 48.430 121.520 50.280 ;
        RECT 130.890 50.200 131.120 50.330 ;
        RECT 131.290 50.040 132.950 60.360 ;
        RECT 133.180 60.040 133.410 60.200 ;
        RECT 133.090 51.555 134.240 60.040 ;
        RECT 133.090 50.565 140.620 51.555 ;
        RECT 133.090 50.350 134.240 50.565 ;
        RECT 133.180 50.200 133.410 50.350 ;
        RECT 131.170 49.810 133.130 50.040 ;
        RECT 131.290 49.780 132.950 49.810 ;
        RECT 131.040 48.480 133.190 49.600 ;
        RECT 139.630 49.190 140.620 50.565 ;
        RECT 147.510 49.190 147.990 49.220 ;
        RECT 139.630 48.710 147.990 49.190 ;
        RECT 110.570 46.650 111.350 47.420 ;
        RECT 112.040 47.390 121.710 48.430 ;
        RECT 131.610 47.770 132.610 48.480 ;
        RECT 111.880 47.160 121.880 47.390 ;
        RECT 102.650 44.740 109.710 45.740 ;
        RECT 109.850 45.580 111.350 46.650 ;
        RECT 110.570 44.820 111.350 45.580 ;
        RECT 111.490 45.150 111.720 47.110 ;
        RECT 112.040 47.030 121.710 47.160 ;
        RECT 122.040 46.960 122.270 47.110 ;
        RECT 123.930 46.960 124.690 46.990 ;
        RECT 122.010 45.920 124.690 46.960 ;
        RECT 122.010 45.890 135.380 45.920 ;
        RECT 111.980 45.100 121.770 45.330 ;
        RECT 122.010 45.270 136.060 45.890 ;
        RECT 122.040 45.150 122.270 45.270 ;
        RECT 111.880 44.870 121.880 45.100 ;
        RECT 123.930 45.080 136.060 45.270 ;
        RECT 108.670 43.880 109.710 44.740 ;
        RECT 108.640 42.840 109.740 43.880 ;
        RECT 111.980 43.690 121.770 44.870 ;
        RECT 112.130 42.320 113.110 43.690 ;
        RECT 107.020 41.340 113.110 42.320 ;
        RECT 107.020 40.370 108.000 41.340 ;
        RECT 103.910 39.370 108.000 40.370 ;
        RECT 108.640 39.610 113.100 40.650 ;
        RECT 112.060 39.430 113.100 39.610 ;
        RECT 103.910 37.110 104.910 39.370 ;
        RECT 98.280 33.230 99.140 33.250 ;
        RECT 98.240 32.940 102.340 33.230 ;
        RECT 107.020 33.120 108.000 39.370 ;
        RECT 110.620 37.750 111.350 38.490 ;
        RECT 112.040 38.430 121.810 39.430 ;
        RECT 111.880 38.200 121.880 38.430 ;
        RECT 109.710 36.690 111.350 37.750 ;
        RECT 110.620 35.850 111.350 36.690 ;
        RECT 111.490 36.190 111.720 38.150 ;
        RECT 112.040 38.010 121.810 38.200 ;
        RECT 122.040 38.000 122.270 38.150 ;
        RECT 123.930 38.000 124.690 45.080 ;
        RECT 129.750 43.250 130.030 43.270 ;
        RECT 112.080 36.140 121.760 36.350 ;
        RECT 122.010 36.300 124.690 38.000 ;
        RECT 128.060 43.210 130.030 43.250 ;
        RECT 128.060 42.930 133.270 43.210 ;
        RECT 128.060 42.760 130.030 42.930 ;
        RECT 128.060 37.825 128.640 42.760 ;
        RECT 128.930 41.320 129.410 42.340 ;
        RECT 129.750 41.700 130.030 42.760 ;
        RECT 128.930 40.960 129.450 41.320 ;
        RECT 128.950 40.580 129.450 40.960 ;
        RECT 128.930 40.120 129.450 40.580 ;
        RECT 128.950 39.160 129.450 40.120 ;
        RECT 129.010 39.110 129.450 39.160 ;
        RECT 130.520 38.660 130.860 41.680 ;
        RECT 131.650 39.870 132.130 42.340 ;
        RECT 131.640 39.320 132.130 39.870 ;
        RECT 132.990 39.380 133.270 42.930 ;
        RECT 134.940 42.340 135.410 43.910 ;
        RECT 134.930 40.960 135.410 42.340 ;
        RECT 135.720 41.710 136.050 45.080 ;
        RECT 137.650 41.880 138.130 42.340 ;
        RECT 134.940 40.580 135.410 40.960 ;
        RECT 134.930 40.120 135.410 40.580 ;
        RECT 134.940 40.110 135.410 40.120 ;
        RECT 136.580 39.380 136.860 41.600 ;
        RECT 137.650 40.960 138.140 41.880 ;
        RECT 137.660 40.580 138.140 40.960 ;
        RECT 137.650 40.120 138.140 40.580 ;
        RECT 131.640 39.270 132.120 39.320 ;
        RECT 132.990 39.100 136.860 39.380 ;
        RECT 137.660 39.240 138.140 40.120 ;
        RECT 139.630 41.875 140.620 48.710 ;
        RECT 147.510 48.680 147.990 48.710 ;
        RECT 144.500 47.040 146.070 47.060 ;
        RECT 146.780 47.040 148.350 47.060 ;
        RECT 149.060 47.040 150.630 47.060 ;
        RECT 151.370 47.040 152.940 47.070 ;
        RECT 144.300 46.810 146.260 47.040 ;
        RECT 146.590 46.810 148.550 47.040 ;
        RECT 148.880 46.810 150.840 47.040 ;
        RECT 151.170 46.810 153.130 47.040 ;
        RECT 144.020 46.540 144.250 46.650 ;
        RECT 142.950 41.875 144.320 46.540 ;
        RECT 139.630 40.885 144.320 41.875 ;
        RECT 137.660 39.180 138.130 39.240 ;
        RECT 130.420 38.410 131.000 38.660 ;
        RECT 131.180 38.590 131.650 38.640 ;
        RECT 122.040 36.190 122.270 36.300 ;
        RECT 123.930 36.290 124.690 36.300 ;
        RECT 111.880 35.910 121.880 36.140 ;
        RECT 112.080 34.700 121.760 35.910 ;
        RECT 98.240 32.350 102.585 32.940 ;
        RECT 98.240 32.120 102.340 32.350 ;
        RECT 103.140 32.170 108.010 33.120 ;
        RECT 120.780 32.980 121.760 34.700 ;
        RECT 127.035 33.715 128.785 37.825 ;
        RECT 130.340 37.750 131.000 38.410 ;
        RECT 130.420 37.480 131.000 37.750 ;
        RECT 131.170 37.630 131.650 38.590 ;
        RECT 131.180 37.590 131.650 37.630 ;
        RECT 130.420 37.230 131.040 37.480 ;
        RECT 130.210 36.230 131.210 37.230 ;
        RECT 131.560 35.170 132.480 35.660 ;
        RECT 130.860 33.640 133.180 35.170 ;
        RECT 131.170 33.260 133.130 33.490 ;
        RECT 130.890 32.980 131.120 33.100 ;
        RECT 103.830 30.520 105.270 32.030 ;
        RECT 104.180 30.110 105.030 30.520 ;
        RECT 107.020 24.740 108.000 32.170 ;
        RECT 120.780 32.020 131.180 32.980 ;
        RECT 120.780 30.690 121.760 32.020 ;
        RECT 112.060 30.330 121.760 30.690 ;
        RECT 112.060 29.470 121.730 30.330 ;
        RECT 110.630 28.690 111.330 29.470 ;
        RECT 111.880 29.240 121.880 29.470 ;
        RECT 109.720 27.720 111.330 28.690 ;
        RECT 110.630 26.980 111.330 27.720 ;
        RECT 111.490 27.230 111.720 29.190 ;
        RECT 112.060 29.090 121.730 29.240 ;
        RECT 122.040 29.080 122.270 29.190 ;
        RECT 123.100 29.080 124.850 31.155 ;
        RECT 112.030 27.180 121.740 27.340 ;
        RECT 121.970 27.330 124.850 29.080 ;
        RECT 122.040 27.230 122.270 27.330 ;
        RECT 111.880 26.950 121.880 27.180 ;
        RECT 112.030 25.810 121.740 26.950 ;
        RECT 112.080 24.740 113.060 25.810 ;
        RECT 107.020 23.760 113.060 24.740 ;
        RECT 129.890 23.170 131.180 32.020 ;
        RECT 130.890 23.100 131.120 23.170 ;
        RECT 131.320 22.940 133.020 33.260 ;
        RECT 133.180 32.980 133.410 33.100 ;
        RECT 133.160 32.940 134.270 32.980 ;
        RECT 139.630 32.940 140.620 40.885 ;
        RECT 142.950 36.830 144.320 40.885 ;
        RECT 144.500 46.370 146.070 46.810 ;
        RECT 144.500 36.910 145.870 46.370 ;
        RECT 146.310 46.220 146.540 46.650 ;
        RECT 146.780 46.420 148.350 46.810 ;
        RECT 146.780 46.370 148.060 46.420 ;
        RECT 146.120 42.000 146.740 46.220 ;
        RECT 146.100 40.380 146.740 42.000 ;
        RECT 146.120 37.250 146.740 40.380 ;
        RECT 144.020 36.650 144.250 36.830 ;
        RECT 144.500 36.490 146.070 36.910 ;
        RECT 146.310 36.650 146.540 37.250 ;
        RECT 147.060 36.910 148.060 46.370 ;
        RECT 148.600 46.210 148.830 46.650 ;
        RECT 149.060 46.420 150.630 46.810 ;
        RECT 149.290 46.410 150.630 46.420 ;
        RECT 148.430 44.750 149.010 46.210 ;
        RECT 148.430 42.900 149.020 44.750 ;
        RECT 148.430 37.200 149.010 42.900 ;
        RECT 146.780 36.830 148.060 36.910 ;
        RECT 146.780 36.490 148.350 36.830 ;
        RECT 148.600 36.650 148.830 37.200 ;
        RECT 149.290 36.910 150.310 46.410 ;
        RECT 150.890 46.120 151.120 46.650 ;
        RECT 151.370 46.410 152.940 46.810 ;
        RECT 151.720 46.400 152.940 46.410 ;
        RECT 150.690 42.020 151.350 46.120 ;
        RECT 150.650 40.360 151.350 42.020 ;
        RECT 150.690 37.270 151.350 40.360 ;
        RECT 149.290 36.830 150.630 36.910 ;
        RECT 149.060 36.490 150.630 36.830 ;
        RECT 150.890 36.650 151.120 37.270 ;
        RECT 151.720 36.910 152.740 46.400 ;
        RECT 153.180 46.170 153.410 46.650 ;
        RECT 153.010 37.280 153.480 46.170 ;
        RECT 153.620 40.270 154.250 42.130 ;
        RECT 151.370 36.850 152.740 36.910 ;
        RECT 151.370 36.490 152.940 36.850 ;
        RECT 153.180 36.650 153.410 37.280 ;
        RECT 144.300 36.260 146.260 36.490 ;
        RECT 146.590 36.260 148.550 36.490 ;
        RECT 148.880 36.260 150.840 36.490 ;
        RECT 151.170 36.260 153.130 36.490 ;
        RECT 144.500 35.120 146.070 36.260 ;
        RECT 146.780 35.120 148.350 36.260 ;
        RECT 149.060 35.120 150.630 36.260 ;
        RECT 151.370 35.130 152.940 36.260 ;
        RECT 145.035 34.015 145.745 35.120 ;
        RECT 147.205 34.015 147.915 35.120 ;
        RECT 149.425 34.015 150.135 35.120 ;
        RECT 151.795 34.015 152.505 35.130 ;
        RECT 145.035 33.305 152.505 34.015 ;
        RECT 133.160 31.950 140.620 32.940 ;
        RECT 133.160 23.210 134.270 31.950 ;
        RECT 133.180 23.100 133.410 23.210 ;
        RECT 131.170 22.710 133.130 22.940 ;
        RECT 142.740 22.885 143.450 22.900 ;
        RECT 146.650 22.885 147.150 22.910 ;
        RECT 150.305 22.890 151.015 33.305 ;
        RECT 150.305 22.885 151.020 22.890 ;
        RECT 131.320 22.680 133.020 22.710 ;
        RECT 132.100 21.050 132.880 22.680 ;
        RECT 139.155 22.330 151.020 22.885 ;
        RECT 139.155 22.175 151.015 22.330 ;
        RECT 131.860 20.050 135.170 21.050 ;
        RECT 113.660 19.080 114.700 19.440 ;
        RECT 110.590 17.590 111.550 18.210 ;
        RECT 113.590 17.830 115.020 19.080 ;
        RECT 139.155 17.670 139.865 22.175 ;
        RECT 142.740 21.230 143.450 22.175 ;
        RECT 142.740 20.220 144.210 21.230 ;
        RECT 145.125 21.220 145.835 22.175 ;
        RECT 146.650 22.130 147.150 22.175 ;
        RECT 144.980 20.410 146.630 21.220 ;
        RECT 147.425 21.210 148.135 22.175 ;
        RECT 145.170 20.220 146.630 20.410 ;
        RECT 147.420 20.220 148.730 21.210 ;
        RECT 150.305 21.200 151.015 22.175 ;
        RECT 149.520 20.220 151.230 21.200 ;
        RECT 142.530 19.990 144.490 20.220 ;
        RECT 144.820 19.990 146.780 20.220 ;
        RECT 147.110 19.990 149.070 20.220 ;
        RECT 149.400 19.990 151.360 20.220 ;
        RECT 142.250 19.670 142.480 19.830 ;
        RECT 141.350 17.670 142.550 19.670 ;
        RECT 110.590 17.070 114.990 17.590 ;
        RECT 134.850 17.480 142.550 17.670 ;
        RECT 134.795 17.230 142.550 17.480 ;
        RECT 110.590 16.470 111.550 17.070 ;
        RECT 134.850 17.050 142.550 17.230 ;
        RECT 141.350 14.970 142.550 17.050 ;
        RECT 142.740 19.620 144.210 19.990 ;
        RECT 142.740 15.090 144.200 19.620 ;
        RECT 144.540 19.310 144.770 19.830 ;
        RECT 145.170 19.720 146.630 19.990 ;
        RECT 146.830 19.720 147.060 19.830 ;
        RECT 144.390 15.380 144.920 19.310 ;
        RECT 142.250 14.830 142.480 14.970 ;
        RECT 142.740 14.670 144.370 15.090 ;
        RECT 144.540 14.830 144.770 15.380 ;
        RECT 145.170 15.090 146.480 19.720 ;
        RECT 146.820 19.550 147.070 19.720 ;
        RECT 147.420 19.700 148.730 19.990 ;
        RECT 146.670 15.160 147.110 19.550 ;
        RECT 144.980 14.930 146.480 15.090 ;
        RECT 146.820 15.000 147.070 15.160 ;
        RECT 147.380 15.070 148.730 19.700 ;
        RECT 149.120 19.310 149.350 19.830 ;
        RECT 149.520 19.790 151.230 19.990 ;
        RECT 149.520 19.630 151.020 19.790 ;
        RECT 148.970 17.920 149.540 19.310 ;
        RECT 148.950 16.790 149.540 17.920 ;
        RECT 148.970 15.410 149.540 16.790 ;
        RECT 144.980 14.670 146.630 14.930 ;
        RECT 146.830 14.830 147.060 15.000 ;
        RECT 147.380 14.960 148.910 15.070 ;
        RECT 147.230 14.670 148.910 14.960 ;
        RECT 149.120 14.830 149.350 15.410 ;
        RECT 149.710 15.070 151.020 19.630 ;
        RECT 151.410 19.610 151.640 19.830 ;
        RECT 151.290 15.070 151.730 19.610 ;
        RECT 149.520 14.870 151.020 15.070 ;
        RECT 149.520 14.670 151.230 14.870 ;
        RECT 151.410 14.830 151.640 15.070 ;
        RECT 151.870 14.850 152.480 18.430 ;
        RECT 142.530 14.440 144.490 14.670 ;
        RECT 144.820 14.440 146.780 14.670 ;
        RECT 147.110 14.440 149.070 14.670 ;
        RECT 149.400 14.440 151.360 14.670 ;
        RECT 142.740 14.420 144.370 14.440 ;
        RECT 144.980 14.410 146.630 14.440 ;
        RECT 147.230 14.410 148.910 14.440 ;
        RECT 149.520 14.410 151.230 14.440 ;
        RECT 154.170 11.520 155.170 13.490 ;
        RECT 128.580 7.150 129.580 9.120 ;
      LAYER met2 ;
        RECT 124.975 78.055 125.365 78.070 ;
        RECT 124.975 77.785 126.565 78.055 ;
        RECT 124.975 77.770 125.365 77.785 ;
        RECT 109.220 63.790 110.090 65.460 ;
        RECT 111.460 62.760 112.010 63.310 ;
        RECT 109.850 55.240 110.690 56.480 ;
        RECT 104.140 53.270 104.650 53.750 ;
        RECT 98.090 51.340 99.170 52.320 ;
        RECT 102.680 45.740 103.680 45.770 ;
        RECT 101.465 44.740 103.680 45.740 ;
        RECT 109.800 45.630 110.790 46.600 ;
        RECT 102.680 44.710 103.680 44.740 ;
        RECT 108.670 39.580 109.710 43.910 ;
        RECT 103.910 38.140 104.910 38.185 ;
        RECT 103.880 37.140 104.940 38.140 ;
        RECT 103.910 37.095 104.910 37.140 ;
        RECT 109.660 36.740 110.850 37.700 ;
        RECT 123.100 35.495 124.850 53.945 ;
        RECT 126.295 37.005 126.565 77.785 ;
        RECT 149.630 64.310 151.050 64.980 ;
        RECT 151.760 64.330 152.440 64.980 ;
        RECT 148.440 49.190 149.090 49.230 ;
        RECT 153.040 49.190 153.520 49.230 ;
        RECT 131.560 47.820 132.660 48.880 ;
        RECT 147.480 48.710 153.520 49.190 ;
        RECT 148.440 44.700 149.090 48.710 ;
        RECT 153.040 44.780 153.520 48.710 ;
        RECT 134.890 43.220 135.460 43.860 ;
        RECT 148.390 42.960 149.090 44.700 ;
        RECT 152.980 42.990 153.530 44.780 ;
        RECT 148.390 42.950 149.070 42.960 ;
        RECT 146.050 40.430 146.790 41.950 ;
        RECT 150.600 40.410 151.360 41.970 ;
        RECT 153.520 40.320 154.300 42.080 ;
        RECT 128.960 39.160 129.500 39.790 ;
        RECT 131.590 39.320 132.170 39.820 ;
        RECT 137.610 39.230 138.180 39.760 ;
        RECT 131.130 37.640 131.700 38.590 ;
        RECT 130.585 37.005 130.855 37.055 ;
        RECT 126.295 36.735 130.855 37.005 ;
        RECT 130.585 36.685 130.855 36.735 ;
        RECT 123.100 33.745 128.815 35.495 ;
        RECT 131.510 34.820 132.530 35.610 ;
        RECT 98.230 32.230 99.190 33.200 ;
        RECT 123.100 31.125 124.850 33.745 ;
        RECT 104.130 30.160 105.080 31.020 ;
        RECT 123.070 29.375 124.880 31.125 ;
        RECT 109.670 27.770 110.810 28.640 ;
        RECT 146.640 22.860 147.150 22.900 ;
        RECT 146.600 22.180 147.200 22.860 ;
        RECT 150.490 22.360 151.770 22.860 ;
        RECT 134.140 21.050 135.140 21.080 ;
        RECT 134.140 20.050 136.355 21.050 ;
        RECT 134.140 20.020 135.140 20.050 ;
        RECT 113.610 18.520 114.750 19.390 ;
        RECT 146.640 19.250 147.150 22.180 ;
        RECT 146.620 18.530 147.150 19.250 ;
        RECT 151.270 19.130 151.770 22.360 ;
        RECT 151.240 18.490 151.780 19.130 ;
        RECT 110.540 16.520 111.600 18.160 ;
        RECT 144.360 16.820 144.940 17.850 ;
        RECT 148.900 16.840 149.540 17.870 ;
        RECT 151.840 16.300 152.460 17.010 ;
        RECT 154.170 13.460 155.170 14.605 ;
        RECT 154.140 12.460 155.200 13.460 ;
        RECT 128.580 9.090 129.580 9.975 ;
        RECT 128.550 8.090 129.610 9.090 ;
      LAYER met3 ;
        RECT 118.030 209.370 118.410 209.690 ;
        RECT 118.070 206.830 118.370 209.370 ;
        RECT 118.060 206.450 118.380 206.830 ;
        RECT 118.030 84.160 118.410 84.480 ;
        RECT 118.070 83.140 118.370 84.160 ;
        RECT 118.060 82.760 118.380 83.140 ;
        RECT 123.950 78.070 124.330 78.080 ;
        RECT 124.995 78.070 125.345 78.095 ;
        RECT 123.950 77.770 125.345 78.070 ;
        RECT 123.950 77.760 124.330 77.770 ;
        RECT 124.995 77.745 125.345 77.770 ;
        RECT 109.245 63.740 110.065 65.510 ;
        RECT 149.655 64.260 151.025 65.030 ;
        RECT 151.785 64.280 152.415 65.030 ;
        RECT 111.485 62.710 111.985 63.360 ;
        RECT 109.875 55.190 110.665 56.530 ;
        RECT 104.165 53.220 104.625 53.800 ;
        RECT 98.115 51.290 99.145 52.370 ;
        RECT 131.585 47.770 132.635 48.930 ;
        RECT 101.485 45.740 102.535 45.765 ;
        RECT 95.550 44.740 102.535 45.740 ;
        RECT 109.825 45.580 110.765 46.650 ;
        RECT 42.945 21.390 44.435 21.415 ;
        RECT 42.940 19.890 54.520 21.390 ;
        RECT 42.945 19.865 44.435 19.890 ;
        RECT 95.550 4.650 96.550 44.740 ;
        RECT 101.485 44.715 102.535 44.740 ;
        RECT 134.915 43.170 135.435 43.910 ;
        RECT 146.075 40.380 146.765 42.000 ;
        RECT 150.625 40.360 151.335 42.020 ;
        RECT 153.545 40.270 154.275 42.130 ;
        RECT 128.985 39.110 129.475 39.840 ;
        RECT 131.615 39.270 132.145 39.870 ;
        RECT 137.635 39.180 138.155 39.810 ;
        RECT 103.885 37.115 104.935 38.165 ;
        RECT 103.910 36.610 104.910 37.115 ;
        RECT 109.685 36.690 110.825 37.750 ;
        RECT 131.155 37.590 131.675 38.640 ;
        RECT 101.560 35.610 104.910 36.610 ;
        RECT 98.255 32.180 99.165 33.250 ;
        RECT 101.560 6.440 102.560 35.610 ;
        RECT 131.535 34.770 132.505 35.660 ;
        RECT 104.155 30.110 105.055 31.070 ;
        RECT 109.695 27.720 110.785 28.690 ;
        RECT 135.285 21.050 136.335 21.075 ;
        RECT 135.285 20.050 157.270 21.050 ;
        RECT 135.285 20.025 136.335 20.050 ;
        RECT 113.635 18.470 114.725 19.440 ;
        RECT 110.565 16.470 111.575 18.210 ;
        RECT 144.385 16.770 144.915 17.900 ;
        RECT 148.925 16.790 149.515 17.920 ;
        RECT 151.865 16.250 152.435 17.060 ;
        RECT 154.170 14.585 155.170 15.530 ;
        RECT 154.145 13.535 155.195 14.585 ;
        RECT 128.580 9.955 129.580 10.810 ;
        RECT 128.555 8.905 129.605 9.955 ;
        RECT 101.560 5.780 135.210 6.440 ;
        RECT 101.560 5.440 135.230 5.780 ;
        RECT 95.550 3.650 113.300 4.650 ;
        RECT 134.210 4.370 135.230 5.440 ;
        RECT 112.250 3.440 113.300 3.650 ;
        RECT 112.250 2.665 113.150 3.440 ;
        RECT 134.330 3.225 135.230 4.370 ;
        RECT 112.225 1.775 113.175 2.665 ;
        RECT 134.305 2.335 135.255 3.225 ;
        RECT 156.270 2.720 157.270 20.050 ;
        RECT 134.330 2.330 135.230 2.335 ;
        RECT 112.250 1.770 113.150 1.775 ;
      LAYER met4 ;
        RECT 3.980 224.760 3.990 225.250 ;
        RECT 3.980 223.750 4.280 224.760 ;
        RECT 7.670 223.750 7.970 224.760 ;
        RECT 11.350 223.750 11.650 224.760 ;
        RECT 15.030 223.750 15.330 224.760 ;
        RECT 18.710 223.750 19.010 224.760 ;
        RECT 22.390 223.750 22.690 224.760 ;
        RECT 26.070 223.750 26.370 224.760 ;
        RECT 29.750 223.750 30.050 224.760 ;
        RECT 33.430 223.750 33.730 224.760 ;
        RECT 37.110 223.750 37.410 224.760 ;
        RECT 40.790 223.750 41.090 224.760 ;
        RECT 44.470 223.750 44.770 224.760 ;
        RECT 48.150 223.750 48.450 224.760 ;
        RECT 51.830 223.750 52.130 224.760 ;
        RECT 55.510 223.750 55.810 224.760 ;
        RECT 59.190 223.750 59.490 224.760 ;
        RECT 62.870 223.750 63.170 224.760 ;
        RECT 66.550 223.750 66.850 224.760 ;
        RECT 70.230 223.750 70.530 224.760 ;
        RECT 73.910 223.750 74.210 224.760 ;
        RECT 77.590 223.750 77.890 224.760 ;
        RECT 81.270 223.750 81.570 224.760 ;
        RECT 84.950 223.750 85.250 224.760 ;
        RECT 88.630 223.750 88.930 224.760 ;
        RECT 3.980 223.450 88.930 223.750 ;
        RECT 5.480 223.420 6.980 223.450 ;
        RECT 15.030 223.410 15.330 223.450 ;
        RECT 18.710 223.440 22.710 223.450 ;
        RECT 26.070 223.420 26.370 223.450 ;
        RECT 29.750 223.400 30.050 223.450 ;
        RECT 44.470 223.420 44.770 223.450 ;
        RECT 2.500 219.050 2.520 220.550 ;
        RECT 45.230 220.110 45.530 223.450 ;
        RECT 51.830 223.420 52.130 223.450 ;
        RECT 55.510 223.440 55.810 223.450 ;
        RECT 59.190 223.440 59.490 223.450 ;
        RECT 62.870 223.390 63.170 223.450 ;
        RECT 45.230 219.810 49.000 220.110 ;
        RECT 84.950 218.190 85.250 223.450 ;
        RECT 118.070 209.695 118.370 224.760 ;
        RECT 118.055 209.365 118.385 209.695 ;
        RECT 118.055 206.475 118.385 206.805 ;
        RECT 118.070 84.485 118.370 206.475 ;
        RECT 118.055 84.155 118.385 84.485 ;
        RECT 118.055 82.785 118.385 83.115 ;
        RECT 118.070 78.070 118.370 82.785 ;
        RECT 123.975 78.070 124.305 78.085 ;
        RECT 117.980 77.770 124.305 78.070 ;
        RECT 118.070 77.250 118.370 77.770 ;
        RECT 123.975 77.755 124.305 77.770 ;
        RECT 50.500 71.880 149.390 71.980 ;
        RECT 50.500 70.940 149.400 71.880 ;
        RECT 50.500 70.480 149.390 70.940 ;
        RECT 109.265 65.450 110.045 65.465 ;
        RECT 97.830 63.810 110.045 65.450 ;
        RECT 52.985 21.390 54.495 21.395 ;
        RECT 97.830 21.390 99.470 63.810 ;
        RECT 109.265 63.785 110.045 63.810 ;
        RECT 147.890 65.370 149.390 70.480 ;
        RECT 147.890 63.870 153.360 65.370 ;
        RECT 110.720 60.810 112.220 63.340 ;
        RECT 109.270 60.100 132.930 60.810 ;
        RECT 147.890 60.100 150.680 63.870 ;
        RECT 109.270 59.310 150.680 60.100 ;
        RECT 109.270 54.550 110.770 59.310 ;
        RECT 103.400 53.050 110.770 54.550 ;
        RECT 109.270 37.705 110.770 53.050 ;
        RECT 131.430 58.600 150.680 59.310 ;
        RECT 131.430 48.340 132.930 58.600 ;
        RECT 131.430 46.840 138.710 48.340 ;
        RECT 127.890 42.720 135.990 44.360 ;
        RECT 109.270 36.735 110.805 37.705 ;
        RECT 109.270 31.370 110.770 36.735 ;
        RECT 103.940 29.870 110.770 31.370 ;
        RECT 2.500 19.890 44.440 21.390 ;
        RECT 52.985 19.890 99.470 21.390 ;
        RECT 109.270 21.650 110.770 29.870 ;
        RECT 109.270 20.150 114.800 21.650 ;
        RECT 52.985 19.885 54.495 19.890 ;
        RECT 93.510 19.690 95.010 19.890 ;
        RECT 97.830 18.150 99.470 19.890 ;
        RECT 113.300 18.900 114.800 20.150 ;
        RECT 113.655 18.515 114.705 18.900 ;
        RECT 110.585 18.150 111.555 18.165 ;
        RECT 97.830 16.515 111.555 18.150 ;
        RECT 97.830 16.510 111.420 16.515 ;
        RECT 107.700 12.980 109.340 16.510 ;
        RECT 127.890 12.980 129.530 42.720 ;
        RECT 131.570 39.270 132.590 39.880 ;
        RECT 131.590 38.595 132.590 39.270 ;
        RECT 131.175 37.635 132.590 38.595 ;
        RECT 131.570 36.140 132.590 37.635 ;
        RECT 137.210 36.140 138.710 46.840 ;
        RECT 149.180 41.975 150.680 58.600 ;
        RECT 146.095 41.660 146.745 41.955 ;
        RECT 149.180 41.660 151.315 41.975 ;
        RECT 153.565 41.660 154.255 42.085 ;
        RECT 144.840 40.160 155.170 41.660 ;
        RECT 131.000 34.640 138.710 36.140 ;
        RECT 144.405 17.670 144.895 17.855 ;
        RECT 148.945 17.670 149.495 17.875 ;
        RECT 153.670 17.670 155.170 40.160 ;
        RECT 143.440 16.170 155.170 17.670 ;
        RECT 154.170 15.505 155.170 16.170 ;
        RECT 154.165 14.495 155.175 15.505 ;
        RECT 107.700 12.470 129.530 12.980 ;
        RECT 107.700 11.340 129.580 12.470 ;
        RECT 128.580 10.785 129.580 11.340 ;
        RECT 128.575 9.775 129.585 10.785 ;
        RECT 112.250 1.000 113.150 2.670 ;
        RECT 134.330 1.000 135.230 3.230 ;
        RECT 156.265 2.745 157.275 3.755 ;
        RECT 156.270 1.000 157.270 2.745 ;
        RECT 156.270 0.030 156.410 1.000 ;
  END
END tt_um_brucemack_sb_mixer
END LIBRARY

