VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_devinatkin_dual_oscillator
  CLASS BLOCK ;
  FOREIGN tt_um_devinatkin_dual_oscillator ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.000000 ;
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 108.000000 ;
    ANTENNADIFFAREA 225.588425 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  OBS
      LAYER pwell ;
        RECT 89.360 152.840 131.460 155.800 ;
        RECT 89.350 150.850 107.310 152.840 ;
        RECT 89.370 16.065 93.150 146.860 ;
      LAYER nwell ;
        RECT 93.150 56.490 102.050 146.860 ;
      LAYER pwell ;
        RECT 102.050 56.490 105.830 146.860 ;
        RECT 105.850 146.610 115.070 146.860 ;
        RECT 105.850 132.990 131.240 146.610 ;
      LAYER nwell ;
        RECT 131.250 132.990 148.350 146.860 ;
      LAYER pwell ;
        RECT 115.070 132.980 148.350 132.990 ;
        RECT 105.850 126.210 112.950 132.980 ;
      LAYER nwell ;
        RECT 112.950 130.520 125.300 132.980 ;
      LAYER pwell ;
        RECT 125.300 130.520 148.350 132.980 ;
      LAYER nwell ;
        RECT 112.950 126.210 125.290 130.520 ;
      LAYER pwell ;
        RECT 105.840 108.940 114.040 126.210 ;
      LAYER nwell ;
        RECT 114.040 108.940 125.290 126.210 ;
      LAYER pwell ;
        RECT 125.290 108.950 148.350 130.520 ;
        RECT 105.850 108.690 115.070 108.940 ;
        RECT 105.850 95.070 131.240 108.690 ;
      LAYER nwell ;
        RECT 131.250 95.070 148.350 108.940 ;
      LAYER pwell ;
        RECT 115.070 95.060 148.350 95.070 ;
        RECT 105.850 88.290 112.950 95.060 ;
      LAYER nwell ;
        RECT 112.950 92.600 125.300 95.060 ;
      LAYER pwell ;
        RECT 125.300 92.600 148.350 95.060 ;
      LAYER nwell ;
        RECT 112.950 88.290 125.290 92.600 ;
      LAYER pwell ;
        RECT 105.840 71.020 114.040 88.290 ;
      LAYER nwell ;
        RECT 114.040 71.020 125.290 88.290 ;
      LAYER pwell ;
        RECT 125.290 71.030 148.350 92.600 ;
      LAYER nwell ;
        RECT 93.150 16.065 97.600 56.490 ;
      LAYER li1 ;
        RECT 89.540 155.450 131.280 155.620 ;
        RECT 89.540 153.190 89.710 155.450 ;
        RECT 90.390 154.880 130.430 155.050 ;
        RECT 90.050 153.820 90.220 154.820 ;
        RECT 130.600 153.820 130.770 154.820 ;
        RECT 90.390 153.590 130.430 153.760 ;
        RECT 131.110 153.190 131.280 155.450 ;
        RECT 89.540 153.020 131.280 153.190 ;
        RECT 89.530 152.490 107.130 152.660 ;
        RECT 89.530 152.270 89.700 152.490 ;
        RECT 89.530 151.580 89.710 152.270 ;
        RECT 90.260 151.930 90.430 152.010 ;
        RECT 106.230 151.930 106.400 152.010 ;
        RECT 90.260 151.760 92.245 151.930 ;
        RECT 104.415 151.760 106.400 151.930 ;
        RECT 90.260 151.680 90.430 151.760 ;
        RECT 106.230 151.680 106.400 151.760 ;
        RECT 89.530 151.200 89.700 151.580 ;
        RECT 106.960 151.200 107.130 152.490 ;
        RECT 89.530 151.030 107.130 151.200 ;
        RECT 93.440 146.680 94.240 146.690 ;
        RECT 100.960 146.680 101.760 146.690 ;
        RECT 89.480 146.510 92.980 146.680 ;
        RECT 89.470 146.500 92.980 146.510 ;
        RECT 89.470 145.400 89.650 146.500 ;
        RECT 89.480 142.680 89.650 145.400 ;
        RECT 90.050 145.210 91.050 145.380 ;
        RECT 91.340 145.210 92.340 145.380 ;
        RECT 89.820 144.000 89.990 145.040 ;
        RECT 91.110 144.000 91.280 145.040 ;
        RECT 92.400 144.000 92.570 145.040 ;
        RECT 90.050 143.660 91.050 143.830 ;
        RECT 91.340 143.660 92.340 143.830 ;
        RECT 92.810 142.680 92.980 146.500 ;
        RECT 89.480 142.510 92.980 142.680 ;
        RECT 89.470 142.410 92.980 142.510 ;
        RECT 89.470 141.400 89.650 142.410 ;
        RECT 89.480 138.620 89.650 141.400 ;
        RECT 90.050 141.210 91.050 141.380 ;
        RECT 91.340 141.210 92.340 141.380 ;
        RECT 89.820 140.000 89.990 141.040 ;
        RECT 91.110 140.000 91.280 141.040 ;
        RECT 92.400 140.000 92.570 141.040 ;
        RECT 90.050 139.660 91.050 139.830 ;
        RECT 91.340 139.660 92.340 139.830 ;
        RECT 92.810 138.620 92.980 142.410 ;
        RECT 89.480 138.410 92.980 138.620 ;
        RECT 89.470 138.400 92.980 138.410 ;
        RECT 89.470 137.300 89.650 138.400 ;
        RECT 89.480 134.530 89.650 137.300 ;
        RECT 90.050 137.110 91.050 137.280 ;
        RECT 91.340 137.110 92.340 137.280 ;
        RECT 89.820 135.900 89.990 136.940 ;
        RECT 91.110 135.900 91.280 136.940 ;
        RECT 92.400 135.900 92.570 136.940 ;
        RECT 90.050 135.560 91.050 135.730 ;
        RECT 91.340 135.560 92.340 135.730 ;
        RECT 92.810 134.530 92.980 138.400 ;
        RECT 89.480 134.360 92.980 134.530 ;
        RECT 89.470 134.310 92.980 134.360 ;
        RECT 89.470 133.250 89.650 134.310 ;
        RECT 89.480 130.480 89.650 133.250 ;
        RECT 90.050 133.060 91.050 133.230 ;
        RECT 91.340 133.060 92.340 133.230 ;
        RECT 89.820 131.850 89.990 132.890 ;
        RECT 91.110 131.850 91.280 132.890 ;
        RECT 92.400 131.850 92.570 132.890 ;
        RECT 90.050 131.510 91.050 131.680 ;
        RECT 91.340 131.510 92.340 131.680 ;
        RECT 92.810 130.480 92.980 134.310 ;
        RECT 89.480 130.310 92.980 130.480 ;
        RECT 89.470 130.260 92.980 130.310 ;
        RECT 89.470 129.200 89.650 130.260 ;
        RECT 89.480 126.430 89.650 129.200 ;
        RECT 90.050 129.010 91.050 129.180 ;
        RECT 91.340 129.010 92.340 129.180 ;
        RECT 89.820 127.800 89.990 128.840 ;
        RECT 91.110 127.800 91.280 128.840 ;
        RECT 92.400 127.800 92.570 128.840 ;
        RECT 90.050 127.460 91.050 127.630 ;
        RECT 91.340 127.460 92.340 127.630 ;
        RECT 92.810 126.430 92.980 130.260 ;
        RECT 89.480 126.260 92.980 126.430 ;
        RECT 89.470 126.210 92.980 126.260 ;
        RECT 89.470 125.150 89.650 126.210 ;
        RECT 89.480 122.380 89.650 125.150 ;
        RECT 90.050 124.960 91.050 125.130 ;
        RECT 91.340 124.960 92.340 125.130 ;
        RECT 89.820 123.750 89.990 124.790 ;
        RECT 91.110 123.750 91.280 124.790 ;
        RECT 92.400 123.750 92.570 124.790 ;
        RECT 90.050 123.410 91.050 123.580 ;
        RECT 91.340 123.410 92.340 123.580 ;
        RECT 92.810 122.380 92.980 126.210 ;
        RECT 89.480 122.210 92.980 122.380 ;
        RECT 89.470 122.160 92.980 122.210 ;
        RECT 89.470 121.100 89.650 122.160 ;
        RECT 89.480 118.330 89.650 121.100 ;
        RECT 90.050 120.910 91.050 121.080 ;
        RECT 91.340 120.910 92.340 121.080 ;
        RECT 89.820 119.700 89.990 120.740 ;
        RECT 91.110 119.700 91.280 120.740 ;
        RECT 92.400 119.700 92.570 120.740 ;
        RECT 90.050 119.360 91.050 119.530 ;
        RECT 91.340 119.360 92.340 119.530 ;
        RECT 92.810 118.330 92.980 122.160 ;
        RECT 89.480 118.160 92.980 118.330 ;
        RECT 89.470 118.110 92.980 118.160 ;
        RECT 89.470 117.050 89.650 118.110 ;
        RECT 89.480 114.280 89.650 117.050 ;
        RECT 90.050 116.860 91.050 117.030 ;
        RECT 91.340 116.860 92.340 117.030 ;
        RECT 89.820 115.650 89.990 116.690 ;
        RECT 91.110 115.650 91.280 116.690 ;
        RECT 92.400 115.650 92.570 116.690 ;
        RECT 90.050 115.310 91.050 115.480 ;
        RECT 91.340 115.310 92.340 115.480 ;
        RECT 92.810 114.280 92.980 118.110 ;
        RECT 89.480 114.110 92.980 114.280 ;
        RECT 89.470 114.060 92.980 114.110 ;
        RECT 89.470 113.000 89.650 114.060 ;
        RECT 89.480 110.230 89.650 113.000 ;
        RECT 90.050 112.810 91.050 112.980 ;
        RECT 91.340 112.810 92.340 112.980 ;
        RECT 89.820 111.600 89.990 112.640 ;
        RECT 91.110 111.600 91.280 112.640 ;
        RECT 92.400 111.600 92.570 112.640 ;
        RECT 90.050 111.260 91.050 111.430 ;
        RECT 91.340 111.260 92.340 111.430 ;
        RECT 92.810 110.230 92.980 114.060 ;
        RECT 89.480 110.060 92.980 110.230 ;
        RECT 89.470 110.010 92.980 110.060 ;
        RECT 89.470 108.950 89.650 110.010 ;
        RECT 89.480 106.180 89.650 108.950 ;
        RECT 90.050 108.760 91.050 108.930 ;
        RECT 91.340 108.760 92.340 108.930 ;
        RECT 89.820 107.550 89.990 108.590 ;
        RECT 91.110 107.550 91.280 108.590 ;
        RECT 92.400 107.550 92.570 108.590 ;
        RECT 90.050 107.210 91.050 107.380 ;
        RECT 91.340 107.210 92.340 107.380 ;
        RECT 92.810 106.180 92.980 110.010 ;
        RECT 89.480 106.010 92.980 106.180 ;
        RECT 89.470 105.960 92.980 106.010 ;
        RECT 89.470 104.900 89.650 105.960 ;
        RECT 89.480 102.130 89.650 104.900 ;
        RECT 90.050 104.710 91.050 104.880 ;
        RECT 91.340 104.710 92.340 104.880 ;
        RECT 89.820 103.500 89.990 104.540 ;
        RECT 91.110 103.500 91.280 104.540 ;
        RECT 92.400 103.500 92.570 104.540 ;
        RECT 90.050 103.160 91.050 103.330 ;
        RECT 91.340 103.160 92.340 103.330 ;
        RECT 92.810 102.130 92.980 105.960 ;
        RECT 89.480 101.960 92.980 102.130 ;
        RECT 89.470 101.910 92.980 101.960 ;
        RECT 89.470 100.850 89.650 101.910 ;
        RECT 89.480 98.080 89.650 100.850 ;
        RECT 90.050 100.660 91.050 100.830 ;
        RECT 91.340 100.660 92.340 100.830 ;
        RECT 89.820 99.450 89.990 100.490 ;
        RECT 91.110 99.450 91.280 100.490 ;
        RECT 92.400 99.450 92.570 100.490 ;
        RECT 90.050 99.110 91.050 99.280 ;
        RECT 91.340 99.110 92.340 99.280 ;
        RECT 92.810 98.080 92.980 101.910 ;
        RECT 89.480 97.910 92.980 98.080 ;
        RECT 89.470 97.860 92.980 97.910 ;
        RECT 89.470 96.800 89.650 97.860 ;
        RECT 89.480 94.030 89.650 96.800 ;
        RECT 90.050 96.610 91.050 96.780 ;
        RECT 91.340 96.610 92.340 96.780 ;
        RECT 89.820 95.400 89.990 96.440 ;
        RECT 91.110 95.400 91.280 96.440 ;
        RECT 92.400 95.400 92.570 96.440 ;
        RECT 90.050 95.060 91.050 95.230 ;
        RECT 91.340 95.060 92.340 95.230 ;
        RECT 92.810 94.030 92.980 97.860 ;
        RECT 89.480 93.860 92.980 94.030 ;
        RECT 89.470 93.810 92.980 93.860 ;
        RECT 89.470 92.750 89.650 93.810 ;
        RECT 89.480 89.980 89.650 92.750 ;
        RECT 90.050 92.560 91.050 92.730 ;
        RECT 91.340 92.560 92.340 92.730 ;
        RECT 89.820 91.350 89.990 92.390 ;
        RECT 91.110 91.350 91.280 92.390 ;
        RECT 92.400 91.350 92.570 92.390 ;
        RECT 90.050 91.010 91.050 91.180 ;
        RECT 91.340 91.010 92.340 91.180 ;
        RECT 92.810 89.980 92.980 93.810 ;
        RECT 89.480 89.810 92.980 89.980 ;
        RECT 89.470 89.760 92.980 89.810 ;
        RECT 89.470 88.700 89.650 89.760 ;
        RECT 89.480 85.930 89.650 88.700 ;
        RECT 90.050 88.510 91.050 88.680 ;
        RECT 91.340 88.510 92.340 88.680 ;
        RECT 89.820 87.300 89.990 88.340 ;
        RECT 91.110 87.300 91.280 88.340 ;
        RECT 92.400 87.300 92.570 88.340 ;
        RECT 90.050 86.960 91.050 87.130 ;
        RECT 91.340 86.960 92.340 87.130 ;
        RECT 92.810 85.930 92.980 89.760 ;
        RECT 89.480 85.760 92.980 85.930 ;
        RECT 89.470 85.710 92.980 85.760 ;
        RECT 89.470 84.650 89.650 85.710 ;
        RECT 89.480 81.880 89.650 84.650 ;
        RECT 90.050 84.460 91.050 84.630 ;
        RECT 91.340 84.460 92.340 84.630 ;
        RECT 89.820 83.250 89.990 84.290 ;
        RECT 91.110 83.250 91.280 84.290 ;
        RECT 92.400 83.250 92.570 84.290 ;
        RECT 90.050 82.910 91.050 83.080 ;
        RECT 91.340 82.910 92.340 83.080 ;
        RECT 92.810 81.880 92.980 85.710 ;
        RECT 89.480 81.710 92.980 81.880 ;
        RECT 89.470 81.660 92.980 81.710 ;
        RECT 89.470 80.600 89.650 81.660 ;
        RECT 89.480 77.830 89.650 80.600 ;
        RECT 90.050 80.410 91.050 80.580 ;
        RECT 91.340 80.410 92.340 80.580 ;
        RECT 89.820 79.200 89.990 80.240 ;
        RECT 91.110 79.200 91.280 80.240 ;
        RECT 92.400 79.200 92.570 80.240 ;
        RECT 90.050 78.860 91.050 79.030 ;
        RECT 91.340 78.860 92.340 79.030 ;
        RECT 92.810 77.830 92.980 81.660 ;
        RECT 89.480 77.660 92.980 77.830 ;
        RECT 89.470 77.610 92.980 77.660 ;
        RECT 89.470 76.550 89.650 77.610 ;
        RECT 89.480 73.780 89.650 76.550 ;
        RECT 90.050 76.360 91.050 76.530 ;
        RECT 91.340 76.360 92.340 76.530 ;
        RECT 89.820 75.150 89.990 76.190 ;
        RECT 91.110 75.150 91.280 76.190 ;
        RECT 92.400 75.150 92.570 76.190 ;
        RECT 90.050 74.810 91.050 74.980 ;
        RECT 91.340 74.810 92.340 74.980 ;
        RECT 92.810 73.780 92.980 77.610 ;
        RECT 89.480 73.610 92.980 73.780 ;
        RECT 89.470 73.560 92.980 73.610 ;
        RECT 89.470 72.500 89.650 73.560 ;
        RECT 89.480 69.730 89.650 72.500 ;
        RECT 90.050 72.310 91.050 72.480 ;
        RECT 91.340 72.310 92.340 72.480 ;
        RECT 89.820 71.100 89.990 72.140 ;
        RECT 91.110 71.100 91.280 72.140 ;
        RECT 92.400 71.100 92.570 72.140 ;
        RECT 90.050 70.760 91.050 70.930 ;
        RECT 91.340 70.760 92.340 70.930 ;
        RECT 92.810 69.730 92.980 73.560 ;
        RECT 89.480 69.560 92.980 69.730 ;
        RECT 89.470 69.510 92.980 69.560 ;
        RECT 89.470 68.450 89.650 69.510 ;
        RECT 89.480 65.680 89.650 68.450 ;
        RECT 90.050 68.260 91.050 68.430 ;
        RECT 91.340 68.260 92.340 68.430 ;
        RECT 89.820 67.050 89.990 68.090 ;
        RECT 91.110 67.050 91.280 68.090 ;
        RECT 92.400 67.050 92.570 68.090 ;
        RECT 90.050 66.710 91.050 66.880 ;
        RECT 91.340 66.710 92.340 66.880 ;
        RECT 92.810 65.680 92.980 69.510 ;
        RECT 89.480 65.510 92.980 65.680 ;
        RECT 89.470 65.460 92.980 65.510 ;
        RECT 89.470 64.400 89.650 65.460 ;
        RECT 89.480 61.630 89.650 64.400 ;
        RECT 90.050 64.210 91.050 64.380 ;
        RECT 91.340 64.210 92.340 64.380 ;
        RECT 89.820 63.000 89.990 64.040 ;
        RECT 91.110 63.000 91.280 64.040 ;
        RECT 92.400 63.000 92.570 64.040 ;
        RECT 90.050 62.660 91.050 62.830 ;
        RECT 91.340 62.660 92.340 62.830 ;
        RECT 92.810 61.630 92.980 65.460 ;
        RECT 89.480 61.460 92.980 61.630 ;
        RECT 89.470 61.410 92.980 61.460 ;
        RECT 89.470 60.350 89.650 61.410 ;
        RECT 89.480 57.580 89.650 60.350 ;
        RECT 90.050 60.160 91.050 60.330 ;
        RECT 91.340 60.160 92.340 60.330 ;
        RECT 89.820 58.950 89.990 59.990 ;
        RECT 91.110 58.950 91.280 59.990 ;
        RECT 92.400 58.950 92.570 59.990 ;
        RECT 90.050 58.610 91.050 58.780 ;
        RECT 91.340 58.610 92.340 58.780 ;
        RECT 92.810 57.580 92.980 61.410 ;
        RECT 89.480 57.410 92.980 57.580 ;
        RECT 89.470 57.360 92.980 57.410 ;
        RECT 89.470 56.300 89.650 57.360 ;
        RECT 89.480 53.530 89.650 56.300 ;
        RECT 90.050 56.110 91.050 56.280 ;
        RECT 91.340 56.110 92.340 56.280 ;
        RECT 89.820 54.900 89.990 55.940 ;
        RECT 91.110 54.900 91.280 55.940 ;
        RECT 92.400 54.900 92.570 55.940 ;
        RECT 90.050 54.560 91.050 54.730 ;
        RECT 91.340 54.560 92.340 54.730 ;
        RECT 92.810 53.530 92.980 57.360 ;
        RECT 89.480 53.360 92.980 53.530 ;
        RECT 89.470 53.310 92.980 53.360 ;
        RECT 89.470 52.250 89.650 53.310 ;
        RECT 89.480 49.480 89.650 52.250 ;
        RECT 90.050 52.060 91.050 52.230 ;
        RECT 91.340 52.060 92.340 52.230 ;
        RECT 89.820 50.850 89.990 51.890 ;
        RECT 91.110 50.850 91.280 51.890 ;
        RECT 92.400 50.850 92.570 51.890 ;
        RECT 90.050 50.510 91.050 50.680 ;
        RECT 91.340 50.510 92.340 50.680 ;
        RECT 92.810 49.480 92.980 53.310 ;
        RECT 89.480 49.310 92.980 49.480 ;
        RECT 89.470 49.260 92.980 49.310 ;
        RECT 89.470 48.200 89.650 49.260 ;
        RECT 89.480 45.430 89.650 48.200 ;
        RECT 90.050 48.010 91.050 48.180 ;
        RECT 91.340 48.010 92.340 48.180 ;
        RECT 89.820 46.800 89.990 47.840 ;
        RECT 91.110 46.800 91.280 47.840 ;
        RECT 92.400 46.800 92.570 47.840 ;
        RECT 90.050 46.460 91.050 46.630 ;
        RECT 91.340 46.460 92.340 46.630 ;
        RECT 92.810 45.430 92.980 49.260 ;
        RECT 89.480 45.260 92.980 45.430 ;
        RECT 89.470 45.210 92.980 45.260 ;
        RECT 89.470 44.150 89.650 45.210 ;
        RECT 89.480 41.380 89.650 44.150 ;
        RECT 90.050 43.960 91.050 44.130 ;
        RECT 91.340 43.960 92.340 44.130 ;
        RECT 89.820 42.750 89.990 43.790 ;
        RECT 91.110 42.750 91.280 43.790 ;
        RECT 92.400 42.750 92.570 43.790 ;
        RECT 90.050 42.410 91.050 42.580 ;
        RECT 91.340 42.410 92.340 42.580 ;
        RECT 92.810 41.380 92.980 45.210 ;
        RECT 89.480 41.210 92.980 41.380 ;
        RECT 89.470 41.160 92.980 41.210 ;
        RECT 89.470 40.100 89.650 41.160 ;
        RECT 89.480 37.330 89.650 40.100 ;
        RECT 90.050 39.910 91.050 40.080 ;
        RECT 91.340 39.910 92.340 40.080 ;
        RECT 89.820 38.700 89.990 39.740 ;
        RECT 91.110 38.700 91.280 39.740 ;
        RECT 92.400 38.700 92.570 39.740 ;
        RECT 90.050 38.360 91.050 38.530 ;
        RECT 91.340 38.360 92.340 38.530 ;
        RECT 92.810 37.330 92.980 41.160 ;
        RECT 89.480 37.160 92.980 37.330 ;
        RECT 89.470 37.110 92.980 37.160 ;
        RECT 89.470 36.050 89.650 37.110 ;
        RECT 89.480 33.280 89.650 36.050 ;
        RECT 90.050 35.860 91.050 36.030 ;
        RECT 91.340 35.860 92.340 36.030 ;
        RECT 89.820 34.650 89.990 35.690 ;
        RECT 91.110 34.650 91.280 35.690 ;
        RECT 92.400 34.650 92.570 35.690 ;
        RECT 90.050 34.310 91.050 34.480 ;
        RECT 91.340 34.310 92.340 34.480 ;
        RECT 92.810 33.280 92.980 37.110 ;
        RECT 89.480 33.110 92.980 33.280 ;
        RECT 89.470 33.060 92.980 33.110 ;
        RECT 89.470 32.000 89.650 33.060 ;
        RECT 89.480 29.220 89.650 32.000 ;
        RECT 90.050 31.810 91.050 31.980 ;
        RECT 91.340 31.810 92.340 31.980 ;
        RECT 89.820 30.600 89.990 31.640 ;
        RECT 91.110 30.600 91.280 31.640 ;
        RECT 92.400 30.600 92.570 31.640 ;
        RECT 90.050 30.260 91.050 30.430 ;
        RECT 91.340 30.260 92.340 30.430 ;
        RECT 92.810 29.220 92.980 33.060 ;
        RECT 89.480 29.025 92.980 29.220 ;
        RECT 89.470 29.010 92.980 29.025 ;
        RECT 89.470 27.915 89.650 29.010 ;
        RECT 89.480 25.135 89.650 27.915 ;
        RECT 90.050 27.725 91.050 27.895 ;
        RECT 91.340 27.725 92.340 27.895 ;
        RECT 89.820 26.515 89.990 27.555 ;
        RECT 91.110 26.515 91.280 27.555 ;
        RECT 92.400 26.515 92.570 27.555 ;
        RECT 90.050 26.175 91.050 26.345 ;
        RECT 91.340 26.175 92.340 26.345 ;
        RECT 92.810 25.135 92.980 29.010 ;
        RECT 89.480 24.900 92.980 25.135 ;
        RECT 89.470 24.890 92.980 24.900 ;
        RECT 89.470 23.790 89.650 24.890 ;
        RECT 89.480 21.010 89.650 23.790 ;
        RECT 90.050 23.600 91.050 23.770 ;
        RECT 91.340 23.600 92.340 23.770 ;
        RECT 89.820 22.390 89.990 23.430 ;
        RECT 91.110 22.390 91.280 23.430 ;
        RECT 92.400 22.390 92.570 23.430 ;
        RECT 90.050 22.050 91.050 22.220 ;
        RECT 91.340 22.050 92.340 22.220 ;
        RECT 92.810 21.010 92.980 24.890 ;
        RECT 89.480 20.800 92.980 21.010 ;
        RECT 93.330 146.510 97.430 146.680 ;
        RECT 93.330 142.690 93.500 146.510 ;
        RECT 94.240 145.685 95.240 145.855 ;
        RECT 95.530 145.685 96.530 145.855 ;
        RECT 94.010 143.430 94.180 145.470 ;
        RECT 95.300 143.430 95.470 145.470 ;
        RECT 96.590 143.430 96.760 145.470 ;
        RECT 94.240 143.045 95.240 143.215 ;
        RECT 95.530 143.045 96.530 143.215 ;
        RECT 93.330 142.680 94.240 142.690 ;
        RECT 97.250 142.680 97.430 146.510 ;
        RECT 93.330 142.410 97.430 142.680 ;
        RECT 93.330 138.620 93.500 142.410 ;
        RECT 94.240 141.685 95.240 141.855 ;
        RECT 95.530 141.685 96.530 141.855 ;
        RECT 94.010 139.430 94.180 141.470 ;
        RECT 95.300 139.430 95.470 141.470 ;
        RECT 96.590 139.430 96.760 141.470 ;
        RECT 94.240 139.045 95.240 139.215 ;
        RECT 95.530 139.045 96.530 139.215 ;
        RECT 97.250 138.620 97.430 142.410 ;
        RECT 93.330 138.410 97.430 138.620 ;
        RECT 93.330 134.540 93.500 138.410 ;
        RECT 94.240 137.585 95.240 137.755 ;
        RECT 95.530 137.585 96.530 137.755 ;
        RECT 94.010 135.330 94.180 137.370 ;
        RECT 95.300 135.330 95.470 137.370 ;
        RECT 96.590 135.330 96.760 137.370 ;
        RECT 94.240 134.945 95.240 135.115 ;
        RECT 95.530 134.945 96.530 135.115 ;
        RECT 93.330 134.530 94.240 134.540 ;
        RECT 97.250 134.530 97.430 138.410 ;
        RECT 93.330 134.310 97.430 134.530 ;
        RECT 93.330 130.490 93.500 134.310 ;
        RECT 94.240 133.535 95.240 133.705 ;
        RECT 95.530 133.535 96.530 133.705 ;
        RECT 94.010 131.280 94.180 133.320 ;
        RECT 95.300 131.280 95.470 133.320 ;
        RECT 96.590 131.280 96.760 133.320 ;
        RECT 94.240 130.895 95.240 131.065 ;
        RECT 95.530 130.895 96.530 131.065 ;
        RECT 93.330 130.480 94.240 130.490 ;
        RECT 97.250 130.480 97.430 134.310 ;
        RECT 93.330 130.260 97.430 130.480 ;
        RECT 93.330 126.440 93.500 130.260 ;
        RECT 94.240 129.485 95.240 129.655 ;
        RECT 95.530 129.485 96.530 129.655 ;
        RECT 94.010 127.230 94.180 129.270 ;
        RECT 95.300 127.230 95.470 129.270 ;
        RECT 96.590 127.230 96.760 129.270 ;
        RECT 94.240 126.845 95.240 127.015 ;
        RECT 95.530 126.845 96.530 127.015 ;
        RECT 93.330 126.430 94.240 126.440 ;
        RECT 97.250 126.430 97.430 130.260 ;
        RECT 93.330 126.210 97.430 126.430 ;
        RECT 93.330 122.390 93.500 126.210 ;
        RECT 94.240 125.435 95.240 125.605 ;
        RECT 95.530 125.435 96.530 125.605 ;
        RECT 94.010 123.180 94.180 125.220 ;
        RECT 95.300 123.180 95.470 125.220 ;
        RECT 96.590 123.180 96.760 125.220 ;
        RECT 94.240 122.795 95.240 122.965 ;
        RECT 95.530 122.795 96.530 122.965 ;
        RECT 93.330 122.380 94.240 122.390 ;
        RECT 97.250 122.380 97.430 126.210 ;
        RECT 93.330 122.160 97.430 122.380 ;
        RECT 93.330 118.340 93.500 122.160 ;
        RECT 94.240 121.385 95.240 121.555 ;
        RECT 95.530 121.385 96.530 121.555 ;
        RECT 94.010 119.130 94.180 121.170 ;
        RECT 95.300 119.130 95.470 121.170 ;
        RECT 96.590 119.130 96.760 121.170 ;
        RECT 94.240 118.745 95.240 118.915 ;
        RECT 95.530 118.745 96.530 118.915 ;
        RECT 93.330 118.330 94.240 118.340 ;
        RECT 97.250 118.330 97.430 122.160 ;
        RECT 93.330 118.110 97.430 118.330 ;
        RECT 93.330 114.290 93.500 118.110 ;
        RECT 94.240 117.335 95.240 117.505 ;
        RECT 95.530 117.335 96.530 117.505 ;
        RECT 94.010 115.080 94.180 117.120 ;
        RECT 95.300 115.080 95.470 117.120 ;
        RECT 96.590 115.080 96.760 117.120 ;
        RECT 94.240 114.695 95.240 114.865 ;
        RECT 95.530 114.695 96.530 114.865 ;
        RECT 93.330 114.280 94.240 114.290 ;
        RECT 97.250 114.280 97.430 118.110 ;
        RECT 93.330 114.060 97.430 114.280 ;
        RECT 93.330 110.240 93.500 114.060 ;
        RECT 94.240 113.285 95.240 113.455 ;
        RECT 95.530 113.285 96.530 113.455 ;
        RECT 94.010 111.030 94.180 113.070 ;
        RECT 95.300 111.030 95.470 113.070 ;
        RECT 96.590 111.030 96.760 113.070 ;
        RECT 94.240 110.645 95.240 110.815 ;
        RECT 95.530 110.645 96.530 110.815 ;
        RECT 93.330 110.230 94.240 110.240 ;
        RECT 97.250 110.230 97.430 114.060 ;
        RECT 93.330 110.010 97.430 110.230 ;
        RECT 93.330 106.190 93.500 110.010 ;
        RECT 94.240 109.235 95.240 109.405 ;
        RECT 95.530 109.235 96.530 109.405 ;
        RECT 94.010 106.980 94.180 109.020 ;
        RECT 95.300 106.980 95.470 109.020 ;
        RECT 96.590 106.980 96.760 109.020 ;
        RECT 94.240 106.595 95.240 106.765 ;
        RECT 95.530 106.595 96.530 106.765 ;
        RECT 93.330 106.180 94.240 106.190 ;
        RECT 97.250 106.180 97.430 110.010 ;
        RECT 93.330 105.960 97.430 106.180 ;
        RECT 93.330 102.140 93.500 105.960 ;
        RECT 94.240 105.185 95.240 105.355 ;
        RECT 95.530 105.185 96.530 105.355 ;
        RECT 94.010 102.930 94.180 104.970 ;
        RECT 95.300 102.930 95.470 104.970 ;
        RECT 96.590 102.930 96.760 104.970 ;
        RECT 94.240 102.545 95.240 102.715 ;
        RECT 95.530 102.545 96.530 102.715 ;
        RECT 93.330 102.130 94.240 102.140 ;
        RECT 97.250 102.130 97.430 105.960 ;
        RECT 93.330 101.910 97.430 102.130 ;
        RECT 93.330 98.090 93.500 101.910 ;
        RECT 94.240 101.135 95.240 101.305 ;
        RECT 95.530 101.135 96.530 101.305 ;
        RECT 94.010 98.880 94.180 100.920 ;
        RECT 95.300 98.880 95.470 100.920 ;
        RECT 96.590 98.880 96.760 100.920 ;
        RECT 94.240 98.495 95.240 98.665 ;
        RECT 95.530 98.495 96.530 98.665 ;
        RECT 93.330 98.080 94.240 98.090 ;
        RECT 97.250 98.080 97.430 101.910 ;
        RECT 93.330 97.860 97.430 98.080 ;
        RECT 93.330 94.040 93.500 97.860 ;
        RECT 94.240 97.085 95.240 97.255 ;
        RECT 95.530 97.085 96.530 97.255 ;
        RECT 94.010 94.830 94.180 96.870 ;
        RECT 95.300 94.830 95.470 96.870 ;
        RECT 96.590 94.830 96.760 96.870 ;
        RECT 94.240 94.445 95.240 94.615 ;
        RECT 95.530 94.445 96.530 94.615 ;
        RECT 93.330 94.030 94.240 94.040 ;
        RECT 97.250 94.030 97.430 97.860 ;
        RECT 93.330 93.810 97.430 94.030 ;
        RECT 93.330 89.990 93.500 93.810 ;
        RECT 94.240 93.035 95.240 93.205 ;
        RECT 95.530 93.035 96.530 93.205 ;
        RECT 94.010 90.780 94.180 92.820 ;
        RECT 95.300 90.780 95.470 92.820 ;
        RECT 96.590 90.780 96.760 92.820 ;
        RECT 94.240 90.395 95.240 90.565 ;
        RECT 95.530 90.395 96.530 90.565 ;
        RECT 93.330 89.980 94.240 89.990 ;
        RECT 97.250 89.980 97.430 93.810 ;
        RECT 93.330 89.760 97.430 89.980 ;
        RECT 93.330 85.940 93.500 89.760 ;
        RECT 94.240 88.985 95.240 89.155 ;
        RECT 95.530 88.985 96.530 89.155 ;
        RECT 94.010 86.730 94.180 88.770 ;
        RECT 95.300 86.730 95.470 88.770 ;
        RECT 96.590 86.730 96.760 88.770 ;
        RECT 94.240 86.345 95.240 86.515 ;
        RECT 95.530 86.345 96.530 86.515 ;
        RECT 93.330 85.930 94.240 85.940 ;
        RECT 97.250 85.930 97.430 89.760 ;
        RECT 93.330 85.710 97.430 85.930 ;
        RECT 93.330 81.890 93.500 85.710 ;
        RECT 94.240 84.935 95.240 85.105 ;
        RECT 95.530 84.935 96.530 85.105 ;
        RECT 94.010 82.680 94.180 84.720 ;
        RECT 95.300 82.680 95.470 84.720 ;
        RECT 96.590 82.680 96.760 84.720 ;
        RECT 94.240 82.295 95.240 82.465 ;
        RECT 95.530 82.295 96.530 82.465 ;
        RECT 93.330 81.880 94.240 81.890 ;
        RECT 97.250 81.880 97.430 85.710 ;
        RECT 93.330 81.660 97.430 81.880 ;
        RECT 93.330 77.840 93.500 81.660 ;
        RECT 94.240 80.885 95.240 81.055 ;
        RECT 95.530 80.885 96.530 81.055 ;
        RECT 94.010 78.630 94.180 80.670 ;
        RECT 95.300 78.630 95.470 80.670 ;
        RECT 96.590 78.630 96.760 80.670 ;
        RECT 94.240 78.245 95.240 78.415 ;
        RECT 95.530 78.245 96.530 78.415 ;
        RECT 93.330 77.830 94.240 77.840 ;
        RECT 97.250 77.830 97.430 81.660 ;
        RECT 93.330 77.610 97.430 77.830 ;
        RECT 93.330 73.790 93.500 77.610 ;
        RECT 94.240 76.835 95.240 77.005 ;
        RECT 95.530 76.835 96.530 77.005 ;
        RECT 94.010 74.580 94.180 76.620 ;
        RECT 95.300 74.580 95.470 76.620 ;
        RECT 96.590 74.580 96.760 76.620 ;
        RECT 94.240 74.195 95.240 74.365 ;
        RECT 95.530 74.195 96.530 74.365 ;
        RECT 93.330 73.780 94.240 73.790 ;
        RECT 97.250 73.780 97.430 77.610 ;
        RECT 93.330 73.560 97.430 73.780 ;
        RECT 93.330 69.740 93.500 73.560 ;
        RECT 94.240 72.785 95.240 72.955 ;
        RECT 95.530 72.785 96.530 72.955 ;
        RECT 94.010 70.530 94.180 72.570 ;
        RECT 95.300 70.530 95.470 72.570 ;
        RECT 96.590 70.530 96.760 72.570 ;
        RECT 94.240 70.145 95.240 70.315 ;
        RECT 95.530 70.145 96.530 70.315 ;
        RECT 93.330 69.730 94.240 69.740 ;
        RECT 97.250 69.730 97.430 73.560 ;
        RECT 93.330 69.510 97.430 69.730 ;
        RECT 93.330 65.690 93.500 69.510 ;
        RECT 94.240 68.735 95.240 68.905 ;
        RECT 95.530 68.735 96.530 68.905 ;
        RECT 94.010 66.480 94.180 68.520 ;
        RECT 95.300 66.480 95.470 68.520 ;
        RECT 96.590 66.480 96.760 68.520 ;
        RECT 94.240 66.095 95.240 66.265 ;
        RECT 95.530 66.095 96.530 66.265 ;
        RECT 93.330 65.680 94.240 65.690 ;
        RECT 97.250 65.680 97.430 69.510 ;
        RECT 93.330 65.460 97.430 65.680 ;
        RECT 93.330 61.640 93.500 65.460 ;
        RECT 94.240 64.685 95.240 64.855 ;
        RECT 95.530 64.685 96.530 64.855 ;
        RECT 94.010 62.430 94.180 64.470 ;
        RECT 95.300 62.430 95.470 64.470 ;
        RECT 96.590 62.430 96.760 64.470 ;
        RECT 94.240 62.045 95.240 62.215 ;
        RECT 95.530 62.045 96.530 62.215 ;
        RECT 93.330 61.630 94.240 61.640 ;
        RECT 97.250 61.630 97.430 65.460 ;
        RECT 93.330 61.410 97.430 61.630 ;
        RECT 93.330 57.590 93.500 61.410 ;
        RECT 94.240 60.635 95.240 60.805 ;
        RECT 95.530 60.635 96.530 60.805 ;
        RECT 94.010 58.380 94.180 60.420 ;
        RECT 95.300 58.380 95.470 60.420 ;
        RECT 96.590 58.380 96.760 60.420 ;
        RECT 94.240 57.995 95.240 58.165 ;
        RECT 95.530 57.995 96.530 58.165 ;
        RECT 93.330 57.580 94.240 57.590 ;
        RECT 97.250 57.580 97.430 61.410 ;
        RECT 97.770 146.510 101.870 146.680 ;
        RECT 97.770 142.620 97.950 146.510 ;
        RECT 98.670 145.685 99.670 145.855 ;
        RECT 99.960 145.685 100.960 145.855 ;
        RECT 98.440 143.430 98.610 145.470 ;
        RECT 99.730 143.430 99.900 145.470 ;
        RECT 101.020 143.430 101.190 145.470 ;
        RECT 98.670 143.045 99.670 143.215 ;
        RECT 99.960 143.045 100.960 143.215 ;
        RECT 101.700 142.630 101.870 146.510 ;
        RECT 100.960 142.620 101.870 142.630 ;
        RECT 97.770 142.410 101.870 142.620 ;
        RECT 97.770 138.560 97.950 142.410 ;
        RECT 98.670 141.625 99.670 141.795 ;
        RECT 99.960 141.625 100.960 141.795 ;
        RECT 98.440 139.370 98.610 141.410 ;
        RECT 99.730 139.370 99.900 141.410 ;
        RECT 101.020 139.370 101.190 141.410 ;
        RECT 98.670 138.985 99.670 139.155 ;
        RECT 99.960 138.985 100.960 139.155 ;
        RECT 101.700 138.570 101.870 142.410 ;
        RECT 100.960 138.560 101.870 138.570 ;
        RECT 97.770 138.350 101.870 138.560 ;
        RECT 97.770 134.500 97.950 138.350 ;
        RECT 98.670 137.565 99.670 137.735 ;
        RECT 99.960 137.565 100.960 137.735 ;
        RECT 98.440 135.310 98.610 137.350 ;
        RECT 99.730 135.310 99.900 137.350 ;
        RECT 101.020 135.310 101.190 137.350 ;
        RECT 98.670 134.925 99.670 135.095 ;
        RECT 99.960 134.925 100.960 135.095 ;
        RECT 101.700 134.510 101.870 138.350 ;
        RECT 100.960 134.500 101.870 134.510 ;
        RECT 97.770 134.290 101.870 134.500 ;
        RECT 97.770 130.440 97.950 134.290 ;
        RECT 98.670 133.505 99.670 133.675 ;
        RECT 99.960 133.505 100.960 133.675 ;
        RECT 98.440 131.250 98.610 133.290 ;
        RECT 99.730 131.250 99.900 133.290 ;
        RECT 101.020 131.250 101.190 133.290 ;
        RECT 98.670 130.865 99.670 131.035 ;
        RECT 99.960 130.865 100.960 131.035 ;
        RECT 101.700 130.450 101.870 134.290 ;
        RECT 100.960 130.440 101.870 130.450 ;
        RECT 97.770 130.230 101.870 130.440 ;
        RECT 97.770 126.380 97.950 130.230 ;
        RECT 98.670 129.445 99.670 129.615 ;
        RECT 99.960 129.445 100.960 129.615 ;
        RECT 98.440 127.190 98.610 129.230 ;
        RECT 99.730 127.190 99.900 129.230 ;
        RECT 101.020 127.190 101.190 129.230 ;
        RECT 98.670 126.805 99.670 126.975 ;
        RECT 99.960 126.805 100.960 126.975 ;
        RECT 101.700 126.390 101.870 130.230 ;
        RECT 100.960 126.380 101.870 126.390 ;
        RECT 97.770 126.170 101.870 126.380 ;
        RECT 97.770 122.320 97.950 126.170 ;
        RECT 98.670 125.385 99.670 125.555 ;
        RECT 99.960 125.385 100.960 125.555 ;
        RECT 98.440 123.130 98.610 125.170 ;
        RECT 99.730 123.130 99.900 125.170 ;
        RECT 101.020 123.130 101.190 125.170 ;
        RECT 98.670 122.745 99.670 122.915 ;
        RECT 99.960 122.745 100.960 122.915 ;
        RECT 101.700 122.330 101.870 126.170 ;
        RECT 100.960 122.320 101.870 122.330 ;
        RECT 97.770 122.110 101.870 122.320 ;
        RECT 97.770 118.260 97.950 122.110 ;
        RECT 98.670 121.325 99.670 121.495 ;
        RECT 99.960 121.325 100.960 121.495 ;
        RECT 98.440 119.070 98.610 121.110 ;
        RECT 99.730 119.070 99.900 121.110 ;
        RECT 101.020 119.070 101.190 121.110 ;
        RECT 98.670 118.685 99.670 118.855 ;
        RECT 99.960 118.685 100.960 118.855 ;
        RECT 101.700 118.270 101.870 122.110 ;
        RECT 100.960 118.260 101.870 118.270 ;
        RECT 97.770 118.050 101.870 118.260 ;
        RECT 97.770 114.200 97.950 118.050 ;
        RECT 98.670 117.265 99.670 117.435 ;
        RECT 99.960 117.265 100.960 117.435 ;
        RECT 98.440 115.010 98.610 117.050 ;
        RECT 99.730 115.010 99.900 117.050 ;
        RECT 101.020 115.010 101.190 117.050 ;
        RECT 98.670 114.625 99.670 114.795 ;
        RECT 99.960 114.625 100.960 114.795 ;
        RECT 101.700 114.210 101.870 118.050 ;
        RECT 100.960 114.200 101.870 114.210 ;
        RECT 97.770 113.990 101.870 114.200 ;
        RECT 97.770 110.140 97.950 113.990 ;
        RECT 98.670 113.205 99.670 113.375 ;
        RECT 99.960 113.205 100.960 113.375 ;
        RECT 98.440 110.950 98.610 112.990 ;
        RECT 99.730 110.950 99.900 112.990 ;
        RECT 101.020 110.950 101.190 112.990 ;
        RECT 98.670 110.565 99.670 110.735 ;
        RECT 99.960 110.565 100.960 110.735 ;
        RECT 101.700 110.150 101.870 113.990 ;
        RECT 100.960 110.140 101.870 110.150 ;
        RECT 97.770 109.930 101.870 110.140 ;
        RECT 97.770 106.080 97.950 109.930 ;
        RECT 98.670 109.145 99.670 109.315 ;
        RECT 99.960 109.145 100.960 109.315 ;
        RECT 98.440 106.890 98.610 108.930 ;
        RECT 99.730 106.890 99.900 108.930 ;
        RECT 101.020 106.890 101.190 108.930 ;
        RECT 98.670 106.505 99.670 106.675 ;
        RECT 99.960 106.505 100.960 106.675 ;
        RECT 101.700 106.090 101.870 109.930 ;
        RECT 100.960 106.080 101.870 106.090 ;
        RECT 97.770 105.870 101.870 106.080 ;
        RECT 97.770 102.020 97.950 105.870 ;
        RECT 98.670 105.085 99.670 105.255 ;
        RECT 99.960 105.085 100.960 105.255 ;
        RECT 98.440 102.830 98.610 104.870 ;
        RECT 99.730 102.830 99.900 104.870 ;
        RECT 101.020 102.830 101.190 104.870 ;
        RECT 98.670 102.445 99.670 102.615 ;
        RECT 99.960 102.445 100.960 102.615 ;
        RECT 101.700 102.030 101.870 105.870 ;
        RECT 100.960 102.020 101.870 102.030 ;
        RECT 97.770 101.810 101.870 102.020 ;
        RECT 97.770 97.960 97.950 101.810 ;
        RECT 98.670 101.025 99.670 101.195 ;
        RECT 99.960 101.025 100.960 101.195 ;
        RECT 98.440 98.770 98.610 100.810 ;
        RECT 99.730 98.770 99.900 100.810 ;
        RECT 101.020 98.770 101.190 100.810 ;
        RECT 98.670 98.385 99.670 98.555 ;
        RECT 99.960 98.385 100.960 98.555 ;
        RECT 101.700 97.970 101.870 101.810 ;
        RECT 100.960 97.960 101.870 97.970 ;
        RECT 97.770 97.750 101.870 97.960 ;
        RECT 97.770 93.900 97.950 97.750 ;
        RECT 98.670 96.965 99.670 97.135 ;
        RECT 99.960 96.965 100.960 97.135 ;
        RECT 98.440 94.710 98.610 96.750 ;
        RECT 99.730 94.710 99.900 96.750 ;
        RECT 101.020 94.710 101.190 96.750 ;
        RECT 98.670 94.325 99.670 94.495 ;
        RECT 99.960 94.325 100.960 94.495 ;
        RECT 101.700 93.910 101.870 97.750 ;
        RECT 100.960 93.900 101.870 93.910 ;
        RECT 97.770 93.690 101.870 93.900 ;
        RECT 97.770 89.840 97.950 93.690 ;
        RECT 98.670 92.905 99.670 93.075 ;
        RECT 99.960 92.905 100.960 93.075 ;
        RECT 98.440 90.650 98.610 92.690 ;
        RECT 99.730 90.650 99.900 92.690 ;
        RECT 101.020 90.650 101.190 92.690 ;
        RECT 98.670 90.265 99.670 90.435 ;
        RECT 99.960 90.265 100.960 90.435 ;
        RECT 101.700 89.850 101.870 93.690 ;
        RECT 100.960 89.840 101.870 89.850 ;
        RECT 97.770 89.630 101.870 89.840 ;
        RECT 97.770 85.780 97.950 89.630 ;
        RECT 98.670 88.845 99.670 89.015 ;
        RECT 99.960 88.845 100.960 89.015 ;
        RECT 98.440 86.590 98.610 88.630 ;
        RECT 99.730 86.590 99.900 88.630 ;
        RECT 101.020 86.590 101.190 88.630 ;
        RECT 98.670 86.205 99.670 86.375 ;
        RECT 99.960 86.205 100.960 86.375 ;
        RECT 101.700 85.790 101.870 89.630 ;
        RECT 100.960 85.780 101.870 85.790 ;
        RECT 97.770 85.570 101.870 85.780 ;
        RECT 97.770 81.720 97.950 85.570 ;
        RECT 98.670 84.785 99.670 84.955 ;
        RECT 99.960 84.785 100.960 84.955 ;
        RECT 98.440 82.530 98.610 84.570 ;
        RECT 99.730 82.530 99.900 84.570 ;
        RECT 101.020 82.530 101.190 84.570 ;
        RECT 98.670 82.145 99.670 82.315 ;
        RECT 99.960 82.145 100.960 82.315 ;
        RECT 101.700 81.730 101.870 85.570 ;
        RECT 100.960 81.720 101.870 81.730 ;
        RECT 97.770 81.510 101.870 81.720 ;
        RECT 97.770 77.660 97.950 81.510 ;
        RECT 98.670 80.725 99.670 80.895 ;
        RECT 99.960 80.725 100.960 80.895 ;
        RECT 98.440 78.470 98.610 80.510 ;
        RECT 99.730 78.470 99.900 80.510 ;
        RECT 101.020 78.470 101.190 80.510 ;
        RECT 98.670 78.085 99.670 78.255 ;
        RECT 99.960 78.085 100.960 78.255 ;
        RECT 101.700 77.670 101.870 81.510 ;
        RECT 100.960 77.660 101.870 77.670 ;
        RECT 97.770 77.450 101.870 77.660 ;
        RECT 97.770 73.600 97.950 77.450 ;
        RECT 98.670 76.665 99.670 76.835 ;
        RECT 99.960 76.665 100.960 76.835 ;
        RECT 98.440 74.410 98.610 76.450 ;
        RECT 99.730 74.410 99.900 76.450 ;
        RECT 101.020 74.410 101.190 76.450 ;
        RECT 98.670 74.025 99.670 74.195 ;
        RECT 99.960 74.025 100.960 74.195 ;
        RECT 101.700 73.610 101.870 77.450 ;
        RECT 100.960 73.600 101.870 73.610 ;
        RECT 97.770 73.390 101.870 73.600 ;
        RECT 97.770 69.540 97.950 73.390 ;
        RECT 98.670 72.605 99.670 72.775 ;
        RECT 99.960 72.605 100.960 72.775 ;
        RECT 98.440 70.350 98.610 72.390 ;
        RECT 99.730 70.350 99.900 72.390 ;
        RECT 101.020 70.350 101.190 72.390 ;
        RECT 98.670 69.965 99.670 70.135 ;
        RECT 99.960 69.965 100.960 70.135 ;
        RECT 101.700 69.550 101.870 73.390 ;
        RECT 100.960 69.540 101.870 69.550 ;
        RECT 97.770 69.330 101.870 69.540 ;
        RECT 97.770 65.480 97.950 69.330 ;
        RECT 98.670 68.545 99.670 68.715 ;
        RECT 99.960 68.545 100.960 68.715 ;
        RECT 98.440 66.290 98.610 68.330 ;
        RECT 99.730 66.290 99.900 68.330 ;
        RECT 101.020 66.290 101.190 68.330 ;
        RECT 98.670 65.905 99.670 66.075 ;
        RECT 99.960 65.905 100.960 66.075 ;
        RECT 101.700 65.490 101.870 69.330 ;
        RECT 100.960 65.480 101.870 65.490 ;
        RECT 97.770 65.270 101.870 65.480 ;
        RECT 97.770 61.420 97.950 65.270 ;
        RECT 98.670 64.485 99.670 64.655 ;
        RECT 99.960 64.485 100.960 64.655 ;
        RECT 98.440 62.230 98.610 64.270 ;
        RECT 99.730 62.230 99.900 64.270 ;
        RECT 101.020 62.230 101.190 64.270 ;
        RECT 98.670 61.845 99.670 62.015 ;
        RECT 99.960 61.845 100.960 62.015 ;
        RECT 101.700 61.420 101.870 65.270 ;
        RECT 97.770 61.210 101.870 61.420 ;
        RECT 102.220 146.510 105.720 146.680 ;
        RECT 102.220 146.500 105.730 146.510 ;
        RECT 102.220 142.620 102.390 146.500 ;
        RECT 105.550 145.400 105.730 146.500 ;
        RECT 106.110 146.230 114.510 146.400 ;
        RECT 131.590 146.260 147.700 146.440 ;
        RECT 102.860 145.210 103.860 145.380 ;
        RECT 104.150 145.210 105.150 145.380 ;
        RECT 102.630 144.000 102.800 145.040 ;
        RECT 103.920 144.000 104.090 145.040 ;
        RECT 105.210 144.000 105.380 145.040 ;
        RECT 102.860 143.660 103.860 143.830 ;
        RECT 104.150 143.660 105.150 143.830 ;
        RECT 105.550 142.620 105.720 145.400 ;
        RECT 102.220 142.450 105.720 142.620 ;
        RECT 102.220 142.410 105.730 142.450 ;
        RECT 102.220 138.560 102.390 142.410 ;
        RECT 105.550 141.340 105.730 142.410 ;
        RECT 102.860 141.150 103.860 141.320 ;
        RECT 104.150 141.150 105.150 141.320 ;
        RECT 102.630 139.940 102.800 140.980 ;
        RECT 103.920 139.940 104.090 140.980 ;
        RECT 105.210 139.940 105.380 140.980 ;
        RECT 102.860 139.600 103.860 139.770 ;
        RECT 104.150 139.600 105.150 139.770 ;
        RECT 105.550 138.560 105.720 141.340 ;
        RECT 102.220 138.390 105.720 138.560 ;
        RECT 102.220 138.350 105.730 138.390 ;
        RECT 102.220 134.500 102.390 138.350 ;
        RECT 105.550 137.280 105.730 138.350 ;
        RECT 102.860 137.090 103.860 137.260 ;
        RECT 104.150 137.090 105.150 137.260 ;
        RECT 102.630 135.880 102.800 136.920 ;
        RECT 103.920 135.880 104.090 136.920 ;
        RECT 105.210 135.880 105.380 136.920 ;
        RECT 102.860 135.540 103.860 135.710 ;
        RECT 104.150 135.540 105.150 135.710 ;
        RECT 105.550 134.500 105.720 137.280 ;
        RECT 102.220 134.330 105.720 134.500 ;
        RECT 102.220 134.290 105.730 134.330 ;
        RECT 102.220 130.440 102.390 134.290 ;
        RECT 105.550 133.220 105.730 134.290 ;
        RECT 106.110 133.430 106.280 146.230 ;
        RECT 108.550 144.190 113.590 144.360 ;
        RECT 108.210 143.130 108.380 144.130 ;
        RECT 113.760 143.130 113.930 144.130 ;
        RECT 108.550 142.900 113.590 143.070 ;
        RECT 108.210 141.840 108.380 142.840 ;
        RECT 113.760 141.840 113.930 142.840 ;
        RECT 108.550 141.610 113.590 141.780 ;
        RECT 108.210 140.550 108.380 141.550 ;
        RECT 113.760 140.550 113.930 141.550 ;
        RECT 108.550 140.320 113.590 140.490 ;
        RECT 108.210 139.260 108.380 140.260 ;
        RECT 113.760 139.260 113.930 140.260 ;
        RECT 108.550 139.030 113.590 139.200 ;
        RECT 108.210 137.970 108.380 138.970 ;
        RECT 113.760 137.970 113.930 138.970 ;
        RECT 108.550 137.740 113.590 137.910 ;
        RECT 108.210 136.680 108.380 137.680 ;
        RECT 113.760 136.680 113.930 137.680 ;
        RECT 108.550 136.450 113.590 136.620 ;
        RECT 108.210 135.390 108.380 136.390 ;
        RECT 113.760 135.390 113.930 136.390 ;
        RECT 108.550 135.160 113.590 135.330 ;
        RECT 108.210 134.100 108.380 135.100 ;
        RECT 113.760 134.100 113.930 135.100 ;
        RECT 108.550 133.870 113.590 134.040 ;
        RECT 114.340 133.430 114.510 146.230 ;
        RECT 106.110 133.260 114.510 133.430 ;
        RECT 115.370 146.090 130.930 146.260 ;
        RECT 115.370 133.570 115.540 146.090 ;
        RECT 117.010 144.470 122.050 144.640 ;
        RECT 124.010 144.470 129.050 144.640 ;
        RECT 116.670 143.410 116.840 144.410 ;
        RECT 122.220 143.410 122.390 144.410 ;
        RECT 123.670 143.410 123.840 144.410 ;
        RECT 129.220 143.410 129.390 144.410 ;
        RECT 117.010 143.180 122.050 143.350 ;
        RECT 124.010 143.180 129.050 143.350 ;
        RECT 117.010 142.470 122.050 142.640 ;
        RECT 124.010 142.470 129.050 142.640 ;
        RECT 116.670 141.410 116.840 142.410 ;
        RECT 122.220 141.410 122.390 142.410 ;
        RECT 123.670 141.410 123.840 142.410 ;
        RECT 129.220 141.410 129.390 142.410 ;
        RECT 117.010 141.180 122.050 141.350 ;
        RECT 124.010 141.180 129.050 141.350 ;
        RECT 117.010 138.470 122.050 138.640 ;
        RECT 124.010 138.470 129.050 138.640 ;
        RECT 116.670 137.410 116.840 138.410 ;
        RECT 122.220 137.410 122.390 138.410 ;
        RECT 123.670 137.410 123.840 138.410 ;
        RECT 129.220 137.410 129.390 138.410 ;
        RECT 117.010 137.180 122.050 137.350 ;
        RECT 124.010 137.180 129.050 137.350 ;
        RECT 117.010 136.470 122.050 136.640 ;
        RECT 124.010 136.470 129.050 136.640 ;
        RECT 116.670 135.410 116.840 136.410 ;
        RECT 122.220 135.410 122.390 136.410 ;
        RECT 123.670 135.410 123.840 136.410 ;
        RECT 129.220 135.410 129.390 136.410 ;
        RECT 117.010 135.180 122.050 135.350 ;
        RECT 124.010 135.180 129.050 135.350 ;
        RECT 130.760 133.570 130.930 146.090 ;
        RECT 115.370 133.400 130.930 133.570 ;
        RECT 131.590 133.600 131.770 146.260 ;
        RECT 132.730 145.450 137.770 145.620 ;
        RECT 141.730 145.450 146.770 145.620 ;
        RECT 132.345 144.890 132.515 145.390 ;
        RECT 137.985 144.890 138.155 145.390 ;
        RECT 141.345 144.890 141.515 145.390 ;
        RECT 146.985 144.890 147.155 145.390 ;
        RECT 132.730 144.660 137.770 144.830 ;
        RECT 141.730 144.660 146.770 144.830 ;
        RECT 132.730 140.950 137.770 141.120 ;
        RECT 141.730 140.950 146.770 141.120 ;
        RECT 132.345 140.390 132.515 140.890 ;
        RECT 137.985 140.390 138.155 140.890 ;
        RECT 141.345 140.390 141.515 140.890 ;
        RECT 146.985 140.390 147.155 140.890 ;
        RECT 132.730 140.160 137.770 140.330 ;
        RECT 141.730 140.160 146.770 140.330 ;
        RECT 132.730 136.450 137.770 136.620 ;
        RECT 141.730 136.450 146.770 136.620 ;
        RECT 132.345 135.890 132.515 136.390 ;
        RECT 137.985 135.890 138.155 136.390 ;
        RECT 141.345 135.890 141.515 136.390 ;
        RECT 146.985 135.890 147.155 136.390 ;
        RECT 132.730 135.660 137.770 135.830 ;
        RECT 141.730 135.660 146.770 135.830 ;
        RECT 147.520 133.600 147.700 146.260 ;
        RECT 131.590 133.420 147.700 133.600 ;
        RECT 102.860 133.030 103.860 133.200 ;
        RECT 104.150 133.030 105.150 133.200 ;
        RECT 102.630 131.820 102.800 132.860 ;
        RECT 103.920 131.820 104.090 132.860 ;
        RECT 105.210 131.820 105.380 132.860 ;
        RECT 102.860 131.480 103.860 131.650 ;
        RECT 104.150 131.480 105.150 131.650 ;
        RECT 105.550 130.440 105.720 133.220 ;
        RECT 106.510 132.795 107.150 132.800 ;
        RECT 108.160 132.795 108.800 132.800 ;
        RECT 109.560 132.795 110.200 132.800 ;
        RECT 110.740 132.795 111.380 132.800 ;
        RECT 102.220 130.270 105.720 130.440 ;
        RECT 106.030 132.625 112.770 132.795 ;
        RECT 106.030 130.365 106.200 132.625 ;
        RECT 106.880 132.055 111.920 132.225 ;
        RECT 106.540 130.995 106.710 131.995 ;
        RECT 112.090 130.995 112.260 131.995 ;
        RECT 106.880 130.765 111.920 130.935 ;
        RECT 112.600 130.365 112.770 132.625 ;
        RECT 113.130 132.630 125.120 132.800 ;
        RECT 113.130 130.870 113.300 132.630 ;
        RECT 114.025 132.060 115.065 132.230 ;
        RECT 113.640 131.500 113.810 132.000 ;
        RECT 115.280 131.500 115.450 132.000 ;
        RECT 114.025 131.270 115.065 131.440 ;
        RECT 115.790 130.870 115.960 132.630 ;
        RECT 116.685 132.060 124.225 132.230 ;
        RECT 116.300 131.500 116.470 132.000 ;
        RECT 124.440 131.500 124.610 132.000 ;
        RECT 116.685 131.270 124.225 131.440 ;
        RECT 124.950 130.870 125.120 132.630 ;
        RECT 113.130 130.700 125.120 130.870 ;
        RECT 117.020 130.425 121.970 130.430 ;
        RECT 102.220 130.230 105.730 130.270 ;
        RECT 102.220 126.380 102.390 130.230 ;
        RECT 105.550 129.160 105.730 130.230 ;
        RECT 106.030 130.195 112.770 130.365 ;
        RECT 115.795 130.255 124.625 130.425 ;
        RECT 102.860 128.970 103.860 129.140 ;
        RECT 104.150 128.970 105.150 129.140 ;
        RECT 102.630 127.760 102.800 128.800 ;
        RECT 103.920 127.760 104.090 128.800 ;
        RECT 105.210 127.760 105.380 128.800 ;
        RECT 102.860 127.420 103.860 127.590 ;
        RECT 104.150 127.420 105.150 127.590 ;
        RECT 105.550 126.380 105.720 129.160 ;
        RECT 115.795 128.495 115.965 130.255 ;
        RECT 124.455 129.950 124.625 130.255 ;
        RECT 116.690 129.685 123.730 129.855 ;
        RECT 116.305 129.125 116.475 129.625 ;
        RECT 123.945 129.125 124.115 129.625 ;
        RECT 116.690 128.895 123.730 129.065 ;
        RECT 124.450 128.810 124.625 129.950 ;
        RECT 124.455 128.495 124.625 128.810 ;
        RECT 115.795 128.325 124.625 128.495 ;
        RECT 115.795 126.565 115.965 128.325 ;
        RECT 124.455 128.020 124.625 128.325 ;
        RECT 116.690 127.755 123.730 127.925 ;
        RECT 116.305 127.195 116.475 127.695 ;
        RECT 123.945 127.195 124.115 127.695 ;
        RECT 116.690 126.965 123.730 127.135 ;
        RECT 124.450 126.880 124.625 128.020 ;
        RECT 124.455 126.565 124.625 126.880 ;
        RECT 115.795 126.395 124.625 126.565 ;
        RECT 102.220 126.210 105.720 126.380 ;
        RECT 102.220 126.170 105.730 126.210 ;
        RECT 102.220 122.320 102.390 126.170 ;
        RECT 105.550 125.100 105.730 126.170 ;
        RECT 106.140 125.570 113.450 125.750 ;
        RECT 102.860 124.910 103.860 125.080 ;
        RECT 104.150 124.910 105.150 125.080 ;
        RECT 102.630 123.700 102.800 124.740 ;
        RECT 103.920 123.700 104.090 124.740 ;
        RECT 105.210 123.700 105.380 124.740 ;
        RECT 102.860 123.360 103.860 123.530 ;
        RECT 104.150 123.360 105.150 123.530 ;
        RECT 105.550 122.320 105.720 125.100 ;
        RECT 102.220 122.150 105.720 122.320 ;
        RECT 102.220 122.110 105.730 122.150 ;
        RECT 102.220 118.260 102.390 122.110 ;
        RECT 105.550 121.040 105.730 122.110 ;
        RECT 102.860 120.850 103.860 121.020 ;
        RECT 104.150 120.850 105.150 121.020 ;
        RECT 102.630 119.640 102.800 120.680 ;
        RECT 103.920 119.640 104.090 120.680 ;
        RECT 105.210 119.640 105.380 120.680 ;
        RECT 102.860 119.300 103.860 119.470 ;
        RECT 104.150 119.300 105.150 119.470 ;
        RECT 105.550 118.260 105.720 121.040 ;
        RECT 102.220 118.090 105.720 118.260 ;
        RECT 102.220 118.050 105.730 118.090 ;
        RECT 102.220 114.200 102.390 118.050 ;
        RECT 105.550 116.980 105.730 118.050 ;
        RECT 102.860 116.790 103.860 116.960 ;
        RECT 104.150 116.790 105.150 116.960 ;
        RECT 102.630 115.580 102.800 116.620 ;
        RECT 103.920 115.580 104.090 116.620 ;
        RECT 105.210 115.580 105.380 116.620 ;
        RECT 102.860 115.240 103.860 115.410 ;
        RECT 104.150 115.240 105.150 115.410 ;
        RECT 105.550 114.200 105.720 116.980 ;
        RECT 102.220 114.030 105.720 114.200 ;
        RECT 102.220 113.990 105.730 114.030 ;
        RECT 102.220 110.140 102.390 113.990 ;
        RECT 105.550 112.920 105.730 113.990 ;
        RECT 102.860 112.730 103.860 112.900 ;
        RECT 104.150 112.730 105.150 112.900 ;
        RECT 102.630 111.520 102.800 112.560 ;
        RECT 103.920 111.520 104.090 112.560 ;
        RECT 105.210 111.520 105.380 112.560 ;
        RECT 102.860 111.180 103.860 111.350 ;
        RECT 104.150 111.180 105.150 111.350 ;
        RECT 105.550 110.140 105.720 112.920 ;
        RECT 102.220 109.970 105.720 110.140 ;
        RECT 102.220 109.930 105.730 109.970 ;
        RECT 102.220 106.080 102.390 109.930 ;
        RECT 105.550 108.860 105.730 109.930 ;
        RECT 106.140 109.440 106.310 125.570 ;
        RECT 107.080 124.840 112.120 125.010 ;
        RECT 106.740 124.280 106.910 124.780 ;
        RECT 112.290 124.280 112.460 124.780 ;
        RECT 107.080 124.050 112.120 124.220 ;
        RECT 106.740 123.490 106.910 123.990 ;
        RECT 112.290 123.490 112.460 123.990 ;
        RECT 107.080 123.260 112.120 123.430 ;
        RECT 106.740 122.700 106.910 123.200 ;
        RECT 112.290 122.700 112.460 123.200 ;
        RECT 107.080 122.470 112.120 122.640 ;
        RECT 106.740 121.910 106.910 122.410 ;
        RECT 112.290 121.910 112.460 122.410 ;
        RECT 107.080 121.680 112.120 121.850 ;
        RECT 106.740 121.120 106.910 121.620 ;
        RECT 112.290 121.120 112.460 121.620 ;
        RECT 107.080 120.890 112.120 121.060 ;
        RECT 106.740 120.330 106.910 120.830 ;
        RECT 112.290 120.330 112.460 120.830 ;
        RECT 107.080 120.100 112.120 120.270 ;
        RECT 106.740 119.540 106.910 120.040 ;
        RECT 112.290 119.540 112.460 120.040 ;
        RECT 107.080 119.310 112.120 119.480 ;
        RECT 106.740 118.750 106.910 119.250 ;
        RECT 112.290 118.750 112.460 119.250 ;
        RECT 107.080 118.520 112.120 118.690 ;
        RECT 106.740 117.960 106.910 118.460 ;
        RECT 112.290 117.960 112.460 118.460 ;
        RECT 107.080 117.730 112.120 117.900 ;
        RECT 106.740 117.170 106.910 117.670 ;
        RECT 112.290 117.170 112.460 117.670 ;
        RECT 107.080 116.940 112.120 117.110 ;
        RECT 106.740 116.380 106.910 116.880 ;
        RECT 112.290 116.380 112.460 116.880 ;
        RECT 107.080 116.150 112.120 116.320 ;
        RECT 106.740 115.590 106.910 116.090 ;
        RECT 112.290 115.590 112.460 116.090 ;
        RECT 107.080 115.360 112.120 115.530 ;
        RECT 106.740 114.800 106.910 115.300 ;
        RECT 112.290 114.800 112.460 115.300 ;
        RECT 107.080 114.570 112.120 114.740 ;
        RECT 106.740 114.010 106.910 114.510 ;
        RECT 112.290 114.010 112.460 114.510 ;
        RECT 107.080 113.780 112.120 113.950 ;
        RECT 106.740 113.220 106.910 113.720 ;
        RECT 112.290 113.220 112.460 113.720 ;
        RECT 107.080 112.990 112.120 113.160 ;
        RECT 106.740 112.430 106.910 112.930 ;
        RECT 112.290 112.430 112.460 112.930 ;
        RECT 107.080 112.200 112.120 112.370 ;
        RECT 106.740 111.640 106.910 112.140 ;
        RECT 112.290 111.640 112.460 112.140 ;
        RECT 107.080 111.410 112.120 111.580 ;
        RECT 106.740 110.850 106.910 111.350 ;
        RECT 112.290 110.850 112.460 111.350 ;
        RECT 107.080 110.620 112.120 110.790 ;
        RECT 106.740 110.060 106.910 110.560 ;
        RECT 112.290 110.060 112.460 110.560 ;
        RECT 107.080 109.830 112.120 110.000 ;
        RECT 113.280 109.440 113.450 125.570 ;
        RECT 114.260 125.580 121.030 125.750 ;
        RECT 114.260 112.820 114.430 125.580 ;
        RECT 115.140 124.660 120.180 124.830 ;
        RECT 114.755 124.100 114.925 124.600 ;
        RECT 120.395 124.100 120.565 124.600 ;
        RECT 115.140 123.870 120.180 124.040 ;
        RECT 114.755 123.310 114.925 123.810 ;
        RECT 120.395 123.310 120.565 123.810 ;
        RECT 115.140 123.080 120.180 123.250 ;
        RECT 114.755 122.520 114.925 123.020 ;
        RECT 120.395 122.520 120.565 123.020 ;
        RECT 115.140 122.290 120.180 122.460 ;
        RECT 114.755 121.730 114.925 122.230 ;
        RECT 120.395 121.730 120.565 122.230 ;
        RECT 115.140 121.500 120.180 121.670 ;
        RECT 114.755 120.940 114.925 121.440 ;
        RECT 120.395 120.940 120.565 121.440 ;
        RECT 115.140 120.710 120.180 120.880 ;
        RECT 114.755 120.150 114.925 120.650 ;
        RECT 120.395 120.150 120.565 120.650 ;
        RECT 115.140 119.920 120.180 120.090 ;
        RECT 114.755 119.360 114.925 119.860 ;
        RECT 120.395 119.360 120.565 119.860 ;
        RECT 115.140 119.130 120.180 119.300 ;
        RECT 114.755 118.570 114.925 119.070 ;
        RECT 120.395 118.570 120.565 119.070 ;
        RECT 115.140 118.340 120.180 118.510 ;
        RECT 114.755 117.780 114.925 118.280 ;
        RECT 120.395 117.780 120.565 118.280 ;
        RECT 115.140 117.550 120.180 117.720 ;
        RECT 114.755 116.990 114.925 117.490 ;
        RECT 120.395 116.990 120.565 117.490 ;
        RECT 115.140 116.760 120.180 116.930 ;
        RECT 114.755 116.200 114.925 116.700 ;
        RECT 120.395 116.200 120.565 116.700 ;
        RECT 115.140 115.970 120.180 116.140 ;
        RECT 114.755 115.410 114.925 115.910 ;
        RECT 120.395 115.410 120.565 115.910 ;
        RECT 115.140 115.180 120.180 115.350 ;
        RECT 114.755 114.620 114.925 115.120 ;
        RECT 120.395 114.620 120.565 115.120 ;
        RECT 115.140 114.390 120.180 114.560 ;
        RECT 114.755 113.830 114.925 114.330 ;
        RECT 120.395 113.830 120.565 114.330 ;
        RECT 115.140 113.600 120.180 113.770 ;
        RECT 120.860 112.820 121.030 125.580 ;
        RECT 114.260 112.650 121.030 112.820 ;
        RECT 106.140 109.260 113.450 109.440 ;
        RECT 102.860 108.670 103.860 108.840 ;
        RECT 104.150 108.670 105.150 108.840 ;
        RECT 102.630 107.460 102.800 108.500 ;
        RECT 103.920 107.460 104.090 108.500 ;
        RECT 105.210 107.460 105.380 108.500 ;
        RECT 102.860 107.120 103.860 107.290 ;
        RECT 104.150 107.120 105.150 107.290 ;
        RECT 105.550 106.080 105.720 108.860 ;
        RECT 102.220 105.910 105.720 106.080 ;
        RECT 106.110 108.310 114.510 108.480 ;
        RECT 131.590 108.340 147.700 108.520 ;
        RECT 102.220 105.870 105.730 105.910 ;
        RECT 102.220 102.020 102.390 105.870 ;
        RECT 105.550 104.800 105.730 105.870 ;
        RECT 102.860 104.610 103.860 104.780 ;
        RECT 104.150 104.610 105.150 104.780 ;
        RECT 102.630 103.400 102.800 104.440 ;
        RECT 103.920 103.400 104.090 104.440 ;
        RECT 105.210 103.400 105.380 104.440 ;
        RECT 102.860 103.060 103.860 103.230 ;
        RECT 104.150 103.060 105.150 103.230 ;
        RECT 105.550 102.020 105.720 104.800 ;
        RECT 102.220 101.850 105.720 102.020 ;
        RECT 102.220 101.810 105.730 101.850 ;
        RECT 102.220 97.960 102.390 101.810 ;
        RECT 105.550 100.740 105.730 101.810 ;
        RECT 102.860 100.550 103.860 100.720 ;
        RECT 104.150 100.550 105.150 100.720 ;
        RECT 102.630 99.340 102.800 100.380 ;
        RECT 103.920 99.340 104.090 100.380 ;
        RECT 105.210 99.340 105.380 100.380 ;
        RECT 102.860 99.000 103.860 99.170 ;
        RECT 104.150 99.000 105.150 99.170 ;
        RECT 105.550 97.960 105.720 100.740 ;
        RECT 102.220 97.790 105.720 97.960 ;
        RECT 102.220 97.750 105.730 97.790 ;
        RECT 102.220 93.900 102.390 97.750 ;
        RECT 105.550 96.680 105.730 97.750 ;
        RECT 102.860 96.490 103.860 96.660 ;
        RECT 104.150 96.490 105.150 96.660 ;
        RECT 102.630 95.280 102.800 96.320 ;
        RECT 103.920 95.280 104.090 96.320 ;
        RECT 105.210 95.280 105.380 96.320 ;
        RECT 102.860 94.940 103.860 95.110 ;
        RECT 104.150 94.940 105.150 95.110 ;
        RECT 105.550 93.900 105.720 96.680 ;
        RECT 106.110 95.510 106.280 108.310 ;
        RECT 108.550 106.270 113.590 106.440 ;
        RECT 108.210 105.210 108.380 106.210 ;
        RECT 113.760 105.210 113.930 106.210 ;
        RECT 108.550 104.980 113.590 105.150 ;
        RECT 108.210 103.920 108.380 104.920 ;
        RECT 113.760 103.920 113.930 104.920 ;
        RECT 108.550 103.690 113.590 103.860 ;
        RECT 108.210 102.630 108.380 103.630 ;
        RECT 113.760 102.630 113.930 103.630 ;
        RECT 108.550 102.400 113.590 102.570 ;
        RECT 108.210 101.340 108.380 102.340 ;
        RECT 113.760 101.340 113.930 102.340 ;
        RECT 108.550 101.110 113.590 101.280 ;
        RECT 108.210 100.050 108.380 101.050 ;
        RECT 113.760 100.050 113.930 101.050 ;
        RECT 108.550 99.820 113.590 99.990 ;
        RECT 108.210 98.760 108.380 99.760 ;
        RECT 113.760 98.760 113.930 99.760 ;
        RECT 108.550 98.530 113.590 98.700 ;
        RECT 108.210 97.470 108.380 98.470 ;
        RECT 113.760 97.470 113.930 98.470 ;
        RECT 108.550 97.240 113.590 97.410 ;
        RECT 108.210 96.180 108.380 97.180 ;
        RECT 113.760 96.180 113.930 97.180 ;
        RECT 108.550 95.950 113.590 96.120 ;
        RECT 114.340 95.510 114.510 108.310 ;
        RECT 106.110 95.340 114.510 95.510 ;
        RECT 115.370 108.170 130.930 108.340 ;
        RECT 115.370 95.650 115.540 108.170 ;
        RECT 117.010 106.550 122.050 106.720 ;
        RECT 124.010 106.550 129.050 106.720 ;
        RECT 116.670 105.490 116.840 106.490 ;
        RECT 122.220 105.490 122.390 106.490 ;
        RECT 123.670 105.490 123.840 106.490 ;
        RECT 129.220 105.490 129.390 106.490 ;
        RECT 117.010 105.260 122.050 105.430 ;
        RECT 124.010 105.260 129.050 105.430 ;
        RECT 117.010 104.550 122.050 104.720 ;
        RECT 124.010 104.550 129.050 104.720 ;
        RECT 116.670 103.490 116.840 104.490 ;
        RECT 122.220 103.490 122.390 104.490 ;
        RECT 123.670 103.490 123.840 104.490 ;
        RECT 129.220 103.490 129.390 104.490 ;
        RECT 117.010 103.260 122.050 103.430 ;
        RECT 124.010 103.260 129.050 103.430 ;
        RECT 117.010 100.550 122.050 100.720 ;
        RECT 124.010 100.550 129.050 100.720 ;
        RECT 116.670 99.490 116.840 100.490 ;
        RECT 122.220 99.490 122.390 100.490 ;
        RECT 123.670 99.490 123.840 100.490 ;
        RECT 129.220 99.490 129.390 100.490 ;
        RECT 117.010 99.260 122.050 99.430 ;
        RECT 124.010 99.260 129.050 99.430 ;
        RECT 117.010 98.550 122.050 98.720 ;
        RECT 124.010 98.550 129.050 98.720 ;
        RECT 116.670 97.490 116.840 98.490 ;
        RECT 122.220 97.490 122.390 98.490 ;
        RECT 123.670 97.490 123.840 98.490 ;
        RECT 129.220 97.490 129.390 98.490 ;
        RECT 117.010 97.260 122.050 97.430 ;
        RECT 124.010 97.260 129.050 97.430 ;
        RECT 130.760 95.650 130.930 108.170 ;
        RECT 115.370 95.480 130.930 95.650 ;
        RECT 131.590 95.680 131.770 108.340 ;
        RECT 132.730 107.530 137.770 107.700 ;
        RECT 141.730 107.530 146.770 107.700 ;
        RECT 132.345 106.970 132.515 107.470 ;
        RECT 137.985 106.970 138.155 107.470 ;
        RECT 141.345 106.970 141.515 107.470 ;
        RECT 146.985 106.970 147.155 107.470 ;
        RECT 132.730 106.740 137.770 106.910 ;
        RECT 141.730 106.740 146.770 106.910 ;
        RECT 132.730 103.030 137.770 103.200 ;
        RECT 141.730 103.030 146.770 103.200 ;
        RECT 132.345 102.470 132.515 102.970 ;
        RECT 137.985 102.470 138.155 102.970 ;
        RECT 141.345 102.470 141.515 102.970 ;
        RECT 146.985 102.470 147.155 102.970 ;
        RECT 132.730 102.240 137.770 102.410 ;
        RECT 141.730 102.240 146.770 102.410 ;
        RECT 132.730 98.530 137.770 98.700 ;
        RECT 141.730 98.530 146.770 98.700 ;
        RECT 132.345 97.970 132.515 98.470 ;
        RECT 137.985 97.970 138.155 98.470 ;
        RECT 141.345 97.970 141.515 98.470 ;
        RECT 146.985 97.970 147.155 98.470 ;
        RECT 132.730 97.740 137.770 97.910 ;
        RECT 141.730 97.740 146.770 97.910 ;
        RECT 147.520 95.680 147.700 108.340 ;
        RECT 131.590 95.500 147.700 95.680 ;
        RECT 106.510 94.875 107.150 94.880 ;
        RECT 108.160 94.875 108.800 94.880 ;
        RECT 109.560 94.875 110.200 94.880 ;
        RECT 110.740 94.875 111.380 94.880 ;
        RECT 102.220 93.730 105.720 93.900 ;
        RECT 106.030 94.705 112.770 94.875 ;
        RECT 102.220 93.690 105.730 93.730 ;
        RECT 102.220 89.840 102.390 93.690 ;
        RECT 105.550 92.620 105.730 93.690 ;
        RECT 102.860 92.430 103.860 92.600 ;
        RECT 104.150 92.430 105.150 92.600 ;
        RECT 102.630 91.220 102.800 92.260 ;
        RECT 103.920 91.220 104.090 92.260 ;
        RECT 105.210 91.220 105.380 92.260 ;
        RECT 102.860 90.880 103.860 91.050 ;
        RECT 104.150 90.880 105.150 91.050 ;
        RECT 105.550 89.840 105.720 92.620 ;
        RECT 106.030 92.445 106.200 94.705 ;
        RECT 106.880 94.135 111.920 94.305 ;
        RECT 106.540 93.075 106.710 94.075 ;
        RECT 112.090 93.075 112.260 94.075 ;
        RECT 106.880 92.845 111.920 93.015 ;
        RECT 112.600 92.445 112.770 94.705 ;
        RECT 113.130 94.710 125.120 94.880 ;
        RECT 113.130 92.950 113.300 94.710 ;
        RECT 114.025 94.140 115.065 94.310 ;
        RECT 113.640 93.580 113.810 94.080 ;
        RECT 115.280 93.580 115.450 94.080 ;
        RECT 114.025 93.350 115.065 93.520 ;
        RECT 115.790 92.950 115.960 94.710 ;
        RECT 116.685 94.140 124.225 94.310 ;
        RECT 116.300 93.580 116.470 94.080 ;
        RECT 124.440 93.580 124.610 94.080 ;
        RECT 116.685 93.350 124.225 93.520 ;
        RECT 124.950 92.950 125.120 94.710 ;
        RECT 113.130 92.780 125.120 92.950 ;
        RECT 117.020 92.505 121.970 92.510 ;
        RECT 106.030 92.275 112.770 92.445 ;
        RECT 115.795 92.335 124.625 92.505 ;
        RECT 102.220 89.670 105.720 89.840 ;
        RECT 115.795 90.575 115.965 92.335 ;
        RECT 124.455 92.030 124.625 92.335 ;
        RECT 116.690 91.765 123.730 91.935 ;
        RECT 116.305 91.205 116.475 91.705 ;
        RECT 123.945 91.205 124.115 91.705 ;
        RECT 116.690 90.975 123.730 91.145 ;
        RECT 124.450 90.890 124.625 92.030 ;
        RECT 124.455 90.575 124.625 90.890 ;
        RECT 115.795 90.405 124.625 90.575 ;
        RECT 102.220 89.630 105.730 89.670 ;
        RECT 102.220 85.780 102.390 89.630 ;
        RECT 105.550 88.560 105.730 89.630 ;
        RECT 115.795 88.645 115.965 90.405 ;
        RECT 124.455 90.100 124.625 90.405 ;
        RECT 116.690 89.835 123.730 90.005 ;
        RECT 116.305 89.275 116.475 89.775 ;
        RECT 123.945 89.275 124.115 89.775 ;
        RECT 116.690 89.045 123.730 89.215 ;
        RECT 124.450 88.960 124.625 90.100 ;
        RECT 124.455 88.645 124.625 88.960 ;
        RECT 102.860 88.370 103.860 88.540 ;
        RECT 104.150 88.370 105.150 88.540 ;
        RECT 102.630 87.160 102.800 88.200 ;
        RECT 103.920 87.160 104.090 88.200 ;
        RECT 105.210 87.160 105.380 88.200 ;
        RECT 102.860 86.820 103.860 86.990 ;
        RECT 104.150 86.820 105.150 86.990 ;
        RECT 105.550 85.780 105.720 88.560 ;
        RECT 115.795 88.475 124.625 88.645 ;
        RECT 102.220 85.610 105.720 85.780 ;
        RECT 106.140 87.650 113.450 87.830 ;
        RECT 102.220 85.570 105.730 85.610 ;
        RECT 102.220 81.720 102.390 85.570 ;
        RECT 105.550 84.500 105.730 85.570 ;
        RECT 102.860 84.310 103.860 84.480 ;
        RECT 104.150 84.310 105.150 84.480 ;
        RECT 102.630 83.100 102.800 84.140 ;
        RECT 103.920 83.100 104.090 84.140 ;
        RECT 105.210 83.100 105.380 84.140 ;
        RECT 102.860 82.760 103.860 82.930 ;
        RECT 104.150 82.760 105.150 82.930 ;
        RECT 105.550 81.720 105.720 84.500 ;
        RECT 102.220 81.550 105.720 81.720 ;
        RECT 102.220 81.510 105.730 81.550 ;
        RECT 102.220 77.660 102.390 81.510 ;
        RECT 105.550 80.440 105.730 81.510 ;
        RECT 102.860 80.250 103.860 80.420 ;
        RECT 104.150 80.250 105.150 80.420 ;
        RECT 102.630 79.040 102.800 80.080 ;
        RECT 103.920 79.040 104.090 80.080 ;
        RECT 105.210 79.040 105.380 80.080 ;
        RECT 102.860 78.700 103.860 78.870 ;
        RECT 104.150 78.700 105.150 78.870 ;
        RECT 105.550 77.660 105.720 80.440 ;
        RECT 102.220 77.490 105.720 77.660 ;
        RECT 102.220 77.450 105.730 77.490 ;
        RECT 102.220 73.600 102.390 77.450 ;
        RECT 105.550 76.380 105.730 77.450 ;
        RECT 102.860 76.190 103.860 76.360 ;
        RECT 104.150 76.190 105.150 76.360 ;
        RECT 102.630 74.980 102.800 76.020 ;
        RECT 103.920 74.980 104.090 76.020 ;
        RECT 105.210 74.980 105.380 76.020 ;
        RECT 102.860 74.640 103.860 74.810 ;
        RECT 104.150 74.640 105.150 74.810 ;
        RECT 105.550 73.600 105.720 76.380 ;
        RECT 102.220 73.430 105.720 73.600 ;
        RECT 102.220 73.390 105.730 73.430 ;
        RECT 102.220 69.540 102.390 73.390 ;
        RECT 105.550 72.320 105.730 73.390 ;
        RECT 102.860 72.130 103.860 72.300 ;
        RECT 104.150 72.130 105.150 72.300 ;
        RECT 102.630 70.920 102.800 71.960 ;
        RECT 103.920 70.920 104.090 71.960 ;
        RECT 105.210 70.920 105.380 71.960 ;
        RECT 102.860 70.580 103.860 70.750 ;
        RECT 104.150 70.580 105.150 70.750 ;
        RECT 105.550 69.540 105.720 72.320 ;
        RECT 106.140 71.520 106.310 87.650 ;
        RECT 107.080 86.920 112.120 87.090 ;
        RECT 106.740 86.360 106.910 86.860 ;
        RECT 112.290 86.360 112.460 86.860 ;
        RECT 107.080 86.130 112.120 86.300 ;
        RECT 106.740 85.570 106.910 86.070 ;
        RECT 112.290 85.570 112.460 86.070 ;
        RECT 107.080 85.340 112.120 85.510 ;
        RECT 106.740 84.780 106.910 85.280 ;
        RECT 112.290 84.780 112.460 85.280 ;
        RECT 107.080 84.550 112.120 84.720 ;
        RECT 106.740 83.990 106.910 84.490 ;
        RECT 112.290 83.990 112.460 84.490 ;
        RECT 107.080 83.760 112.120 83.930 ;
        RECT 106.740 83.200 106.910 83.700 ;
        RECT 112.290 83.200 112.460 83.700 ;
        RECT 107.080 82.970 112.120 83.140 ;
        RECT 106.740 82.410 106.910 82.910 ;
        RECT 112.290 82.410 112.460 82.910 ;
        RECT 107.080 82.180 112.120 82.350 ;
        RECT 106.740 81.620 106.910 82.120 ;
        RECT 112.290 81.620 112.460 82.120 ;
        RECT 107.080 81.390 112.120 81.560 ;
        RECT 106.740 80.830 106.910 81.330 ;
        RECT 112.290 80.830 112.460 81.330 ;
        RECT 107.080 80.600 112.120 80.770 ;
        RECT 106.740 80.040 106.910 80.540 ;
        RECT 112.290 80.040 112.460 80.540 ;
        RECT 107.080 79.810 112.120 79.980 ;
        RECT 106.740 79.250 106.910 79.750 ;
        RECT 112.290 79.250 112.460 79.750 ;
        RECT 107.080 79.020 112.120 79.190 ;
        RECT 106.740 78.460 106.910 78.960 ;
        RECT 112.290 78.460 112.460 78.960 ;
        RECT 107.080 78.230 112.120 78.400 ;
        RECT 106.740 77.670 106.910 78.170 ;
        RECT 112.290 77.670 112.460 78.170 ;
        RECT 107.080 77.440 112.120 77.610 ;
        RECT 106.740 76.880 106.910 77.380 ;
        RECT 112.290 76.880 112.460 77.380 ;
        RECT 107.080 76.650 112.120 76.820 ;
        RECT 106.740 76.090 106.910 76.590 ;
        RECT 112.290 76.090 112.460 76.590 ;
        RECT 107.080 75.860 112.120 76.030 ;
        RECT 106.740 75.300 106.910 75.800 ;
        RECT 112.290 75.300 112.460 75.800 ;
        RECT 107.080 75.070 112.120 75.240 ;
        RECT 106.740 74.510 106.910 75.010 ;
        RECT 112.290 74.510 112.460 75.010 ;
        RECT 107.080 74.280 112.120 74.450 ;
        RECT 106.740 73.720 106.910 74.220 ;
        RECT 112.290 73.720 112.460 74.220 ;
        RECT 107.080 73.490 112.120 73.660 ;
        RECT 106.740 72.930 106.910 73.430 ;
        RECT 112.290 72.930 112.460 73.430 ;
        RECT 107.080 72.700 112.120 72.870 ;
        RECT 106.740 72.140 106.910 72.640 ;
        RECT 112.290 72.140 112.460 72.640 ;
        RECT 107.080 71.910 112.120 72.080 ;
        RECT 113.280 71.520 113.450 87.650 ;
        RECT 114.260 87.660 121.030 87.830 ;
        RECT 114.260 74.900 114.430 87.660 ;
        RECT 115.140 86.740 120.180 86.910 ;
        RECT 114.755 86.180 114.925 86.680 ;
        RECT 120.395 86.180 120.565 86.680 ;
        RECT 115.140 85.950 120.180 86.120 ;
        RECT 114.755 85.390 114.925 85.890 ;
        RECT 120.395 85.390 120.565 85.890 ;
        RECT 115.140 85.160 120.180 85.330 ;
        RECT 114.755 84.600 114.925 85.100 ;
        RECT 120.395 84.600 120.565 85.100 ;
        RECT 115.140 84.370 120.180 84.540 ;
        RECT 114.755 83.810 114.925 84.310 ;
        RECT 120.395 83.810 120.565 84.310 ;
        RECT 115.140 83.580 120.180 83.750 ;
        RECT 114.755 83.020 114.925 83.520 ;
        RECT 120.395 83.020 120.565 83.520 ;
        RECT 115.140 82.790 120.180 82.960 ;
        RECT 114.755 82.230 114.925 82.730 ;
        RECT 120.395 82.230 120.565 82.730 ;
        RECT 115.140 82.000 120.180 82.170 ;
        RECT 114.755 81.440 114.925 81.940 ;
        RECT 120.395 81.440 120.565 81.940 ;
        RECT 115.140 81.210 120.180 81.380 ;
        RECT 114.755 80.650 114.925 81.150 ;
        RECT 120.395 80.650 120.565 81.150 ;
        RECT 115.140 80.420 120.180 80.590 ;
        RECT 114.755 79.860 114.925 80.360 ;
        RECT 120.395 79.860 120.565 80.360 ;
        RECT 115.140 79.630 120.180 79.800 ;
        RECT 114.755 79.070 114.925 79.570 ;
        RECT 120.395 79.070 120.565 79.570 ;
        RECT 115.140 78.840 120.180 79.010 ;
        RECT 114.755 78.280 114.925 78.780 ;
        RECT 120.395 78.280 120.565 78.780 ;
        RECT 115.140 78.050 120.180 78.220 ;
        RECT 114.755 77.490 114.925 77.990 ;
        RECT 120.395 77.490 120.565 77.990 ;
        RECT 115.140 77.260 120.180 77.430 ;
        RECT 114.755 76.700 114.925 77.200 ;
        RECT 120.395 76.700 120.565 77.200 ;
        RECT 115.140 76.470 120.180 76.640 ;
        RECT 114.755 75.910 114.925 76.410 ;
        RECT 120.395 75.910 120.565 76.410 ;
        RECT 115.140 75.680 120.180 75.850 ;
        RECT 120.860 74.900 121.030 87.660 ;
        RECT 114.260 74.730 121.030 74.900 ;
        RECT 106.140 71.340 113.450 71.520 ;
        RECT 102.220 69.370 105.720 69.540 ;
        RECT 102.220 69.330 105.730 69.370 ;
        RECT 102.220 65.480 102.390 69.330 ;
        RECT 105.550 68.260 105.730 69.330 ;
        RECT 102.860 68.070 103.860 68.240 ;
        RECT 104.150 68.070 105.150 68.240 ;
        RECT 102.630 66.860 102.800 67.900 ;
        RECT 103.920 66.860 104.090 67.900 ;
        RECT 105.210 66.860 105.380 67.900 ;
        RECT 102.860 66.520 103.860 66.690 ;
        RECT 104.150 66.520 105.150 66.690 ;
        RECT 105.550 65.480 105.720 68.260 ;
        RECT 102.220 65.310 105.720 65.480 ;
        RECT 102.220 65.270 105.730 65.310 ;
        RECT 102.220 61.420 102.390 65.270 ;
        RECT 105.550 64.200 105.730 65.270 ;
        RECT 102.860 64.010 103.860 64.180 ;
        RECT 104.150 64.010 105.150 64.180 ;
        RECT 102.630 62.800 102.800 63.840 ;
        RECT 103.920 62.800 104.090 63.840 ;
        RECT 105.210 62.800 105.380 63.840 ;
        RECT 102.860 62.460 103.860 62.630 ;
        RECT 104.150 62.460 105.150 62.630 ;
        RECT 105.550 61.420 105.720 64.200 ;
        RECT 102.220 61.210 105.720 61.420 ;
        RECT 100.960 60.940 101.760 60.950 ;
        RECT 93.330 57.360 97.430 57.580 ;
        RECT 93.330 53.540 93.500 57.360 ;
        RECT 94.240 56.585 95.240 56.755 ;
        RECT 95.530 56.585 96.530 56.755 ;
        RECT 94.010 54.330 94.180 56.370 ;
        RECT 95.300 54.330 95.470 56.370 ;
        RECT 96.590 54.330 96.760 56.370 ;
        RECT 94.240 53.945 95.240 54.115 ;
        RECT 95.530 53.945 96.530 54.115 ;
        RECT 93.330 53.530 94.240 53.540 ;
        RECT 97.250 53.530 97.430 57.360 ;
        RECT 97.770 60.770 101.870 60.940 ;
        RECT 97.770 56.880 97.950 60.770 ;
        RECT 98.670 59.945 99.670 60.115 ;
        RECT 99.960 59.945 100.960 60.115 ;
        RECT 98.440 57.690 98.610 59.730 ;
        RECT 99.730 57.690 99.900 59.730 ;
        RECT 101.020 57.690 101.190 59.730 ;
        RECT 98.670 57.305 99.670 57.475 ;
        RECT 99.960 57.305 100.960 57.475 ;
        RECT 101.700 56.880 101.870 60.770 ;
        RECT 97.770 56.670 101.870 56.880 ;
        RECT 102.220 60.770 105.720 60.940 ;
        RECT 102.220 60.760 105.730 60.770 ;
        RECT 102.220 56.880 102.390 60.760 ;
        RECT 105.550 59.660 105.730 60.760 ;
        RECT 102.860 59.470 103.860 59.640 ;
        RECT 104.150 59.470 105.150 59.640 ;
        RECT 102.630 58.260 102.800 59.300 ;
        RECT 103.920 58.260 104.090 59.300 ;
        RECT 105.210 58.260 105.380 59.300 ;
        RECT 102.860 57.920 103.860 58.090 ;
        RECT 104.150 57.920 105.150 58.090 ;
        RECT 105.550 56.880 105.720 59.660 ;
        RECT 102.220 56.670 105.720 56.880 ;
        RECT 93.330 53.310 97.430 53.530 ;
        RECT 93.330 49.490 93.500 53.310 ;
        RECT 94.240 52.535 95.240 52.705 ;
        RECT 95.530 52.535 96.530 52.705 ;
        RECT 94.010 50.280 94.180 52.320 ;
        RECT 95.300 50.280 95.470 52.320 ;
        RECT 96.590 50.280 96.760 52.320 ;
        RECT 94.240 49.895 95.240 50.065 ;
        RECT 95.530 49.895 96.530 50.065 ;
        RECT 93.330 49.480 94.240 49.490 ;
        RECT 97.250 49.480 97.430 53.310 ;
        RECT 93.330 49.260 97.430 49.480 ;
        RECT 93.330 45.440 93.500 49.260 ;
        RECT 94.240 48.485 95.240 48.655 ;
        RECT 95.530 48.485 96.530 48.655 ;
        RECT 94.010 46.230 94.180 48.270 ;
        RECT 95.300 46.230 95.470 48.270 ;
        RECT 96.590 46.230 96.760 48.270 ;
        RECT 94.240 45.845 95.240 46.015 ;
        RECT 95.530 45.845 96.530 46.015 ;
        RECT 93.330 45.430 94.240 45.440 ;
        RECT 97.250 45.430 97.430 49.260 ;
        RECT 93.330 45.210 97.430 45.430 ;
        RECT 93.330 41.390 93.500 45.210 ;
        RECT 94.240 44.435 95.240 44.605 ;
        RECT 95.530 44.435 96.530 44.605 ;
        RECT 94.010 42.180 94.180 44.220 ;
        RECT 95.300 42.180 95.470 44.220 ;
        RECT 96.590 42.180 96.760 44.220 ;
        RECT 94.240 41.795 95.240 41.965 ;
        RECT 95.530 41.795 96.530 41.965 ;
        RECT 93.330 41.380 94.240 41.390 ;
        RECT 97.250 41.380 97.430 45.210 ;
        RECT 93.330 41.160 97.430 41.380 ;
        RECT 93.330 37.340 93.500 41.160 ;
        RECT 94.240 40.385 95.240 40.555 ;
        RECT 95.530 40.385 96.530 40.555 ;
        RECT 94.010 38.130 94.180 40.170 ;
        RECT 95.300 38.130 95.470 40.170 ;
        RECT 96.590 38.130 96.760 40.170 ;
        RECT 94.240 37.745 95.240 37.915 ;
        RECT 95.530 37.745 96.530 37.915 ;
        RECT 93.330 37.330 94.240 37.340 ;
        RECT 97.250 37.330 97.430 41.160 ;
        RECT 93.330 37.110 97.430 37.330 ;
        RECT 93.330 33.290 93.500 37.110 ;
        RECT 94.240 36.335 95.240 36.505 ;
        RECT 95.530 36.335 96.530 36.505 ;
        RECT 94.010 34.080 94.180 36.120 ;
        RECT 95.300 34.080 95.470 36.120 ;
        RECT 96.590 34.080 96.760 36.120 ;
        RECT 94.240 33.695 95.240 33.865 ;
        RECT 95.530 33.695 96.530 33.865 ;
        RECT 93.330 33.280 94.240 33.290 ;
        RECT 97.250 33.280 97.430 37.110 ;
        RECT 93.330 33.060 97.430 33.280 ;
        RECT 93.330 29.220 93.500 33.060 ;
        RECT 94.240 32.285 95.240 32.455 ;
        RECT 95.530 32.285 96.530 32.455 ;
        RECT 94.010 30.030 94.180 32.070 ;
        RECT 95.300 30.030 95.470 32.070 ;
        RECT 96.590 30.030 96.760 32.070 ;
        RECT 94.240 29.645 95.240 29.815 ;
        RECT 95.530 29.645 96.530 29.815 ;
        RECT 97.250 29.220 97.430 33.060 ;
        RECT 93.330 29.010 97.430 29.220 ;
        RECT 93.330 25.135 93.500 29.010 ;
        RECT 94.240 28.200 95.240 28.370 ;
        RECT 95.530 28.200 96.530 28.370 ;
        RECT 94.010 25.945 94.180 27.985 ;
        RECT 95.300 25.945 95.470 27.985 ;
        RECT 96.590 25.945 96.760 27.985 ;
        RECT 94.240 25.560 95.240 25.730 ;
        RECT 95.530 25.560 96.530 25.730 ;
        RECT 97.250 25.135 97.430 29.010 ;
        RECT 93.330 24.900 97.430 25.135 ;
        RECT 93.330 21.010 93.500 24.900 ;
        RECT 94.240 24.075 95.240 24.245 ;
        RECT 95.530 24.075 96.530 24.245 ;
        RECT 94.010 21.820 94.180 23.860 ;
        RECT 95.300 21.820 95.470 23.860 ;
        RECT 96.590 21.820 96.760 23.860 ;
        RECT 94.240 21.435 95.240 21.605 ;
        RECT 95.530 21.435 96.530 21.605 ;
        RECT 97.250 21.010 97.430 24.900 ;
        RECT 93.330 20.800 97.430 21.010 ;
        RECT 93.440 20.515 94.240 20.525 ;
        RECT 89.480 20.345 92.980 20.515 ;
        RECT 89.470 20.335 92.980 20.345 ;
        RECT 89.470 19.235 89.650 20.335 ;
        RECT 89.480 16.455 89.650 19.235 ;
        RECT 90.050 19.045 91.050 19.215 ;
        RECT 91.340 19.045 92.340 19.215 ;
        RECT 89.820 17.835 89.990 18.875 ;
        RECT 91.110 17.835 91.280 18.875 ;
        RECT 92.400 17.835 92.570 18.875 ;
        RECT 90.050 17.495 91.050 17.665 ;
        RECT 91.340 17.495 92.340 17.665 ;
        RECT 92.810 16.455 92.980 20.335 ;
        RECT 89.480 16.245 92.980 16.455 ;
        RECT 93.330 20.345 97.430 20.515 ;
        RECT 93.330 16.455 93.500 20.345 ;
        RECT 94.240 19.520 95.240 19.690 ;
        RECT 95.530 19.520 96.530 19.690 ;
        RECT 94.010 17.265 94.180 19.305 ;
        RECT 95.300 17.265 95.470 19.305 ;
        RECT 96.590 17.265 96.760 19.305 ;
        RECT 94.240 16.880 95.240 17.050 ;
        RECT 95.530 16.880 96.530 17.050 ;
        RECT 97.250 16.455 97.430 20.345 ;
        RECT 93.330 16.245 97.430 16.455 ;
      LAYER mcon ;
        RECT 90.020 155.450 129.900 155.620 ;
        RECT 89.540 153.500 89.710 155.140 ;
        RECT 90.470 154.880 130.350 155.050 ;
        RECT 90.050 153.900 90.220 154.740 ;
        RECT 130.600 153.900 130.770 154.740 ;
        RECT 90.470 153.590 130.350 153.760 ;
        RECT 89.540 151.580 89.710 152.270 ;
        RECT 90.260 151.760 92.245 151.930 ;
        RECT 104.415 151.760 106.400 151.930 ;
        RECT 90.130 145.210 90.970 145.380 ;
        RECT 91.420 145.210 92.260 145.380 ;
        RECT 89.820 144.080 89.990 144.960 ;
        RECT 91.110 144.080 91.280 144.960 ;
        RECT 92.400 144.080 92.570 144.960 ;
        RECT 90.130 143.660 90.970 143.830 ;
        RECT 91.420 143.660 92.260 143.830 ;
        RECT 89.480 142.750 89.650 143.190 ;
        RECT 90.130 141.210 90.970 141.380 ;
        RECT 91.420 141.210 92.260 141.380 ;
        RECT 89.820 140.080 89.990 140.960 ;
        RECT 91.110 140.080 91.280 140.960 ;
        RECT 92.400 140.080 92.570 140.960 ;
        RECT 90.130 139.660 90.970 139.830 ;
        RECT 91.420 139.660 92.260 139.830 ;
        RECT 89.480 138.750 89.650 139.190 ;
        RECT 90.130 137.110 90.970 137.280 ;
        RECT 91.420 137.110 92.260 137.280 ;
        RECT 89.820 135.980 89.990 136.860 ;
        RECT 91.110 135.980 91.280 136.860 ;
        RECT 92.400 135.980 92.570 136.860 ;
        RECT 90.130 135.560 90.970 135.730 ;
        RECT 91.420 135.560 92.260 135.730 ;
        RECT 89.480 134.650 89.650 135.090 ;
        RECT 90.130 133.060 90.970 133.230 ;
        RECT 91.420 133.060 92.260 133.230 ;
        RECT 89.820 131.930 89.990 132.810 ;
        RECT 91.110 131.930 91.280 132.810 ;
        RECT 92.400 131.930 92.570 132.810 ;
        RECT 90.130 131.510 90.970 131.680 ;
        RECT 91.420 131.510 92.260 131.680 ;
        RECT 89.480 130.600 89.650 131.040 ;
        RECT 90.130 129.010 90.970 129.180 ;
        RECT 91.420 129.010 92.260 129.180 ;
        RECT 89.820 127.880 89.990 128.760 ;
        RECT 91.110 127.880 91.280 128.760 ;
        RECT 92.400 127.880 92.570 128.760 ;
        RECT 90.130 127.460 90.970 127.630 ;
        RECT 91.420 127.460 92.260 127.630 ;
        RECT 89.480 126.550 89.650 126.990 ;
        RECT 90.130 124.960 90.970 125.130 ;
        RECT 91.420 124.960 92.260 125.130 ;
        RECT 89.820 123.830 89.990 124.710 ;
        RECT 91.110 123.830 91.280 124.710 ;
        RECT 92.400 123.830 92.570 124.710 ;
        RECT 90.130 123.410 90.970 123.580 ;
        RECT 91.420 123.410 92.260 123.580 ;
        RECT 89.480 122.500 89.650 122.940 ;
        RECT 90.130 120.910 90.970 121.080 ;
        RECT 91.420 120.910 92.260 121.080 ;
        RECT 89.820 119.780 89.990 120.660 ;
        RECT 91.110 119.780 91.280 120.660 ;
        RECT 92.400 119.780 92.570 120.660 ;
        RECT 90.130 119.360 90.970 119.530 ;
        RECT 91.420 119.360 92.260 119.530 ;
        RECT 89.480 118.450 89.650 118.890 ;
        RECT 90.130 116.860 90.970 117.030 ;
        RECT 91.420 116.860 92.260 117.030 ;
        RECT 89.820 115.730 89.990 116.610 ;
        RECT 91.110 115.730 91.280 116.610 ;
        RECT 92.400 115.730 92.570 116.610 ;
        RECT 90.130 115.310 90.970 115.480 ;
        RECT 91.420 115.310 92.260 115.480 ;
        RECT 89.480 114.400 89.650 114.840 ;
        RECT 90.130 112.810 90.970 112.980 ;
        RECT 91.420 112.810 92.260 112.980 ;
        RECT 89.820 111.680 89.990 112.560 ;
        RECT 91.110 111.680 91.280 112.560 ;
        RECT 92.400 111.680 92.570 112.560 ;
        RECT 90.130 111.260 90.970 111.430 ;
        RECT 91.420 111.260 92.260 111.430 ;
        RECT 89.480 110.350 89.650 110.790 ;
        RECT 90.130 108.760 90.970 108.930 ;
        RECT 91.420 108.760 92.260 108.930 ;
        RECT 89.820 107.630 89.990 108.510 ;
        RECT 91.110 107.630 91.280 108.510 ;
        RECT 92.400 107.630 92.570 108.510 ;
        RECT 90.130 107.210 90.970 107.380 ;
        RECT 91.420 107.210 92.260 107.380 ;
        RECT 89.480 106.300 89.650 106.740 ;
        RECT 90.130 104.710 90.970 104.880 ;
        RECT 91.420 104.710 92.260 104.880 ;
        RECT 89.820 103.580 89.990 104.460 ;
        RECT 91.110 103.580 91.280 104.460 ;
        RECT 92.400 103.580 92.570 104.460 ;
        RECT 90.130 103.160 90.970 103.330 ;
        RECT 91.420 103.160 92.260 103.330 ;
        RECT 89.480 102.250 89.650 102.690 ;
        RECT 90.130 100.660 90.970 100.830 ;
        RECT 91.420 100.660 92.260 100.830 ;
        RECT 89.820 99.530 89.990 100.410 ;
        RECT 91.110 99.530 91.280 100.410 ;
        RECT 92.400 99.530 92.570 100.410 ;
        RECT 90.130 99.110 90.970 99.280 ;
        RECT 91.420 99.110 92.260 99.280 ;
        RECT 89.480 98.200 89.650 98.640 ;
        RECT 90.130 96.610 90.970 96.780 ;
        RECT 91.420 96.610 92.260 96.780 ;
        RECT 89.820 95.480 89.990 96.360 ;
        RECT 91.110 95.480 91.280 96.360 ;
        RECT 92.400 95.480 92.570 96.360 ;
        RECT 90.130 95.060 90.970 95.230 ;
        RECT 91.420 95.060 92.260 95.230 ;
        RECT 89.480 94.150 89.650 94.590 ;
        RECT 90.130 92.560 90.970 92.730 ;
        RECT 91.420 92.560 92.260 92.730 ;
        RECT 89.820 91.430 89.990 92.310 ;
        RECT 91.110 91.430 91.280 92.310 ;
        RECT 92.400 91.430 92.570 92.310 ;
        RECT 90.130 91.010 90.970 91.180 ;
        RECT 91.420 91.010 92.260 91.180 ;
        RECT 89.480 90.100 89.650 90.540 ;
        RECT 90.130 88.510 90.970 88.680 ;
        RECT 91.420 88.510 92.260 88.680 ;
        RECT 89.820 87.380 89.990 88.260 ;
        RECT 91.110 87.380 91.280 88.260 ;
        RECT 92.400 87.380 92.570 88.260 ;
        RECT 90.130 86.960 90.970 87.130 ;
        RECT 91.420 86.960 92.260 87.130 ;
        RECT 89.480 86.050 89.650 86.490 ;
        RECT 90.130 84.460 90.970 84.630 ;
        RECT 91.420 84.460 92.260 84.630 ;
        RECT 89.820 83.330 89.990 84.210 ;
        RECT 91.110 83.330 91.280 84.210 ;
        RECT 92.400 83.330 92.570 84.210 ;
        RECT 90.130 82.910 90.970 83.080 ;
        RECT 91.420 82.910 92.260 83.080 ;
        RECT 89.480 82.000 89.650 82.440 ;
        RECT 90.130 80.410 90.970 80.580 ;
        RECT 91.420 80.410 92.260 80.580 ;
        RECT 89.820 79.280 89.990 80.160 ;
        RECT 91.110 79.280 91.280 80.160 ;
        RECT 92.400 79.280 92.570 80.160 ;
        RECT 90.130 78.860 90.970 79.030 ;
        RECT 91.420 78.860 92.260 79.030 ;
        RECT 89.480 77.950 89.650 78.390 ;
        RECT 90.130 76.360 90.970 76.530 ;
        RECT 91.420 76.360 92.260 76.530 ;
        RECT 89.820 75.230 89.990 76.110 ;
        RECT 91.110 75.230 91.280 76.110 ;
        RECT 92.400 75.230 92.570 76.110 ;
        RECT 90.130 74.810 90.970 74.980 ;
        RECT 91.420 74.810 92.260 74.980 ;
        RECT 89.480 73.900 89.650 74.340 ;
        RECT 90.130 72.310 90.970 72.480 ;
        RECT 91.420 72.310 92.260 72.480 ;
        RECT 89.820 71.180 89.990 72.060 ;
        RECT 91.110 71.180 91.280 72.060 ;
        RECT 92.400 71.180 92.570 72.060 ;
        RECT 90.130 70.760 90.970 70.930 ;
        RECT 91.420 70.760 92.260 70.930 ;
        RECT 89.480 69.850 89.650 70.290 ;
        RECT 90.130 68.260 90.970 68.430 ;
        RECT 91.420 68.260 92.260 68.430 ;
        RECT 89.820 67.130 89.990 68.010 ;
        RECT 91.110 67.130 91.280 68.010 ;
        RECT 92.400 67.130 92.570 68.010 ;
        RECT 90.130 66.710 90.970 66.880 ;
        RECT 91.420 66.710 92.260 66.880 ;
        RECT 89.480 65.800 89.650 66.240 ;
        RECT 90.130 64.210 90.970 64.380 ;
        RECT 91.420 64.210 92.260 64.380 ;
        RECT 89.820 63.080 89.990 63.960 ;
        RECT 91.110 63.080 91.280 63.960 ;
        RECT 92.400 63.080 92.570 63.960 ;
        RECT 90.130 62.660 90.970 62.830 ;
        RECT 91.420 62.660 92.260 62.830 ;
        RECT 89.480 61.750 89.650 62.190 ;
        RECT 90.130 60.160 90.970 60.330 ;
        RECT 91.420 60.160 92.260 60.330 ;
        RECT 89.820 59.030 89.990 59.910 ;
        RECT 91.110 59.030 91.280 59.910 ;
        RECT 92.400 59.030 92.570 59.910 ;
        RECT 90.130 58.610 90.970 58.780 ;
        RECT 91.420 58.610 92.260 58.780 ;
        RECT 89.480 57.700 89.650 58.140 ;
        RECT 90.130 56.110 90.970 56.280 ;
        RECT 91.420 56.110 92.260 56.280 ;
        RECT 89.820 54.980 89.990 55.860 ;
        RECT 91.110 54.980 91.280 55.860 ;
        RECT 92.400 54.980 92.570 55.860 ;
        RECT 90.130 54.560 90.970 54.730 ;
        RECT 91.420 54.560 92.260 54.730 ;
        RECT 89.480 53.650 89.650 54.090 ;
        RECT 90.130 52.060 90.970 52.230 ;
        RECT 91.420 52.060 92.260 52.230 ;
        RECT 89.820 50.930 89.990 51.810 ;
        RECT 91.110 50.930 91.280 51.810 ;
        RECT 92.400 50.930 92.570 51.810 ;
        RECT 90.130 50.510 90.970 50.680 ;
        RECT 91.420 50.510 92.260 50.680 ;
        RECT 89.480 49.600 89.650 50.040 ;
        RECT 90.130 48.010 90.970 48.180 ;
        RECT 91.420 48.010 92.260 48.180 ;
        RECT 89.820 46.880 89.990 47.760 ;
        RECT 91.110 46.880 91.280 47.760 ;
        RECT 92.400 46.880 92.570 47.760 ;
        RECT 90.130 46.460 90.970 46.630 ;
        RECT 91.420 46.460 92.260 46.630 ;
        RECT 89.480 45.550 89.650 45.990 ;
        RECT 90.130 43.960 90.970 44.130 ;
        RECT 91.420 43.960 92.260 44.130 ;
        RECT 89.820 42.830 89.990 43.710 ;
        RECT 91.110 42.830 91.280 43.710 ;
        RECT 92.400 42.830 92.570 43.710 ;
        RECT 90.130 42.410 90.970 42.580 ;
        RECT 91.420 42.410 92.260 42.580 ;
        RECT 89.480 41.500 89.650 41.940 ;
        RECT 90.130 39.910 90.970 40.080 ;
        RECT 91.420 39.910 92.260 40.080 ;
        RECT 89.820 38.780 89.990 39.660 ;
        RECT 91.110 38.780 91.280 39.660 ;
        RECT 92.400 38.780 92.570 39.660 ;
        RECT 90.130 38.360 90.970 38.530 ;
        RECT 91.420 38.360 92.260 38.530 ;
        RECT 89.480 37.450 89.650 37.890 ;
        RECT 90.130 35.860 90.970 36.030 ;
        RECT 91.420 35.860 92.260 36.030 ;
        RECT 89.820 34.730 89.990 35.610 ;
        RECT 91.110 34.730 91.280 35.610 ;
        RECT 92.400 34.730 92.570 35.610 ;
        RECT 90.130 34.310 90.970 34.480 ;
        RECT 91.420 34.310 92.260 34.480 ;
        RECT 89.480 33.400 89.650 33.840 ;
        RECT 90.130 31.810 90.970 31.980 ;
        RECT 91.420 31.810 92.260 31.980 ;
        RECT 89.820 30.680 89.990 31.560 ;
        RECT 91.110 30.680 91.280 31.560 ;
        RECT 92.400 30.680 92.570 31.560 ;
        RECT 90.130 30.260 90.970 30.430 ;
        RECT 91.420 30.260 92.260 30.430 ;
        RECT 89.480 29.350 89.650 29.790 ;
        RECT 90.130 27.725 90.970 27.895 ;
        RECT 91.420 27.725 92.260 27.895 ;
        RECT 89.820 26.595 89.990 27.475 ;
        RECT 91.110 26.595 91.280 27.475 ;
        RECT 92.400 26.595 92.570 27.475 ;
        RECT 90.130 26.175 90.970 26.345 ;
        RECT 91.420 26.175 92.260 26.345 ;
        RECT 89.480 25.265 89.650 25.705 ;
        RECT 90.130 23.600 90.970 23.770 ;
        RECT 91.420 23.600 92.260 23.770 ;
        RECT 89.820 22.470 89.990 23.350 ;
        RECT 91.110 22.470 91.280 23.350 ;
        RECT 92.400 22.470 92.570 23.350 ;
        RECT 90.130 22.050 90.970 22.220 ;
        RECT 91.420 22.050 92.260 22.220 ;
        RECT 89.480 21.140 89.650 21.580 ;
        RECT 94.320 145.685 95.160 145.855 ;
        RECT 95.610 145.685 96.450 145.855 ;
        RECT 94.010 143.510 94.180 145.390 ;
        RECT 95.300 143.510 95.470 145.390 ;
        RECT 96.590 143.510 96.760 145.390 ;
        RECT 94.320 143.045 95.160 143.215 ;
        RECT 95.610 143.045 96.450 143.215 ;
        RECT 97.250 142.710 97.430 146.380 ;
        RECT 94.320 141.685 95.160 141.855 ;
        RECT 95.610 141.685 96.450 141.855 ;
        RECT 94.010 139.510 94.180 141.390 ;
        RECT 95.300 139.510 95.470 141.390 ;
        RECT 96.590 139.510 96.760 141.390 ;
        RECT 94.320 139.045 95.160 139.215 ;
        RECT 95.610 139.045 96.450 139.215 ;
        RECT 97.250 138.710 97.430 142.380 ;
        RECT 94.320 137.585 95.160 137.755 ;
        RECT 95.610 137.585 96.450 137.755 ;
        RECT 94.010 135.410 94.180 137.290 ;
        RECT 95.300 135.410 95.470 137.290 ;
        RECT 96.590 135.410 96.760 137.290 ;
        RECT 94.320 134.945 95.160 135.115 ;
        RECT 95.610 134.945 96.450 135.115 ;
        RECT 97.250 134.610 97.430 138.280 ;
        RECT 94.320 133.535 95.160 133.705 ;
        RECT 95.610 133.535 96.450 133.705 ;
        RECT 94.010 131.360 94.180 133.240 ;
        RECT 95.300 131.360 95.470 133.240 ;
        RECT 96.590 131.360 96.760 133.240 ;
        RECT 94.320 130.895 95.160 131.065 ;
        RECT 95.610 130.895 96.450 131.065 ;
        RECT 97.250 130.560 97.430 134.230 ;
        RECT 94.320 129.485 95.160 129.655 ;
        RECT 95.610 129.485 96.450 129.655 ;
        RECT 94.010 127.310 94.180 129.190 ;
        RECT 95.300 127.310 95.470 129.190 ;
        RECT 96.590 127.310 96.760 129.190 ;
        RECT 94.320 126.845 95.160 127.015 ;
        RECT 95.610 126.845 96.450 127.015 ;
        RECT 97.250 126.510 97.430 130.180 ;
        RECT 94.320 125.435 95.160 125.605 ;
        RECT 95.610 125.435 96.450 125.605 ;
        RECT 94.010 123.260 94.180 125.140 ;
        RECT 95.300 123.260 95.470 125.140 ;
        RECT 96.590 123.260 96.760 125.140 ;
        RECT 94.320 122.795 95.160 122.965 ;
        RECT 95.610 122.795 96.450 122.965 ;
        RECT 97.250 122.460 97.430 126.130 ;
        RECT 94.320 121.385 95.160 121.555 ;
        RECT 95.610 121.385 96.450 121.555 ;
        RECT 94.010 119.210 94.180 121.090 ;
        RECT 95.300 119.210 95.470 121.090 ;
        RECT 96.590 119.210 96.760 121.090 ;
        RECT 94.320 118.745 95.160 118.915 ;
        RECT 95.610 118.745 96.450 118.915 ;
        RECT 97.250 118.410 97.430 122.080 ;
        RECT 94.320 117.335 95.160 117.505 ;
        RECT 95.610 117.335 96.450 117.505 ;
        RECT 94.010 115.160 94.180 117.040 ;
        RECT 95.300 115.160 95.470 117.040 ;
        RECT 96.590 115.160 96.760 117.040 ;
        RECT 94.320 114.695 95.160 114.865 ;
        RECT 95.610 114.695 96.450 114.865 ;
        RECT 97.250 114.360 97.430 118.030 ;
        RECT 94.320 113.285 95.160 113.455 ;
        RECT 95.610 113.285 96.450 113.455 ;
        RECT 94.010 111.110 94.180 112.990 ;
        RECT 95.300 111.110 95.470 112.990 ;
        RECT 96.590 111.110 96.760 112.990 ;
        RECT 94.320 110.645 95.160 110.815 ;
        RECT 95.610 110.645 96.450 110.815 ;
        RECT 97.250 110.310 97.430 113.980 ;
        RECT 94.320 109.235 95.160 109.405 ;
        RECT 95.610 109.235 96.450 109.405 ;
        RECT 94.010 107.060 94.180 108.940 ;
        RECT 95.300 107.060 95.470 108.940 ;
        RECT 96.590 107.060 96.760 108.940 ;
        RECT 94.320 106.595 95.160 106.765 ;
        RECT 95.610 106.595 96.450 106.765 ;
        RECT 97.250 106.260 97.430 109.930 ;
        RECT 94.320 105.185 95.160 105.355 ;
        RECT 95.610 105.185 96.450 105.355 ;
        RECT 94.010 103.010 94.180 104.890 ;
        RECT 95.300 103.010 95.470 104.890 ;
        RECT 96.590 103.010 96.760 104.890 ;
        RECT 94.320 102.545 95.160 102.715 ;
        RECT 95.610 102.545 96.450 102.715 ;
        RECT 97.250 102.210 97.430 105.880 ;
        RECT 94.320 101.135 95.160 101.305 ;
        RECT 95.610 101.135 96.450 101.305 ;
        RECT 94.010 98.960 94.180 100.840 ;
        RECT 95.300 98.960 95.470 100.840 ;
        RECT 96.590 98.960 96.760 100.840 ;
        RECT 94.320 98.495 95.160 98.665 ;
        RECT 95.610 98.495 96.450 98.665 ;
        RECT 97.250 98.160 97.430 101.830 ;
        RECT 94.320 97.085 95.160 97.255 ;
        RECT 95.610 97.085 96.450 97.255 ;
        RECT 94.010 94.910 94.180 96.790 ;
        RECT 95.300 94.910 95.470 96.790 ;
        RECT 96.590 94.910 96.760 96.790 ;
        RECT 94.320 94.445 95.160 94.615 ;
        RECT 95.610 94.445 96.450 94.615 ;
        RECT 97.250 94.110 97.430 97.780 ;
        RECT 94.320 93.035 95.160 93.205 ;
        RECT 95.610 93.035 96.450 93.205 ;
        RECT 94.010 90.860 94.180 92.740 ;
        RECT 95.300 90.860 95.470 92.740 ;
        RECT 96.590 90.860 96.760 92.740 ;
        RECT 94.320 90.395 95.160 90.565 ;
        RECT 95.610 90.395 96.450 90.565 ;
        RECT 97.250 90.060 97.430 93.730 ;
        RECT 94.320 88.985 95.160 89.155 ;
        RECT 95.610 88.985 96.450 89.155 ;
        RECT 94.010 86.810 94.180 88.690 ;
        RECT 95.300 86.810 95.470 88.690 ;
        RECT 96.590 86.810 96.760 88.690 ;
        RECT 94.320 86.345 95.160 86.515 ;
        RECT 95.610 86.345 96.450 86.515 ;
        RECT 97.250 86.010 97.430 89.680 ;
        RECT 94.320 84.935 95.160 85.105 ;
        RECT 95.610 84.935 96.450 85.105 ;
        RECT 94.010 82.760 94.180 84.640 ;
        RECT 95.300 82.760 95.470 84.640 ;
        RECT 96.590 82.760 96.760 84.640 ;
        RECT 94.320 82.295 95.160 82.465 ;
        RECT 95.610 82.295 96.450 82.465 ;
        RECT 97.250 81.960 97.430 85.630 ;
        RECT 94.320 80.885 95.160 81.055 ;
        RECT 95.610 80.885 96.450 81.055 ;
        RECT 94.010 78.710 94.180 80.590 ;
        RECT 95.300 78.710 95.470 80.590 ;
        RECT 96.590 78.710 96.760 80.590 ;
        RECT 94.320 78.245 95.160 78.415 ;
        RECT 95.610 78.245 96.450 78.415 ;
        RECT 97.250 77.910 97.430 81.580 ;
        RECT 94.320 76.835 95.160 77.005 ;
        RECT 95.610 76.835 96.450 77.005 ;
        RECT 94.010 74.660 94.180 76.540 ;
        RECT 95.300 74.660 95.470 76.540 ;
        RECT 96.590 74.660 96.760 76.540 ;
        RECT 94.320 74.195 95.160 74.365 ;
        RECT 95.610 74.195 96.450 74.365 ;
        RECT 97.250 73.860 97.430 77.530 ;
        RECT 94.320 72.785 95.160 72.955 ;
        RECT 95.610 72.785 96.450 72.955 ;
        RECT 94.010 70.610 94.180 72.490 ;
        RECT 95.300 70.610 95.470 72.490 ;
        RECT 96.590 70.610 96.760 72.490 ;
        RECT 94.320 70.145 95.160 70.315 ;
        RECT 95.610 70.145 96.450 70.315 ;
        RECT 97.250 69.810 97.430 73.480 ;
        RECT 94.320 68.735 95.160 68.905 ;
        RECT 95.610 68.735 96.450 68.905 ;
        RECT 94.010 66.560 94.180 68.440 ;
        RECT 95.300 66.560 95.470 68.440 ;
        RECT 96.590 66.560 96.760 68.440 ;
        RECT 94.320 66.095 95.160 66.265 ;
        RECT 95.610 66.095 96.450 66.265 ;
        RECT 97.250 65.760 97.430 69.430 ;
        RECT 94.320 64.685 95.160 64.855 ;
        RECT 95.610 64.685 96.450 64.855 ;
        RECT 94.010 62.510 94.180 64.390 ;
        RECT 95.300 62.510 95.470 64.390 ;
        RECT 96.590 62.510 96.760 64.390 ;
        RECT 94.320 62.045 95.160 62.215 ;
        RECT 95.610 62.045 96.450 62.215 ;
        RECT 97.250 61.710 97.430 65.380 ;
        RECT 94.320 60.635 95.160 60.805 ;
        RECT 95.610 60.635 96.450 60.805 ;
        RECT 94.010 58.460 94.180 60.340 ;
        RECT 95.300 58.460 95.470 60.340 ;
        RECT 96.590 58.460 96.760 60.340 ;
        RECT 94.320 57.995 95.160 58.165 ;
        RECT 95.610 57.995 96.450 58.165 ;
        RECT 97.250 57.660 97.430 61.330 ;
        RECT 97.770 142.710 97.950 146.380 ;
        RECT 98.750 145.685 99.590 145.855 ;
        RECT 100.040 145.685 100.880 145.855 ;
        RECT 98.440 143.510 98.610 145.390 ;
        RECT 99.730 143.510 99.900 145.390 ;
        RECT 101.020 143.510 101.190 145.390 ;
        RECT 98.750 143.045 99.590 143.215 ;
        RECT 100.040 143.045 100.880 143.215 ;
        RECT 97.770 138.650 97.950 142.320 ;
        RECT 98.750 141.625 99.590 141.795 ;
        RECT 100.040 141.625 100.880 141.795 ;
        RECT 98.440 139.450 98.610 141.330 ;
        RECT 99.730 139.450 99.900 141.330 ;
        RECT 101.020 139.450 101.190 141.330 ;
        RECT 98.750 138.985 99.590 139.155 ;
        RECT 100.040 138.985 100.880 139.155 ;
        RECT 97.770 134.590 97.950 138.260 ;
        RECT 98.750 137.565 99.590 137.735 ;
        RECT 100.040 137.565 100.880 137.735 ;
        RECT 98.440 135.390 98.610 137.270 ;
        RECT 99.730 135.390 99.900 137.270 ;
        RECT 101.020 135.390 101.190 137.270 ;
        RECT 98.750 134.925 99.590 135.095 ;
        RECT 100.040 134.925 100.880 135.095 ;
        RECT 97.770 130.530 97.950 134.200 ;
        RECT 98.750 133.505 99.590 133.675 ;
        RECT 100.040 133.505 100.880 133.675 ;
        RECT 98.440 131.330 98.610 133.210 ;
        RECT 99.730 131.330 99.900 133.210 ;
        RECT 101.020 131.330 101.190 133.210 ;
        RECT 98.750 130.865 99.590 131.035 ;
        RECT 100.040 130.865 100.880 131.035 ;
        RECT 97.770 126.470 97.950 130.140 ;
        RECT 98.750 129.445 99.590 129.615 ;
        RECT 100.040 129.445 100.880 129.615 ;
        RECT 98.440 127.270 98.610 129.150 ;
        RECT 99.730 127.270 99.900 129.150 ;
        RECT 101.020 127.270 101.190 129.150 ;
        RECT 98.750 126.805 99.590 126.975 ;
        RECT 100.040 126.805 100.880 126.975 ;
        RECT 97.770 122.410 97.950 126.080 ;
        RECT 98.750 125.385 99.590 125.555 ;
        RECT 100.040 125.385 100.880 125.555 ;
        RECT 98.440 123.210 98.610 125.090 ;
        RECT 99.730 123.210 99.900 125.090 ;
        RECT 101.020 123.210 101.190 125.090 ;
        RECT 98.750 122.745 99.590 122.915 ;
        RECT 100.040 122.745 100.880 122.915 ;
        RECT 97.770 118.350 97.950 122.020 ;
        RECT 98.750 121.325 99.590 121.495 ;
        RECT 100.040 121.325 100.880 121.495 ;
        RECT 98.440 119.150 98.610 121.030 ;
        RECT 99.730 119.150 99.900 121.030 ;
        RECT 101.020 119.150 101.190 121.030 ;
        RECT 98.750 118.685 99.590 118.855 ;
        RECT 100.040 118.685 100.880 118.855 ;
        RECT 97.770 114.290 97.950 117.960 ;
        RECT 98.750 117.265 99.590 117.435 ;
        RECT 100.040 117.265 100.880 117.435 ;
        RECT 98.440 115.090 98.610 116.970 ;
        RECT 99.730 115.090 99.900 116.970 ;
        RECT 101.020 115.090 101.190 116.970 ;
        RECT 98.750 114.625 99.590 114.795 ;
        RECT 100.040 114.625 100.880 114.795 ;
        RECT 97.770 110.230 97.950 113.900 ;
        RECT 98.750 113.205 99.590 113.375 ;
        RECT 100.040 113.205 100.880 113.375 ;
        RECT 98.440 111.030 98.610 112.910 ;
        RECT 99.730 111.030 99.900 112.910 ;
        RECT 101.020 111.030 101.190 112.910 ;
        RECT 98.750 110.565 99.590 110.735 ;
        RECT 100.040 110.565 100.880 110.735 ;
        RECT 97.770 106.170 97.950 109.840 ;
        RECT 98.750 109.145 99.590 109.315 ;
        RECT 100.040 109.145 100.880 109.315 ;
        RECT 98.440 106.970 98.610 108.850 ;
        RECT 99.730 106.970 99.900 108.850 ;
        RECT 101.020 106.970 101.190 108.850 ;
        RECT 98.750 106.505 99.590 106.675 ;
        RECT 100.040 106.505 100.880 106.675 ;
        RECT 97.770 102.110 97.950 105.780 ;
        RECT 98.750 105.085 99.590 105.255 ;
        RECT 100.040 105.085 100.880 105.255 ;
        RECT 98.440 102.910 98.610 104.790 ;
        RECT 99.730 102.910 99.900 104.790 ;
        RECT 101.020 102.910 101.190 104.790 ;
        RECT 98.750 102.445 99.590 102.615 ;
        RECT 100.040 102.445 100.880 102.615 ;
        RECT 97.770 98.050 97.950 101.720 ;
        RECT 98.750 101.025 99.590 101.195 ;
        RECT 100.040 101.025 100.880 101.195 ;
        RECT 98.440 98.850 98.610 100.730 ;
        RECT 99.730 98.850 99.900 100.730 ;
        RECT 101.020 98.850 101.190 100.730 ;
        RECT 98.750 98.385 99.590 98.555 ;
        RECT 100.040 98.385 100.880 98.555 ;
        RECT 97.770 93.990 97.950 97.660 ;
        RECT 98.750 96.965 99.590 97.135 ;
        RECT 100.040 96.965 100.880 97.135 ;
        RECT 98.440 94.790 98.610 96.670 ;
        RECT 99.730 94.790 99.900 96.670 ;
        RECT 101.020 94.790 101.190 96.670 ;
        RECT 98.750 94.325 99.590 94.495 ;
        RECT 100.040 94.325 100.880 94.495 ;
        RECT 97.770 89.930 97.950 93.600 ;
        RECT 98.750 92.905 99.590 93.075 ;
        RECT 100.040 92.905 100.880 93.075 ;
        RECT 98.440 90.730 98.610 92.610 ;
        RECT 99.730 90.730 99.900 92.610 ;
        RECT 101.020 90.730 101.190 92.610 ;
        RECT 98.750 90.265 99.590 90.435 ;
        RECT 100.040 90.265 100.880 90.435 ;
        RECT 97.770 85.870 97.950 89.540 ;
        RECT 98.750 88.845 99.590 89.015 ;
        RECT 100.040 88.845 100.880 89.015 ;
        RECT 98.440 86.670 98.610 88.550 ;
        RECT 99.730 86.670 99.900 88.550 ;
        RECT 101.020 86.670 101.190 88.550 ;
        RECT 98.750 86.205 99.590 86.375 ;
        RECT 100.040 86.205 100.880 86.375 ;
        RECT 97.770 81.810 97.950 85.480 ;
        RECT 98.750 84.785 99.590 84.955 ;
        RECT 100.040 84.785 100.880 84.955 ;
        RECT 98.440 82.610 98.610 84.490 ;
        RECT 99.730 82.610 99.900 84.490 ;
        RECT 101.020 82.610 101.190 84.490 ;
        RECT 98.750 82.145 99.590 82.315 ;
        RECT 100.040 82.145 100.880 82.315 ;
        RECT 97.770 77.750 97.950 81.420 ;
        RECT 98.750 80.725 99.590 80.895 ;
        RECT 100.040 80.725 100.880 80.895 ;
        RECT 98.440 78.550 98.610 80.430 ;
        RECT 99.730 78.550 99.900 80.430 ;
        RECT 101.020 78.550 101.190 80.430 ;
        RECT 98.750 78.085 99.590 78.255 ;
        RECT 100.040 78.085 100.880 78.255 ;
        RECT 97.770 73.690 97.950 77.360 ;
        RECT 98.750 76.665 99.590 76.835 ;
        RECT 100.040 76.665 100.880 76.835 ;
        RECT 98.440 74.490 98.610 76.370 ;
        RECT 99.730 74.490 99.900 76.370 ;
        RECT 101.020 74.490 101.190 76.370 ;
        RECT 98.750 74.025 99.590 74.195 ;
        RECT 100.040 74.025 100.880 74.195 ;
        RECT 97.770 69.630 97.950 73.300 ;
        RECT 98.750 72.605 99.590 72.775 ;
        RECT 100.040 72.605 100.880 72.775 ;
        RECT 98.440 70.430 98.610 72.310 ;
        RECT 99.730 70.430 99.900 72.310 ;
        RECT 101.020 70.430 101.190 72.310 ;
        RECT 98.750 69.965 99.590 70.135 ;
        RECT 100.040 69.965 100.880 70.135 ;
        RECT 97.770 65.570 97.950 69.240 ;
        RECT 98.750 68.545 99.590 68.715 ;
        RECT 100.040 68.545 100.880 68.715 ;
        RECT 98.440 66.370 98.610 68.250 ;
        RECT 99.730 66.370 99.900 68.250 ;
        RECT 101.020 66.370 101.190 68.250 ;
        RECT 98.750 65.905 99.590 66.075 ;
        RECT 100.040 65.905 100.880 66.075 ;
        RECT 97.770 61.510 97.950 65.180 ;
        RECT 98.750 64.485 99.590 64.655 ;
        RECT 100.040 64.485 100.880 64.655 ;
        RECT 98.440 62.310 98.610 64.190 ;
        RECT 99.730 62.310 99.900 64.190 ;
        RECT 101.020 62.310 101.190 64.190 ;
        RECT 98.750 61.845 99.590 62.015 ;
        RECT 100.040 61.845 100.880 62.015 ;
        RECT 138.520 146.260 139.140 146.440 ;
        RECT 102.940 145.210 103.780 145.380 ;
        RECT 104.230 145.210 105.070 145.380 ;
        RECT 102.630 144.080 102.800 144.960 ;
        RECT 103.920 144.080 104.090 144.960 ;
        RECT 105.210 144.080 105.380 144.960 ;
        RECT 102.940 143.660 103.780 143.830 ;
        RECT 104.230 143.660 105.070 143.830 ;
        RECT 105.550 142.750 105.720 143.190 ;
        RECT 102.940 141.150 103.780 141.320 ;
        RECT 104.230 141.150 105.070 141.320 ;
        RECT 102.630 140.020 102.800 140.900 ;
        RECT 103.920 140.020 104.090 140.900 ;
        RECT 105.210 140.020 105.380 140.900 ;
        RECT 102.940 139.600 103.780 139.770 ;
        RECT 104.230 139.600 105.070 139.770 ;
        RECT 105.550 138.690 105.720 139.130 ;
        RECT 102.940 137.090 103.780 137.260 ;
        RECT 104.230 137.090 105.070 137.260 ;
        RECT 102.630 135.960 102.800 136.840 ;
        RECT 103.920 135.960 104.090 136.840 ;
        RECT 105.210 135.960 105.380 136.840 ;
        RECT 102.940 135.540 103.780 135.710 ;
        RECT 104.230 135.540 105.070 135.710 ;
        RECT 105.550 134.630 105.720 135.070 ;
        RECT 106.110 134.780 106.280 144.490 ;
        RECT 108.630 144.190 113.510 144.360 ;
        RECT 108.210 143.210 108.380 144.050 ;
        RECT 113.760 143.210 113.930 144.050 ;
        RECT 108.630 142.900 113.510 143.070 ;
        RECT 108.210 141.920 108.380 142.760 ;
        RECT 113.760 141.920 113.930 142.760 ;
        RECT 108.630 141.610 113.510 141.780 ;
        RECT 108.210 140.630 108.380 141.470 ;
        RECT 113.760 140.630 113.930 141.470 ;
        RECT 108.630 140.320 113.510 140.490 ;
        RECT 108.210 139.340 108.380 140.180 ;
        RECT 113.760 139.340 113.930 140.180 ;
        RECT 108.630 139.030 113.510 139.200 ;
        RECT 108.210 138.050 108.380 138.890 ;
        RECT 113.760 138.050 113.930 138.890 ;
        RECT 108.630 137.740 113.510 137.910 ;
        RECT 108.210 136.760 108.380 137.600 ;
        RECT 113.760 136.760 113.930 137.600 ;
        RECT 108.630 136.450 113.510 136.620 ;
        RECT 108.210 135.470 108.380 136.310 ;
        RECT 113.760 135.470 113.930 136.310 ;
        RECT 108.630 135.160 113.510 135.330 ;
        RECT 108.210 134.180 108.380 135.020 ;
        RECT 113.760 134.180 113.930 135.020 ;
        RECT 108.630 133.870 113.510 134.040 ;
        RECT 115.370 143.420 115.540 145.630 ;
        RECT 117.090 144.470 121.970 144.640 ;
        RECT 124.090 144.470 128.970 144.640 ;
        RECT 116.670 143.490 116.840 144.330 ;
        RECT 122.220 143.490 122.390 144.330 ;
        RECT 123.670 143.490 123.840 144.330 ;
        RECT 129.220 143.490 129.390 144.330 ;
        RECT 117.090 143.180 121.970 143.350 ;
        RECT 124.090 143.180 128.970 143.350 ;
        RECT 117.090 142.470 121.970 142.640 ;
        RECT 124.090 142.470 128.970 142.640 ;
        RECT 116.670 141.490 116.840 142.330 ;
        RECT 122.220 141.490 122.390 142.330 ;
        RECT 123.670 141.490 123.840 142.330 ;
        RECT 129.220 141.490 129.390 142.330 ;
        RECT 117.090 141.180 121.970 141.350 ;
        RECT 124.090 141.180 128.970 141.350 ;
        RECT 117.090 138.470 121.970 138.640 ;
        RECT 124.090 138.470 128.970 138.640 ;
        RECT 116.670 137.490 116.840 138.330 ;
        RECT 122.220 137.490 122.390 138.330 ;
        RECT 123.670 137.490 123.840 138.330 ;
        RECT 129.220 137.490 129.390 138.330 ;
        RECT 117.090 137.180 121.970 137.350 ;
        RECT 124.090 137.180 128.970 137.350 ;
        RECT 117.090 136.470 121.970 136.640 ;
        RECT 124.090 136.470 128.970 136.640 ;
        RECT 116.670 135.490 116.840 136.330 ;
        RECT 122.220 135.490 122.390 136.330 ;
        RECT 123.670 135.490 123.840 136.330 ;
        RECT 129.220 135.490 129.390 136.330 ;
        RECT 117.090 135.180 121.970 135.350 ;
        RECT 124.090 135.180 128.970 135.350 ;
        RECT 132.810 145.450 137.690 145.620 ;
        RECT 141.810 145.450 146.690 145.620 ;
        RECT 132.345 144.970 132.515 145.310 ;
        RECT 137.985 144.970 138.155 145.310 ;
        RECT 141.345 144.970 141.515 145.310 ;
        RECT 146.985 144.970 147.155 145.310 ;
        RECT 132.810 144.660 137.690 144.830 ;
        RECT 141.810 144.660 146.690 144.830 ;
        RECT 132.810 140.950 137.690 141.120 ;
        RECT 141.810 140.950 146.690 141.120 ;
        RECT 132.345 140.470 132.515 140.810 ;
        RECT 137.985 140.470 138.155 140.810 ;
        RECT 141.345 140.470 141.515 140.810 ;
        RECT 146.985 140.470 147.155 140.810 ;
        RECT 132.810 140.160 137.690 140.330 ;
        RECT 141.810 140.160 146.690 140.330 ;
        RECT 132.810 136.450 137.690 136.620 ;
        RECT 141.810 136.450 146.690 136.620 ;
        RECT 132.345 135.970 132.515 136.310 ;
        RECT 137.985 135.970 138.155 136.310 ;
        RECT 141.345 135.970 141.515 136.310 ;
        RECT 146.985 135.970 147.155 136.310 ;
        RECT 132.810 135.660 137.690 135.830 ;
        RECT 141.810 135.660 146.690 135.830 ;
        RECT 147.520 134.160 147.700 145.830 ;
        RECT 138.410 133.420 139.470 133.600 ;
        RECT 102.940 133.030 103.780 133.200 ;
        RECT 104.230 133.030 105.070 133.200 ;
        RECT 102.630 131.900 102.800 132.780 ;
        RECT 103.920 131.900 104.090 132.780 ;
        RECT 105.210 131.900 105.380 132.780 ;
        RECT 102.940 131.480 103.780 131.650 ;
        RECT 104.230 131.480 105.070 131.650 ;
        RECT 105.550 130.570 105.720 131.010 ;
        RECT 106.510 132.630 107.150 132.800 ;
        RECT 108.160 132.630 108.800 132.800 ;
        RECT 109.560 132.630 110.200 132.800 ;
        RECT 110.740 132.630 111.380 132.800 ;
        RECT 106.030 130.680 106.200 132.320 ;
        RECT 106.960 132.055 111.840 132.225 ;
        RECT 106.540 131.075 106.710 131.915 ;
        RECT 112.090 131.075 112.260 131.915 ;
        RECT 106.960 130.765 111.840 130.935 ;
        RECT 123.660 132.630 124.230 132.800 ;
        RECT 114.105 132.060 114.985 132.230 ;
        RECT 113.640 131.580 113.810 131.920 ;
        RECT 115.280 131.580 115.450 131.920 ;
        RECT 114.105 131.270 114.985 131.440 ;
        RECT 116.765 132.060 124.145 132.230 ;
        RECT 116.300 131.580 116.470 131.920 ;
        RECT 124.440 131.580 124.610 131.920 ;
        RECT 116.765 131.270 124.145 131.440 ;
        RECT 124.950 131.180 125.120 132.320 ;
        RECT 117.020 130.700 121.970 130.870 ;
        RECT 122.800 130.700 123.940 130.870 ;
        RECT 117.020 130.260 121.970 130.430 ;
        RECT 102.940 128.970 103.780 129.140 ;
        RECT 104.230 128.970 105.070 129.140 ;
        RECT 102.630 127.840 102.800 128.720 ;
        RECT 103.920 127.840 104.090 128.720 ;
        RECT 105.210 127.840 105.380 128.720 ;
        RECT 102.940 127.420 103.780 127.590 ;
        RECT 104.230 127.420 105.070 127.590 ;
        RECT 105.550 126.510 105.720 126.950 ;
        RECT 116.770 129.685 123.650 129.855 ;
        RECT 116.305 129.205 116.475 129.545 ;
        RECT 123.945 129.205 124.115 129.545 ;
        RECT 116.770 128.895 123.650 129.065 ;
        RECT 124.450 128.810 124.620 129.950 ;
        RECT 116.770 127.755 123.650 127.925 ;
        RECT 116.305 127.275 116.475 127.615 ;
        RECT 123.945 127.275 124.115 127.615 ;
        RECT 116.770 126.965 123.650 127.135 ;
        RECT 124.450 126.880 124.620 128.020 ;
        RECT 102.940 124.910 103.780 125.080 ;
        RECT 104.230 124.910 105.070 125.080 ;
        RECT 102.630 123.780 102.800 124.660 ;
        RECT 103.920 123.780 104.090 124.660 ;
        RECT 105.210 123.780 105.380 124.660 ;
        RECT 102.940 123.360 103.780 123.530 ;
        RECT 104.230 123.360 105.070 123.530 ;
        RECT 105.550 122.450 105.720 122.890 ;
        RECT 107.160 124.840 112.040 125.010 ;
        RECT 106.140 122.900 106.310 124.370 ;
        RECT 106.740 124.360 106.910 124.700 ;
        RECT 112.290 124.360 112.460 124.700 ;
        RECT 107.160 124.050 112.040 124.220 ;
        RECT 106.740 123.570 106.910 123.910 ;
        RECT 112.290 123.570 112.460 123.910 ;
        RECT 107.160 123.260 112.040 123.430 ;
        RECT 106.740 122.780 106.910 123.120 ;
        RECT 112.290 122.780 112.460 123.120 ;
        RECT 107.160 122.470 112.040 122.640 ;
        RECT 106.740 121.990 106.910 122.330 ;
        RECT 112.290 121.990 112.460 122.330 ;
        RECT 107.160 121.680 112.040 121.850 ;
        RECT 102.940 120.850 103.780 121.020 ;
        RECT 104.230 120.850 105.070 121.020 ;
        RECT 102.630 119.720 102.800 120.600 ;
        RECT 103.920 119.720 104.090 120.600 ;
        RECT 105.210 119.720 105.380 120.600 ;
        RECT 102.940 119.300 103.780 119.470 ;
        RECT 104.230 119.300 105.070 119.470 ;
        RECT 105.550 118.390 105.720 118.830 ;
        RECT 106.140 120.070 106.310 121.540 ;
        RECT 106.740 121.200 106.910 121.540 ;
        RECT 112.290 121.200 112.460 121.540 ;
        RECT 107.160 120.890 112.040 121.060 ;
        RECT 106.740 120.410 106.910 120.750 ;
        RECT 112.290 120.410 112.460 120.750 ;
        RECT 107.160 120.100 112.040 120.270 ;
        RECT 106.740 119.620 106.910 119.960 ;
        RECT 112.290 119.620 112.460 119.960 ;
        RECT 107.160 119.310 112.040 119.480 ;
        RECT 106.140 117.720 106.310 119.190 ;
        RECT 106.740 118.830 106.910 119.170 ;
        RECT 112.290 118.830 112.460 119.170 ;
        RECT 107.160 118.520 112.040 118.690 ;
        RECT 106.740 118.040 106.910 118.380 ;
        RECT 112.290 118.040 112.460 118.380 ;
        RECT 107.160 117.730 112.040 117.900 ;
        RECT 102.940 116.790 103.780 116.960 ;
        RECT 104.230 116.790 105.070 116.960 ;
        RECT 102.630 115.660 102.800 116.540 ;
        RECT 103.920 115.660 104.090 116.540 ;
        RECT 105.210 115.660 105.380 116.540 ;
        RECT 102.940 115.240 103.780 115.410 ;
        RECT 104.230 115.240 105.070 115.410 ;
        RECT 105.550 114.330 105.720 114.770 ;
        RECT 106.740 117.250 106.910 117.590 ;
        RECT 112.290 117.250 112.460 117.590 ;
        RECT 107.160 116.940 112.040 117.110 ;
        RECT 106.140 115.200 106.310 116.670 ;
        RECT 106.740 116.460 106.910 116.800 ;
        RECT 112.290 116.460 112.460 116.800 ;
        RECT 107.160 116.150 112.040 116.320 ;
        RECT 106.740 115.670 106.910 116.010 ;
        RECT 112.290 115.670 112.460 116.010 ;
        RECT 107.160 115.360 112.040 115.530 ;
        RECT 106.740 114.880 106.910 115.220 ;
        RECT 112.290 114.880 112.460 115.220 ;
        RECT 107.160 114.570 112.040 114.740 ;
        RECT 102.940 112.730 103.780 112.900 ;
        RECT 104.230 112.730 105.070 112.900 ;
        RECT 102.630 111.600 102.800 112.480 ;
        RECT 103.920 111.600 104.090 112.480 ;
        RECT 105.210 111.600 105.380 112.480 ;
        RECT 102.940 111.180 103.780 111.350 ;
        RECT 104.230 111.180 105.070 111.350 ;
        RECT 105.550 110.270 105.720 110.710 ;
        RECT 106.140 112.620 106.310 114.090 ;
        RECT 106.740 114.090 106.910 114.430 ;
        RECT 112.290 114.090 112.460 114.430 ;
        RECT 107.160 113.780 112.040 113.950 ;
        RECT 106.740 113.300 106.910 113.640 ;
        RECT 112.290 113.300 112.460 113.640 ;
        RECT 107.160 112.990 112.040 113.160 ;
        RECT 106.740 112.510 106.910 112.850 ;
        RECT 112.290 112.510 112.460 112.850 ;
        RECT 107.160 112.200 112.040 112.370 ;
        RECT 106.740 111.720 106.910 112.060 ;
        RECT 112.290 111.720 112.460 112.060 ;
        RECT 106.140 110.050 106.310 111.520 ;
        RECT 107.160 111.410 112.040 111.580 ;
        RECT 106.740 110.930 106.910 111.270 ;
        RECT 112.290 110.930 112.460 111.270 ;
        RECT 107.160 110.620 112.040 110.790 ;
        RECT 106.740 110.140 106.910 110.480 ;
        RECT 112.290 110.140 112.460 110.480 ;
        RECT 107.160 109.830 112.040 110.000 ;
        RECT 115.220 124.660 120.100 124.830 ;
        RECT 114.755 124.180 114.925 124.520 ;
        RECT 120.395 124.180 120.565 124.520 ;
        RECT 115.220 123.870 120.100 124.040 ;
        RECT 114.755 123.390 114.925 123.730 ;
        RECT 120.395 123.390 120.565 123.730 ;
        RECT 115.220 123.080 120.100 123.250 ;
        RECT 120.860 123.170 121.030 124.310 ;
        RECT 114.755 122.600 114.925 122.940 ;
        RECT 120.395 122.600 120.565 122.940 ;
        RECT 115.220 122.290 120.100 122.460 ;
        RECT 114.755 121.810 114.925 122.150 ;
        RECT 120.395 121.810 120.565 122.150 ;
        RECT 115.220 121.500 120.100 121.670 ;
        RECT 114.755 121.020 114.925 121.360 ;
        RECT 120.395 121.020 120.565 121.360 ;
        RECT 120.860 120.930 121.030 122.070 ;
        RECT 115.220 120.710 120.100 120.880 ;
        RECT 114.755 120.230 114.925 120.570 ;
        RECT 120.395 120.230 120.565 120.570 ;
        RECT 115.220 119.920 120.100 120.090 ;
        RECT 114.755 119.440 114.925 119.780 ;
        RECT 120.395 119.440 120.565 119.780 ;
        RECT 115.220 119.130 120.100 119.300 ;
        RECT 114.755 118.650 114.925 118.990 ;
        RECT 120.395 118.650 120.565 118.990 ;
        RECT 120.860 118.630 121.030 119.770 ;
        RECT 115.220 118.340 120.100 118.510 ;
        RECT 114.755 117.860 114.925 118.200 ;
        RECT 120.395 117.860 120.565 118.200 ;
        RECT 115.220 117.550 120.100 117.720 ;
        RECT 114.755 117.070 114.925 117.410 ;
        RECT 120.395 117.070 120.565 117.410 ;
        RECT 115.220 116.760 120.100 116.930 ;
        RECT 114.755 116.280 114.925 116.620 ;
        RECT 120.395 116.280 120.565 116.620 ;
        RECT 120.860 116.190 121.030 117.330 ;
        RECT 115.220 115.970 120.100 116.140 ;
        RECT 114.755 115.490 114.925 115.830 ;
        RECT 120.395 115.490 120.565 115.830 ;
        RECT 115.220 115.180 120.100 115.350 ;
        RECT 114.755 114.700 114.925 115.040 ;
        RECT 120.395 114.700 120.565 115.040 ;
        RECT 115.220 114.390 120.100 114.560 ;
        RECT 114.755 113.910 114.925 114.250 ;
        RECT 120.395 113.910 120.565 114.250 ;
        RECT 120.860 113.790 121.030 114.930 ;
        RECT 115.220 113.600 120.100 113.770 ;
        RECT 102.940 108.670 103.780 108.840 ;
        RECT 104.230 108.670 105.070 108.840 ;
        RECT 102.630 107.540 102.800 108.420 ;
        RECT 103.920 107.540 104.090 108.420 ;
        RECT 105.210 107.540 105.380 108.420 ;
        RECT 102.940 107.120 103.780 107.290 ;
        RECT 104.230 107.120 105.070 107.290 ;
        RECT 105.550 106.210 105.720 106.650 ;
        RECT 138.520 108.340 139.140 108.520 ;
        RECT 102.940 104.610 103.780 104.780 ;
        RECT 104.230 104.610 105.070 104.780 ;
        RECT 102.630 103.480 102.800 104.360 ;
        RECT 103.920 103.480 104.090 104.360 ;
        RECT 105.210 103.480 105.380 104.360 ;
        RECT 102.940 103.060 103.780 103.230 ;
        RECT 104.230 103.060 105.070 103.230 ;
        RECT 105.550 102.150 105.720 102.590 ;
        RECT 102.940 100.550 103.780 100.720 ;
        RECT 104.230 100.550 105.070 100.720 ;
        RECT 102.630 99.420 102.800 100.300 ;
        RECT 103.920 99.420 104.090 100.300 ;
        RECT 105.210 99.420 105.380 100.300 ;
        RECT 102.940 99.000 103.780 99.170 ;
        RECT 104.230 99.000 105.070 99.170 ;
        RECT 105.550 98.090 105.720 98.530 ;
        RECT 106.110 96.860 106.280 106.570 ;
        RECT 108.630 106.270 113.510 106.440 ;
        RECT 108.210 105.290 108.380 106.130 ;
        RECT 113.760 105.290 113.930 106.130 ;
        RECT 108.630 104.980 113.510 105.150 ;
        RECT 108.210 104.000 108.380 104.840 ;
        RECT 113.760 104.000 113.930 104.840 ;
        RECT 108.630 103.690 113.510 103.860 ;
        RECT 108.210 102.710 108.380 103.550 ;
        RECT 113.760 102.710 113.930 103.550 ;
        RECT 108.630 102.400 113.510 102.570 ;
        RECT 108.210 101.420 108.380 102.260 ;
        RECT 113.760 101.420 113.930 102.260 ;
        RECT 108.630 101.110 113.510 101.280 ;
        RECT 108.210 100.130 108.380 100.970 ;
        RECT 113.760 100.130 113.930 100.970 ;
        RECT 108.630 99.820 113.510 99.990 ;
        RECT 108.210 98.840 108.380 99.680 ;
        RECT 113.760 98.840 113.930 99.680 ;
        RECT 108.630 98.530 113.510 98.700 ;
        RECT 108.210 97.550 108.380 98.390 ;
        RECT 113.760 97.550 113.930 98.390 ;
        RECT 108.630 97.240 113.510 97.410 ;
        RECT 102.940 96.490 103.780 96.660 ;
        RECT 104.230 96.490 105.070 96.660 ;
        RECT 102.630 95.360 102.800 96.240 ;
        RECT 103.920 95.360 104.090 96.240 ;
        RECT 105.210 95.360 105.380 96.240 ;
        RECT 102.940 94.940 103.780 95.110 ;
        RECT 104.230 94.940 105.070 95.110 ;
        RECT 108.210 96.260 108.380 97.100 ;
        RECT 113.760 96.260 113.930 97.100 ;
        RECT 108.630 95.950 113.510 96.120 ;
        RECT 115.370 105.500 115.540 107.710 ;
        RECT 117.090 106.550 121.970 106.720 ;
        RECT 124.090 106.550 128.970 106.720 ;
        RECT 116.670 105.570 116.840 106.410 ;
        RECT 122.220 105.570 122.390 106.410 ;
        RECT 123.670 105.570 123.840 106.410 ;
        RECT 129.220 105.570 129.390 106.410 ;
        RECT 117.090 105.260 121.970 105.430 ;
        RECT 124.090 105.260 128.970 105.430 ;
        RECT 117.090 104.550 121.970 104.720 ;
        RECT 124.090 104.550 128.970 104.720 ;
        RECT 116.670 103.570 116.840 104.410 ;
        RECT 122.220 103.570 122.390 104.410 ;
        RECT 123.670 103.570 123.840 104.410 ;
        RECT 129.220 103.570 129.390 104.410 ;
        RECT 117.090 103.260 121.970 103.430 ;
        RECT 124.090 103.260 128.970 103.430 ;
        RECT 117.090 100.550 121.970 100.720 ;
        RECT 124.090 100.550 128.970 100.720 ;
        RECT 116.670 99.570 116.840 100.410 ;
        RECT 122.220 99.570 122.390 100.410 ;
        RECT 123.670 99.570 123.840 100.410 ;
        RECT 129.220 99.570 129.390 100.410 ;
        RECT 117.090 99.260 121.970 99.430 ;
        RECT 124.090 99.260 128.970 99.430 ;
        RECT 117.090 98.550 121.970 98.720 ;
        RECT 124.090 98.550 128.970 98.720 ;
        RECT 116.670 97.570 116.840 98.410 ;
        RECT 122.220 97.570 122.390 98.410 ;
        RECT 123.670 97.570 123.840 98.410 ;
        RECT 129.220 97.570 129.390 98.410 ;
        RECT 117.090 97.260 121.970 97.430 ;
        RECT 124.090 97.260 128.970 97.430 ;
        RECT 132.810 107.530 137.690 107.700 ;
        RECT 141.810 107.530 146.690 107.700 ;
        RECT 132.345 107.050 132.515 107.390 ;
        RECT 137.985 107.050 138.155 107.390 ;
        RECT 141.345 107.050 141.515 107.390 ;
        RECT 146.985 107.050 147.155 107.390 ;
        RECT 132.810 106.740 137.690 106.910 ;
        RECT 141.810 106.740 146.690 106.910 ;
        RECT 132.810 103.030 137.690 103.200 ;
        RECT 141.810 103.030 146.690 103.200 ;
        RECT 132.345 102.550 132.515 102.890 ;
        RECT 137.985 102.550 138.155 102.890 ;
        RECT 141.345 102.550 141.515 102.890 ;
        RECT 146.985 102.550 147.155 102.890 ;
        RECT 132.810 102.240 137.690 102.410 ;
        RECT 141.810 102.240 146.690 102.410 ;
        RECT 132.810 98.530 137.690 98.700 ;
        RECT 141.810 98.530 146.690 98.700 ;
        RECT 132.345 98.050 132.515 98.390 ;
        RECT 137.985 98.050 138.155 98.390 ;
        RECT 141.345 98.050 141.515 98.390 ;
        RECT 146.985 98.050 147.155 98.390 ;
        RECT 132.810 97.740 137.690 97.910 ;
        RECT 141.810 97.740 146.690 97.910 ;
        RECT 147.520 96.240 147.700 107.910 ;
        RECT 138.410 95.500 139.470 95.680 ;
        RECT 105.550 94.030 105.720 94.470 ;
        RECT 106.510 94.710 107.150 94.880 ;
        RECT 108.160 94.710 108.800 94.880 ;
        RECT 109.560 94.710 110.200 94.880 ;
        RECT 110.740 94.710 111.380 94.880 ;
        RECT 106.030 92.760 106.200 94.400 ;
        RECT 106.960 94.135 111.840 94.305 ;
        RECT 106.540 93.155 106.710 93.995 ;
        RECT 112.090 93.155 112.260 93.995 ;
        RECT 106.960 92.845 111.840 93.015 ;
        RECT 102.940 92.430 103.780 92.600 ;
        RECT 104.230 92.430 105.070 92.600 ;
        RECT 102.630 91.300 102.800 92.180 ;
        RECT 103.920 91.300 104.090 92.180 ;
        RECT 105.210 91.300 105.380 92.180 ;
        RECT 102.940 90.880 103.780 91.050 ;
        RECT 104.230 90.880 105.070 91.050 ;
        RECT 123.660 94.710 124.230 94.880 ;
        RECT 114.105 94.140 114.985 94.310 ;
        RECT 113.640 93.660 113.810 94.000 ;
        RECT 115.280 93.660 115.450 94.000 ;
        RECT 114.105 93.350 114.985 93.520 ;
        RECT 116.765 94.140 124.145 94.310 ;
        RECT 116.300 93.660 116.470 94.000 ;
        RECT 124.440 93.660 124.610 94.000 ;
        RECT 116.765 93.350 124.145 93.520 ;
        RECT 124.950 93.260 125.120 94.400 ;
        RECT 117.020 92.780 121.970 92.950 ;
        RECT 122.800 92.780 123.940 92.950 ;
        RECT 117.020 92.340 121.970 92.510 ;
        RECT 105.550 89.970 105.720 90.410 ;
        RECT 116.770 91.765 123.650 91.935 ;
        RECT 116.305 91.285 116.475 91.625 ;
        RECT 123.945 91.285 124.115 91.625 ;
        RECT 116.770 90.975 123.650 91.145 ;
        RECT 124.450 90.890 124.620 92.030 ;
        RECT 116.770 89.835 123.650 90.005 ;
        RECT 116.305 89.355 116.475 89.695 ;
        RECT 123.945 89.355 124.115 89.695 ;
        RECT 116.770 89.045 123.650 89.215 ;
        RECT 124.450 88.960 124.620 90.100 ;
        RECT 102.940 88.370 103.780 88.540 ;
        RECT 104.230 88.370 105.070 88.540 ;
        RECT 102.630 87.240 102.800 88.120 ;
        RECT 103.920 87.240 104.090 88.120 ;
        RECT 105.210 87.240 105.380 88.120 ;
        RECT 102.940 86.820 103.780 86.990 ;
        RECT 104.230 86.820 105.070 86.990 ;
        RECT 105.550 85.910 105.720 86.350 ;
        RECT 107.160 86.920 112.040 87.090 ;
        RECT 106.140 84.980 106.310 86.450 ;
        RECT 106.740 86.440 106.910 86.780 ;
        RECT 112.290 86.440 112.460 86.780 ;
        RECT 107.160 86.130 112.040 86.300 ;
        RECT 106.740 85.650 106.910 85.990 ;
        RECT 112.290 85.650 112.460 85.990 ;
        RECT 107.160 85.340 112.040 85.510 ;
        RECT 102.940 84.310 103.780 84.480 ;
        RECT 104.230 84.310 105.070 84.480 ;
        RECT 102.630 83.180 102.800 84.060 ;
        RECT 103.920 83.180 104.090 84.060 ;
        RECT 105.210 83.180 105.380 84.060 ;
        RECT 102.940 82.760 103.780 82.930 ;
        RECT 104.230 82.760 105.070 82.930 ;
        RECT 105.550 81.850 105.720 82.290 ;
        RECT 106.740 84.860 106.910 85.200 ;
        RECT 112.290 84.860 112.460 85.200 ;
        RECT 107.160 84.550 112.040 84.720 ;
        RECT 106.740 84.070 106.910 84.410 ;
        RECT 112.290 84.070 112.460 84.410 ;
        RECT 107.160 83.760 112.040 83.930 ;
        RECT 106.140 82.150 106.310 83.620 ;
        RECT 106.740 83.280 106.910 83.620 ;
        RECT 112.290 83.280 112.460 83.620 ;
        RECT 107.160 82.970 112.040 83.140 ;
        RECT 106.740 82.490 106.910 82.830 ;
        RECT 112.290 82.490 112.460 82.830 ;
        RECT 107.160 82.180 112.040 82.350 ;
        RECT 106.740 81.700 106.910 82.040 ;
        RECT 112.290 81.700 112.460 82.040 ;
        RECT 107.160 81.390 112.040 81.560 ;
        RECT 102.940 80.250 103.780 80.420 ;
        RECT 104.230 80.250 105.070 80.420 ;
        RECT 102.630 79.120 102.800 80.000 ;
        RECT 103.920 79.120 104.090 80.000 ;
        RECT 105.210 79.120 105.380 80.000 ;
        RECT 102.940 78.700 103.780 78.870 ;
        RECT 104.230 78.700 105.070 78.870 ;
        RECT 105.550 77.790 105.720 78.230 ;
        RECT 106.140 79.800 106.310 81.270 ;
        RECT 106.740 80.910 106.910 81.250 ;
        RECT 112.290 80.910 112.460 81.250 ;
        RECT 107.160 80.600 112.040 80.770 ;
        RECT 106.740 80.120 106.910 80.460 ;
        RECT 112.290 80.120 112.460 80.460 ;
        RECT 107.160 79.810 112.040 79.980 ;
        RECT 106.740 79.330 106.910 79.670 ;
        RECT 112.290 79.330 112.460 79.670 ;
        RECT 107.160 79.020 112.040 79.190 ;
        RECT 106.140 77.280 106.310 78.750 ;
        RECT 106.740 78.540 106.910 78.880 ;
        RECT 112.290 78.540 112.460 78.880 ;
        RECT 107.160 78.230 112.040 78.400 ;
        RECT 106.740 77.750 106.910 78.090 ;
        RECT 112.290 77.750 112.460 78.090 ;
        RECT 107.160 77.440 112.040 77.610 ;
        RECT 102.940 76.190 103.780 76.360 ;
        RECT 104.230 76.190 105.070 76.360 ;
        RECT 102.630 75.060 102.800 75.940 ;
        RECT 103.920 75.060 104.090 75.940 ;
        RECT 105.210 75.060 105.380 75.940 ;
        RECT 102.940 74.640 103.780 74.810 ;
        RECT 104.230 74.640 105.070 74.810 ;
        RECT 105.550 73.730 105.720 74.170 ;
        RECT 106.740 76.960 106.910 77.300 ;
        RECT 112.290 76.960 112.460 77.300 ;
        RECT 107.160 76.650 112.040 76.820 ;
        RECT 106.140 74.700 106.310 76.170 ;
        RECT 106.740 76.170 106.910 76.510 ;
        RECT 112.290 76.170 112.460 76.510 ;
        RECT 107.160 75.860 112.040 76.030 ;
        RECT 106.740 75.380 106.910 75.720 ;
        RECT 112.290 75.380 112.460 75.720 ;
        RECT 107.160 75.070 112.040 75.240 ;
        RECT 106.740 74.590 106.910 74.930 ;
        RECT 112.290 74.590 112.460 74.930 ;
        RECT 107.160 74.280 112.040 74.450 ;
        RECT 106.740 73.800 106.910 74.140 ;
        RECT 112.290 73.800 112.460 74.140 ;
        RECT 102.940 72.130 103.780 72.300 ;
        RECT 104.230 72.130 105.070 72.300 ;
        RECT 102.630 71.000 102.800 71.880 ;
        RECT 103.920 71.000 104.090 71.880 ;
        RECT 105.210 71.000 105.380 71.880 ;
        RECT 102.940 70.580 103.780 70.750 ;
        RECT 104.230 70.580 105.070 70.750 ;
        RECT 106.140 72.130 106.310 73.600 ;
        RECT 107.160 73.490 112.040 73.660 ;
        RECT 106.740 73.010 106.910 73.350 ;
        RECT 112.290 73.010 112.460 73.350 ;
        RECT 107.160 72.700 112.040 72.870 ;
        RECT 106.740 72.220 106.910 72.560 ;
        RECT 112.290 72.220 112.460 72.560 ;
        RECT 107.160 71.910 112.040 72.080 ;
        RECT 115.220 86.740 120.100 86.910 ;
        RECT 114.755 86.260 114.925 86.600 ;
        RECT 120.395 86.260 120.565 86.600 ;
        RECT 115.220 85.950 120.100 86.120 ;
        RECT 114.755 85.470 114.925 85.810 ;
        RECT 120.395 85.470 120.565 85.810 ;
        RECT 115.220 85.160 120.100 85.330 ;
        RECT 120.860 85.250 121.030 86.390 ;
        RECT 114.755 84.680 114.925 85.020 ;
        RECT 120.395 84.680 120.565 85.020 ;
        RECT 115.220 84.370 120.100 84.540 ;
        RECT 114.755 83.890 114.925 84.230 ;
        RECT 120.395 83.890 120.565 84.230 ;
        RECT 115.220 83.580 120.100 83.750 ;
        RECT 114.755 83.100 114.925 83.440 ;
        RECT 120.395 83.100 120.565 83.440 ;
        RECT 120.860 83.010 121.030 84.150 ;
        RECT 115.220 82.790 120.100 82.960 ;
        RECT 114.755 82.310 114.925 82.650 ;
        RECT 120.395 82.310 120.565 82.650 ;
        RECT 115.220 82.000 120.100 82.170 ;
        RECT 114.755 81.520 114.925 81.860 ;
        RECT 120.395 81.520 120.565 81.860 ;
        RECT 115.220 81.210 120.100 81.380 ;
        RECT 114.755 80.730 114.925 81.070 ;
        RECT 120.395 80.730 120.565 81.070 ;
        RECT 120.860 80.710 121.030 81.850 ;
        RECT 115.220 80.420 120.100 80.590 ;
        RECT 114.755 79.940 114.925 80.280 ;
        RECT 120.395 79.940 120.565 80.280 ;
        RECT 115.220 79.630 120.100 79.800 ;
        RECT 114.755 79.150 114.925 79.490 ;
        RECT 120.395 79.150 120.565 79.490 ;
        RECT 115.220 78.840 120.100 79.010 ;
        RECT 114.755 78.360 114.925 78.700 ;
        RECT 120.395 78.360 120.565 78.700 ;
        RECT 120.860 78.270 121.030 79.410 ;
        RECT 115.220 78.050 120.100 78.220 ;
        RECT 114.755 77.570 114.925 77.910 ;
        RECT 120.395 77.570 120.565 77.910 ;
        RECT 115.220 77.260 120.100 77.430 ;
        RECT 114.755 76.780 114.925 77.120 ;
        RECT 120.395 76.780 120.565 77.120 ;
        RECT 115.220 76.470 120.100 76.640 ;
        RECT 114.755 75.990 114.925 76.330 ;
        RECT 120.395 75.990 120.565 76.330 ;
        RECT 120.860 75.870 121.030 77.010 ;
        RECT 115.220 75.680 120.100 75.850 ;
        RECT 105.550 69.670 105.720 70.110 ;
        RECT 102.940 68.070 103.780 68.240 ;
        RECT 104.230 68.070 105.070 68.240 ;
        RECT 102.630 66.940 102.800 67.820 ;
        RECT 103.920 66.940 104.090 67.820 ;
        RECT 105.210 66.940 105.380 67.820 ;
        RECT 102.940 66.520 103.780 66.690 ;
        RECT 104.230 66.520 105.070 66.690 ;
        RECT 105.550 65.610 105.720 66.050 ;
        RECT 102.940 64.010 103.780 64.180 ;
        RECT 104.230 64.010 105.070 64.180 ;
        RECT 102.630 62.880 102.800 63.760 ;
        RECT 103.920 62.880 104.090 63.760 ;
        RECT 105.210 62.880 105.380 63.760 ;
        RECT 102.940 62.460 103.780 62.630 ;
        RECT 104.230 62.460 105.070 62.630 ;
        RECT 105.550 61.550 105.720 61.990 ;
        RECT 94.320 56.585 95.160 56.755 ;
        RECT 95.610 56.585 96.450 56.755 ;
        RECT 94.010 54.410 94.180 56.290 ;
        RECT 95.300 54.410 95.470 56.290 ;
        RECT 96.590 54.410 96.760 56.290 ;
        RECT 94.320 53.945 95.160 54.115 ;
        RECT 95.610 53.945 96.450 54.115 ;
        RECT 97.250 53.610 97.430 57.280 ;
        RECT 97.770 56.970 97.950 60.640 ;
        RECT 98.750 59.945 99.590 60.115 ;
        RECT 100.040 59.945 100.880 60.115 ;
        RECT 98.440 57.770 98.610 59.650 ;
        RECT 99.730 57.770 99.900 59.650 ;
        RECT 101.020 57.770 101.190 59.650 ;
        RECT 98.750 57.305 99.590 57.475 ;
        RECT 100.040 57.305 100.880 57.475 ;
        RECT 102.940 59.470 103.780 59.640 ;
        RECT 104.230 59.470 105.070 59.640 ;
        RECT 102.630 58.340 102.800 59.220 ;
        RECT 103.920 58.340 104.090 59.220 ;
        RECT 105.210 58.340 105.380 59.220 ;
        RECT 102.940 57.920 103.780 58.090 ;
        RECT 104.230 57.920 105.070 58.090 ;
        RECT 105.550 57.010 105.720 57.450 ;
        RECT 94.320 52.535 95.160 52.705 ;
        RECT 95.610 52.535 96.450 52.705 ;
        RECT 94.010 50.360 94.180 52.240 ;
        RECT 95.300 50.360 95.470 52.240 ;
        RECT 96.590 50.360 96.760 52.240 ;
        RECT 94.320 49.895 95.160 50.065 ;
        RECT 95.610 49.895 96.450 50.065 ;
        RECT 97.250 49.560 97.430 53.230 ;
        RECT 94.320 48.485 95.160 48.655 ;
        RECT 95.610 48.485 96.450 48.655 ;
        RECT 94.010 46.310 94.180 48.190 ;
        RECT 95.300 46.310 95.470 48.190 ;
        RECT 96.590 46.310 96.760 48.190 ;
        RECT 94.320 45.845 95.160 46.015 ;
        RECT 95.610 45.845 96.450 46.015 ;
        RECT 97.250 45.510 97.430 49.180 ;
        RECT 94.320 44.435 95.160 44.605 ;
        RECT 95.610 44.435 96.450 44.605 ;
        RECT 94.010 42.260 94.180 44.140 ;
        RECT 95.300 42.260 95.470 44.140 ;
        RECT 96.590 42.260 96.760 44.140 ;
        RECT 94.320 41.795 95.160 41.965 ;
        RECT 95.610 41.795 96.450 41.965 ;
        RECT 97.250 41.460 97.430 45.130 ;
        RECT 94.320 40.385 95.160 40.555 ;
        RECT 95.610 40.385 96.450 40.555 ;
        RECT 94.010 38.210 94.180 40.090 ;
        RECT 95.300 38.210 95.470 40.090 ;
        RECT 96.590 38.210 96.760 40.090 ;
        RECT 94.320 37.745 95.160 37.915 ;
        RECT 95.610 37.745 96.450 37.915 ;
        RECT 97.250 37.410 97.430 41.080 ;
        RECT 94.320 36.335 95.160 36.505 ;
        RECT 95.610 36.335 96.450 36.505 ;
        RECT 94.010 34.160 94.180 36.040 ;
        RECT 95.300 34.160 95.470 36.040 ;
        RECT 96.590 34.160 96.760 36.040 ;
        RECT 94.320 33.695 95.160 33.865 ;
        RECT 95.610 33.695 96.450 33.865 ;
        RECT 97.250 33.360 97.430 37.030 ;
        RECT 94.320 32.285 95.160 32.455 ;
        RECT 95.610 32.285 96.450 32.455 ;
        RECT 94.010 30.110 94.180 31.990 ;
        RECT 95.300 30.110 95.470 31.990 ;
        RECT 96.590 30.110 96.760 31.990 ;
        RECT 94.320 29.645 95.160 29.815 ;
        RECT 95.610 29.645 96.450 29.815 ;
        RECT 97.250 29.310 97.430 32.980 ;
        RECT 94.320 28.200 95.160 28.370 ;
        RECT 95.610 28.200 96.450 28.370 ;
        RECT 94.010 26.025 94.180 27.905 ;
        RECT 95.300 26.025 95.470 27.905 ;
        RECT 96.590 26.025 96.760 27.905 ;
        RECT 94.320 25.560 95.160 25.730 ;
        RECT 95.610 25.560 96.450 25.730 ;
        RECT 97.250 25.225 97.430 28.895 ;
        RECT 94.320 24.075 95.160 24.245 ;
        RECT 95.610 24.075 96.450 24.245 ;
        RECT 94.010 21.900 94.180 23.780 ;
        RECT 95.300 21.900 95.470 23.780 ;
        RECT 96.590 21.900 96.760 23.780 ;
        RECT 94.320 21.435 95.160 21.605 ;
        RECT 95.610 21.435 96.450 21.605 ;
        RECT 97.250 21.100 97.430 24.770 ;
        RECT 90.130 19.045 90.970 19.215 ;
        RECT 91.420 19.045 92.260 19.215 ;
        RECT 89.820 17.915 89.990 18.795 ;
        RECT 91.110 17.915 91.280 18.795 ;
        RECT 92.400 17.915 92.570 18.795 ;
        RECT 90.130 17.495 90.970 17.665 ;
        RECT 91.420 17.495 92.260 17.665 ;
        RECT 89.480 16.585 89.650 17.025 ;
        RECT 94.320 19.520 95.160 19.690 ;
        RECT 95.610 19.520 96.450 19.690 ;
        RECT 94.010 17.345 94.180 19.225 ;
        RECT 95.300 17.345 95.470 19.225 ;
        RECT 96.590 17.345 96.760 19.225 ;
        RECT 94.320 16.880 95.160 17.050 ;
        RECT 95.610 16.880 96.450 17.050 ;
        RECT 97.250 16.545 97.430 20.215 ;
      LAYER met1 ;
        RECT 89.360 155.700 89.930 155.800 ;
        RECT 89.360 155.620 130.350 155.700 ;
        RECT 89.360 155.450 130.800 155.620 ;
        RECT 89.360 155.300 130.350 155.450 ;
        RECT 89.360 155.060 89.930 155.300 ;
        RECT 90.470 155.080 130.350 155.300 ;
        RECT 89.360 151.550 89.810 155.060 ;
        RECT 90.410 154.850 130.410 155.080 ;
        RECT 90.020 154.740 90.250 154.800 ;
        RECT 90.020 154.680 90.260 154.740 ;
        RECT 90.020 153.840 90.430 154.680 ;
        RECT 90.040 153.790 90.430 153.840 ;
        RECT 130.570 153.790 130.800 154.800 ;
        RECT 90.040 153.560 130.800 153.790 ;
        RECT 90.040 151.750 92.350 153.560 ;
        RECT 90.200 151.730 92.305 151.750 ;
        RECT 89.360 146.860 89.930 151.550 ;
        RECT 96.530 150.210 99.090 150.790 ;
        RECT 104.270 150.210 107.140 152.670 ;
        RECT 96.530 149.635 107.740 150.210 ;
        RECT 96.530 148.985 108.805 149.635 ;
        RECT 96.530 148.410 107.740 148.985 ;
        RECT 96.530 147.980 99.090 148.410 ;
        RECT 87.680 145.770 89.930 146.860 ;
        RECT 92.810 145.860 93.500 146.640 ;
        RECT 94.260 145.860 95.220 145.885 ;
        RECT 87.680 145.020 89.910 145.770 ;
        RECT 91.420 145.690 95.220 145.860 ;
        RECT 91.420 145.410 92.260 145.690 ;
        RECT 94.260 145.655 95.220 145.690 ;
        RECT 95.550 145.655 96.510 145.885 ;
        RECT 92.470 145.450 94.190 145.470 ;
        RECT 90.070 145.180 91.030 145.410 ;
        RECT 91.360 145.180 92.320 145.410 ;
        RECT 87.680 144.020 90.020 145.020 ;
        RECT 87.680 143.490 89.910 144.020 ;
        RECT 90.290 143.860 90.810 145.180 ;
        RECT 91.080 144.020 91.310 145.020 ;
        RECT 91.560 143.860 92.080 145.180 ;
        RECT 92.470 145.020 94.210 145.450 ;
        RECT 92.370 144.020 94.210 145.020 ;
        RECT 90.070 143.630 91.030 143.860 ;
        RECT 91.360 143.630 92.320 143.860 ;
        RECT 87.680 143.370 89.920 143.490 ;
        RECT 92.470 143.450 94.210 144.020 ;
        RECT 92.470 143.430 94.190 143.450 ;
        RECT 87.680 143.020 89.930 143.370 ;
        RECT 89.370 142.230 89.930 143.020 ;
        RECT 92.810 143.020 93.500 143.430 ;
        RECT 94.490 143.245 95.010 145.655 ;
        RECT 95.270 143.450 95.500 145.450 ;
        RECT 95.820 143.245 96.340 145.655 ;
        RECT 96.700 145.450 98.500 147.980 ;
        RECT 98.690 145.655 99.650 145.885 ;
        RECT 99.980 145.860 100.940 145.885 ;
        RECT 101.700 145.860 102.390 146.640 ;
        RECT 105.290 146.400 105.830 146.860 ;
        RECT 108.155 146.665 108.805 148.985 ;
        RECT 138.220 146.685 139.170 146.730 ;
        RECT 134.855 146.670 139.170 146.685 ;
        RECT 118.350 146.665 139.170 146.670 ;
        RECT 99.980 145.690 103.780 145.860 ;
        RECT 99.980 145.655 100.940 145.690 ;
        RECT 96.560 143.450 98.640 145.450 ;
        RECT 92.810 142.400 93.510 143.020 ;
        RECT 94.260 143.015 95.220 143.245 ;
        RECT 95.550 143.015 96.510 143.245 ;
        RECT 89.370 141.020 89.910 142.230 ;
        RECT 92.810 141.860 93.500 142.400 ;
        RECT 94.260 141.860 95.220 141.885 ;
        RECT 91.420 141.690 95.220 141.860 ;
        RECT 91.420 141.410 92.260 141.690 ;
        RECT 94.260 141.655 95.220 141.690 ;
        RECT 95.550 141.655 96.510 141.885 ;
        RECT 92.470 141.450 94.190 141.470 ;
        RECT 90.070 141.180 91.030 141.410 ;
        RECT 91.360 141.180 92.320 141.410 ;
        RECT 89.370 140.020 90.020 141.020 ;
        RECT 89.370 139.490 89.910 140.020 ;
        RECT 90.290 139.860 90.810 141.180 ;
        RECT 91.080 140.020 91.310 141.020 ;
        RECT 91.560 139.860 92.080 141.180 ;
        RECT 92.470 141.020 94.210 141.450 ;
        RECT 92.370 140.020 94.210 141.020 ;
        RECT 90.070 139.630 91.030 139.860 ;
        RECT 91.360 139.630 92.320 139.860 ;
        RECT 89.370 139.370 89.920 139.490 ;
        RECT 92.470 139.450 94.210 140.020 ;
        RECT 92.470 139.430 94.190 139.450 ;
        RECT 89.370 138.230 89.930 139.370 ;
        RECT 92.810 139.020 93.500 139.430 ;
        RECT 94.490 139.245 95.010 141.655 ;
        RECT 95.270 139.450 95.500 141.450 ;
        RECT 95.820 139.245 96.340 141.655 ;
        RECT 96.700 141.450 98.500 143.450 ;
        RECT 98.860 143.245 99.380 145.655 ;
        RECT 99.700 143.450 99.930 145.450 ;
        RECT 100.190 143.245 100.710 145.655 ;
        RECT 101.010 145.450 102.730 145.470 ;
        RECT 100.990 145.020 102.730 145.450 ;
        RECT 102.940 145.410 103.780 145.690 ;
        RECT 105.290 145.830 106.460 146.400 ;
        RECT 108.155 146.170 139.170 146.665 ;
        RECT 108.155 146.165 108.805 146.170 ;
        RECT 134.855 146.155 139.170 146.170 ;
        RECT 138.220 146.110 139.170 146.155 ;
        RECT 102.880 145.180 103.840 145.410 ;
        RECT 104.170 145.180 105.130 145.410 ;
        RECT 100.990 144.020 102.830 145.020 ;
        RECT 100.990 143.450 102.730 144.020 ;
        RECT 103.120 143.860 103.640 145.180 ;
        RECT 103.890 144.020 104.120 145.020 ;
        RECT 104.390 143.860 104.910 145.180 ;
        RECT 105.290 145.020 115.760 145.830 ;
        RECT 136.890 145.650 137.610 145.850 ;
        RECT 132.750 145.420 137.750 145.650 ;
        RECT 105.180 144.970 115.760 145.020 ;
        RECT 105.180 144.020 106.460 144.970 ;
        RECT 102.880 143.630 103.840 143.860 ;
        RECT 104.170 143.630 105.130 143.860 ;
        RECT 105.290 143.490 106.460 144.020 ;
        RECT 107.250 144.110 108.400 144.780 ;
        RECT 112.650 144.390 113.570 144.460 ;
        RECT 108.550 144.160 113.570 144.390 ;
        RECT 107.250 143.600 108.410 144.110 ;
        RECT 112.650 144.040 113.570 144.160 ;
        RECT 101.010 143.430 102.730 143.450 ;
        RECT 98.690 143.015 99.650 143.245 ;
        RECT 99.980 143.015 100.940 143.245 ;
        RECT 101.700 143.020 102.390 143.430 ;
        RECT 105.280 143.370 106.460 143.490 ;
        RECT 101.690 142.400 102.390 143.020 ;
        RECT 98.690 141.595 99.650 141.825 ;
        RECT 99.980 141.800 100.940 141.825 ;
        RECT 101.700 141.800 102.390 142.400 ;
        RECT 105.270 143.300 106.460 143.370 ;
        RECT 105.270 142.640 106.630 143.300 ;
        RECT 107.990 143.150 108.410 143.600 ;
        RECT 107.990 142.820 108.380 143.150 ;
        RECT 108.550 143.100 109.650 143.300 ;
        RECT 108.550 142.870 113.570 143.100 ;
        RECT 105.270 142.230 106.460 142.640 ;
        RECT 105.280 141.800 106.460 142.230 ;
        RECT 99.980 141.630 103.780 141.800 ;
        RECT 99.980 141.595 100.940 141.630 ;
        RECT 96.560 141.390 98.500 141.450 ;
        RECT 96.560 139.450 98.640 141.390 ;
        RECT 96.700 139.390 98.640 139.450 ;
        RECT 92.810 138.400 93.510 139.020 ;
        RECT 94.260 139.015 95.220 139.245 ;
        RECT 95.550 139.015 96.510 139.245 ;
        RECT 89.370 136.920 89.910 138.230 ;
        RECT 92.810 137.760 93.500 138.400 ;
        RECT 94.260 137.760 95.220 137.785 ;
        RECT 91.420 137.590 95.220 137.760 ;
        RECT 91.420 137.310 92.260 137.590 ;
        RECT 94.260 137.555 95.220 137.590 ;
        RECT 95.550 137.555 96.510 137.785 ;
        RECT 92.470 137.350 94.190 137.370 ;
        RECT 90.070 137.080 91.030 137.310 ;
        RECT 91.360 137.080 92.320 137.310 ;
        RECT 89.370 135.920 90.020 136.920 ;
        RECT 89.370 135.390 89.910 135.920 ;
        RECT 90.290 135.760 90.810 137.080 ;
        RECT 91.080 135.920 91.310 136.920 ;
        RECT 91.560 135.760 92.080 137.080 ;
        RECT 92.470 136.920 94.210 137.350 ;
        RECT 92.370 135.920 94.210 136.920 ;
        RECT 90.070 135.530 91.030 135.760 ;
        RECT 91.360 135.530 92.320 135.760 ;
        RECT 89.370 135.270 89.920 135.390 ;
        RECT 92.470 135.350 94.210 135.920 ;
        RECT 92.470 135.330 94.190 135.350 ;
        RECT 89.370 134.130 89.930 135.270 ;
        RECT 92.810 134.920 93.500 135.330 ;
        RECT 94.490 135.145 95.010 137.555 ;
        RECT 95.270 135.350 95.500 137.350 ;
        RECT 95.820 135.145 96.340 137.555 ;
        RECT 96.700 137.350 98.500 139.390 ;
        RECT 98.860 139.185 99.380 141.595 ;
        RECT 99.700 139.390 99.930 141.390 ;
        RECT 100.190 139.185 100.710 141.595 ;
        RECT 101.010 141.390 102.730 141.410 ;
        RECT 100.990 140.960 102.730 141.390 ;
        RECT 102.940 141.350 103.780 141.630 ;
        RECT 102.880 141.120 103.840 141.350 ;
        RECT 104.170 141.120 105.130 141.350 ;
        RECT 100.990 139.960 102.830 140.960 ;
        RECT 100.990 139.390 102.730 139.960 ;
        RECT 103.120 139.800 103.640 141.120 ;
        RECT 103.890 139.960 104.120 140.960 ;
        RECT 104.390 139.800 104.910 141.120 ;
        RECT 105.290 140.960 106.460 141.800 ;
        RECT 105.180 139.960 106.460 140.960 ;
        RECT 102.880 139.570 103.840 139.800 ;
        RECT 104.170 139.570 105.130 139.800 ;
        RECT 105.290 139.430 106.460 139.960 ;
        RECT 101.010 139.370 102.730 139.390 ;
        RECT 98.690 138.955 99.650 139.185 ;
        RECT 99.980 138.955 100.940 139.185 ;
        RECT 101.700 138.960 102.390 139.370 ;
        RECT 105.280 139.310 106.460 139.430 ;
        RECT 101.690 138.340 102.390 138.960 ;
        RECT 98.690 137.535 99.650 137.765 ;
        RECT 99.980 137.740 100.940 137.765 ;
        RECT 101.700 137.740 102.390 138.340 ;
        RECT 105.270 138.170 106.460 139.310 ;
        RECT 99.980 137.570 103.780 137.740 ;
        RECT 99.980 137.535 100.940 137.570 ;
        RECT 96.560 137.330 98.500 137.350 ;
        RECT 96.560 135.350 98.640 137.330 ;
        RECT 96.700 135.330 98.640 135.350 ;
        RECT 92.810 134.300 93.510 134.920 ;
        RECT 94.260 134.915 95.220 135.145 ;
        RECT 95.550 134.915 96.510 135.145 ;
        RECT 89.370 132.870 89.910 134.130 ;
        RECT 92.810 133.710 93.500 134.300 ;
        RECT 94.260 133.710 95.220 133.735 ;
        RECT 91.420 133.540 95.220 133.710 ;
        RECT 91.420 133.260 92.260 133.540 ;
        RECT 94.260 133.505 95.220 133.540 ;
        RECT 95.550 133.505 96.510 133.735 ;
        RECT 92.470 133.300 94.190 133.320 ;
        RECT 90.070 133.030 91.030 133.260 ;
        RECT 91.360 133.030 92.320 133.260 ;
        RECT 89.370 131.870 90.020 132.870 ;
        RECT 89.370 131.340 89.910 131.870 ;
        RECT 90.290 131.710 90.810 133.030 ;
        RECT 91.080 131.870 91.310 132.870 ;
        RECT 91.560 131.710 92.080 133.030 ;
        RECT 92.470 132.870 94.210 133.300 ;
        RECT 92.370 131.870 94.210 132.870 ;
        RECT 90.070 131.480 91.030 131.710 ;
        RECT 91.360 131.480 92.320 131.710 ;
        RECT 89.370 131.220 89.920 131.340 ;
        RECT 92.470 131.300 94.210 131.870 ;
        RECT 92.470 131.280 94.190 131.300 ;
        RECT 89.370 130.080 89.930 131.220 ;
        RECT 92.810 130.870 93.500 131.280 ;
        RECT 94.490 131.095 95.010 133.505 ;
        RECT 95.270 131.300 95.500 133.300 ;
        RECT 95.820 131.095 96.340 133.505 ;
        RECT 96.700 133.300 98.500 135.330 ;
        RECT 98.860 135.125 99.380 137.535 ;
        RECT 99.700 135.330 99.930 137.330 ;
        RECT 100.190 135.125 100.710 137.535 ;
        RECT 101.010 137.330 102.730 137.350 ;
        RECT 100.990 136.900 102.730 137.330 ;
        RECT 102.940 137.290 103.780 137.570 ;
        RECT 102.880 137.060 103.840 137.290 ;
        RECT 104.170 137.060 105.130 137.290 ;
        RECT 100.990 135.900 102.830 136.900 ;
        RECT 100.990 135.330 102.730 135.900 ;
        RECT 103.120 135.740 103.640 137.060 ;
        RECT 103.890 135.900 104.120 136.900 ;
        RECT 104.390 135.740 104.910 137.060 ;
        RECT 105.290 136.900 106.460 138.170 ;
        RECT 105.180 135.900 106.460 136.900 ;
        RECT 102.880 135.510 103.840 135.740 ;
        RECT 104.170 135.510 105.130 135.740 ;
        RECT 105.290 135.370 106.460 135.900 ;
        RECT 101.010 135.310 102.730 135.330 ;
        RECT 98.690 134.895 99.650 135.125 ;
        RECT 99.980 134.895 100.940 135.125 ;
        RECT 101.700 134.900 102.390 135.310 ;
        RECT 105.280 135.250 106.460 135.370 ;
        RECT 101.690 134.280 102.390 134.900 ;
        RECT 98.690 133.475 99.650 133.705 ;
        RECT 99.980 133.680 100.940 133.705 ;
        RECT 101.700 133.680 102.390 134.280 ;
        RECT 105.270 134.110 106.460 135.250 ;
        RECT 107.990 141.860 108.410 142.820 ;
        RECT 108.550 142.630 109.650 142.870 ;
        RECT 107.990 141.530 108.380 141.860 ;
        RECT 112.650 141.810 113.570 141.880 ;
        RECT 108.560 141.580 113.570 141.810 ;
        RECT 107.990 140.570 108.410 141.530 ;
        RECT 112.650 141.460 113.570 141.580 ;
        RECT 107.990 140.240 108.380 140.570 ;
        RECT 108.630 140.530 109.570 140.600 ;
        RECT 108.560 140.520 113.520 140.530 ;
        RECT 108.560 140.300 113.570 140.520 ;
        RECT 108.570 140.290 113.570 140.300 ;
        RECT 107.990 139.980 108.410 140.240 ;
        RECT 108.630 140.210 109.570 140.290 ;
        RECT 113.730 139.980 114.010 144.130 ;
        RECT 115.180 143.320 115.760 144.970 ;
        RECT 120.080 144.670 121.600 144.770 ;
        RECT 127.280 144.670 129.000 144.810 ;
        RECT 117.030 144.440 122.030 144.670 ;
        RECT 124.030 144.440 129.030 144.670 ;
        RECT 116.640 143.430 116.870 144.390 ;
        RECT 120.080 144.250 121.600 144.440 ;
        RECT 122.220 144.390 123.080 144.400 ;
        RECT 127.280 144.390 129.000 144.440 ;
        RECT 129.280 144.390 130.870 144.420 ;
        RECT 122.190 143.430 123.090 144.390 ;
        RECT 123.640 143.430 123.870 144.390 ;
        RECT 129.190 143.430 130.870 144.390 ;
        RECT 122.200 143.410 123.090 143.430 ;
        RECT 129.210 143.410 130.870 143.430 ;
        RECT 122.220 143.390 123.090 143.410 ;
        RECT 117.030 143.350 122.030 143.380 ;
        RECT 117.010 142.650 122.060 143.350 ;
        RECT 117.010 142.460 122.050 142.650 ;
        RECT 117.030 142.440 122.030 142.460 ;
        RECT 116.640 141.430 116.870 142.390 ;
        RECT 117.990 141.380 119.510 141.470 ;
        RECT 117.030 141.150 122.030 141.380 ;
        RECT 117.990 140.950 119.510 141.150 ;
        RECT 107.990 139.530 108.460 139.980 ;
        RECT 113.640 139.530 114.010 139.980 ;
        RECT 107.990 139.280 108.410 139.530 ;
        RECT 107.990 138.950 108.380 139.280 ;
        RECT 112.640 139.230 113.570 139.290 ;
        RECT 108.560 139.000 113.570 139.230 ;
        RECT 107.990 137.990 108.410 138.950 ;
        RECT 112.640 138.910 113.570 139.000 ;
        RECT 107.990 137.660 108.380 137.990 ;
        RECT 108.620 137.950 109.570 138.040 ;
        RECT 108.560 137.940 113.520 137.950 ;
        RECT 108.560 137.720 113.570 137.940 ;
        RECT 108.570 137.710 113.570 137.720 ;
        RECT 108.620 137.660 109.570 137.710 ;
        RECT 107.990 136.700 108.410 137.660 ;
        RECT 107.990 136.370 108.380 136.700 ;
        RECT 112.650 136.660 113.570 136.730 ;
        RECT 108.560 136.430 113.570 136.660 ;
        RECT 108.570 136.420 113.570 136.430 ;
        RECT 107.990 135.410 108.410 136.370 ;
        RECT 112.650 136.360 113.570 136.420 ;
        RECT 107.990 135.080 108.380 135.410 ;
        RECT 108.620 135.360 109.570 135.440 ;
        RECT 108.560 135.130 113.570 135.360 ;
        RECT 107.270 134.110 108.420 135.080 ;
        RECT 108.620 135.040 109.570 135.130 ;
        RECT 113.730 134.120 114.010 139.530 ;
        RECT 122.190 140.480 122.470 142.420 ;
        RECT 122.770 142.410 123.090 143.390 ;
        RECT 124.030 143.360 129.030 143.380 ;
        RECT 124.000 142.470 129.050 143.360 ;
        RECT 129.760 143.070 130.870 143.410 ;
        RECT 124.030 142.440 129.030 142.470 ;
        RECT 122.770 142.390 123.830 142.410 ;
        RECT 122.770 141.430 123.870 142.390 ;
        RECT 129.190 141.430 129.420 142.390 ;
        RECT 122.770 141.410 123.830 141.430 ;
        RECT 122.190 139.450 122.580 140.480 ;
        RECT 122.770 138.960 123.090 141.410 ;
        RECT 124.030 141.150 129.030 141.380 ;
        RECT 124.990 140.820 126.720 141.150 ;
        RECT 129.760 140.620 130.080 143.070 ;
        RECT 132.260 142.220 132.590 145.420 ;
        RECT 136.890 145.280 137.610 145.420 ;
        RECT 137.960 145.370 138.290 145.430 ;
        RECT 137.170 144.860 137.790 144.920 ;
        RECT 137.955 144.910 138.290 145.370 ;
        RECT 132.750 144.630 137.790 144.860 ;
        RECT 137.170 144.420 137.790 144.630 ;
        RECT 131.930 141.330 132.590 142.220 ;
        RECT 129.750 138.990 130.080 140.620 ;
        RECT 120.090 138.670 121.610 138.800 ;
        RECT 117.030 138.440 122.030 138.670 ;
        RECT 116.640 137.430 116.870 138.390 ;
        RECT 120.090 138.280 121.610 138.440 ;
        RECT 122.760 138.430 123.100 138.960 ;
        RECT 127.150 138.670 129.040 138.790 ;
        RECT 124.030 138.440 129.040 138.670 ;
        RECT 122.190 137.380 123.100 138.430 ;
        RECT 123.640 137.430 123.870 138.390 ;
        RECT 127.150 138.170 129.040 138.440 ;
        RECT 129.760 138.410 130.080 138.990 ;
        RECT 129.220 138.390 130.080 138.410 ;
        RECT 129.190 137.430 130.080 138.390 ;
        RECT 129.220 137.400 130.080 137.430 ;
        RECT 132.260 140.330 132.590 141.330 ;
        RECT 136.940 141.150 137.660 141.270 ;
        RECT 132.750 140.920 137.750 141.150 ;
        RECT 136.940 140.700 137.660 140.920 ;
        RECT 137.960 140.870 138.290 144.910 ;
        RECT 137.955 140.410 138.290 140.870 ;
        RECT 132.750 140.330 137.750 140.360 ;
        RECT 132.260 140.250 137.750 140.330 ;
        RECT 137.960 140.250 138.290 140.410 ;
        RECT 132.260 140.130 138.290 140.250 ;
        RECT 132.260 140.080 132.920 140.130 ;
        RECT 117.030 137.360 122.030 137.380 ;
        RECT 117.000 137.150 122.030 137.360 ;
        RECT 117.000 136.670 121.820 137.150 ;
        RECT 117.000 136.470 122.030 136.670 ;
        RECT 117.030 136.440 122.030 136.470 ;
        RECT 116.640 135.430 116.870 136.390 ;
        RECT 118.020 135.380 119.540 135.480 ;
        RECT 122.180 135.410 122.530 136.450 ;
        RECT 122.760 136.430 123.100 137.380 ;
        RECT 124.030 137.360 129.030 137.380 ;
        RECT 124.010 136.470 129.060 137.360 ;
        RECT 124.030 136.440 129.030 136.470 ;
        RECT 122.760 136.390 123.840 136.430 ;
        RECT 117.030 135.150 122.030 135.380 ;
        RECT 118.020 134.960 119.540 135.150 ;
        RECT 122.760 134.990 123.870 136.390 ;
        RECT 129.190 135.430 129.420 136.390 ;
        RECT 132.260 135.900 132.590 140.080 ;
        RECT 136.970 139.900 138.290 140.130 ;
        RECT 136.900 136.650 137.720 136.820 ;
        RECT 132.750 136.420 137.750 136.650 ;
        RECT 136.900 136.320 137.720 136.420 ;
        RECT 137.960 136.370 138.290 139.900 ;
        RECT 132.970 135.860 134.770 136.010 ;
        RECT 137.955 135.910 138.290 136.370 ;
        RECT 137.120 135.860 137.780 135.880 ;
        RECT 132.750 135.630 137.780 135.860 ;
        RECT 124.030 135.150 129.030 135.380 ;
        RECT 132.970 135.190 134.770 135.630 ;
        RECT 137.120 135.410 137.780 135.630 ;
        RECT 124.990 134.810 126.720 135.150 ;
        RECT 99.980 133.510 103.780 133.680 ;
        RECT 99.980 133.475 100.940 133.510 ;
        RECT 96.560 133.270 98.500 133.300 ;
        RECT 96.560 131.300 98.640 133.270 ;
        RECT 96.700 131.270 98.640 131.300 ;
        RECT 92.810 130.250 93.510 130.870 ;
        RECT 94.260 130.865 95.220 131.095 ;
        RECT 95.550 130.865 96.510 131.095 ;
        RECT 89.370 128.820 89.910 130.080 ;
        RECT 92.810 129.660 93.500 130.250 ;
        RECT 94.260 129.660 95.220 129.685 ;
        RECT 91.420 129.490 95.220 129.660 ;
        RECT 91.420 129.210 92.260 129.490 ;
        RECT 94.260 129.455 95.220 129.490 ;
        RECT 95.550 129.455 96.510 129.685 ;
        RECT 92.470 129.250 94.190 129.270 ;
        RECT 90.070 128.980 91.030 129.210 ;
        RECT 91.360 128.980 92.320 129.210 ;
        RECT 89.370 127.820 90.020 128.820 ;
        RECT 89.370 127.290 89.910 127.820 ;
        RECT 90.290 127.660 90.810 128.980 ;
        RECT 91.080 127.820 91.310 128.820 ;
        RECT 91.560 127.660 92.080 128.980 ;
        RECT 92.470 128.820 94.210 129.250 ;
        RECT 92.370 127.820 94.210 128.820 ;
        RECT 90.070 127.430 91.030 127.660 ;
        RECT 91.360 127.430 92.320 127.660 ;
        RECT 89.370 127.170 89.920 127.290 ;
        RECT 92.470 127.250 94.210 127.820 ;
        RECT 92.470 127.230 94.190 127.250 ;
        RECT 89.370 126.030 89.930 127.170 ;
        RECT 92.810 126.820 93.500 127.230 ;
        RECT 94.490 127.045 95.010 129.455 ;
        RECT 95.270 127.250 95.500 129.250 ;
        RECT 95.820 127.045 96.340 129.455 ;
        RECT 96.700 129.250 98.500 131.270 ;
        RECT 98.860 131.065 99.380 133.475 ;
        RECT 99.700 131.270 99.930 133.270 ;
        RECT 100.190 131.065 100.710 133.475 ;
        RECT 101.010 133.270 102.730 133.290 ;
        RECT 100.990 132.840 102.730 133.270 ;
        RECT 102.940 133.230 103.780 133.510 ;
        RECT 102.880 133.000 103.840 133.230 ;
        RECT 104.170 133.000 105.130 133.230 ;
        RECT 100.990 131.840 102.830 132.840 ;
        RECT 100.990 131.270 102.730 131.840 ;
        RECT 103.120 131.680 103.640 133.000 ;
        RECT 103.890 131.840 104.120 132.840 ;
        RECT 104.390 131.680 104.910 133.000 ;
        RECT 105.290 132.890 106.460 134.110 ;
        RECT 112.650 134.070 113.580 134.120 ;
        RECT 108.570 133.840 113.580 134.070 ;
        RECT 112.650 133.800 113.580 133.840 ;
        RECT 138.610 133.780 139.000 146.110 ;
        RECT 139.480 135.440 140.120 145.930 ;
        RECT 140.660 135.520 141.050 145.980 ;
        RECT 141.780 145.650 142.730 145.730 ;
        RECT 141.750 145.420 146.750 145.650 ;
        RECT 141.240 144.910 141.570 145.400 ;
        RECT 141.780 145.290 142.730 145.420 ;
        RECT 141.240 144.860 142.530 144.910 ;
        RECT 141.240 144.840 146.750 144.860 ;
        RECT 146.940 144.840 147.270 145.450 ;
        RECT 141.240 144.630 147.270 144.840 ;
        RECT 141.240 144.620 142.530 144.630 ;
        RECT 141.240 135.960 141.570 144.620 ;
        RECT 146.430 144.580 147.270 144.630 ;
        RECT 141.770 141.150 142.710 141.340 ;
        RECT 141.750 140.920 146.750 141.150 ;
        RECT 141.770 140.870 142.710 140.920 ;
        RECT 141.740 140.360 142.710 140.460 ;
        RECT 141.740 140.130 146.750 140.360 ;
        RECT 141.740 139.740 142.710 140.130 ;
        RECT 141.710 136.650 142.710 136.800 ;
        RECT 141.710 136.420 146.750 136.650 ;
        RECT 141.710 136.340 142.710 136.420 ;
        RECT 146.940 136.020 147.270 144.580 ;
        RECT 141.240 135.880 142.540 135.960 ;
        RECT 141.290 135.860 142.540 135.880 ;
        RECT 146.520 135.930 147.270 136.020 ;
        RECT 146.520 135.860 147.240 135.930 ;
        RECT 141.290 135.650 147.240 135.860 ;
        RECT 141.290 135.630 146.750 135.650 ;
        RECT 141.290 135.610 142.540 135.630 ;
        RECT 147.460 134.830 148.020 146.440 ;
        RECT 138.330 132.980 139.560 133.780 ;
        RECT 147.460 132.980 148.030 134.830 ;
        RECT 105.290 132.840 111.920 132.890 ;
        RECT 105.180 132.200 111.920 132.840 ;
        RECT 114.070 132.260 116.495 132.380 ;
        RECT 123.450 132.320 148.030 132.980 ;
        RECT 123.450 132.260 124.230 132.320 ;
        RECT 105.180 132.050 106.350 132.200 ;
        RECT 106.900 132.050 111.920 132.200 ;
        RECT 114.045 132.170 116.495 132.260 ;
        RECT 105.180 131.840 106.330 132.050 ;
        RECT 106.900 132.025 111.900 132.050 ;
        RECT 114.045 132.030 115.045 132.170 ;
        RECT 115.710 132.150 116.495 132.170 ;
        RECT 115.710 132.120 116.090 132.150 ;
        RECT 102.880 131.450 103.840 131.680 ;
        RECT 104.170 131.450 105.130 131.680 ;
        RECT 105.290 131.310 106.330 131.840 ;
        RECT 101.010 131.250 102.730 131.270 ;
        RECT 98.690 130.835 99.650 131.065 ;
        RECT 99.980 130.835 100.940 131.065 ;
        RECT 101.700 130.840 102.390 131.250 ;
        RECT 105.280 131.190 106.330 131.310 ;
        RECT 101.690 130.220 102.390 130.840 ;
        RECT 98.690 129.415 99.650 129.645 ;
        RECT 99.980 129.620 100.940 129.645 ;
        RECT 101.700 129.620 102.390 130.220 ;
        RECT 105.270 130.050 106.330 131.190 ;
        RECT 106.510 131.720 106.740 131.975 ;
        RECT 112.060 131.720 112.290 131.975 ;
        RECT 106.510 131.380 112.290 131.720 ;
        RECT 106.510 131.015 106.740 131.380 ;
        RECT 112.060 131.015 112.290 131.380 ;
        RECT 113.560 131.470 113.850 132.000 ;
        RECT 116.265 131.980 116.495 132.150 ;
        RECT 116.705 132.060 124.230 132.260 ;
        RECT 116.705 132.030 124.205 132.060 ;
        RECT 124.800 131.990 148.030 132.320 ;
        RECT 115.245 131.470 115.635 131.980 ;
        RECT 116.265 131.470 116.500 131.980 ;
        RECT 124.410 131.770 124.640 131.980 ;
        RECT 123.630 131.520 124.640 131.770 ;
        RECT 123.630 131.470 124.610 131.520 ;
        RECT 106.900 130.950 111.900 130.965 ;
        RECT 106.870 130.740 111.900 130.950 ;
        RECT 106.870 130.600 111.905 130.740 ;
        RECT 113.560 130.710 115.960 131.470 ;
        RECT 116.265 131.430 124.610 131.470 ;
        RECT 116.265 131.240 124.205 131.430 ;
        RECT 124.800 131.150 125.290 131.990 ;
        RECT 124.390 130.940 125.290 131.150 ;
        RECT 112.170 130.600 115.960 130.710 ;
        RECT 106.870 130.470 115.960 130.600 ;
        RECT 111.690 130.410 112.390 130.470 ;
        RECT 113.560 130.460 115.960 130.470 ;
        RECT 99.980 129.450 103.780 129.620 ;
        RECT 99.980 129.415 100.940 129.450 ;
        RECT 96.560 129.210 98.500 129.250 ;
        RECT 96.560 127.250 98.640 129.210 ;
        RECT 96.700 127.210 98.640 127.250 ;
        RECT 92.810 126.200 93.510 126.820 ;
        RECT 94.260 126.815 95.220 127.045 ;
        RECT 95.550 126.815 96.510 127.045 ;
        RECT 89.370 124.770 89.910 126.030 ;
        RECT 92.810 125.610 93.500 126.200 ;
        RECT 94.260 125.610 95.220 125.635 ;
        RECT 91.420 125.440 95.220 125.610 ;
        RECT 91.420 125.160 92.260 125.440 ;
        RECT 94.260 125.405 95.220 125.440 ;
        RECT 95.550 125.405 96.510 125.635 ;
        RECT 92.470 125.200 94.190 125.220 ;
        RECT 90.070 124.930 91.030 125.160 ;
        RECT 91.360 124.930 92.320 125.160 ;
        RECT 89.370 123.770 90.020 124.770 ;
        RECT 89.370 123.240 89.910 123.770 ;
        RECT 90.290 123.610 90.810 124.930 ;
        RECT 91.080 123.770 91.310 124.770 ;
        RECT 91.560 123.610 92.080 124.930 ;
        RECT 92.470 124.770 94.210 125.200 ;
        RECT 92.370 123.770 94.210 124.770 ;
        RECT 90.070 123.380 91.030 123.610 ;
        RECT 91.360 123.380 92.320 123.610 ;
        RECT 89.370 123.120 89.920 123.240 ;
        RECT 92.470 123.200 94.210 123.770 ;
        RECT 92.470 123.180 94.190 123.200 ;
        RECT 89.370 121.980 89.930 123.120 ;
        RECT 92.810 122.770 93.500 123.180 ;
        RECT 94.490 122.995 95.010 125.405 ;
        RECT 95.270 123.200 95.500 125.200 ;
        RECT 95.820 122.995 96.340 125.405 ;
        RECT 96.700 125.200 98.500 127.210 ;
        RECT 98.860 127.005 99.380 129.415 ;
        RECT 99.700 127.210 99.930 129.210 ;
        RECT 100.190 127.005 100.710 129.415 ;
        RECT 101.010 129.210 102.730 129.230 ;
        RECT 100.990 128.780 102.730 129.210 ;
        RECT 102.940 129.170 103.780 129.450 ;
        RECT 102.880 128.940 103.840 129.170 ;
        RECT 104.170 128.940 105.130 129.170 ;
        RECT 100.990 127.780 102.830 128.780 ;
        RECT 100.990 127.210 102.730 127.780 ;
        RECT 103.120 127.620 103.640 128.940 ;
        RECT 103.890 127.780 104.120 128.780 ;
        RECT 104.390 127.620 104.910 128.940 ;
        RECT 105.290 128.780 106.330 130.050 ;
        RECT 115.790 129.810 115.960 130.460 ;
        RECT 116.760 130.590 125.290 130.940 ;
        RECT 116.760 130.190 122.380 130.590 ;
        RECT 122.740 129.900 123.650 130.220 ;
        RECT 116.700 129.885 123.670 129.900 ;
        RECT 115.790 129.510 116.510 129.810 ;
        RECT 116.700 129.655 123.710 129.885 ;
        RECT 116.700 129.560 123.670 129.655 ;
        RECT 105.180 127.780 106.330 128.780 ;
        RECT 116.210 128.590 116.510 129.510 ;
        RECT 102.880 127.390 103.840 127.620 ;
        RECT 104.170 127.390 105.130 127.620 ;
        RECT 105.290 127.250 106.330 127.780 ;
        RECT 101.010 127.190 102.730 127.210 ;
        RECT 98.690 126.775 99.650 127.005 ;
        RECT 99.980 126.775 100.940 127.005 ;
        RECT 101.700 126.780 102.390 127.190 ;
        RECT 105.280 127.130 106.330 127.250 ;
        RECT 101.690 126.160 102.390 126.780 ;
        RECT 98.690 125.355 99.650 125.585 ;
        RECT 99.980 125.560 100.940 125.585 ;
        RECT 101.700 125.560 102.390 126.160 ;
        RECT 105.270 125.990 106.330 127.130 ;
        RECT 105.290 125.750 106.330 125.990 ;
        RECT 99.980 125.390 103.780 125.560 ;
        RECT 99.980 125.355 100.940 125.390 ;
        RECT 96.560 125.150 98.500 125.200 ;
        RECT 96.560 123.200 98.640 125.150 ;
        RECT 96.700 123.150 98.640 123.200 ;
        RECT 92.810 122.150 93.510 122.770 ;
        RECT 94.260 122.765 95.220 122.995 ;
        RECT 95.550 122.765 96.510 122.995 ;
        RECT 89.370 120.720 89.910 121.980 ;
        RECT 92.810 121.560 93.500 122.150 ;
        RECT 94.260 121.560 95.220 121.585 ;
        RECT 91.420 121.390 95.220 121.560 ;
        RECT 91.420 121.110 92.260 121.390 ;
        RECT 94.260 121.355 95.220 121.390 ;
        RECT 95.550 121.355 96.510 121.585 ;
        RECT 92.470 121.150 94.190 121.170 ;
        RECT 90.070 120.880 91.030 121.110 ;
        RECT 91.360 120.880 92.320 121.110 ;
        RECT 89.370 119.720 90.020 120.720 ;
        RECT 89.370 119.190 89.910 119.720 ;
        RECT 90.290 119.560 90.810 120.880 ;
        RECT 91.080 119.720 91.310 120.720 ;
        RECT 91.560 119.560 92.080 120.880 ;
        RECT 92.470 120.720 94.210 121.150 ;
        RECT 92.370 119.720 94.210 120.720 ;
        RECT 90.070 119.330 91.030 119.560 ;
        RECT 91.360 119.330 92.320 119.560 ;
        RECT 89.370 119.070 89.920 119.190 ;
        RECT 92.470 119.150 94.210 119.720 ;
        RECT 92.470 119.130 94.190 119.150 ;
        RECT 89.370 117.930 89.930 119.070 ;
        RECT 92.810 118.720 93.500 119.130 ;
        RECT 94.490 118.945 95.010 121.355 ;
        RECT 95.270 119.150 95.500 121.150 ;
        RECT 95.820 118.945 96.340 121.355 ;
        RECT 96.700 121.150 98.500 123.150 ;
        RECT 98.860 122.945 99.380 125.355 ;
        RECT 99.700 123.150 99.930 125.150 ;
        RECT 100.190 122.945 100.710 125.355 ;
        RECT 101.010 125.150 102.730 125.170 ;
        RECT 100.990 124.720 102.730 125.150 ;
        RECT 102.940 125.110 103.780 125.390 ;
        RECT 102.880 124.880 103.840 125.110 ;
        RECT 104.170 124.880 105.130 125.110 ;
        RECT 100.990 123.720 102.830 124.720 ;
        RECT 100.990 123.150 102.730 123.720 ;
        RECT 103.120 123.560 103.640 124.880 ;
        RECT 103.890 123.720 104.120 124.720 ;
        RECT 104.390 123.560 104.910 124.880 ;
        RECT 105.290 124.720 106.450 125.750 ;
        RECT 107.120 125.040 111.960 125.100 ;
        RECT 107.100 124.810 112.100 125.040 ;
        RECT 105.180 123.720 106.450 124.720 ;
        RECT 102.880 123.330 103.840 123.560 ;
        RECT 104.170 123.330 105.130 123.560 ;
        RECT 105.290 123.190 106.450 123.720 ;
        RECT 101.010 123.130 102.730 123.150 ;
        RECT 98.690 122.715 99.650 122.945 ;
        RECT 99.980 122.715 100.940 122.945 ;
        RECT 101.700 122.720 102.390 123.130 ;
        RECT 105.280 123.070 106.450 123.190 ;
        RECT 101.690 122.100 102.390 122.720 ;
        RECT 98.690 121.295 99.650 121.525 ;
        RECT 99.980 121.500 100.940 121.525 ;
        RECT 101.700 121.500 102.390 122.100 ;
        RECT 105.270 121.930 106.450 123.070 ;
        RECT 99.980 121.330 103.780 121.500 ;
        RECT 99.980 121.295 100.940 121.330 ;
        RECT 96.560 121.090 98.500 121.150 ;
        RECT 96.560 119.150 98.640 121.090 ;
        RECT 96.700 119.090 98.640 119.150 ;
        RECT 92.810 118.100 93.510 118.720 ;
        RECT 94.260 118.715 95.220 118.945 ;
        RECT 95.550 118.715 96.510 118.945 ;
        RECT 89.370 116.670 89.910 117.930 ;
        RECT 92.810 117.510 93.500 118.100 ;
        RECT 94.260 117.510 95.220 117.535 ;
        RECT 91.420 117.340 95.220 117.510 ;
        RECT 91.420 117.060 92.260 117.340 ;
        RECT 94.260 117.305 95.220 117.340 ;
        RECT 95.550 117.305 96.510 117.535 ;
        RECT 92.470 117.100 94.190 117.120 ;
        RECT 90.070 116.830 91.030 117.060 ;
        RECT 91.360 116.830 92.320 117.060 ;
        RECT 89.370 115.670 90.020 116.670 ;
        RECT 89.370 115.140 89.910 115.670 ;
        RECT 90.290 115.510 90.810 116.830 ;
        RECT 91.080 115.670 91.310 116.670 ;
        RECT 91.560 115.510 92.080 116.830 ;
        RECT 92.470 116.670 94.210 117.100 ;
        RECT 92.370 115.670 94.210 116.670 ;
        RECT 90.070 115.280 91.030 115.510 ;
        RECT 91.360 115.280 92.320 115.510 ;
        RECT 89.370 115.020 89.920 115.140 ;
        RECT 92.470 115.100 94.210 115.670 ;
        RECT 92.470 115.080 94.190 115.100 ;
        RECT 89.370 113.880 89.930 115.020 ;
        RECT 92.810 114.670 93.500 115.080 ;
        RECT 94.490 114.895 95.010 117.305 ;
        RECT 95.270 115.100 95.500 117.100 ;
        RECT 95.820 114.895 96.340 117.305 ;
        RECT 96.700 117.100 98.500 119.090 ;
        RECT 98.860 118.885 99.380 121.295 ;
        RECT 99.700 119.090 99.930 121.090 ;
        RECT 100.190 118.885 100.710 121.295 ;
        RECT 101.010 121.090 102.730 121.110 ;
        RECT 100.990 120.660 102.730 121.090 ;
        RECT 102.940 121.050 103.780 121.330 ;
        RECT 102.880 120.820 103.840 121.050 ;
        RECT 104.170 120.820 105.130 121.050 ;
        RECT 100.990 119.660 102.830 120.660 ;
        RECT 100.990 119.090 102.730 119.660 ;
        RECT 103.120 119.500 103.640 120.820 ;
        RECT 103.890 119.660 104.120 120.660 ;
        RECT 104.390 119.500 104.910 120.820 ;
        RECT 105.290 120.660 106.450 121.930 ;
        RECT 105.180 119.660 106.450 120.660 ;
        RECT 102.880 119.270 103.840 119.500 ;
        RECT 104.170 119.270 105.130 119.500 ;
        RECT 105.290 119.130 106.450 119.660 ;
        RECT 101.010 119.070 102.730 119.090 ;
        RECT 98.690 118.655 99.650 118.885 ;
        RECT 99.980 118.655 100.940 118.885 ;
        RECT 101.700 118.660 102.390 119.070 ;
        RECT 105.280 119.010 106.450 119.130 ;
        RECT 101.690 118.040 102.390 118.660 ;
        RECT 98.690 117.235 99.650 117.465 ;
        RECT 99.980 117.440 100.940 117.465 ;
        RECT 101.700 117.440 102.390 118.040 ;
        RECT 105.270 117.870 106.450 119.010 ;
        RECT 99.980 117.270 103.780 117.440 ;
        RECT 99.980 117.235 100.940 117.270 ;
        RECT 96.560 117.030 98.500 117.100 ;
        RECT 96.560 115.100 98.640 117.030 ;
        RECT 96.700 115.030 98.640 115.100 ;
        RECT 92.810 114.050 93.510 114.670 ;
        RECT 94.260 114.665 95.220 114.895 ;
        RECT 95.550 114.665 96.510 114.895 ;
        RECT 89.370 112.620 89.910 113.880 ;
        RECT 92.810 113.460 93.500 114.050 ;
        RECT 94.260 113.460 95.220 113.485 ;
        RECT 91.420 113.290 95.220 113.460 ;
        RECT 91.420 113.010 92.260 113.290 ;
        RECT 94.260 113.255 95.220 113.290 ;
        RECT 95.550 113.255 96.510 113.485 ;
        RECT 92.470 113.050 94.190 113.070 ;
        RECT 90.070 112.780 91.030 113.010 ;
        RECT 91.360 112.780 92.320 113.010 ;
        RECT 89.370 111.620 90.020 112.620 ;
        RECT 89.370 111.090 89.910 111.620 ;
        RECT 90.290 111.460 90.810 112.780 ;
        RECT 91.080 111.620 91.310 112.620 ;
        RECT 91.560 111.460 92.080 112.780 ;
        RECT 92.470 112.620 94.210 113.050 ;
        RECT 92.370 111.620 94.210 112.620 ;
        RECT 90.070 111.230 91.030 111.460 ;
        RECT 91.360 111.230 92.320 111.460 ;
        RECT 89.370 110.970 89.920 111.090 ;
        RECT 92.470 111.050 94.210 111.620 ;
        RECT 92.470 111.030 94.190 111.050 ;
        RECT 89.370 109.830 89.930 110.970 ;
        RECT 92.810 110.620 93.500 111.030 ;
        RECT 94.490 110.845 95.010 113.255 ;
        RECT 95.270 111.050 95.500 113.050 ;
        RECT 95.820 110.845 96.340 113.255 ;
        RECT 96.700 113.050 98.500 115.030 ;
        RECT 98.860 114.825 99.380 117.235 ;
        RECT 99.700 115.030 99.930 117.030 ;
        RECT 100.190 114.825 100.710 117.235 ;
        RECT 101.010 117.030 102.730 117.050 ;
        RECT 100.990 116.600 102.730 117.030 ;
        RECT 102.940 116.990 103.780 117.270 ;
        RECT 102.880 116.760 103.840 116.990 ;
        RECT 104.170 116.760 105.130 116.990 ;
        RECT 100.990 115.600 102.830 116.600 ;
        RECT 100.990 115.030 102.730 115.600 ;
        RECT 103.120 115.440 103.640 116.760 ;
        RECT 103.890 115.600 104.120 116.600 ;
        RECT 104.390 115.440 104.910 116.760 ;
        RECT 105.290 116.600 106.450 117.870 ;
        RECT 105.180 115.600 106.450 116.600 ;
        RECT 102.880 115.210 103.840 115.440 ;
        RECT 104.170 115.210 105.130 115.440 ;
        RECT 105.290 115.070 106.450 115.600 ;
        RECT 101.010 115.010 102.730 115.030 ;
        RECT 98.690 114.595 99.650 114.825 ;
        RECT 99.980 114.595 100.940 114.825 ;
        RECT 101.700 114.600 102.390 115.010 ;
        RECT 105.280 114.950 106.450 115.070 ;
        RECT 101.690 113.980 102.390 114.600 ;
        RECT 98.690 113.175 99.650 113.405 ;
        RECT 99.980 113.380 100.940 113.405 ;
        RECT 101.700 113.380 102.390 113.980 ;
        RECT 105.270 113.810 106.450 114.950 ;
        RECT 99.980 113.210 103.780 113.380 ;
        RECT 99.980 113.175 100.940 113.210 ;
        RECT 96.560 112.970 98.500 113.050 ;
        RECT 96.560 111.050 98.640 112.970 ;
        RECT 96.700 110.970 98.640 111.050 ;
        RECT 92.810 110.000 93.510 110.620 ;
        RECT 94.260 110.615 95.220 110.845 ;
        RECT 95.550 110.615 96.510 110.845 ;
        RECT 89.370 108.570 89.910 109.830 ;
        RECT 92.810 109.410 93.500 110.000 ;
        RECT 94.260 109.410 95.220 109.435 ;
        RECT 91.420 109.240 95.220 109.410 ;
        RECT 91.420 108.960 92.260 109.240 ;
        RECT 94.260 109.205 95.220 109.240 ;
        RECT 95.550 109.205 96.510 109.435 ;
        RECT 92.470 109.000 94.190 109.020 ;
        RECT 90.070 108.730 91.030 108.960 ;
        RECT 91.360 108.730 92.320 108.960 ;
        RECT 89.370 107.570 90.020 108.570 ;
        RECT 89.370 107.040 89.910 107.570 ;
        RECT 90.290 107.410 90.810 108.730 ;
        RECT 91.080 107.570 91.310 108.570 ;
        RECT 91.560 107.410 92.080 108.730 ;
        RECT 92.470 108.570 94.210 109.000 ;
        RECT 92.370 107.570 94.210 108.570 ;
        RECT 90.070 107.180 91.030 107.410 ;
        RECT 91.360 107.180 92.320 107.410 ;
        RECT 89.370 106.920 89.920 107.040 ;
        RECT 92.470 107.000 94.210 107.570 ;
        RECT 92.470 106.980 94.190 107.000 ;
        RECT 89.370 105.780 89.930 106.920 ;
        RECT 92.810 106.570 93.500 106.980 ;
        RECT 94.490 106.795 95.010 109.205 ;
        RECT 95.270 107.000 95.500 109.000 ;
        RECT 95.820 106.795 96.340 109.205 ;
        RECT 96.700 109.000 98.500 110.970 ;
        RECT 98.860 110.765 99.380 113.175 ;
        RECT 99.700 110.970 99.930 112.970 ;
        RECT 100.190 110.765 100.710 113.175 ;
        RECT 101.010 112.970 102.730 112.990 ;
        RECT 100.990 112.540 102.730 112.970 ;
        RECT 102.940 112.930 103.780 113.210 ;
        RECT 102.880 112.700 103.840 112.930 ;
        RECT 104.170 112.700 105.130 112.930 ;
        RECT 100.990 111.540 102.830 112.540 ;
        RECT 100.990 110.970 102.730 111.540 ;
        RECT 103.120 111.380 103.640 112.700 ;
        RECT 103.890 111.540 104.120 112.540 ;
        RECT 104.390 111.380 104.910 112.700 ;
        RECT 105.290 112.540 106.450 113.810 ;
        RECT 105.180 111.540 106.450 112.540 ;
        RECT 102.880 111.150 103.840 111.380 ;
        RECT 104.170 111.150 105.130 111.380 ;
        RECT 105.290 111.010 106.450 111.540 ;
        RECT 101.010 110.950 102.730 110.970 ;
        RECT 98.690 110.535 99.650 110.765 ;
        RECT 99.980 110.535 100.940 110.765 ;
        RECT 101.700 110.540 102.390 110.950 ;
        RECT 105.280 110.890 106.450 111.010 ;
        RECT 101.690 109.920 102.390 110.540 ;
        RECT 98.690 109.115 99.650 109.345 ;
        RECT 99.980 109.320 100.940 109.345 ;
        RECT 101.700 109.320 102.390 109.920 ;
        RECT 105.270 109.750 106.450 110.890 ;
        RECT 106.620 124.760 106.930 124.810 ;
        RECT 107.120 124.760 111.960 124.810 ;
        RECT 106.620 124.300 106.940 124.760 ;
        RECT 110.810 124.330 112.020 124.340 ;
        RECT 106.620 123.970 106.930 124.300 ;
        RECT 110.800 124.250 112.020 124.330 ;
        RECT 107.100 124.020 112.100 124.250 ;
        RECT 110.800 123.970 112.020 124.020 ;
        RECT 106.620 123.510 106.940 123.970 ;
        RECT 110.810 123.940 112.020 123.970 ;
        RECT 112.260 123.920 113.130 128.380 ;
        RECT 116.220 127.200 116.510 128.590 ;
        RECT 116.680 127.740 123.720 129.100 ;
        RECT 116.710 127.725 123.710 127.740 ;
        RECT 122.740 127.230 123.650 127.250 ;
        RECT 116.700 127.165 123.670 127.230 ;
        RECT 123.900 127.200 124.190 129.630 ;
        RECT 116.700 126.935 123.710 127.165 ;
        RECT 116.700 126.890 123.670 126.935 ;
        RECT 122.740 126.690 123.650 126.890 ;
        RECT 124.390 125.750 125.290 130.590 ;
        RECT 141.710 130.490 147.190 130.750 ;
        RECT 141.710 130.160 147.290 130.490 ;
        RECT 141.710 130.070 142.380 130.160 ;
        RECT 141.690 128.110 142.380 130.070 ;
        RECT 146.820 128.460 147.290 130.160 ;
        RECT 146.820 128.110 147.320 128.460 ;
        RECT 141.690 127.520 147.320 128.110 ;
        RECT 141.830 127.480 147.320 127.520 ;
        RECT 141.710 126.680 147.360 127.190 ;
        RECT 112.260 123.870 113.110 123.920 ;
        RECT 106.620 123.180 106.930 123.510 ;
        RECT 107.290 123.460 108.570 123.550 ;
        RECT 112.260 123.510 112.590 123.870 ;
        RECT 113.820 123.700 115.000 125.200 ;
        RECT 120.790 124.920 125.290 125.750 ;
        RECT 144.700 125.930 145.240 126.680 ;
        RECT 146.750 125.930 147.340 126.680 ;
        RECT 144.700 125.620 147.340 125.930 ;
        RECT 144.870 125.580 147.340 125.620 ;
        RECT 115.320 124.860 116.580 124.920 ;
        RECT 115.160 124.630 120.160 124.860 ;
        RECT 115.320 124.570 116.580 124.630 ;
        RECT 118.910 124.070 120.030 124.090 ;
        RECT 115.160 123.840 120.160 124.070 ;
        RECT 118.910 123.740 120.030 123.840 ;
        RECT 114.040 123.690 115.000 123.700 ;
        RECT 107.100 123.230 112.100 123.460 ;
        RECT 106.620 122.720 106.940 123.180 ;
        RECT 107.290 123.150 108.570 123.230 ;
        RECT 112.280 123.180 112.590 123.510 ;
        RECT 112.260 122.720 112.590 123.180 ;
        RECT 106.620 122.390 106.930 122.720 ;
        RECT 110.800 122.670 112.020 122.710 ;
        RECT 107.100 122.440 112.100 122.670 ;
        RECT 106.620 121.930 106.940 122.390 ;
        RECT 110.800 122.350 112.020 122.440 ;
        RECT 112.280 122.390 112.590 122.720 ;
        RECT 106.620 121.600 106.930 121.930 ;
        RECT 107.290 121.880 108.570 121.950 ;
        RECT 112.260 121.930 112.590 122.390 ;
        RECT 107.100 121.650 112.100 121.880 ;
        RECT 106.620 121.140 106.940 121.600 ;
        RECT 107.290 121.550 108.570 121.650 ;
        RECT 112.280 121.600 112.590 121.930 ;
        RECT 112.260 121.140 112.590 121.600 ;
        RECT 106.620 120.810 106.930 121.140 ;
        RECT 110.800 121.090 112.040 121.140 ;
        RECT 107.100 120.860 112.100 121.090 ;
        RECT 106.620 120.350 106.940 120.810 ;
        RECT 110.800 120.790 112.040 120.860 ;
        RECT 112.280 120.810 112.590 121.140 ;
        RECT 106.620 120.020 106.930 120.350 ;
        RECT 107.250 120.300 108.580 120.360 ;
        RECT 112.260 120.350 112.590 120.810 ;
        RECT 107.100 120.070 112.100 120.300 ;
        RECT 106.620 119.560 106.940 120.020 ;
        RECT 107.250 119.960 108.580 120.070 ;
        RECT 112.280 120.020 112.590 120.350 ;
        RECT 112.260 119.560 112.590 120.020 ;
        RECT 106.620 119.230 106.930 119.560 ;
        RECT 110.790 119.510 111.940 119.530 ;
        RECT 107.100 119.280 112.100 119.510 ;
        RECT 106.620 118.770 106.940 119.230 ;
        RECT 110.790 119.170 111.940 119.280 ;
        RECT 112.280 119.230 112.590 119.560 ;
        RECT 106.620 118.440 106.930 118.770 ;
        RECT 107.300 118.720 108.560 118.830 ;
        RECT 112.260 118.770 112.590 119.230 ;
        RECT 107.100 118.490 112.100 118.720 ;
        RECT 106.620 117.980 106.940 118.440 ;
        RECT 107.300 118.380 108.560 118.490 ;
        RECT 112.280 118.440 112.590 118.770 ;
        RECT 112.260 117.980 112.590 118.440 ;
        RECT 106.620 117.650 106.930 117.980 ;
        RECT 110.800 117.930 111.920 117.970 ;
        RECT 107.100 117.700 112.100 117.930 ;
        RECT 106.620 117.190 106.940 117.650 ;
        RECT 110.800 117.630 111.920 117.700 ;
        RECT 112.280 117.650 112.590 117.980 ;
        RECT 112.260 117.190 112.590 117.650 ;
        RECT 106.620 116.860 106.930 117.190 ;
        RECT 107.310 117.140 108.570 117.180 ;
        RECT 107.100 116.910 112.100 117.140 ;
        RECT 106.620 116.400 106.940 116.860 ;
        RECT 107.310 116.830 108.570 116.910 ;
        RECT 112.280 116.860 112.590 117.190 ;
        RECT 112.260 116.400 112.590 116.860 ;
        RECT 106.620 116.070 106.930 116.400 ;
        RECT 110.800 116.350 111.950 116.380 ;
        RECT 107.100 116.120 112.100 116.350 ;
        RECT 106.620 115.610 106.940 116.070 ;
        RECT 110.800 116.030 111.950 116.120 ;
        RECT 112.280 116.070 112.590 116.400 ;
        RECT 106.620 115.280 106.930 115.610 ;
        RECT 107.300 115.560 108.570 115.620 ;
        RECT 112.260 115.610 112.590 116.070 ;
        RECT 107.100 115.330 112.100 115.560 ;
        RECT 106.620 114.820 106.940 115.280 ;
        RECT 107.300 115.260 108.570 115.330 ;
        RECT 112.280 115.280 112.590 115.610 ;
        RECT 112.260 114.820 112.590 115.280 ;
        RECT 106.620 114.490 106.930 114.820 ;
        RECT 110.800 114.770 111.990 114.810 ;
        RECT 107.100 114.540 112.100 114.770 ;
        RECT 106.620 114.030 106.940 114.490 ;
        RECT 110.800 114.450 111.990 114.540 ;
        RECT 112.280 114.490 112.590 114.820 ;
        RECT 112.260 114.030 112.590 114.490 ;
        RECT 106.620 113.700 106.930 114.030 ;
        RECT 107.290 113.980 108.570 114.020 ;
        RECT 107.100 113.750 112.100 113.980 ;
        RECT 106.620 113.240 106.940 113.700 ;
        RECT 107.290 113.660 108.570 113.750 ;
        RECT 112.280 113.700 112.590 114.030 ;
        RECT 112.260 113.240 112.590 113.700 ;
        RECT 114.700 113.680 115.000 123.690 ;
        RECT 115.310 123.280 116.570 123.360 ;
        RECT 115.160 123.050 120.160 123.280 ;
        RECT 115.310 123.000 116.570 123.050 ;
        RECT 118.920 122.490 120.040 122.520 ;
        RECT 115.160 122.260 120.160 122.490 ;
        RECT 118.920 122.180 120.040 122.260 ;
        RECT 115.320 121.700 116.580 121.770 ;
        RECT 115.160 121.470 120.160 121.700 ;
        RECT 115.320 121.410 116.580 121.470 ;
        RECT 118.920 120.910 120.010 120.940 ;
        RECT 115.160 120.680 120.160 120.910 ;
        RECT 118.920 120.580 120.010 120.680 ;
        RECT 115.320 120.120 116.580 120.170 ;
        RECT 115.160 119.890 120.160 120.120 ;
        RECT 115.320 119.810 116.580 119.890 ;
        RECT 118.920 119.330 120.080 119.400 ;
        RECT 115.160 119.100 120.160 119.330 ;
        RECT 118.920 118.980 120.080 119.100 ;
        RECT 115.320 118.540 116.580 118.570 ;
        RECT 115.160 118.310 120.160 118.540 ;
        RECT 115.320 118.230 116.580 118.310 ;
        RECT 118.920 117.750 120.070 117.850 ;
        RECT 115.160 117.520 120.160 117.750 ;
        RECT 118.920 117.390 120.070 117.520 ;
        RECT 115.320 116.960 116.580 117.040 ;
        RECT 115.160 116.730 120.160 116.960 ;
        RECT 115.320 116.700 116.580 116.730 ;
        RECT 118.920 116.170 120.020 116.250 ;
        RECT 115.160 115.940 120.160 116.170 ;
        RECT 118.920 115.830 120.020 115.940 ;
        RECT 115.320 115.380 116.580 115.410 ;
        RECT 115.160 115.150 120.160 115.380 ;
        RECT 115.320 115.070 116.580 115.150 ;
        RECT 118.920 114.590 120.000 114.680 ;
        RECT 115.160 114.360 120.160 114.590 ;
        RECT 118.920 114.250 120.000 114.360 ;
        RECT 115.320 113.800 116.580 113.830 ;
        RECT 115.160 113.570 120.160 113.800 ;
        RECT 120.350 113.700 120.650 124.650 ;
        RECT 115.320 113.480 116.580 113.570 ;
        RECT 106.620 112.910 106.930 113.240 ;
        RECT 110.800 113.190 111.950 113.220 ;
        RECT 107.100 112.960 112.100 113.190 ;
        RECT 106.620 112.450 106.940 112.910 ;
        RECT 110.800 112.870 111.950 112.960 ;
        RECT 112.280 112.910 112.590 113.240 ;
        RECT 112.260 112.450 112.590 112.910 ;
        RECT 106.620 112.120 106.930 112.450 ;
        RECT 107.300 112.400 108.570 112.430 ;
        RECT 107.100 112.170 112.100 112.400 ;
        RECT 106.620 111.660 106.940 112.120 ;
        RECT 107.300 112.040 108.570 112.170 ;
        RECT 112.280 112.120 112.590 112.450 ;
        RECT 110.810 111.660 111.990 111.710 ;
        RECT 112.260 111.660 112.590 112.120 ;
        RECT 120.790 112.110 121.210 124.920 ;
        RECT 141.690 124.250 147.380 124.760 ;
        RECT 141.690 123.730 145.170 124.250 ;
        RECT 144.660 122.940 145.170 123.730 ;
        RECT 144.670 122.380 145.170 122.940 ;
        RECT 141.710 122.350 145.170 122.380 ;
        RECT 146.850 123.730 147.380 124.250 ;
        RECT 146.850 122.690 147.320 123.730 ;
        RECT 146.850 122.350 147.400 122.690 ;
        RECT 141.710 121.660 147.400 122.350 ;
        RECT 141.730 119.260 147.420 119.860 ;
        RECT 141.730 118.820 147.440 119.260 ;
        RECT 146.580 117.480 147.440 118.820 ;
        RECT 141.790 116.450 147.480 117.480 ;
        RECT 146.580 115.070 147.440 116.450 ;
        RECT 141.850 114.030 147.540 115.070 ;
        RECT 141.770 112.410 147.460 112.600 ;
        RECT 106.620 111.330 106.930 111.660 ;
        RECT 110.800 111.610 111.990 111.660 ;
        RECT 107.100 111.380 112.100 111.610 ;
        RECT 106.620 110.870 106.940 111.330 ;
        RECT 110.800 111.320 111.990 111.380 ;
        RECT 112.280 111.330 112.590 111.660 ;
        RECT 141.770 111.910 147.550 112.410 ;
        RECT 141.770 111.560 144.700 111.910 ;
        RECT 110.810 111.290 111.990 111.320 ;
        RECT 112.260 110.870 112.590 111.330 ;
        RECT 106.620 110.540 106.930 110.870 ;
        RECT 107.300 110.820 108.580 110.850 ;
        RECT 107.100 110.590 112.100 110.820 ;
        RECT 106.620 110.080 106.940 110.540 ;
        RECT 107.300 110.490 108.580 110.590 ;
        RECT 112.280 110.540 112.590 110.870 ;
        RECT 112.260 110.080 112.590 110.540 ;
        RECT 106.620 109.970 106.930 110.080 ;
        RECT 110.790 110.030 111.990 110.060 ;
        RECT 107.100 109.800 112.100 110.030 ;
        RECT 112.280 109.980 112.590 110.080 ;
        RECT 144.200 110.520 144.700 111.560 ;
        RECT 146.850 110.520 147.550 111.910 ;
        RECT 144.200 110.210 147.550 110.520 ;
        RECT 144.200 109.960 147.540 110.210 ;
        RECT 99.980 109.150 103.780 109.320 ;
        RECT 99.980 109.115 100.940 109.150 ;
        RECT 96.560 108.910 98.500 109.000 ;
        RECT 96.560 107.000 98.640 108.910 ;
        RECT 96.700 106.910 98.640 107.000 ;
        RECT 92.810 105.950 93.510 106.570 ;
        RECT 94.260 106.565 95.220 106.795 ;
        RECT 95.550 106.565 96.510 106.795 ;
        RECT 89.370 104.520 89.910 105.780 ;
        RECT 92.810 105.360 93.500 105.950 ;
        RECT 94.260 105.360 95.220 105.385 ;
        RECT 91.420 105.190 95.220 105.360 ;
        RECT 91.420 104.910 92.260 105.190 ;
        RECT 94.260 105.155 95.220 105.190 ;
        RECT 95.550 105.155 96.510 105.385 ;
        RECT 92.470 104.950 94.190 104.970 ;
        RECT 90.070 104.680 91.030 104.910 ;
        RECT 91.360 104.680 92.320 104.910 ;
        RECT 89.370 103.520 90.020 104.520 ;
        RECT 89.370 102.990 89.910 103.520 ;
        RECT 90.290 103.360 90.810 104.680 ;
        RECT 91.080 103.520 91.310 104.520 ;
        RECT 91.560 103.360 92.080 104.680 ;
        RECT 92.470 104.520 94.210 104.950 ;
        RECT 92.370 103.520 94.210 104.520 ;
        RECT 90.070 103.130 91.030 103.360 ;
        RECT 91.360 103.130 92.320 103.360 ;
        RECT 89.370 102.870 89.920 102.990 ;
        RECT 92.470 102.950 94.210 103.520 ;
        RECT 92.470 102.930 94.190 102.950 ;
        RECT 89.370 101.730 89.930 102.870 ;
        RECT 92.810 102.520 93.500 102.930 ;
        RECT 94.490 102.745 95.010 105.155 ;
        RECT 95.270 102.950 95.500 104.950 ;
        RECT 95.820 102.745 96.340 105.155 ;
        RECT 96.700 104.950 98.500 106.910 ;
        RECT 98.860 106.705 99.380 109.115 ;
        RECT 99.700 106.910 99.930 108.910 ;
        RECT 100.190 106.705 100.710 109.115 ;
        RECT 101.010 108.910 102.730 108.930 ;
        RECT 100.990 108.480 102.730 108.910 ;
        RECT 102.940 108.870 103.780 109.150 ;
        RECT 105.290 109.260 106.450 109.750 ;
        RECT 110.790 109.700 111.990 109.800 ;
        RECT 102.880 108.640 103.840 108.870 ;
        RECT 104.170 108.640 105.130 108.870 ;
        RECT 100.990 107.480 102.830 108.480 ;
        RECT 100.990 106.910 102.730 107.480 ;
        RECT 103.120 107.320 103.640 108.640 ;
        RECT 103.890 107.480 104.120 108.480 ;
        RECT 104.390 107.320 104.910 108.640 ;
        RECT 105.290 108.480 106.110 109.260 ;
        RECT 109.605 108.670 139.000 108.855 ;
        RECT 105.180 107.910 106.460 108.480 ;
        RECT 109.605 108.465 139.170 108.670 ;
        RECT 138.490 108.190 139.170 108.465 ;
        RECT 105.180 107.480 115.760 107.910 ;
        RECT 136.890 107.730 137.610 107.930 ;
        RECT 102.880 107.090 103.840 107.320 ;
        RECT 104.170 107.090 105.130 107.320 ;
        RECT 105.290 107.050 115.760 107.480 ;
        RECT 130.090 107.285 130.540 107.675 ;
        RECT 132.750 107.500 137.750 107.730 ;
        RECT 105.290 106.950 106.460 107.050 ;
        RECT 101.010 106.890 102.730 106.910 ;
        RECT 98.690 106.475 99.650 106.705 ;
        RECT 99.980 106.475 100.940 106.705 ;
        RECT 101.700 106.480 102.390 106.890 ;
        RECT 105.280 106.830 106.460 106.950 ;
        RECT 101.690 105.860 102.390 106.480 ;
        RECT 98.690 105.055 99.650 105.285 ;
        RECT 99.980 105.260 100.940 105.285 ;
        RECT 101.700 105.260 102.390 105.860 ;
        RECT 105.270 105.690 106.460 106.830 ;
        RECT 112.650 106.470 113.570 106.540 ;
        RECT 108.550 106.240 113.570 106.470 ;
        RECT 105.290 105.380 106.460 105.690 ;
        RECT 107.990 106.190 108.380 106.210 ;
        RECT 99.980 105.090 103.780 105.260 ;
        RECT 99.980 105.055 100.940 105.090 ;
        RECT 96.560 104.850 98.500 104.950 ;
        RECT 96.560 102.950 98.640 104.850 ;
        RECT 96.700 102.850 98.640 102.950 ;
        RECT 92.810 101.900 93.510 102.520 ;
        RECT 94.260 102.515 95.220 102.745 ;
        RECT 95.550 102.515 96.510 102.745 ;
        RECT 89.370 100.470 89.910 101.730 ;
        RECT 92.810 101.310 93.500 101.900 ;
        RECT 94.260 101.310 95.220 101.335 ;
        RECT 91.420 101.140 95.220 101.310 ;
        RECT 91.420 100.860 92.260 101.140 ;
        RECT 94.260 101.105 95.220 101.140 ;
        RECT 95.550 101.105 96.510 101.335 ;
        RECT 92.470 100.900 94.190 100.920 ;
        RECT 90.070 100.630 91.030 100.860 ;
        RECT 91.360 100.630 92.320 100.860 ;
        RECT 89.370 99.470 90.020 100.470 ;
        RECT 89.370 98.940 89.910 99.470 ;
        RECT 90.290 99.310 90.810 100.630 ;
        RECT 91.080 99.470 91.310 100.470 ;
        RECT 91.560 99.310 92.080 100.630 ;
        RECT 92.470 100.470 94.210 100.900 ;
        RECT 92.370 99.470 94.210 100.470 ;
        RECT 90.070 99.080 91.030 99.310 ;
        RECT 91.360 99.080 92.320 99.310 ;
        RECT 89.370 98.820 89.920 98.940 ;
        RECT 92.470 98.900 94.210 99.470 ;
        RECT 92.470 98.880 94.190 98.900 ;
        RECT 89.370 97.680 89.930 98.820 ;
        RECT 92.810 98.470 93.500 98.880 ;
        RECT 94.490 98.695 95.010 101.105 ;
        RECT 95.270 98.900 95.500 100.900 ;
        RECT 95.820 98.695 96.340 101.105 ;
        RECT 96.700 100.900 98.500 102.850 ;
        RECT 98.860 102.645 99.380 105.055 ;
        RECT 99.700 102.850 99.930 104.850 ;
        RECT 100.190 102.645 100.710 105.055 ;
        RECT 101.010 104.850 102.730 104.870 ;
        RECT 100.990 104.420 102.730 104.850 ;
        RECT 102.940 104.810 103.780 105.090 ;
        RECT 102.880 104.580 103.840 104.810 ;
        RECT 104.170 104.580 105.130 104.810 ;
        RECT 105.290 104.720 106.630 105.380 ;
        RECT 107.990 105.230 108.410 106.190 ;
        RECT 112.650 106.120 113.570 106.240 ;
        RECT 107.990 104.900 108.380 105.230 ;
        RECT 108.550 105.180 109.650 105.380 ;
        RECT 108.550 104.950 113.570 105.180 ;
        RECT 100.990 103.420 102.830 104.420 ;
        RECT 100.990 102.850 102.730 103.420 ;
        RECT 103.120 103.260 103.640 104.580 ;
        RECT 103.890 103.420 104.120 104.420 ;
        RECT 104.390 103.260 104.910 104.580 ;
        RECT 105.290 104.420 106.460 104.720 ;
        RECT 105.180 103.420 106.460 104.420 ;
        RECT 102.880 103.030 103.840 103.260 ;
        RECT 104.170 103.030 105.130 103.260 ;
        RECT 105.290 102.890 106.460 103.420 ;
        RECT 101.010 102.830 102.730 102.850 ;
        RECT 98.690 102.415 99.650 102.645 ;
        RECT 99.980 102.415 100.940 102.645 ;
        RECT 101.700 102.420 102.390 102.830 ;
        RECT 105.280 102.770 106.460 102.890 ;
        RECT 101.690 101.800 102.390 102.420 ;
        RECT 98.690 100.995 99.650 101.225 ;
        RECT 99.980 101.200 100.940 101.225 ;
        RECT 101.700 101.200 102.390 101.800 ;
        RECT 105.270 101.630 106.460 102.770 ;
        RECT 107.990 103.940 108.410 104.900 ;
        RECT 108.550 104.710 109.650 104.950 ;
        RECT 107.990 103.610 108.380 103.940 ;
        RECT 112.650 103.890 113.570 103.960 ;
        RECT 108.560 103.660 113.570 103.890 ;
        RECT 107.990 102.650 108.410 103.610 ;
        RECT 112.650 103.540 113.570 103.660 ;
        RECT 107.990 102.580 108.380 102.650 ;
        RECT 108.630 102.610 109.570 102.680 ;
        RECT 99.980 101.030 103.780 101.200 ;
        RECT 99.980 100.995 100.940 101.030 ;
        RECT 96.560 100.790 98.500 100.900 ;
        RECT 96.560 98.900 98.640 100.790 ;
        RECT 96.700 98.790 98.640 98.900 ;
        RECT 92.810 97.850 93.510 98.470 ;
        RECT 94.260 98.465 95.220 98.695 ;
        RECT 95.550 98.465 96.510 98.695 ;
        RECT 89.370 96.420 89.910 97.680 ;
        RECT 92.810 97.260 93.500 97.850 ;
        RECT 94.260 97.260 95.220 97.285 ;
        RECT 91.420 97.090 95.220 97.260 ;
        RECT 91.420 96.810 92.260 97.090 ;
        RECT 94.260 97.055 95.220 97.090 ;
        RECT 95.550 97.055 96.510 97.285 ;
        RECT 92.470 96.850 94.190 96.870 ;
        RECT 90.070 96.580 91.030 96.810 ;
        RECT 91.360 96.580 92.320 96.810 ;
        RECT 89.370 95.420 90.020 96.420 ;
        RECT 89.370 94.890 89.910 95.420 ;
        RECT 90.290 95.260 90.810 96.580 ;
        RECT 91.080 95.420 91.310 96.420 ;
        RECT 91.560 95.260 92.080 96.580 ;
        RECT 92.470 96.420 94.210 96.850 ;
        RECT 92.370 95.420 94.210 96.420 ;
        RECT 90.070 95.030 91.030 95.260 ;
        RECT 91.360 95.030 92.320 95.260 ;
        RECT 89.370 94.770 89.920 94.890 ;
        RECT 92.470 94.850 94.210 95.420 ;
        RECT 92.470 94.830 94.190 94.850 ;
        RECT 89.370 93.630 89.930 94.770 ;
        RECT 92.810 94.420 93.500 94.830 ;
        RECT 94.490 94.645 95.010 97.055 ;
        RECT 95.270 94.850 95.500 96.850 ;
        RECT 95.820 94.645 96.340 97.055 ;
        RECT 96.700 96.850 98.500 98.790 ;
        RECT 98.860 98.585 99.380 100.995 ;
        RECT 99.700 98.790 99.930 100.790 ;
        RECT 100.190 98.585 100.710 100.995 ;
        RECT 101.010 100.790 102.730 100.810 ;
        RECT 100.990 100.360 102.730 100.790 ;
        RECT 102.940 100.750 103.780 101.030 ;
        RECT 102.880 100.520 103.840 100.750 ;
        RECT 104.170 100.520 105.130 100.750 ;
        RECT 100.990 99.360 102.830 100.360 ;
        RECT 100.990 98.790 102.730 99.360 ;
        RECT 103.120 99.200 103.640 100.520 ;
        RECT 103.890 99.360 104.120 100.360 ;
        RECT 104.390 99.200 104.910 100.520 ;
        RECT 105.290 100.360 106.460 101.630 ;
        RECT 107.100 102.320 108.380 102.580 ;
        RECT 108.560 102.600 113.520 102.610 ;
        RECT 108.560 102.380 113.570 102.600 ;
        RECT 108.570 102.370 113.570 102.380 ;
        RECT 107.100 102.060 108.410 102.320 ;
        RECT 108.630 102.290 109.570 102.370 ;
        RECT 113.730 102.060 114.010 106.210 ;
        RECT 115.180 105.400 115.760 107.050 ;
        RECT 120.080 106.750 121.600 106.850 ;
        RECT 127.280 106.750 129.000 106.890 ;
        RECT 117.030 106.520 122.030 106.750 ;
        RECT 124.030 106.520 129.030 106.750 ;
        RECT 116.640 105.510 116.870 106.470 ;
        RECT 120.080 106.330 121.600 106.520 ;
        RECT 122.220 106.470 123.080 106.480 ;
        RECT 127.280 106.470 129.000 106.520 ;
        RECT 130.120 106.500 130.510 107.285 ;
        RECT 129.280 106.470 130.870 106.500 ;
        RECT 122.190 105.510 123.090 106.470 ;
        RECT 123.640 105.510 123.870 106.470 ;
        RECT 129.190 105.510 130.870 106.470 ;
        RECT 122.200 105.490 123.090 105.510 ;
        RECT 129.210 105.490 130.870 105.510 ;
        RECT 122.220 105.470 123.090 105.490 ;
        RECT 117.030 105.430 122.030 105.460 ;
        RECT 117.010 104.730 122.060 105.430 ;
        RECT 117.010 104.540 122.050 104.730 ;
        RECT 117.030 104.520 122.030 104.540 ;
        RECT 116.640 103.510 116.870 104.470 ;
        RECT 117.990 103.460 119.510 103.550 ;
        RECT 117.030 103.230 122.030 103.460 ;
        RECT 117.990 103.030 119.510 103.230 ;
        RECT 107.100 101.610 108.460 102.060 ;
        RECT 113.640 101.610 114.010 102.060 ;
        RECT 107.100 101.360 108.410 101.610 ;
        RECT 107.100 101.220 108.380 101.360 ;
        RECT 112.640 101.310 113.570 101.370 ;
        RECT 105.180 99.360 106.460 100.360 ;
        RECT 102.880 98.970 103.840 99.200 ;
        RECT 104.170 98.970 105.130 99.200 ;
        RECT 105.290 98.830 106.460 99.360 ;
        RECT 101.010 98.770 102.730 98.790 ;
        RECT 98.690 98.355 99.650 98.585 ;
        RECT 99.980 98.355 100.940 98.585 ;
        RECT 101.700 98.360 102.390 98.770 ;
        RECT 105.280 98.710 106.460 98.830 ;
        RECT 101.690 97.740 102.390 98.360 ;
        RECT 98.690 96.935 99.650 97.165 ;
        RECT 99.980 97.140 100.940 97.165 ;
        RECT 101.700 97.140 102.390 97.740 ;
        RECT 105.270 97.570 106.460 98.710 ;
        RECT 99.980 96.970 103.780 97.140 ;
        RECT 99.980 96.935 100.940 96.970 ;
        RECT 96.560 96.730 98.500 96.850 ;
        RECT 96.560 94.850 98.640 96.730 ;
        RECT 96.700 94.730 98.640 94.850 ;
        RECT 92.810 93.800 93.510 94.420 ;
        RECT 94.260 94.415 95.220 94.645 ;
        RECT 95.550 94.415 96.510 94.645 ;
        RECT 89.370 92.370 89.910 93.630 ;
        RECT 92.810 93.210 93.500 93.800 ;
        RECT 94.260 93.210 95.220 93.235 ;
        RECT 91.420 93.040 95.220 93.210 ;
        RECT 91.420 92.760 92.260 93.040 ;
        RECT 94.260 93.005 95.220 93.040 ;
        RECT 95.550 93.005 96.510 93.235 ;
        RECT 92.470 92.800 94.190 92.820 ;
        RECT 90.070 92.530 91.030 92.760 ;
        RECT 91.360 92.530 92.320 92.760 ;
        RECT 89.370 91.370 90.020 92.370 ;
        RECT 89.370 90.840 89.910 91.370 ;
        RECT 90.290 91.210 90.810 92.530 ;
        RECT 91.080 91.370 91.310 92.370 ;
        RECT 91.560 91.210 92.080 92.530 ;
        RECT 92.470 92.370 94.210 92.800 ;
        RECT 92.370 91.370 94.210 92.370 ;
        RECT 90.070 90.980 91.030 91.210 ;
        RECT 91.360 90.980 92.320 91.210 ;
        RECT 89.370 90.720 89.920 90.840 ;
        RECT 92.470 90.800 94.210 91.370 ;
        RECT 92.470 90.780 94.190 90.800 ;
        RECT 89.370 89.580 89.930 90.720 ;
        RECT 92.810 90.370 93.500 90.780 ;
        RECT 94.490 90.595 95.010 93.005 ;
        RECT 95.270 90.800 95.500 92.800 ;
        RECT 95.820 90.595 96.340 93.005 ;
        RECT 96.700 92.800 98.500 94.730 ;
        RECT 98.860 94.525 99.380 96.935 ;
        RECT 99.700 94.730 99.930 96.730 ;
        RECT 100.190 94.525 100.710 96.935 ;
        RECT 101.010 96.730 102.730 96.750 ;
        RECT 100.990 96.300 102.730 96.730 ;
        RECT 102.940 96.690 103.780 96.970 ;
        RECT 102.880 96.460 103.840 96.690 ;
        RECT 104.170 96.460 105.130 96.690 ;
        RECT 100.990 95.300 102.830 96.300 ;
        RECT 100.990 94.730 102.730 95.300 ;
        RECT 103.120 95.140 103.640 96.460 ;
        RECT 103.890 95.300 104.120 96.300 ;
        RECT 104.390 95.140 104.910 96.460 ;
        RECT 105.290 96.300 106.460 97.570 ;
        RECT 107.990 101.030 108.380 101.220 ;
        RECT 108.560 101.080 113.570 101.310 ;
        RECT 107.990 100.070 108.410 101.030 ;
        RECT 112.640 100.990 113.570 101.080 ;
        RECT 107.990 99.740 108.380 100.070 ;
        RECT 108.620 100.030 109.570 100.120 ;
        RECT 108.560 100.020 113.520 100.030 ;
        RECT 108.560 99.800 113.570 100.020 ;
        RECT 108.570 99.790 113.570 99.800 ;
        RECT 108.620 99.740 109.570 99.790 ;
        RECT 107.990 98.780 108.410 99.740 ;
        RECT 107.990 98.450 108.380 98.780 ;
        RECT 112.650 98.740 113.570 98.810 ;
        RECT 108.560 98.510 113.570 98.740 ;
        RECT 108.570 98.500 113.570 98.510 ;
        RECT 107.990 97.490 108.410 98.450 ;
        RECT 112.650 98.440 113.570 98.500 ;
        RECT 107.990 97.160 108.380 97.490 ;
        RECT 108.620 97.440 109.570 97.520 ;
        RECT 108.560 97.210 113.570 97.440 ;
        RECT 105.180 95.300 106.460 96.300 ;
        RECT 107.270 96.190 108.420 97.160 ;
        RECT 108.620 97.120 109.570 97.210 ;
        RECT 113.730 96.200 114.010 101.610 ;
        RECT 122.190 102.560 122.470 104.500 ;
        RECT 122.770 104.490 123.090 105.470 ;
        RECT 124.030 105.440 129.030 105.460 ;
        RECT 124.000 104.550 129.050 105.440 ;
        RECT 129.760 105.150 130.870 105.490 ;
        RECT 124.030 104.520 129.030 104.550 ;
        RECT 122.770 104.470 123.830 104.490 ;
        RECT 122.770 103.510 123.870 104.470 ;
        RECT 129.190 103.510 129.420 104.470 ;
        RECT 122.770 103.490 123.830 103.510 ;
        RECT 122.190 101.530 122.580 102.560 ;
        RECT 122.770 101.040 123.090 103.490 ;
        RECT 124.030 103.230 129.030 103.460 ;
        RECT 124.990 102.900 126.720 103.230 ;
        RECT 129.760 102.700 130.080 105.150 ;
        RECT 132.260 104.300 132.590 107.500 ;
        RECT 136.890 107.360 137.610 107.500 ;
        RECT 137.960 107.450 138.290 107.510 ;
        RECT 137.170 106.940 137.790 107.000 ;
        RECT 137.955 106.990 138.290 107.450 ;
        RECT 132.750 106.710 137.790 106.940 ;
        RECT 137.170 106.500 137.790 106.710 ;
        RECT 131.930 103.410 132.590 104.300 ;
        RECT 129.750 101.070 130.080 102.700 ;
        RECT 120.090 100.750 121.610 100.880 ;
        RECT 117.030 100.520 122.030 100.750 ;
        RECT 116.640 99.510 116.870 100.470 ;
        RECT 120.090 100.360 121.610 100.520 ;
        RECT 122.760 100.510 123.100 101.040 ;
        RECT 127.150 100.750 129.040 100.870 ;
        RECT 124.030 100.520 129.040 100.750 ;
        RECT 122.190 99.460 123.100 100.510 ;
        RECT 123.640 99.510 123.870 100.470 ;
        RECT 127.150 100.250 129.040 100.520 ;
        RECT 129.760 100.490 130.080 101.070 ;
        RECT 129.220 100.470 130.080 100.490 ;
        RECT 129.190 99.510 130.080 100.470 ;
        RECT 129.220 99.480 130.080 99.510 ;
        RECT 132.260 102.410 132.590 103.410 ;
        RECT 136.940 103.230 137.660 103.350 ;
        RECT 132.750 103.000 137.750 103.230 ;
        RECT 136.940 102.780 137.660 103.000 ;
        RECT 137.960 102.950 138.290 106.990 ;
        RECT 137.955 102.490 138.290 102.950 ;
        RECT 132.750 102.410 137.750 102.440 ;
        RECT 132.260 102.330 137.750 102.410 ;
        RECT 137.960 102.330 138.290 102.490 ;
        RECT 132.260 102.210 138.290 102.330 ;
        RECT 132.260 102.160 132.920 102.210 ;
        RECT 117.030 99.440 122.030 99.460 ;
        RECT 117.000 99.230 122.030 99.440 ;
        RECT 117.000 98.750 121.820 99.230 ;
        RECT 117.000 98.550 122.030 98.750 ;
        RECT 117.030 98.520 122.030 98.550 ;
        RECT 116.640 97.510 116.870 98.470 ;
        RECT 118.020 97.460 119.540 97.560 ;
        RECT 122.180 97.490 122.530 98.530 ;
        RECT 122.760 98.510 123.100 99.460 ;
        RECT 124.030 99.440 129.030 99.460 ;
        RECT 124.010 98.550 129.060 99.440 ;
        RECT 124.030 98.520 129.030 98.550 ;
        RECT 122.760 98.470 123.840 98.510 ;
        RECT 117.030 97.230 122.030 97.460 ;
        RECT 118.020 97.040 119.540 97.230 ;
        RECT 122.760 97.070 123.870 98.470 ;
        RECT 129.190 97.510 129.420 98.470 ;
        RECT 132.260 97.980 132.590 102.160 ;
        RECT 136.970 101.980 138.290 102.210 ;
        RECT 136.900 98.730 137.720 98.900 ;
        RECT 132.750 98.500 137.750 98.730 ;
        RECT 136.900 98.400 137.720 98.500 ;
        RECT 137.960 98.450 138.290 101.980 ;
        RECT 132.970 97.940 134.770 98.090 ;
        RECT 137.955 97.990 138.290 98.450 ;
        RECT 137.120 97.940 137.780 97.960 ;
        RECT 132.750 97.710 137.780 97.940 ;
        RECT 124.030 97.230 129.030 97.460 ;
        RECT 132.970 97.270 134.770 97.710 ;
        RECT 137.120 97.490 137.780 97.710 ;
        RECT 124.990 96.890 126.720 97.230 ;
        RECT 112.650 96.150 113.580 96.200 ;
        RECT 108.570 95.920 113.580 96.150 ;
        RECT 112.650 95.880 113.580 95.920 ;
        RECT 138.610 95.860 139.000 108.190 ;
        RECT 139.480 97.520 140.120 108.010 ;
        RECT 140.660 97.600 141.050 108.060 ;
        RECT 141.780 107.730 142.730 107.810 ;
        RECT 141.750 107.500 146.750 107.730 ;
        RECT 141.240 106.990 141.570 107.480 ;
        RECT 141.780 107.370 142.730 107.500 ;
        RECT 141.240 106.940 142.530 106.990 ;
        RECT 141.240 106.920 146.750 106.940 ;
        RECT 146.940 106.920 147.270 107.530 ;
        RECT 141.240 106.710 147.270 106.920 ;
        RECT 141.240 106.700 142.530 106.710 ;
        RECT 141.240 98.040 141.570 106.700 ;
        RECT 146.430 106.660 147.270 106.710 ;
        RECT 141.770 103.230 142.710 103.420 ;
        RECT 141.750 103.000 146.750 103.230 ;
        RECT 141.770 102.950 142.710 103.000 ;
        RECT 141.740 102.440 142.710 102.540 ;
        RECT 141.740 102.210 146.750 102.440 ;
        RECT 141.740 101.820 142.710 102.210 ;
        RECT 141.710 98.730 142.710 98.880 ;
        RECT 141.710 98.500 146.750 98.730 ;
        RECT 141.710 98.420 142.710 98.500 ;
        RECT 146.940 98.100 147.270 106.660 ;
        RECT 141.240 97.960 142.540 98.040 ;
        RECT 141.290 97.940 142.540 97.960 ;
        RECT 146.520 98.010 147.270 98.100 ;
        RECT 146.520 97.940 147.240 98.010 ;
        RECT 141.290 97.730 147.240 97.940 ;
        RECT 141.290 97.710 146.750 97.730 ;
        RECT 141.290 97.690 142.540 97.710 ;
        RECT 147.460 96.910 148.020 108.520 ;
        RECT 102.880 94.910 103.840 95.140 ;
        RECT 104.170 94.910 105.130 95.140 ;
        RECT 105.290 94.970 106.460 95.300 ;
        RECT 138.330 95.060 139.560 95.860 ;
        RECT 147.460 95.060 148.030 96.910 ;
        RECT 105.290 94.770 111.920 94.970 ;
        RECT 101.010 94.710 102.730 94.730 ;
        RECT 98.690 94.295 99.650 94.525 ;
        RECT 99.980 94.295 100.940 94.525 ;
        RECT 101.700 94.300 102.390 94.710 ;
        RECT 105.280 94.650 111.920 94.770 ;
        RECT 101.690 93.680 102.390 94.300 ;
        RECT 98.690 92.875 99.650 93.105 ;
        RECT 99.980 93.080 100.940 93.105 ;
        RECT 101.700 93.080 102.390 93.680 ;
        RECT 105.270 94.280 111.920 94.650 ;
        RECT 114.070 94.340 116.495 94.460 ;
        RECT 123.450 94.400 148.030 95.060 ;
        RECT 123.450 94.340 124.230 94.400 ;
        RECT 105.270 94.130 106.350 94.280 ;
        RECT 106.900 94.130 111.920 94.280 ;
        RECT 114.045 94.250 116.495 94.340 ;
        RECT 105.270 93.510 106.330 94.130 ;
        RECT 106.900 94.105 111.900 94.130 ;
        RECT 114.045 94.110 115.045 94.250 ;
        RECT 115.710 94.230 116.495 94.250 ;
        RECT 115.710 94.200 116.090 94.230 ;
        RECT 99.980 92.910 103.780 93.080 ;
        RECT 99.980 92.875 100.940 92.910 ;
        RECT 96.560 92.670 98.500 92.800 ;
        RECT 96.560 90.800 98.640 92.670 ;
        RECT 96.700 90.670 98.640 90.800 ;
        RECT 92.810 89.750 93.510 90.370 ;
        RECT 94.260 90.365 95.220 90.595 ;
        RECT 95.550 90.365 96.510 90.595 ;
        RECT 89.370 88.320 89.910 89.580 ;
        RECT 92.810 89.160 93.500 89.750 ;
        RECT 94.260 89.160 95.220 89.185 ;
        RECT 91.420 88.990 95.220 89.160 ;
        RECT 91.420 88.710 92.260 88.990 ;
        RECT 94.260 88.955 95.220 88.990 ;
        RECT 95.550 88.955 96.510 89.185 ;
        RECT 92.470 88.750 94.190 88.770 ;
        RECT 90.070 88.480 91.030 88.710 ;
        RECT 91.360 88.480 92.320 88.710 ;
        RECT 89.370 87.320 90.020 88.320 ;
        RECT 89.370 86.790 89.910 87.320 ;
        RECT 90.290 87.160 90.810 88.480 ;
        RECT 91.080 87.320 91.310 88.320 ;
        RECT 91.560 87.160 92.080 88.480 ;
        RECT 92.470 88.320 94.210 88.750 ;
        RECT 92.370 87.320 94.210 88.320 ;
        RECT 90.070 86.930 91.030 87.160 ;
        RECT 91.360 86.930 92.320 87.160 ;
        RECT 89.370 86.670 89.920 86.790 ;
        RECT 92.470 86.750 94.210 87.320 ;
        RECT 92.470 86.730 94.190 86.750 ;
        RECT 89.370 85.530 89.930 86.670 ;
        RECT 92.810 86.320 93.500 86.730 ;
        RECT 94.490 86.545 95.010 88.955 ;
        RECT 95.270 86.750 95.500 88.750 ;
        RECT 95.820 86.545 96.340 88.955 ;
        RECT 96.700 88.750 98.500 90.670 ;
        RECT 98.860 90.465 99.380 92.875 ;
        RECT 99.700 90.670 99.930 92.670 ;
        RECT 100.190 90.465 100.710 92.875 ;
        RECT 101.010 92.670 102.730 92.690 ;
        RECT 100.990 92.240 102.730 92.670 ;
        RECT 102.940 92.630 103.780 92.910 ;
        RECT 102.880 92.400 103.840 92.630 ;
        RECT 104.170 92.400 105.130 92.630 ;
        RECT 100.990 91.240 102.830 92.240 ;
        RECT 100.990 90.670 102.730 91.240 ;
        RECT 103.120 91.080 103.640 92.400 ;
        RECT 103.890 91.240 104.120 92.240 ;
        RECT 104.390 91.080 104.910 92.400 ;
        RECT 105.290 92.240 106.330 93.510 ;
        RECT 106.510 93.800 106.740 94.055 ;
        RECT 112.060 93.800 112.290 94.055 ;
        RECT 106.510 93.460 112.290 93.800 ;
        RECT 106.510 93.095 106.740 93.460 ;
        RECT 112.060 93.095 112.290 93.460 ;
        RECT 113.560 93.550 113.850 94.080 ;
        RECT 116.265 94.060 116.495 94.230 ;
        RECT 116.705 94.140 124.230 94.340 ;
        RECT 116.705 94.110 124.205 94.140 ;
        RECT 124.800 94.070 148.030 94.400 ;
        RECT 115.245 93.550 115.635 94.060 ;
        RECT 116.265 93.550 116.500 94.060 ;
        RECT 124.410 93.850 124.640 94.060 ;
        RECT 123.630 93.600 124.640 93.850 ;
        RECT 123.630 93.550 124.610 93.600 ;
        RECT 106.900 93.030 111.900 93.045 ;
        RECT 106.870 92.820 111.900 93.030 ;
        RECT 106.870 92.680 111.905 92.820 ;
        RECT 113.560 92.790 115.960 93.550 ;
        RECT 116.265 93.510 124.610 93.550 ;
        RECT 116.265 93.320 124.205 93.510 ;
        RECT 124.800 93.230 125.290 94.070 ;
        RECT 124.390 93.020 125.290 93.230 ;
        RECT 112.170 92.680 115.960 92.790 ;
        RECT 106.870 92.550 115.960 92.680 ;
        RECT 111.690 92.490 112.390 92.550 ;
        RECT 113.560 92.540 115.960 92.550 ;
        RECT 105.180 91.240 106.330 92.240 ;
        RECT 115.790 91.890 115.960 92.540 ;
        RECT 116.760 92.670 125.290 93.020 ;
        RECT 116.760 92.270 122.380 92.670 ;
        RECT 122.740 91.980 123.650 92.300 ;
        RECT 116.700 91.965 123.670 91.980 ;
        RECT 115.790 91.590 116.510 91.890 ;
        RECT 116.700 91.735 123.710 91.965 ;
        RECT 116.700 91.640 123.670 91.735 ;
        RECT 102.880 90.850 103.840 91.080 ;
        RECT 104.170 90.850 105.130 91.080 ;
        RECT 105.290 90.710 106.330 91.240 ;
        RECT 101.010 90.650 102.730 90.670 ;
        RECT 98.690 90.235 99.650 90.465 ;
        RECT 99.980 90.235 100.940 90.465 ;
        RECT 101.700 90.240 102.390 90.650 ;
        RECT 105.280 90.590 106.330 90.710 ;
        RECT 116.210 90.670 116.510 91.590 ;
        RECT 101.690 89.620 102.390 90.240 ;
        RECT 98.690 88.815 99.650 89.045 ;
        RECT 99.980 89.020 100.940 89.045 ;
        RECT 101.700 89.020 102.390 89.620 ;
        RECT 105.270 89.450 106.330 90.590 ;
        RECT 99.980 88.850 103.780 89.020 ;
        RECT 99.980 88.815 100.940 88.850 ;
        RECT 96.560 88.610 98.500 88.750 ;
        RECT 96.560 86.750 98.640 88.610 ;
        RECT 96.700 86.610 98.640 86.750 ;
        RECT 92.810 85.700 93.510 86.320 ;
        RECT 94.260 86.315 95.220 86.545 ;
        RECT 95.550 86.315 96.510 86.545 ;
        RECT 89.370 84.270 89.910 85.530 ;
        RECT 92.810 85.110 93.500 85.700 ;
        RECT 94.260 85.110 95.220 85.135 ;
        RECT 91.420 84.940 95.220 85.110 ;
        RECT 91.420 84.660 92.260 84.940 ;
        RECT 94.260 84.905 95.220 84.940 ;
        RECT 95.550 84.905 96.510 85.135 ;
        RECT 92.470 84.700 94.190 84.720 ;
        RECT 90.070 84.430 91.030 84.660 ;
        RECT 91.360 84.430 92.320 84.660 ;
        RECT 89.370 83.270 90.020 84.270 ;
        RECT 89.370 82.740 89.910 83.270 ;
        RECT 90.290 83.110 90.810 84.430 ;
        RECT 91.080 83.270 91.310 84.270 ;
        RECT 91.560 83.110 92.080 84.430 ;
        RECT 92.470 84.270 94.210 84.700 ;
        RECT 92.370 83.270 94.210 84.270 ;
        RECT 90.070 82.880 91.030 83.110 ;
        RECT 91.360 82.880 92.320 83.110 ;
        RECT 89.370 82.620 89.920 82.740 ;
        RECT 92.470 82.700 94.210 83.270 ;
        RECT 92.470 82.680 94.190 82.700 ;
        RECT 89.370 81.480 89.930 82.620 ;
        RECT 92.810 82.270 93.500 82.680 ;
        RECT 94.490 82.495 95.010 84.905 ;
        RECT 95.270 82.700 95.500 84.700 ;
        RECT 95.820 82.495 96.340 84.905 ;
        RECT 96.700 84.700 98.500 86.610 ;
        RECT 98.860 86.405 99.380 88.815 ;
        RECT 99.700 86.610 99.930 88.610 ;
        RECT 100.190 86.405 100.710 88.815 ;
        RECT 101.010 88.610 102.730 88.630 ;
        RECT 100.990 88.180 102.730 88.610 ;
        RECT 102.940 88.570 103.780 88.850 ;
        RECT 102.880 88.340 103.840 88.570 ;
        RECT 104.170 88.340 105.130 88.570 ;
        RECT 100.990 87.180 102.830 88.180 ;
        RECT 100.990 86.610 102.730 87.180 ;
        RECT 103.120 87.020 103.640 88.340 ;
        RECT 103.890 87.180 104.120 88.180 ;
        RECT 104.390 87.020 104.910 88.340 ;
        RECT 105.290 88.180 106.330 89.450 ;
        RECT 105.180 87.830 106.330 88.180 ;
        RECT 105.180 87.180 106.450 87.830 ;
        RECT 102.880 86.790 103.840 87.020 ;
        RECT 104.170 86.790 105.130 87.020 ;
        RECT 105.290 86.650 106.450 87.180 ;
        RECT 107.120 87.120 111.960 87.180 ;
        RECT 107.100 86.890 112.100 87.120 ;
        RECT 101.010 86.590 102.730 86.610 ;
        RECT 98.690 86.175 99.650 86.405 ;
        RECT 99.980 86.175 100.940 86.405 ;
        RECT 101.700 86.180 102.390 86.590 ;
        RECT 105.280 86.530 106.450 86.650 ;
        RECT 101.690 85.560 102.390 86.180 ;
        RECT 98.690 84.755 99.650 84.985 ;
        RECT 99.980 84.960 100.940 84.985 ;
        RECT 101.700 84.960 102.390 85.560 ;
        RECT 105.270 85.390 106.450 86.530 ;
        RECT 99.980 84.790 103.780 84.960 ;
        RECT 99.980 84.755 100.940 84.790 ;
        RECT 96.560 84.550 98.500 84.700 ;
        RECT 96.560 82.700 98.640 84.550 ;
        RECT 96.700 82.550 98.640 82.700 ;
        RECT 92.810 81.650 93.510 82.270 ;
        RECT 94.260 82.265 95.220 82.495 ;
        RECT 95.550 82.265 96.510 82.495 ;
        RECT 89.370 80.220 89.910 81.480 ;
        RECT 92.810 81.060 93.500 81.650 ;
        RECT 94.260 81.060 95.220 81.085 ;
        RECT 91.420 80.890 95.220 81.060 ;
        RECT 91.420 80.610 92.260 80.890 ;
        RECT 94.260 80.855 95.220 80.890 ;
        RECT 95.550 80.855 96.510 81.085 ;
        RECT 92.470 80.650 94.190 80.670 ;
        RECT 90.070 80.380 91.030 80.610 ;
        RECT 91.360 80.380 92.320 80.610 ;
        RECT 89.370 79.220 90.020 80.220 ;
        RECT 89.370 78.690 89.910 79.220 ;
        RECT 90.290 79.060 90.810 80.380 ;
        RECT 91.080 79.220 91.310 80.220 ;
        RECT 91.560 79.060 92.080 80.380 ;
        RECT 92.470 80.220 94.210 80.650 ;
        RECT 92.370 79.220 94.210 80.220 ;
        RECT 90.070 78.830 91.030 79.060 ;
        RECT 91.360 78.830 92.320 79.060 ;
        RECT 89.370 78.570 89.920 78.690 ;
        RECT 92.470 78.650 94.210 79.220 ;
        RECT 92.470 78.630 94.190 78.650 ;
        RECT 89.370 77.430 89.930 78.570 ;
        RECT 92.810 78.220 93.500 78.630 ;
        RECT 94.490 78.445 95.010 80.855 ;
        RECT 95.270 78.650 95.500 80.650 ;
        RECT 95.820 78.445 96.340 80.855 ;
        RECT 96.700 80.650 98.500 82.550 ;
        RECT 98.860 82.345 99.380 84.755 ;
        RECT 99.700 82.550 99.930 84.550 ;
        RECT 100.190 82.345 100.710 84.755 ;
        RECT 101.010 84.550 102.730 84.570 ;
        RECT 100.990 84.120 102.730 84.550 ;
        RECT 102.940 84.510 103.780 84.790 ;
        RECT 102.880 84.280 103.840 84.510 ;
        RECT 104.170 84.280 105.130 84.510 ;
        RECT 100.990 83.120 102.830 84.120 ;
        RECT 100.990 82.550 102.730 83.120 ;
        RECT 103.120 82.960 103.640 84.280 ;
        RECT 103.890 83.120 104.120 84.120 ;
        RECT 104.390 82.960 104.910 84.280 ;
        RECT 105.290 84.120 106.450 85.390 ;
        RECT 105.180 83.120 106.450 84.120 ;
        RECT 102.880 82.730 103.840 82.960 ;
        RECT 104.170 82.730 105.130 82.960 ;
        RECT 105.290 82.590 106.450 83.120 ;
        RECT 101.010 82.530 102.730 82.550 ;
        RECT 98.690 82.115 99.650 82.345 ;
        RECT 99.980 82.115 100.940 82.345 ;
        RECT 101.700 82.120 102.390 82.530 ;
        RECT 105.280 82.470 106.450 82.590 ;
        RECT 101.690 81.500 102.390 82.120 ;
        RECT 98.690 80.695 99.650 80.925 ;
        RECT 99.980 80.900 100.940 80.925 ;
        RECT 101.700 80.900 102.390 81.500 ;
        RECT 105.270 81.330 106.450 82.470 ;
        RECT 99.980 80.730 103.780 80.900 ;
        RECT 99.980 80.695 100.940 80.730 ;
        RECT 96.560 80.490 98.500 80.650 ;
        RECT 96.560 78.650 98.640 80.490 ;
        RECT 96.700 78.490 98.640 78.650 ;
        RECT 92.810 77.600 93.510 78.220 ;
        RECT 94.260 78.215 95.220 78.445 ;
        RECT 95.550 78.215 96.510 78.445 ;
        RECT 89.370 76.170 89.910 77.430 ;
        RECT 92.810 77.010 93.500 77.600 ;
        RECT 94.260 77.010 95.220 77.035 ;
        RECT 91.420 76.840 95.220 77.010 ;
        RECT 91.420 76.560 92.260 76.840 ;
        RECT 94.260 76.805 95.220 76.840 ;
        RECT 95.550 76.805 96.510 77.035 ;
        RECT 92.470 76.600 94.190 76.620 ;
        RECT 90.070 76.330 91.030 76.560 ;
        RECT 91.360 76.330 92.320 76.560 ;
        RECT 89.370 75.170 90.020 76.170 ;
        RECT 89.370 74.640 89.910 75.170 ;
        RECT 90.290 75.010 90.810 76.330 ;
        RECT 91.080 75.170 91.310 76.170 ;
        RECT 91.560 75.010 92.080 76.330 ;
        RECT 92.470 76.170 94.210 76.600 ;
        RECT 92.370 75.170 94.210 76.170 ;
        RECT 90.070 74.780 91.030 75.010 ;
        RECT 91.360 74.780 92.320 75.010 ;
        RECT 89.370 74.520 89.920 74.640 ;
        RECT 92.470 74.600 94.210 75.170 ;
        RECT 92.470 74.580 94.190 74.600 ;
        RECT 89.370 73.380 89.930 74.520 ;
        RECT 92.810 74.170 93.500 74.580 ;
        RECT 94.490 74.395 95.010 76.805 ;
        RECT 95.270 74.600 95.500 76.600 ;
        RECT 95.820 74.395 96.340 76.805 ;
        RECT 96.700 76.600 98.500 78.490 ;
        RECT 98.860 78.285 99.380 80.695 ;
        RECT 99.700 78.490 99.930 80.490 ;
        RECT 100.190 78.285 100.710 80.695 ;
        RECT 101.010 80.490 102.730 80.510 ;
        RECT 100.990 80.060 102.730 80.490 ;
        RECT 102.940 80.450 103.780 80.730 ;
        RECT 102.880 80.220 103.840 80.450 ;
        RECT 104.170 80.220 105.130 80.450 ;
        RECT 100.990 79.060 102.830 80.060 ;
        RECT 100.990 78.490 102.730 79.060 ;
        RECT 103.120 78.900 103.640 80.220 ;
        RECT 103.890 79.060 104.120 80.060 ;
        RECT 104.390 78.900 104.910 80.220 ;
        RECT 105.290 80.060 106.450 81.330 ;
        RECT 105.180 79.060 106.450 80.060 ;
        RECT 102.880 78.670 103.840 78.900 ;
        RECT 104.170 78.670 105.130 78.900 ;
        RECT 105.290 78.530 106.450 79.060 ;
        RECT 101.010 78.470 102.730 78.490 ;
        RECT 98.690 78.055 99.650 78.285 ;
        RECT 99.980 78.055 100.940 78.285 ;
        RECT 101.700 78.060 102.390 78.470 ;
        RECT 105.280 78.410 106.450 78.530 ;
        RECT 101.690 77.440 102.390 78.060 ;
        RECT 98.690 76.635 99.650 76.865 ;
        RECT 99.980 76.840 100.940 76.865 ;
        RECT 101.700 76.840 102.390 77.440 ;
        RECT 105.270 77.270 106.450 78.410 ;
        RECT 99.980 76.670 103.780 76.840 ;
        RECT 99.980 76.635 100.940 76.670 ;
        RECT 96.560 76.430 98.500 76.600 ;
        RECT 96.560 74.600 98.640 76.430 ;
        RECT 96.700 74.430 98.640 74.600 ;
        RECT 92.810 73.550 93.510 74.170 ;
        RECT 94.260 74.165 95.220 74.395 ;
        RECT 95.550 74.165 96.510 74.395 ;
        RECT 89.370 72.120 89.910 73.380 ;
        RECT 92.810 72.960 93.500 73.550 ;
        RECT 94.260 72.960 95.220 72.985 ;
        RECT 91.420 72.790 95.220 72.960 ;
        RECT 91.420 72.510 92.260 72.790 ;
        RECT 94.260 72.755 95.220 72.790 ;
        RECT 95.550 72.755 96.510 72.985 ;
        RECT 92.470 72.550 94.190 72.570 ;
        RECT 90.070 72.280 91.030 72.510 ;
        RECT 91.360 72.280 92.320 72.510 ;
        RECT 89.370 71.120 90.020 72.120 ;
        RECT 89.370 70.590 89.910 71.120 ;
        RECT 90.290 70.960 90.810 72.280 ;
        RECT 91.080 71.120 91.310 72.120 ;
        RECT 91.560 70.960 92.080 72.280 ;
        RECT 92.470 72.120 94.210 72.550 ;
        RECT 92.370 71.120 94.210 72.120 ;
        RECT 90.070 70.730 91.030 70.960 ;
        RECT 91.360 70.730 92.320 70.960 ;
        RECT 89.370 70.470 89.920 70.590 ;
        RECT 92.470 70.550 94.210 71.120 ;
        RECT 92.470 70.530 94.190 70.550 ;
        RECT 89.370 69.330 89.930 70.470 ;
        RECT 92.810 70.120 93.500 70.530 ;
        RECT 94.490 70.345 95.010 72.755 ;
        RECT 95.270 70.550 95.500 72.550 ;
        RECT 95.820 70.345 96.340 72.755 ;
        RECT 96.700 72.550 98.500 74.430 ;
        RECT 98.860 74.225 99.380 76.635 ;
        RECT 99.700 74.430 99.930 76.430 ;
        RECT 100.190 74.225 100.710 76.635 ;
        RECT 101.010 76.430 102.730 76.450 ;
        RECT 100.990 76.000 102.730 76.430 ;
        RECT 102.940 76.390 103.780 76.670 ;
        RECT 102.880 76.160 103.840 76.390 ;
        RECT 104.170 76.160 105.130 76.390 ;
        RECT 100.990 75.000 102.830 76.000 ;
        RECT 100.990 74.430 102.730 75.000 ;
        RECT 103.120 74.840 103.640 76.160 ;
        RECT 103.890 75.000 104.120 76.000 ;
        RECT 104.390 74.840 104.910 76.160 ;
        RECT 105.290 76.000 106.450 77.270 ;
        RECT 105.180 75.000 106.450 76.000 ;
        RECT 102.880 74.610 103.840 74.840 ;
        RECT 104.170 74.610 105.130 74.840 ;
        RECT 105.290 74.470 106.450 75.000 ;
        RECT 101.010 74.410 102.730 74.430 ;
        RECT 98.690 73.995 99.650 74.225 ;
        RECT 99.980 73.995 100.940 74.225 ;
        RECT 101.700 74.000 102.390 74.410 ;
        RECT 105.280 74.350 106.450 74.470 ;
        RECT 101.690 73.380 102.390 74.000 ;
        RECT 98.690 72.575 99.650 72.805 ;
        RECT 99.980 72.780 100.940 72.805 ;
        RECT 101.700 72.780 102.390 73.380 ;
        RECT 105.270 73.210 106.450 74.350 ;
        RECT 99.980 72.610 103.780 72.780 ;
        RECT 99.980 72.575 100.940 72.610 ;
        RECT 96.560 72.370 98.500 72.550 ;
        RECT 96.560 70.550 98.640 72.370 ;
        RECT 96.700 70.370 98.640 70.550 ;
        RECT 92.810 69.500 93.510 70.120 ;
        RECT 94.260 70.115 95.220 70.345 ;
        RECT 95.550 70.115 96.510 70.345 ;
        RECT 89.370 68.070 89.910 69.330 ;
        RECT 92.810 68.910 93.500 69.500 ;
        RECT 94.260 68.910 95.220 68.935 ;
        RECT 91.420 68.740 95.220 68.910 ;
        RECT 91.420 68.460 92.260 68.740 ;
        RECT 94.260 68.705 95.220 68.740 ;
        RECT 95.550 68.705 96.510 68.935 ;
        RECT 92.470 68.500 94.190 68.520 ;
        RECT 90.070 68.230 91.030 68.460 ;
        RECT 91.360 68.230 92.320 68.460 ;
        RECT 89.370 67.070 90.020 68.070 ;
        RECT 89.370 66.540 89.910 67.070 ;
        RECT 90.290 66.910 90.810 68.230 ;
        RECT 91.080 67.070 91.310 68.070 ;
        RECT 91.560 66.910 92.080 68.230 ;
        RECT 92.470 68.070 94.210 68.500 ;
        RECT 92.370 67.070 94.210 68.070 ;
        RECT 90.070 66.680 91.030 66.910 ;
        RECT 91.360 66.680 92.320 66.910 ;
        RECT 89.370 66.420 89.920 66.540 ;
        RECT 92.470 66.500 94.210 67.070 ;
        RECT 92.470 66.480 94.190 66.500 ;
        RECT 89.370 65.280 89.930 66.420 ;
        RECT 92.810 66.070 93.500 66.480 ;
        RECT 94.490 66.295 95.010 68.705 ;
        RECT 95.270 66.500 95.500 68.500 ;
        RECT 95.820 66.295 96.340 68.705 ;
        RECT 96.700 68.500 98.500 70.370 ;
        RECT 98.860 70.165 99.380 72.575 ;
        RECT 99.700 70.370 99.930 72.370 ;
        RECT 100.190 70.165 100.710 72.575 ;
        RECT 101.010 72.370 102.730 72.390 ;
        RECT 100.990 71.940 102.730 72.370 ;
        RECT 102.940 72.330 103.780 72.610 ;
        RECT 102.880 72.100 103.840 72.330 ;
        RECT 104.170 72.100 105.130 72.330 ;
        RECT 100.990 70.940 102.830 71.940 ;
        RECT 100.990 70.370 102.730 70.940 ;
        RECT 103.120 70.780 103.640 72.100 ;
        RECT 103.890 70.940 104.120 71.940 ;
        RECT 104.390 70.780 104.910 72.100 ;
        RECT 105.290 71.940 106.450 73.210 ;
        RECT 106.620 86.840 106.930 86.890 ;
        RECT 107.120 86.840 111.960 86.890 ;
        RECT 106.620 86.380 106.940 86.840 ;
        RECT 110.810 86.410 112.020 86.420 ;
        RECT 106.620 86.050 106.930 86.380 ;
        RECT 110.800 86.330 112.020 86.410 ;
        RECT 107.100 86.100 112.100 86.330 ;
        RECT 110.800 86.050 112.020 86.100 ;
        RECT 106.620 85.590 106.940 86.050 ;
        RECT 110.810 86.020 112.020 86.050 ;
        RECT 112.260 86.000 113.130 90.460 ;
        RECT 116.220 89.280 116.510 90.670 ;
        RECT 116.680 89.820 123.720 91.180 ;
        RECT 116.710 89.805 123.710 89.820 ;
        RECT 122.740 89.310 123.650 89.330 ;
        RECT 116.700 89.245 123.670 89.310 ;
        RECT 123.900 89.280 124.190 91.710 ;
        RECT 116.700 89.015 123.710 89.245 ;
        RECT 116.700 88.970 123.670 89.015 ;
        RECT 122.740 88.770 123.650 88.970 ;
        RECT 124.390 87.830 125.290 92.670 ;
        RECT 141.710 92.570 147.190 92.830 ;
        RECT 141.710 92.240 147.290 92.570 ;
        RECT 141.710 92.150 142.380 92.240 ;
        RECT 141.690 90.190 142.380 92.150 ;
        RECT 146.820 90.540 147.290 92.240 ;
        RECT 146.820 90.190 147.320 90.540 ;
        RECT 141.690 89.600 147.320 90.190 ;
        RECT 141.830 89.560 147.320 89.600 ;
        RECT 141.710 88.760 147.360 89.270 ;
        RECT 112.260 85.950 113.110 86.000 ;
        RECT 106.620 85.260 106.930 85.590 ;
        RECT 107.290 85.540 108.570 85.630 ;
        RECT 112.260 85.590 112.590 85.950 ;
        RECT 113.820 85.780 115.000 87.280 ;
        RECT 120.790 87.000 125.290 87.830 ;
        RECT 144.700 88.010 145.240 88.760 ;
        RECT 146.750 88.010 147.340 88.760 ;
        RECT 144.700 87.700 147.340 88.010 ;
        RECT 144.870 87.660 147.340 87.700 ;
        RECT 115.320 86.940 116.580 87.000 ;
        RECT 115.160 86.710 120.160 86.940 ;
        RECT 115.320 86.650 116.580 86.710 ;
        RECT 118.910 86.150 120.030 86.170 ;
        RECT 115.160 85.920 120.160 86.150 ;
        RECT 118.910 85.820 120.030 85.920 ;
        RECT 114.040 85.770 115.000 85.780 ;
        RECT 107.100 85.310 112.100 85.540 ;
        RECT 106.620 84.800 106.940 85.260 ;
        RECT 107.290 85.230 108.570 85.310 ;
        RECT 112.280 85.260 112.590 85.590 ;
        RECT 112.260 84.800 112.590 85.260 ;
        RECT 106.620 84.470 106.930 84.800 ;
        RECT 110.800 84.750 112.020 84.790 ;
        RECT 107.100 84.520 112.100 84.750 ;
        RECT 106.620 84.010 106.940 84.470 ;
        RECT 110.800 84.430 112.020 84.520 ;
        RECT 112.280 84.470 112.590 84.800 ;
        RECT 106.620 83.680 106.930 84.010 ;
        RECT 107.290 83.960 108.570 84.030 ;
        RECT 112.260 84.010 112.590 84.470 ;
        RECT 107.100 83.730 112.100 83.960 ;
        RECT 106.620 83.220 106.940 83.680 ;
        RECT 107.290 83.630 108.570 83.730 ;
        RECT 112.280 83.680 112.590 84.010 ;
        RECT 112.260 83.220 112.590 83.680 ;
        RECT 106.620 82.890 106.930 83.220 ;
        RECT 110.800 83.170 112.040 83.220 ;
        RECT 107.100 82.940 112.100 83.170 ;
        RECT 106.620 82.430 106.940 82.890 ;
        RECT 110.800 82.870 112.040 82.940 ;
        RECT 112.280 82.890 112.590 83.220 ;
        RECT 106.620 82.100 106.930 82.430 ;
        RECT 107.250 82.380 108.580 82.440 ;
        RECT 112.260 82.430 112.590 82.890 ;
        RECT 107.100 82.150 112.100 82.380 ;
        RECT 106.620 81.640 106.940 82.100 ;
        RECT 107.250 82.040 108.580 82.150 ;
        RECT 112.280 82.100 112.590 82.430 ;
        RECT 112.260 81.640 112.590 82.100 ;
        RECT 106.620 81.310 106.930 81.640 ;
        RECT 110.790 81.590 111.940 81.610 ;
        RECT 107.100 81.360 112.100 81.590 ;
        RECT 106.620 80.850 106.940 81.310 ;
        RECT 110.790 81.250 111.940 81.360 ;
        RECT 112.280 81.310 112.590 81.640 ;
        RECT 106.620 80.520 106.930 80.850 ;
        RECT 107.300 80.800 108.560 80.910 ;
        RECT 112.260 80.850 112.590 81.310 ;
        RECT 107.100 80.570 112.100 80.800 ;
        RECT 106.620 80.060 106.940 80.520 ;
        RECT 107.300 80.460 108.560 80.570 ;
        RECT 112.280 80.520 112.590 80.850 ;
        RECT 112.260 80.060 112.590 80.520 ;
        RECT 106.620 79.730 106.930 80.060 ;
        RECT 110.800 80.010 111.920 80.050 ;
        RECT 107.100 79.780 112.100 80.010 ;
        RECT 106.620 79.270 106.940 79.730 ;
        RECT 110.800 79.710 111.920 79.780 ;
        RECT 112.280 79.730 112.590 80.060 ;
        RECT 112.260 79.270 112.590 79.730 ;
        RECT 106.620 78.940 106.930 79.270 ;
        RECT 107.310 79.220 108.570 79.260 ;
        RECT 107.100 78.990 112.100 79.220 ;
        RECT 106.620 78.480 106.940 78.940 ;
        RECT 107.310 78.910 108.570 78.990 ;
        RECT 112.280 78.940 112.590 79.270 ;
        RECT 112.260 78.480 112.590 78.940 ;
        RECT 106.620 78.150 106.930 78.480 ;
        RECT 110.800 78.430 111.950 78.460 ;
        RECT 107.100 78.200 112.100 78.430 ;
        RECT 106.620 77.690 106.940 78.150 ;
        RECT 110.800 78.110 111.950 78.200 ;
        RECT 112.280 78.150 112.590 78.480 ;
        RECT 106.620 77.360 106.930 77.690 ;
        RECT 107.300 77.640 108.570 77.700 ;
        RECT 112.260 77.690 112.590 78.150 ;
        RECT 107.100 77.410 112.100 77.640 ;
        RECT 106.620 76.900 106.940 77.360 ;
        RECT 107.300 77.340 108.570 77.410 ;
        RECT 112.280 77.360 112.590 77.690 ;
        RECT 112.260 76.900 112.590 77.360 ;
        RECT 106.620 76.570 106.930 76.900 ;
        RECT 110.800 76.850 111.990 76.890 ;
        RECT 107.100 76.620 112.100 76.850 ;
        RECT 106.620 76.110 106.940 76.570 ;
        RECT 110.800 76.530 111.990 76.620 ;
        RECT 112.280 76.570 112.590 76.900 ;
        RECT 112.260 76.110 112.590 76.570 ;
        RECT 106.620 75.780 106.930 76.110 ;
        RECT 107.290 76.060 108.570 76.100 ;
        RECT 107.100 75.830 112.100 76.060 ;
        RECT 106.620 75.320 106.940 75.780 ;
        RECT 107.290 75.740 108.570 75.830 ;
        RECT 112.280 75.780 112.590 76.110 ;
        RECT 112.260 75.320 112.590 75.780 ;
        RECT 114.700 75.760 115.000 85.770 ;
        RECT 115.310 85.360 116.570 85.440 ;
        RECT 115.160 85.130 120.160 85.360 ;
        RECT 115.310 85.080 116.570 85.130 ;
        RECT 118.920 84.570 120.040 84.600 ;
        RECT 115.160 84.340 120.160 84.570 ;
        RECT 118.920 84.260 120.040 84.340 ;
        RECT 115.320 83.780 116.580 83.850 ;
        RECT 115.160 83.550 120.160 83.780 ;
        RECT 115.320 83.490 116.580 83.550 ;
        RECT 118.920 82.990 120.010 83.020 ;
        RECT 115.160 82.760 120.160 82.990 ;
        RECT 118.920 82.660 120.010 82.760 ;
        RECT 115.320 82.200 116.580 82.250 ;
        RECT 115.160 81.970 120.160 82.200 ;
        RECT 115.320 81.890 116.580 81.970 ;
        RECT 118.920 81.410 120.080 81.480 ;
        RECT 115.160 81.180 120.160 81.410 ;
        RECT 118.920 81.060 120.080 81.180 ;
        RECT 115.320 80.620 116.580 80.650 ;
        RECT 115.160 80.390 120.160 80.620 ;
        RECT 115.320 80.310 116.580 80.390 ;
        RECT 118.920 79.830 120.070 79.930 ;
        RECT 115.160 79.600 120.160 79.830 ;
        RECT 118.920 79.470 120.070 79.600 ;
        RECT 115.320 79.040 116.580 79.120 ;
        RECT 115.160 78.810 120.160 79.040 ;
        RECT 115.320 78.780 116.580 78.810 ;
        RECT 118.920 78.250 120.020 78.330 ;
        RECT 115.160 78.020 120.160 78.250 ;
        RECT 118.920 77.910 120.020 78.020 ;
        RECT 115.320 77.460 116.580 77.490 ;
        RECT 115.160 77.230 120.160 77.460 ;
        RECT 115.320 77.150 116.580 77.230 ;
        RECT 118.920 76.670 120.000 76.760 ;
        RECT 115.160 76.440 120.160 76.670 ;
        RECT 118.920 76.330 120.000 76.440 ;
        RECT 115.320 75.880 116.580 75.910 ;
        RECT 115.160 75.650 120.160 75.880 ;
        RECT 120.350 75.780 120.650 86.730 ;
        RECT 115.320 75.560 116.580 75.650 ;
        RECT 106.620 74.990 106.930 75.320 ;
        RECT 110.800 75.270 111.950 75.300 ;
        RECT 107.100 75.040 112.100 75.270 ;
        RECT 106.620 74.530 106.940 74.990 ;
        RECT 110.800 74.950 111.950 75.040 ;
        RECT 112.280 74.990 112.590 75.320 ;
        RECT 112.260 74.530 112.590 74.990 ;
        RECT 106.620 74.200 106.930 74.530 ;
        RECT 107.300 74.480 108.570 74.510 ;
        RECT 107.100 74.250 112.100 74.480 ;
        RECT 106.620 73.740 106.940 74.200 ;
        RECT 107.300 74.120 108.570 74.250 ;
        RECT 112.280 74.200 112.590 74.530 ;
        RECT 110.810 73.740 111.990 73.790 ;
        RECT 112.260 73.740 112.590 74.200 ;
        RECT 120.790 74.190 121.210 87.000 ;
        RECT 141.690 86.330 147.380 86.840 ;
        RECT 141.690 85.810 145.170 86.330 ;
        RECT 144.660 85.020 145.170 85.810 ;
        RECT 144.670 84.460 145.170 85.020 ;
        RECT 141.710 84.430 145.170 84.460 ;
        RECT 146.850 85.810 147.380 86.330 ;
        RECT 146.850 84.770 147.320 85.810 ;
        RECT 146.850 84.430 147.400 84.770 ;
        RECT 122.440 82.380 124.340 84.310 ;
        RECT 141.710 83.740 147.400 84.430 ;
        RECT 106.620 73.410 106.930 73.740 ;
        RECT 110.800 73.690 111.990 73.740 ;
        RECT 107.100 73.460 112.100 73.690 ;
        RECT 106.620 72.950 106.940 73.410 ;
        RECT 110.800 73.400 111.990 73.460 ;
        RECT 112.280 73.410 112.590 73.740 ;
        RECT 110.810 73.370 111.990 73.400 ;
        RECT 112.260 72.950 112.590 73.410 ;
        RECT 106.620 72.620 106.930 72.950 ;
        RECT 107.300 72.900 108.580 72.930 ;
        RECT 107.100 72.670 112.100 72.900 ;
        RECT 106.620 72.160 106.940 72.620 ;
        RECT 107.300 72.570 108.580 72.670 ;
        RECT 112.280 72.620 112.590 72.950 ;
        RECT 112.260 72.160 112.590 72.620 ;
        RECT 106.620 72.050 106.930 72.160 ;
        RECT 110.790 72.110 111.990 72.140 ;
        RECT 105.180 71.340 106.450 71.940 ;
        RECT 107.100 71.880 112.100 72.110 ;
        RECT 112.280 72.060 112.590 72.160 ;
        RECT 110.790 71.780 111.990 71.880 ;
        RECT 105.180 70.940 105.830 71.340 ;
        RECT 102.880 70.550 103.840 70.780 ;
        RECT 104.170 70.550 105.130 70.780 ;
        RECT 105.290 70.410 105.830 70.940 ;
        RECT 101.010 70.350 102.730 70.370 ;
        RECT 98.690 69.935 99.650 70.165 ;
        RECT 99.980 69.935 100.940 70.165 ;
        RECT 101.700 69.940 102.390 70.350 ;
        RECT 105.280 70.290 105.830 70.410 ;
        RECT 101.690 69.320 102.390 69.940 ;
        RECT 98.690 68.515 99.650 68.745 ;
        RECT 99.980 68.720 100.940 68.745 ;
        RECT 101.700 68.720 102.390 69.320 ;
        RECT 105.270 69.150 105.830 70.290 ;
        RECT 122.720 70.010 123.660 82.380 ;
        RECT 141.730 81.340 147.420 81.940 ;
        RECT 141.730 80.900 147.440 81.340 ;
        RECT 146.580 79.560 147.440 80.900 ;
        RECT 141.790 78.530 147.480 79.560 ;
        RECT 146.580 77.150 147.440 78.530 ;
        RECT 141.850 76.110 147.540 77.150 ;
        RECT 141.770 74.490 147.460 74.680 ;
        RECT 141.770 73.990 147.550 74.490 ;
        RECT 141.770 73.640 144.700 73.990 ;
        RECT 144.200 72.600 144.700 73.640 ;
        RECT 146.850 72.600 147.550 73.990 ;
        RECT 144.200 72.290 147.550 72.600 ;
        RECT 144.200 72.040 147.540 72.290 ;
        RECT 99.980 68.550 103.780 68.720 ;
        RECT 99.980 68.515 100.940 68.550 ;
        RECT 96.560 68.310 98.500 68.500 ;
        RECT 96.560 66.500 98.640 68.310 ;
        RECT 96.700 66.310 98.640 66.500 ;
        RECT 92.810 65.450 93.510 66.070 ;
        RECT 94.260 66.065 95.220 66.295 ;
        RECT 95.550 66.065 96.510 66.295 ;
        RECT 89.370 64.020 89.910 65.280 ;
        RECT 92.810 64.860 93.500 65.450 ;
        RECT 94.260 64.860 95.220 64.885 ;
        RECT 91.420 64.690 95.220 64.860 ;
        RECT 91.420 64.410 92.260 64.690 ;
        RECT 94.260 64.655 95.220 64.690 ;
        RECT 95.550 64.655 96.510 64.885 ;
        RECT 92.470 64.450 94.190 64.470 ;
        RECT 90.070 64.180 91.030 64.410 ;
        RECT 91.360 64.180 92.320 64.410 ;
        RECT 89.370 63.020 90.020 64.020 ;
        RECT 89.370 62.490 89.910 63.020 ;
        RECT 90.290 62.860 90.810 64.180 ;
        RECT 91.080 63.020 91.310 64.020 ;
        RECT 91.560 62.860 92.080 64.180 ;
        RECT 92.470 64.020 94.210 64.450 ;
        RECT 92.370 63.020 94.210 64.020 ;
        RECT 90.070 62.630 91.030 62.860 ;
        RECT 91.360 62.630 92.320 62.860 ;
        RECT 89.370 62.370 89.920 62.490 ;
        RECT 92.470 62.450 94.210 63.020 ;
        RECT 92.470 62.430 94.190 62.450 ;
        RECT 89.370 61.230 89.930 62.370 ;
        RECT 92.810 62.020 93.500 62.430 ;
        RECT 94.490 62.245 95.010 64.655 ;
        RECT 95.270 62.450 95.500 64.450 ;
        RECT 95.820 62.245 96.340 64.655 ;
        RECT 96.700 64.450 98.500 66.310 ;
        RECT 98.860 66.105 99.380 68.515 ;
        RECT 99.700 66.310 99.930 68.310 ;
        RECT 100.190 66.105 100.710 68.515 ;
        RECT 101.010 68.310 102.730 68.330 ;
        RECT 100.990 67.880 102.730 68.310 ;
        RECT 102.940 68.270 103.780 68.550 ;
        RECT 102.880 68.040 103.840 68.270 ;
        RECT 104.170 68.040 105.130 68.270 ;
        RECT 100.990 66.880 102.830 67.880 ;
        RECT 100.990 66.310 102.730 66.880 ;
        RECT 103.120 66.720 103.640 68.040 ;
        RECT 103.890 66.880 104.120 67.880 ;
        RECT 104.390 66.720 104.910 68.040 ;
        RECT 105.290 67.880 105.830 69.150 ;
        RECT 107.815 69.070 123.660 70.010 ;
        RECT 105.180 66.880 105.830 67.880 ;
        RECT 102.880 66.490 103.840 66.720 ;
        RECT 104.170 66.490 105.130 66.720 ;
        RECT 105.290 66.350 105.830 66.880 ;
        RECT 101.010 66.290 102.730 66.310 ;
        RECT 98.690 65.875 99.650 66.105 ;
        RECT 99.980 65.875 100.940 66.105 ;
        RECT 101.700 65.880 102.390 66.290 ;
        RECT 105.280 66.230 105.830 66.350 ;
        RECT 101.690 65.260 102.390 65.880 ;
        RECT 98.690 64.455 99.650 64.685 ;
        RECT 99.980 64.660 100.940 64.685 ;
        RECT 101.700 64.660 102.390 65.260 ;
        RECT 105.270 65.090 105.830 66.230 ;
        RECT 99.980 64.490 103.780 64.660 ;
        RECT 99.980 64.455 100.940 64.490 ;
        RECT 96.560 64.250 98.500 64.450 ;
        RECT 96.560 62.450 98.640 64.250 ;
        RECT 96.700 62.250 98.640 62.450 ;
        RECT 92.810 61.400 93.510 62.020 ;
        RECT 94.260 62.015 95.220 62.245 ;
        RECT 95.550 62.015 96.510 62.245 ;
        RECT 96.700 61.650 98.500 62.250 ;
        RECT 98.860 62.045 99.380 64.455 ;
        RECT 99.700 62.250 99.930 64.250 ;
        RECT 100.190 62.045 100.710 64.455 ;
        RECT 101.010 64.250 102.730 64.270 ;
        RECT 100.990 63.820 102.730 64.250 ;
        RECT 102.940 64.210 103.780 64.490 ;
        RECT 102.880 63.980 103.840 64.210 ;
        RECT 104.170 63.980 105.130 64.210 ;
        RECT 100.990 62.820 102.830 63.820 ;
        RECT 100.990 62.250 102.730 62.820 ;
        RECT 103.120 62.660 103.640 63.980 ;
        RECT 103.890 62.820 104.120 63.820 ;
        RECT 104.390 62.660 104.910 63.980 ;
        RECT 105.290 63.820 105.830 65.090 ;
        RECT 105.180 62.820 105.830 63.820 ;
        RECT 102.880 62.430 103.840 62.660 ;
        RECT 104.170 62.430 105.130 62.660 ;
        RECT 105.290 62.290 105.830 62.820 ;
        RECT 101.010 62.230 102.730 62.250 ;
        RECT 98.690 61.815 99.650 62.045 ;
        RECT 99.980 61.815 100.940 62.045 ;
        RECT 101.700 61.820 102.390 62.230 ;
        RECT 105.280 62.170 105.830 62.290 ;
        RECT 89.370 59.970 89.910 61.230 ;
        RECT 92.810 60.810 93.500 61.400 ;
        RECT 94.260 60.810 95.220 60.835 ;
        RECT 91.420 60.640 95.220 60.810 ;
        RECT 91.420 60.360 92.260 60.640 ;
        RECT 94.260 60.605 95.220 60.640 ;
        RECT 95.550 60.605 96.510 60.835 ;
        RECT 92.470 60.400 94.190 60.420 ;
        RECT 90.070 60.130 91.030 60.360 ;
        RECT 91.360 60.130 92.320 60.360 ;
        RECT 89.370 58.970 90.020 59.970 ;
        RECT 89.370 58.440 89.910 58.970 ;
        RECT 90.290 58.810 90.810 60.130 ;
        RECT 91.080 58.970 91.310 59.970 ;
        RECT 91.560 58.810 92.080 60.130 ;
        RECT 92.470 59.970 94.210 60.400 ;
        RECT 92.370 58.970 94.210 59.970 ;
        RECT 90.070 58.580 91.030 58.810 ;
        RECT 91.360 58.580 92.320 58.810 ;
        RECT 89.370 58.320 89.920 58.440 ;
        RECT 92.470 58.400 94.210 58.970 ;
        RECT 92.470 58.380 94.190 58.400 ;
        RECT 89.370 57.180 89.930 58.320 ;
        RECT 92.810 57.970 93.500 58.380 ;
        RECT 94.490 58.195 95.010 60.605 ;
        RECT 95.270 58.400 95.500 60.400 ;
        RECT 95.820 58.195 96.340 60.605 ;
        RECT 96.700 60.400 98.505 61.650 ;
        RECT 101.690 61.200 102.390 61.820 ;
        RECT 96.560 59.710 98.505 60.400 ;
        RECT 101.695 60.900 102.385 61.200 ;
        RECT 105.270 61.030 105.830 62.170 ;
        RECT 98.690 59.915 99.650 60.145 ;
        RECT 99.980 60.120 100.940 60.145 ;
        RECT 101.695 60.120 102.390 60.900 ;
        RECT 99.980 59.950 103.780 60.120 ;
        RECT 99.980 59.915 100.940 59.950 ;
        RECT 96.560 58.400 98.640 59.710 ;
        RECT 92.810 57.350 93.510 57.970 ;
        RECT 94.260 57.965 95.220 58.195 ;
        RECT 95.550 57.965 96.510 58.195 ;
        RECT 96.700 57.710 98.640 58.400 ;
        RECT 89.370 55.920 89.910 57.180 ;
        RECT 92.810 56.760 93.500 57.350 ;
        RECT 94.260 56.760 95.220 56.785 ;
        RECT 91.420 56.590 95.220 56.760 ;
        RECT 91.420 56.310 92.260 56.590 ;
        RECT 94.260 56.555 95.220 56.590 ;
        RECT 95.550 56.555 96.510 56.785 ;
        RECT 96.700 56.620 98.505 57.710 ;
        RECT 98.860 57.505 99.380 59.915 ;
        RECT 99.700 57.710 99.930 59.710 ;
        RECT 100.190 57.505 100.710 59.915 ;
        RECT 101.010 59.710 102.730 59.730 ;
        RECT 100.990 59.280 102.730 59.710 ;
        RECT 102.940 59.670 103.780 59.950 ;
        RECT 102.880 59.440 103.840 59.670 ;
        RECT 104.170 59.440 105.130 59.670 ;
        RECT 100.990 58.280 102.830 59.280 ;
        RECT 100.990 57.710 102.730 58.280 ;
        RECT 103.120 58.120 103.640 59.440 ;
        RECT 103.890 58.280 104.120 59.280 ;
        RECT 104.390 58.120 104.910 59.440 ;
        RECT 105.290 59.280 105.830 61.030 ;
        RECT 105.180 58.280 105.830 59.280 ;
        RECT 102.880 57.890 103.840 58.120 ;
        RECT 104.170 57.890 105.130 58.120 ;
        RECT 105.290 57.750 105.830 58.280 ;
        RECT 101.010 57.690 102.730 57.710 ;
        RECT 98.690 57.275 99.650 57.505 ;
        RECT 99.980 57.275 100.940 57.505 ;
        RECT 101.415 57.150 102.390 57.690 ;
        RECT 105.280 57.630 105.830 57.750 ;
        RECT 101.400 56.660 102.390 57.150 ;
        RECT 92.470 56.350 94.190 56.370 ;
        RECT 90.070 56.080 91.030 56.310 ;
        RECT 91.360 56.080 92.320 56.310 ;
        RECT 89.370 54.920 90.020 55.920 ;
        RECT 89.370 54.390 89.910 54.920 ;
        RECT 90.290 54.760 90.810 56.080 ;
        RECT 91.080 54.920 91.310 55.920 ;
        RECT 91.560 54.760 92.080 56.080 ;
        RECT 92.470 55.920 94.210 56.350 ;
        RECT 92.370 54.920 94.210 55.920 ;
        RECT 90.070 54.530 91.030 54.760 ;
        RECT 91.360 54.530 92.320 54.760 ;
        RECT 89.370 54.270 89.920 54.390 ;
        RECT 92.470 54.350 94.210 54.920 ;
        RECT 92.470 54.330 94.190 54.350 ;
        RECT 89.370 53.130 89.930 54.270 ;
        RECT 92.810 53.920 93.500 54.330 ;
        RECT 94.490 54.145 95.010 56.555 ;
        RECT 95.270 54.350 95.500 56.350 ;
        RECT 95.820 54.145 96.340 56.555 ;
        RECT 96.700 56.490 98.500 56.620 ;
        RECT 96.700 56.350 97.600 56.490 ;
        RECT 96.560 54.350 97.600 56.350 ;
        RECT 92.810 53.300 93.510 53.920 ;
        RECT 94.260 53.915 95.220 54.145 ;
        RECT 95.550 53.915 96.510 54.145 ;
        RECT 89.370 51.870 89.910 53.130 ;
        RECT 92.810 52.710 93.500 53.300 ;
        RECT 94.260 52.710 95.220 52.735 ;
        RECT 91.420 52.540 95.220 52.710 ;
        RECT 91.420 52.260 92.260 52.540 ;
        RECT 94.260 52.505 95.220 52.540 ;
        RECT 95.550 52.505 96.510 52.735 ;
        RECT 92.470 52.300 94.190 52.320 ;
        RECT 90.070 52.030 91.030 52.260 ;
        RECT 91.360 52.030 92.320 52.260 ;
        RECT 89.370 50.870 90.020 51.870 ;
        RECT 89.370 50.340 89.910 50.870 ;
        RECT 90.290 50.710 90.810 52.030 ;
        RECT 91.080 50.870 91.310 51.870 ;
        RECT 91.560 50.710 92.080 52.030 ;
        RECT 92.470 51.870 94.210 52.300 ;
        RECT 92.370 50.870 94.210 51.870 ;
        RECT 90.070 50.480 91.030 50.710 ;
        RECT 91.360 50.480 92.320 50.710 ;
        RECT 89.370 50.220 89.920 50.340 ;
        RECT 92.470 50.300 94.210 50.870 ;
        RECT 92.470 50.280 94.190 50.300 ;
        RECT 89.370 49.080 89.930 50.220 ;
        RECT 92.810 49.870 93.500 50.280 ;
        RECT 94.490 50.095 95.010 52.505 ;
        RECT 95.270 50.300 95.500 52.300 ;
        RECT 95.820 50.095 96.340 52.505 ;
        RECT 96.700 52.300 97.600 54.350 ;
        RECT 96.560 50.300 97.600 52.300 ;
        RECT 101.400 53.070 102.380 56.660 ;
        RECT 105.270 56.490 105.830 57.630 ;
        RECT 105.965 53.070 106.945 54.410 ;
        RECT 101.400 52.090 106.950 53.070 ;
        RECT 92.810 49.250 93.510 49.870 ;
        RECT 94.260 49.865 95.220 50.095 ;
        RECT 95.550 49.865 96.510 50.095 ;
        RECT 89.370 47.820 89.910 49.080 ;
        RECT 92.810 48.660 93.500 49.250 ;
        RECT 94.260 48.660 95.220 48.685 ;
        RECT 91.420 48.490 95.220 48.660 ;
        RECT 91.420 48.210 92.260 48.490 ;
        RECT 94.260 48.455 95.220 48.490 ;
        RECT 95.550 48.455 96.510 48.685 ;
        RECT 92.470 48.250 94.190 48.270 ;
        RECT 90.070 47.980 91.030 48.210 ;
        RECT 91.360 47.980 92.320 48.210 ;
        RECT 89.370 46.820 90.020 47.820 ;
        RECT 89.370 46.290 89.910 46.820 ;
        RECT 90.290 46.660 90.810 47.980 ;
        RECT 91.080 46.820 91.310 47.820 ;
        RECT 91.560 46.660 92.080 47.980 ;
        RECT 92.470 47.820 94.210 48.250 ;
        RECT 92.370 46.820 94.210 47.820 ;
        RECT 90.070 46.430 91.030 46.660 ;
        RECT 91.360 46.430 92.320 46.660 ;
        RECT 89.370 46.170 89.920 46.290 ;
        RECT 92.470 46.250 94.210 46.820 ;
        RECT 92.470 46.230 94.190 46.250 ;
        RECT 89.370 45.030 89.930 46.170 ;
        RECT 92.810 45.820 93.500 46.230 ;
        RECT 94.490 46.045 95.010 48.455 ;
        RECT 95.270 46.250 95.500 48.250 ;
        RECT 95.820 46.045 96.340 48.455 ;
        RECT 96.700 48.250 97.600 50.300 ;
        RECT 96.560 46.250 97.600 48.250 ;
        RECT 107.835 47.010 108.740 69.070 ;
        RECT 92.810 45.200 93.510 45.820 ;
        RECT 94.260 45.815 95.220 46.045 ;
        RECT 95.550 45.815 96.510 46.045 ;
        RECT 89.370 43.770 89.910 45.030 ;
        RECT 92.810 44.610 93.500 45.200 ;
        RECT 94.260 44.610 95.220 44.635 ;
        RECT 91.420 44.440 95.220 44.610 ;
        RECT 91.420 44.160 92.260 44.440 ;
        RECT 94.260 44.405 95.220 44.440 ;
        RECT 95.550 44.405 96.510 44.635 ;
        RECT 92.470 44.200 94.190 44.220 ;
        RECT 90.070 43.930 91.030 44.160 ;
        RECT 91.360 43.930 92.320 44.160 ;
        RECT 89.370 42.770 90.020 43.770 ;
        RECT 89.370 42.240 89.910 42.770 ;
        RECT 90.290 42.610 90.810 43.930 ;
        RECT 91.080 42.770 91.310 43.770 ;
        RECT 91.560 42.610 92.080 43.930 ;
        RECT 92.470 43.770 94.210 44.200 ;
        RECT 92.370 42.770 94.210 43.770 ;
        RECT 90.070 42.380 91.030 42.610 ;
        RECT 91.360 42.380 92.320 42.610 ;
        RECT 89.370 42.120 89.920 42.240 ;
        RECT 92.470 42.200 94.210 42.770 ;
        RECT 92.470 42.180 94.190 42.200 ;
        RECT 89.370 40.980 89.930 42.120 ;
        RECT 92.810 41.770 93.500 42.180 ;
        RECT 94.490 41.995 95.010 44.405 ;
        RECT 95.270 42.200 95.500 44.200 ;
        RECT 95.820 41.995 96.340 44.405 ;
        RECT 96.700 44.200 97.600 46.250 ;
        RECT 96.560 42.200 97.600 44.200 ;
        RECT 92.810 41.150 93.510 41.770 ;
        RECT 94.260 41.765 95.220 41.995 ;
        RECT 95.550 41.765 96.510 41.995 ;
        RECT 89.370 39.720 89.910 40.980 ;
        RECT 92.810 40.560 93.500 41.150 ;
        RECT 94.260 40.560 95.220 40.585 ;
        RECT 91.420 40.390 95.220 40.560 ;
        RECT 91.420 40.110 92.260 40.390 ;
        RECT 94.260 40.355 95.220 40.390 ;
        RECT 95.550 40.355 96.510 40.585 ;
        RECT 92.470 40.150 94.190 40.170 ;
        RECT 90.070 39.880 91.030 40.110 ;
        RECT 91.360 39.880 92.320 40.110 ;
        RECT 89.370 38.720 90.020 39.720 ;
        RECT 89.370 38.190 89.910 38.720 ;
        RECT 90.290 38.560 90.810 39.880 ;
        RECT 91.080 38.720 91.310 39.720 ;
        RECT 91.560 38.560 92.080 39.880 ;
        RECT 92.470 39.720 94.210 40.150 ;
        RECT 92.370 38.720 94.210 39.720 ;
        RECT 90.070 38.330 91.030 38.560 ;
        RECT 91.360 38.330 92.320 38.560 ;
        RECT 89.370 38.070 89.920 38.190 ;
        RECT 92.470 38.150 94.210 38.720 ;
        RECT 92.470 38.130 94.190 38.150 ;
        RECT 89.370 36.930 89.930 38.070 ;
        RECT 92.810 37.720 93.500 38.130 ;
        RECT 94.490 37.945 95.010 40.355 ;
        RECT 95.270 38.150 95.500 40.150 ;
        RECT 95.820 37.945 96.340 40.355 ;
        RECT 96.700 40.150 97.600 42.200 ;
        RECT 96.560 38.150 97.600 40.150 ;
        RECT 92.810 37.100 93.510 37.720 ;
        RECT 94.260 37.715 95.220 37.945 ;
        RECT 95.550 37.715 96.510 37.945 ;
        RECT 89.370 35.670 89.910 36.930 ;
        RECT 92.810 36.510 93.500 37.100 ;
        RECT 94.260 36.510 95.220 36.535 ;
        RECT 91.420 36.340 95.220 36.510 ;
        RECT 91.420 36.060 92.260 36.340 ;
        RECT 94.260 36.305 95.220 36.340 ;
        RECT 95.550 36.305 96.510 36.535 ;
        RECT 92.470 36.100 94.190 36.120 ;
        RECT 90.070 35.830 91.030 36.060 ;
        RECT 91.360 35.830 92.320 36.060 ;
        RECT 89.370 34.670 90.020 35.670 ;
        RECT 89.370 34.140 89.910 34.670 ;
        RECT 90.290 34.510 90.810 35.830 ;
        RECT 91.080 34.670 91.310 35.670 ;
        RECT 91.560 34.510 92.080 35.830 ;
        RECT 92.470 35.670 94.210 36.100 ;
        RECT 92.370 34.670 94.210 35.670 ;
        RECT 90.070 34.280 91.030 34.510 ;
        RECT 91.360 34.280 92.320 34.510 ;
        RECT 89.370 34.020 89.920 34.140 ;
        RECT 92.470 34.100 94.210 34.670 ;
        RECT 92.470 34.080 94.190 34.100 ;
        RECT 89.370 32.880 89.930 34.020 ;
        RECT 92.810 33.670 93.500 34.080 ;
        RECT 94.490 33.895 95.010 36.305 ;
        RECT 95.270 34.100 95.500 36.100 ;
        RECT 95.820 33.895 96.340 36.305 ;
        RECT 96.700 36.100 97.600 38.150 ;
        RECT 96.560 34.100 97.600 36.100 ;
        RECT 92.810 33.050 93.510 33.670 ;
        RECT 94.260 33.665 95.220 33.895 ;
        RECT 95.550 33.665 96.510 33.895 ;
        RECT 89.370 31.620 89.910 32.880 ;
        RECT 92.810 32.460 93.500 33.050 ;
        RECT 94.260 32.460 95.220 32.485 ;
        RECT 91.420 32.290 95.220 32.460 ;
        RECT 91.420 32.010 92.260 32.290 ;
        RECT 94.260 32.255 95.220 32.290 ;
        RECT 95.550 32.255 96.510 32.485 ;
        RECT 92.470 32.050 94.190 32.070 ;
        RECT 90.070 31.780 91.030 32.010 ;
        RECT 91.360 31.780 92.320 32.010 ;
        RECT 89.370 30.620 90.020 31.620 ;
        RECT 89.370 30.090 89.910 30.620 ;
        RECT 90.290 30.460 90.810 31.780 ;
        RECT 91.080 30.620 91.310 31.620 ;
        RECT 91.560 30.460 92.080 31.780 ;
        RECT 92.470 31.620 94.210 32.050 ;
        RECT 92.370 30.620 94.210 31.620 ;
        RECT 90.070 30.230 91.030 30.460 ;
        RECT 91.360 30.230 92.320 30.460 ;
        RECT 89.370 29.970 89.920 30.090 ;
        RECT 92.470 30.050 94.210 30.620 ;
        RECT 92.470 30.030 94.190 30.050 ;
        RECT 89.370 28.830 89.930 29.970 ;
        RECT 92.810 29.620 93.500 30.030 ;
        RECT 94.490 29.845 95.010 32.255 ;
        RECT 95.270 30.050 95.500 32.050 ;
        RECT 95.820 29.845 96.340 32.255 ;
        RECT 96.700 32.050 97.600 34.100 ;
        RECT 96.560 30.050 97.600 32.050 ;
        RECT 92.810 29.000 93.510 29.620 ;
        RECT 94.260 29.615 95.220 29.845 ;
        RECT 95.550 29.615 96.510 29.845 ;
        RECT 89.370 27.535 89.910 28.830 ;
        RECT 92.810 28.375 93.500 29.000 ;
        RECT 94.260 28.375 95.220 28.400 ;
        RECT 91.420 28.205 95.220 28.375 ;
        RECT 91.420 27.925 92.260 28.205 ;
        RECT 94.260 28.170 95.220 28.205 ;
        RECT 95.550 28.170 96.510 28.400 ;
        RECT 92.470 27.965 94.190 27.985 ;
        RECT 90.070 27.695 91.030 27.925 ;
        RECT 91.360 27.695 92.320 27.925 ;
        RECT 89.370 26.535 90.020 27.535 ;
        RECT 89.370 26.005 89.910 26.535 ;
        RECT 90.290 26.375 90.810 27.695 ;
        RECT 91.080 26.535 91.310 27.535 ;
        RECT 91.560 26.375 92.080 27.695 ;
        RECT 92.470 27.535 94.210 27.965 ;
        RECT 92.370 26.535 94.210 27.535 ;
        RECT 90.070 26.145 91.030 26.375 ;
        RECT 91.360 26.145 92.320 26.375 ;
        RECT 89.370 25.885 89.920 26.005 ;
        RECT 92.470 25.965 94.210 26.535 ;
        RECT 92.470 25.945 94.190 25.965 ;
        RECT 89.370 24.745 89.930 25.885 ;
        RECT 92.810 25.535 93.500 25.945 ;
        RECT 94.490 25.760 95.010 28.170 ;
        RECT 95.270 25.965 95.500 27.965 ;
        RECT 95.820 25.760 96.340 28.170 ;
        RECT 96.700 27.965 97.600 30.050 ;
        RECT 96.560 25.965 97.600 27.965 ;
        RECT 92.810 24.915 93.510 25.535 ;
        RECT 94.260 25.530 95.220 25.760 ;
        RECT 95.550 25.530 96.510 25.760 ;
        RECT 89.370 23.410 89.910 24.745 ;
        RECT 92.810 24.250 93.500 24.915 ;
        RECT 94.260 24.250 95.220 24.275 ;
        RECT 91.420 24.080 95.220 24.250 ;
        RECT 91.420 23.800 92.260 24.080 ;
        RECT 94.260 24.045 95.220 24.080 ;
        RECT 95.550 24.045 96.510 24.275 ;
        RECT 92.470 23.840 94.190 23.860 ;
        RECT 90.070 23.570 91.030 23.800 ;
        RECT 91.360 23.570 92.320 23.800 ;
        RECT 89.370 22.410 90.020 23.410 ;
        RECT 89.370 21.880 89.910 22.410 ;
        RECT 90.290 22.250 90.810 23.570 ;
        RECT 91.080 22.410 91.310 23.410 ;
        RECT 91.560 22.250 92.080 23.570 ;
        RECT 92.470 23.410 94.210 23.840 ;
        RECT 92.370 22.410 94.210 23.410 ;
        RECT 90.070 22.020 91.030 22.250 ;
        RECT 91.360 22.020 92.320 22.250 ;
        RECT 89.370 21.760 89.920 21.880 ;
        RECT 92.470 21.840 94.210 22.410 ;
        RECT 92.470 21.820 94.190 21.840 ;
        RECT 89.370 20.620 89.930 21.760 ;
        RECT 92.810 21.410 93.500 21.820 ;
        RECT 94.490 21.635 95.010 24.045 ;
        RECT 95.270 21.840 95.500 23.840 ;
        RECT 95.820 21.635 96.340 24.045 ;
        RECT 96.700 23.840 97.600 25.965 ;
        RECT 96.560 21.840 97.600 23.840 ;
        RECT 92.810 20.790 93.510 21.410 ;
        RECT 94.260 21.405 95.220 21.635 ;
        RECT 95.550 21.405 96.510 21.635 ;
        RECT 89.370 18.855 89.910 20.620 ;
        RECT 92.815 20.475 93.505 20.790 ;
        RECT 92.810 19.985 93.505 20.475 ;
        RECT 92.810 19.695 93.500 19.985 ;
        RECT 94.260 19.695 95.220 19.720 ;
        RECT 91.420 19.525 95.220 19.695 ;
        RECT 91.420 19.245 92.260 19.525 ;
        RECT 94.260 19.490 95.220 19.525 ;
        RECT 95.550 19.490 96.510 19.720 ;
        RECT 92.470 19.285 94.190 19.305 ;
        RECT 90.070 19.015 91.030 19.245 ;
        RECT 91.360 19.015 92.320 19.245 ;
        RECT 89.370 17.855 90.020 18.855 ;
        RECT 89.370 17.325 89.910 17.855 ;
        RECT 90.290 17.695 90.810 19.015 ;
        RECT 91.080 17.855 91.310 18.855 ;
        RECT 91.560 17.695 92.080 19.015 ;
        RECT 92.470 18.855 94.210 19.285 ;
        RECT 92.370 17.855 94.210 18.855 ;
        RECT 90.070 17.465 91.030 17.695 ;
        RECT 91.360 17.465 92.320 17.695 ;
        RECT 89.370 17.205 89.920 17.325 ;
        RECT 92.470 17.285 94.210 17.855 ;
        RECT 92.470 17.265 94.190 17.285 ;
        RECT 89.370 16.065 89.930 17.205 ;
        RECT 92.660 15.290 93.670 17.265 ;
        RECT 94.490 17.080 95.010 19.490 ;
        RECT 95.270 17.285 95.500 19.285 ;
        RECT 95.820 17.080 96.340 19.490 ;
        RECT 96.700 19.285 97.600 21.840 ;
        RECT 96.560 17.285 97.600 19.285 ;
        RECT 94.260 16.850 95.220 17.080 ;
        RECT 95.550 16.850 96.510 17.080 ;
        RECT 96.700 16.455 97.600 17.285 ;
        RECT 96.705 16.275 97.600 16.455 ;
        RECT 96.700 16.065 97.600 16.275 ;
        RECT 98.315 46.105 108.740 47.010 ;
        RECT 98.315 15.305 99.220 46.105 ;
        RECT 95.100 15.290 99.220 15.305 ;
        RECT 92.660 14.420 99.220 15.290 ;
        RECT 95.100 14.400 99.220 14.420 ;
      LAYER via ;
        RECT 90.120 151.970 92.150 153.560 ;
        RECT 96.910 148.300 98.670 150.440 ;
        RECT 87.920 143.230 88.630 146.590 ;
        RECT 92.895 145.815 93.445 146.580 ;
        RECT 89.420 144.850 89.870 145.320 ;
        RECT 90.290 144.020 90.810 144.500 ;
        RECT 89.480 142.400 89.860 143.060 ;
        RECT 101.765 145.960 102.325 146.550 ;
        RECT 95.820 144.820 96.340 145.320 ;
        RECT 96.620 144.030 96.890 144.480 ;
        RECT 98.310 144.030 98.580 144.480 ;
        RECT 98.860 144.820 99.380 145.320 ;
        RECT 89.420 140.850 89.870 141.320 ;
        RECT 90.290 140.020 90.810 140.500 ;
        RECT 104.390 144.020 104.910 144.500 ;
        RECT 105.330 144.850 105.780 145.320 ;
        RECT 107.400 143.720 108.240 144.650 ;
        RECT 112.740 144.140 113.510 144.400 ;
        RECT 105.340 142.420 105.690 143.060 ;
        RECT 106.150 142.730 106.540 143.210 ;
        RECT 95.820 140.820 96.340 141.320 ;
        RECT 96.620 140.030 96.890 140.480 ;
        RECT 98.310 139.970 98.580 140.420 ;
        RECT 98.860 140.760 99.380 141.260 ;
        RECT 89.420 136.750 89.870 137.220 ;
        RECT 90.290 135.920 90.810 136.400 ;
        RECT 104.390 139.960 104.910 140.440 ;
        RECT 105.330 140.790 105.780 141.260 ;
        RECT 95.820 136.720 96.340 137.220 ;
        RECT 96.620 135.930 96.890 136.380 ;
        RECT 98.310 135.910 98.580 136.360 ;
        RECT 98.860 136.700 99.380 137.200 ;
        RECT 89.420 132.700 89.870 133.170 ;
        RECT 90.290 131.870 90.810 132.350 ;
        RECT 104.390 135.900 104.910 136.380 ;
        RECT 105.330 136.730 105.780 137.200 ;
        RECT 108.640 142.750 109.530 143.230 ;
        RECT 112.690 141.530 113.510 141.830 ;
        RECT 108.710 140.270 109.510 140.540 ;
        RECT 120.180 144.390 121.510 144.700 ;
        RECT 127.280 144.430 129.000 144.710 ;
        RECT 117.200 142.620 118.350 143.180 ;
        RECT 118.080 141.060 119.410 141.370 ;
        RECT 108.180 139.580 108.440 139.940 ;
        RECT 113.710 139.570 113.970 139.930 ;
        RECT 112.690 138.940 113.530 139.240 ;
        RECT 108.680 137.710 109.520 137.980 ;
        RECT 112.720 136.420 113.520 136.680 ;
        RECT 108.670 135.100 109.520 135.380 ;
        RECT 107.370 134.170 108.000 134.980 ;
        RECT 127.580 142.670 128.730 143.230 ;
        RECT 129.940 143.320 130.720 144.230 ;
        RECT 136.980 145.360 137.550 145.720 ;
        RECT 137.230 144.480 137.730 144.840 ;
        RECT 132.300 143.740 132.570 144.220 ;
        RECT 122.220 139.510 122.490 140.350 ;
        RECT 125.110 140.900 126.630 141.240 ;
        RECT 132.050 141.380 132.540 142.150 ;
        RECT 129.780 139.480 130.050 140.390 ;
        RECT 120.180 138.340 121.510 138.650 ;
        RECT 127.180 138.410 129.010 138.740 ;
        RECT 137.980 143.720 138.250 144.200 ;
        RECT 137.000 140.760 137.570 141.220 ;
        RECT 117.250 136.610 118.400 137.170 ;
        RECT 122.210 135.490 122.470 136.330 ;
        RECT 127.580 136.660 128.730 137.220 ;
        RECT 118.070 135.050 119.400 135.360 ;
        RECT 122.870 135.190 123.720 136.160 ;
        RECT 136.970 136.390 137.660 136.780 ;
        RECT 138.650 145.390 138.940 145.670 ;
        RECT 138.650 140.860 138.940 141.140 ;
        RECT 138.660 136.370 138.950 136.650 ;
        RECT 125.100 134.860 126.600 135.310 ;
        RECT 133.200 135.300 134.620 135.880 ;
        RECT 137.170 135.460 137.750 135.820 ;
        RECT 95.820 132.670 96.340 133.170 ;
        RECT 96.620 131.880 96.890 132.330 ;
        RECT 98.310 131.850 98.580 132.300 ;
        RECT 98.860 132.640 99.380 133.140 ;
        RECT 89.420 128.650 89.870 129.120 ;
        RECT 90.290 127.820 90.810 128.300 ;
        RECT 112.700 133.820 113.510 134.080 ;
        RECT 139.580 144.610 140.050 144.980 ;
        RECT 139.580 139.920 140.040 140.480 ;
        RECT 139.540 135.530 140.030 135.990 ;
        RECT 140.710 145.400 141.000 145.680 ;
        RECT 140.700 140.950 140.990 141.230 ;
        RECT 141.780 145.360 142.680 145.660 ;
        RECT 141.280 143.720 141.550 144.200 ;
        RECT 146.970 143.750 147.240 144.230 ;
        RECT 141.850 140.940 142.640 141.290 ;
        RECT 141.800 139.870 142.540 140.330 ;
        RECT 141.820 136.440 142.610 136.750 ;
        RECT 147.540 145.080 147.940 145.850 ;
        RECT 104.390 131.840 104.910 132.320 ;
        RECT 105.330 132.670 105.780 133.140 ;
        RECT 106.590 131.430 107.880 131.690 ;
        RECT 95.820 128.620 96.340 129.120 ;
        RECT 96.620 127.830 96.890 128.280 ;
        RECT 98.310 127.790 98.580 128.240 ;
        RECT 98.860 128.580 99.380 129.080 ;
        RECT 89.420 124.600 89.870 125.070 ;
        RECT 90.290 123.770 90.810 124.250 ;
        RECT 122.790 129.740 123.600 130.160 ;
        RECT 104.390 127.780 104.910 128.260 ;
        RECT 105.330 128.610 105.780 129.080 ;
        RECT 112.400 127.380 113.010 128.200 ;
        RECT 95.820 124.570 96.340 125.070 ;
        RECT 96.620 123.780 96.890 124.230 ;
        RECT 98.310 123.730 98.580 124.180 ;
        RECT 98.860 124.520 99.380 125.020 ;
        RECT 89.420 120.550 89.870 121.020 ;
        RECT 90.290 119.720 90.810 120.200 ;
        RECT 104.390 123.720 104.910 124.200 ;
        RECT 105.330 124.550 105.780 125.020 ;
        RECT 95.820 120.520 96.340 121.020 ;
        RECT 96.620 119.730 96.890 120.180 ;
        RECT 98.310 119.670 98.580 120.120 ;
        RECT 98.860 120.460 99.380 120.960 ;
        RECT 89.420 116.500 89.870 116.970 ;
        RECT 90.290 115.670 90.810 116.150 ;
        RECT 104.390 119.660 104.910 120.140 ;
        RECT 105.330 120.490 105.780 120.960 ;
        RECT 106.100 118.170 106.410 118.900 ;
        RECT 95.820 116.470 96.340 116.970 ;
        RECT 96.620 115.680 96.890 116.130 ;
        RECT 98.310 115.610 98.580 116.060 ;
        RECT 98.860 116.400 99.380 116.900 ;
        RECT 89.420 112.450 89.870 112.920 ;
        RECT 90.290 111.620 90.810 112.100 ;
        RECT 104.390 115.600 104.910 116.080 ;
        RECT 105.330 116.430 105.780 116.900 ;
        RECT 95.820 112.420 96.340 112.920 ;
        RECT 96.620 111.630 96.890 112.080 ;
        RECT 98.310 111.550 98.580 112.000 ;
        RECT 98.860 112.340 99.380 112.840 ;
        RECT 104.390 111.540 104.910 112.020 ;
        RECT 105.330 112.370 105.780 112.840 ;
        RECT 97.495 109.505 97.885 109.895 ;
        RECT 89.420 108.400 89.870 108.870 ;
        RECT 90.290 107.570 90.810 108.050 ;
        RECT 107.390 124.790 108.430 125.070 ;
        RECT 110.850 124.000 111.960 124.280 ;
        RECT 116.900 127.980 118.420 128.890 ;
        RECT 122.800 126.760 123.610 127.180 ;
        RECT 113.900 123.860 114.820 125.090 ;
        RECT 115.400 124.570 116.530 124.840 ;
        RECT 118.990 123.750 119.960 124.040 ;
        RECT 107.450 123.200 108.490 123.480 ;
        RECT 110.860 122.390 111.930 122.650 ;
        RECT 107.390 121.600 108.500 121.880 ;
        RECT 110.850 120.830 111.980 121.110 ;
        RECT 107.350 120.030 108.480 120.310 ;
        RECT 110.850 119.220 111.890 119.490 ;
        RECT 107.350 118.470 108.500 118.730 ;
        RECT 110.850 117.660 111.860 117.920 ;
        RECT 107.360 116.870 108.520 117.130 ;
        RECT 110.850 116.070 111.870 116.330 ;
        RECT 107.370 115.310 108.510 115.580 ;
        RECT 110.850 114.510 111.870 114.770 ;
        RECT 107.360 113.700 108.530 113.960 ;
        RECT 115.390 123.050 116.530 123.320 ;
        RECT 119.000 122.200 119.980 122.460 ;
        RECT 115.390 121.460 116.530 121.730 ;
        RECT 118.970 120.620 119.970 120.910 ;
        RECT 115.390 119.850 116.530 120.120 ;
        RECT 118.970 119.030 120.020 119.370 ;
        RECT 115.370 118.260 116.540 118.550 ;
        RECT 118.970 117.460 120.000 117.800 ;
        RECT 115.370 116.730 116.540 117.000 ;
        RECT 119.000 115.890 119.960 116.200 ;
        RECT 115.380 115.100 116.540 115.370 ;
        RECT 118.980 114.310 119.940 114.630 ;
        RECT 115.370 113.520 116.530 113.790 ;
        RECT 120.860 119.860 121.150 121.260 ;
        RECT 110.850 112.910 111.870 113.170 ;
        RECT 107.360 112.090 108.520 112.370 ;
        RECT 110.850 111.350 111.910 111.630 ;
        RECT 107.340 110.530 108.520 110.820 ;
        RECT 95.820 108.370 96.340 108.870 ;
        RECT 96.620 107.580 96.890 108.030 ;
        RECT 98.310 107.490 98.580 107.940 ;
        RECT 98.860 108.280 99.380 108.780 ;
        RECT 89.420 104.350 89.870 104.820 ;
        RECT 90.290 103.520 90.810 104.000 ;
        RECT 110.840 109.740 111.910 110.020 ;
        RECT 104.390 107.480 104.910 107.960 ;
        RECT 105.330 108.310 105.780 108.780 ;
        RECT 109.635 108.465 110.025 108.855 ;
        RECT 130.120 107.285 130.510 107.675 ;
        RECT 112.740 106.220 113.510 106.480 ;
        RECT 95.820 104.320 96.340 104.820 ;
        RECT 96.620 103.530 96.890 103.980 ;
        RECT 98.310 103.430 98.580 103.880 ;
        RECT 98.860 104.220 99.380 104.720 ;
        RECT 89.420 100.300 89.870 100.770 ;
        RECT 90.290 99.470 90.810 99.950 ;
        RECT 106.150 104.810 106.540 105.290 ;
        RECT 104.390 103.420 104.910 103.900 ;
        RECT 105.330 104.250 105.780 104.720 ;
        RECT 108.640 104.830 109.530 105.310 ;
        RECT 112.690 103.610 113.510 103.910 ;
        RECT 95.820 100.270 96.340 100.770 ;
        RECT 96.620 99.480 96.890 99.930 ;
        RECT 98.310 99.370 98.580 99.820 ;
        RECT 98.860 100.160 99.380 100.660 ;
        RECT 89.420 96.250 89.870 96.720 ;
        RECT 90.290 95.420 90.810 95.900 ;
        RECT 107.180 101.310 107.630 102.500 ;
        RECT 108.710 102.350 109.510 102.620 ;
        RECT 120.180 106.470 121.510 106.780 ;
        RECT 127.280 106.510 129.000 106.790 ;
        RECT 117.200 104.700 118.350 105.260 ;
        RECT 118.080 103.140 119.410 103.450 ;
        RECT 108.180 101.660 108.440 102.020 ;
        RECT 113.710 101.650 113.970 102.010 ;
        RECT 104.390 99.360 104.910 99.840 ;
        RECT 105.330 100.190 105.780 100.660 ;
        RECT 95.820 96.220 96.340 96.720 ;
        RECT 96.620 95.430 96.890 95.880 ;
        RECT 98.310 95.310 98.580 95.760 ;
        RECT 98.860 96.100 99.380 96.600 ;
        RECT 89.420 92.200 89.870 92.670 ;
        RECT 90.290 91.370 90.810 91.850 ;
        RECT 112.690 101.020 113.530 101.320 ;
        RECT 108.680 99.790 109.520 100.060 ;
        RECT 112.720 98.500 113.520 98.760 ;
        RECT 108.670 97.180 109.520 97.460 ;
        RECT 104.390 95.300 104.910 95.780 ;
        RECT 105.330 96.130 105.780 96.600 ;
        RECT 107.370 96.250 108.000 97.060 ;
        RECT 127.580 104.750 128.730 105.310 ;
        RECT 129.940 105.400 130.720 106.310 ;
        RECT 136.980 107.440 137.550 107.800 ;
        RECT 137.230 106.560 137.730 106.920 ;
        RECT 132.300 105.820 132.570 106.300 ;
        RECT 122.220 101.590 122.490 102.430 ;
        RECT 125.110 102.980 126.630 103.320 ;
        RECT 132.050 103.460 132.540 104.230 ;
        RECT 129.780 101.560 130.050 102.470 ;
        RECT 120.180 100.420 121.510 100.730 ;
        RECT 127.180 100.490 129.010 100.820 ;
        RECT 137.980 105.800 138.250 106.280 ;
        RECT 137.000 102.840 137.570 103.300 ;
        RECT 117.250 98.690 118.400 99.250 ;
        RECT 122.210 97.570 122.470 98.410 ;
        RECT 127.580 98.740 128.730 99.300 ;
        RECT 118.070 97.130 119.400 97.440 ;
        RECT 122.870 97.270 123.720 98.240 ;
        RECT 136.970 98.470 137.660 98.860 ;
        RECT 138.650 107.470 138.940 107.750 ;
        RECT 138.650 102.940 138.940 103.220 ;
        RECT 138.660 98.450 138.950 98.730 ;
        RECT 125.100 96.940 126.600 97.390 ;
        RECT 133.200 97.380 134.620 97.960 ;
        RECT 137.170 97.540 137.750 97.900 ;
        RECT 112.700 95.900 113.510 96.160 ;
        RECT 139.580 106.690 140.050 107.060 ;
        RECT 139.580 102.000 140.040 102.560 ;
        RECT 139.540 97.610 140.030 98.070 ;
        RECT 140.710 107.480 141.000 107.760 ;
        RECT 140.700 103.030 140.990 103.310 ;
        RECT 141.780 107.440 142.680 107.740 ;
        RECT 141.280 105.800 141.550 106.280 ;
        RECT 146.970 105.830 147.240 106.310 ;
        RECT 141.850 103.020 142.640 103.370 ;
        RECT 141.800 101.950 142.540 102.410 ;
        RECT 141.820 98.520 142.610 98.830 ;
        RECT 147.540 107.160 147.940 107.930 ;
        RECT 95.820 92.170 96.340 92.670 ;
        RECT 96.620 91.380 96.890 91.830 ;
        RECT 98.310 91.250 98.580 91.700 ;
        RECT 98.860 92.040 99.380 92.540 ;
        RECT 89.420 88.150 89.870 88.620 ;
        RECT 90.290 87.320 90.810 87.800 ;
        RECT 106.590 93.510 107.880 93.770 ;
        RECT 104.390 91.240 104.910 91.720 ;
        RECT 105.330 92.070 105.780 92.540 ;
        RECT 122.790 91.820 123.600 92.240 ;
        RECT 95.820 88.120 96.340 88.620 ;
        RECT 96.620 87.330 96.890 87.780 ;
        RECT 98.310 87.190 98.580 87.640 ;
        RECT 98.860 87.980 99.380 88.480 ;
        RECT 89.420 84.100 89.870 84.570 ;
        RECT 90.290 83.270 90.810 83.750 ;
        RECT 104.390 87.180 104.910 87.660 ;
        RECT 105.330 88.010 105.780 88.480 ;
        RECT 112.400 89.460 113.010 90.280 ;
        RECT 95.820 84.070 96.340 84.570 ;
        RECT 96.620 83.280 96.890 83.730 ;
        RECT 98.310 83.130 98.580 83.580 ;
        RECT 98.860 83.920 99.380 84.420 ;
        RECT 89.420 80.050 89.870 80.520 ;
        RECT 90.290 79.220 90.810 79.700 ;
        RECT 104.390 83.120 104.910 83.600 ;
        RECT 105.330 83.950 105.780 84.420 ;
        RECT 95.820 80.020 96.340 80.520 ;
        RECT 96.620 79.230 96.890 79.680 ;
        RECT 98.310 79.070 98.580 79.520 ;
        RECT 98.860 79.860 99.380 80.360 ;
        RECT 89.420 76.000 89.870 76.470 ;
        RECT 90.290 75.170 90.810 75.650 ;
        RECT 104.390 79.060 104.910 79.540 ;
        RECT 105.330 79.890 105.780 80.360 ;
        RECT 106.100 80.250 106.410 80.980 ;
        RECT 95.820 75.970 96.340 76.470 ;
        RECT 96.620 75.180 96.890 75.630 ;
        RECT 98.310 75.010 98.580 75.460 ;
        RECT 98.860 75.800 99.380 76.300 ;
        RECT 89.420 71.950 89.870 72.420 ;
        RECT 90.290 71.120 90.810 71.600 ;
        RECT 104.390 75.000 104.910 75.480 ;
        RECT 105.330 75.830 105.780 76.300 ;
        RECT 95.820 71.920 96.340 72.420 ;
        RECT 96.620 71.130 96.890 71.580 ;
        RECT 98.310 70.950 98.580 71.400 ;
        RECT 98.860 71.740 99.380 72.240 ;
        RECT 89.420 67.900 89.870 68.370 ;
        RECT 90.290 67.070 90.810 67.550 ;
        RECT 104.390 70.940 104.910 71.420 ;
        RECT 105.330 71.770 105.780 72.240 ;
        RECT 107.390 86.870 108.430 87.150 ;
        RECT 110.850 86.080 111.960 86.360 ;
        RECT 116.900 90.060 118.420 90.970 ;
        RECT 122.800 88.840 123.610 89.260 ;
        RECT 113.900 85.940 114.820 87.170 ;
        RECT 115.400 86.650 116.530 86.920 ;
        RECT 118.990 85.830 119.960 86.120 ;
        RECT 107.450 85.280 108.490 85.560 ;
        RECT 110.860 84.470 111.930 84.730 ;
        RECT 107.390 83.680 108.500 83.960 ;
        RECT 110.850 82.910 111.980 83.190 ;
        RECT 107.350 82.110 108.480 82.390 ;
        RECT 110.850 81.300 111.890 81.570 ;
        RECT 107.350 80.550 108.500 80.810 ;
        RECT 110.850 79.740 111.860 80.000 ;
        RECT 107.360 78.950 108.520 79.210 ;
        RECT 110.850 78.150 111.870 78.410 ;
        RECT 107.370 77.390 108.510 77.660 ;
        RECT 110.850 76.590 111.870 76.850 ;
        RECT 107.360 75.780 108.530 76.040 ;
        RECT 115.390 85.130 116.530 85.400 ;
        RECT 119.000 84.280 119.980 84.540 ;
        RECT 115.390 83.540 116.530 83.810 ;
        RECT 118.970 82.700 119.970 82.990 ;
        RECT 115.390 81.930 116.530 82.200 ;
        RECT 118.970 81.110 120.020 81.450 ;
        RECT 115.370 80.340 116.540 80.630 ;
        RECT 118.970 79.540 120.000 79.880 ;
        RECT 115.370 78.810 116.540 79.080 ;
        RECT 119.000 77.970 119.960 78.280 ;
        RECT 115.380 77.180 116.540 77.450 ;
        RECT 118.980 76.390 119.940 76.710 ;
        RECT 115.370 75.600 116.530 75.870 ;
        RECT 120.860 81.940 121.150 83.340 ;
        RECT 122.660 82.590 124.190 84.000 ;
        RECT 110.850 74.990 111.870 75.250 ;
        RECT 107.360 74.170 108.520 74.450 ;
        RECT 110.850 73.430 111.910 73.710 ;
        RECT 107.340 72.610 108.520 72.900 ;
        RECT 110.840 71.820 111.910 72.100 ;
        RECT 95.820 67.870 96.340 68.370 ;
        RECT 96.620 67.080 96.890 67.530 ;
        RECT 98.310 66.890 98.580 67.340 ;
        RECT 98.860 67.680 99.380 68.180 ;
        RECT 89.420 63.850 89.870 64.320 ;
        RECT 90.290 63.020 90.810 63.500 ;
        RECT 104.390 66.880 104.910 67.360 ;
        RECT 105.330 67.710 105.780 68.180 ;
        RECT 95.820 63.820 96.340 64.320 ;
        RECT 96.620 63.030 96.890 63.480 ;
        RECT 98.310 62.830 98.580 63.280 ;
        RECT 98.860 63.620 99.380 64.120 ;
        RECT 104.390 62.820 104.910 63.300 ;
        RECT 105.330 63.650 105.780 64.120 ;
        RECT 89.420 59.800 89.870 60.270 ;
        RECT 90.290 58.970 90.810 59.450 ;
        RECT 101.755 61.250 102.325 62.020 ;
        RECT 95.820 59.770 96.340 60.270 ;
        RECT 96.620 58.980 96.890 59.430 ;
        RECT 98.310 58.290 98.580 58.740 ;
        RECT 98.860 59.080 99.380 59.580 ;
        RECT 104.390 58.280 104.910 58.760 ;
        RECT 105.330 59.110 105.780 59.580 ;
        RECT 89.420 55.750 89.870 56.220 ;
        RECT 90.290 54.920 90.810 55.400 ;
        RECT 95.820 55.720 96.340 56.220 ;
        RECT 96.620 54.930 96.890 55.380 ;
        RECT 89.420 51.700 89.870 52.170 ;
        RECT 90.290 50.870 90.810 51.350 ;
        RECT 95.820 51.670 96.340 52.170 ;
        RECT 105.965 53.400 106.945 54.380 ;
        RECT 96.620 50.880 96.890 51.330 ;
        RECT 89.420 47.650 89.870 48.120 ;
        RECT 90.290 46.820 90.810 47.300 ;
        RECT 95.820 47.620 96.340 48.120 ;
        RECT 96.620 46.830 96.890 47.280 ;
        RECT 89.420 43.600 89.870 44.070 ;
        RECT 90.290 42.770 90.810 43.250 ;
        RECT 95.820 43.570 96.340 44.070 ;
        RECT 96.620 42.780 96.890 43.230 ;
        RECT 89.420 39.550 89.870 40.020 ;
        RECT 90.290 38.720 90.810 39.200 ;
        RECT 95.820 39.520 96.340 40.020 ;
        RECT 96.620 38.730 96.890 39.180 ;
        RECT 89.420 35.500 89.870 35.970 ;
        RECT 90.290 34.670 90.810 35.150 ;
        RECT 95.820 35.470 96.340 35.970 ;
        RECT 96.620 34.680 96.890 35.130 ;
        RECT 89.420 31.450 89.870 31.920 ;
        RECT 90.290 30.620 90.810 31.100 ;
        RECT 95.820 31.420 96.340 31.920 ;
        RECT 96.620 30.630 96.890 31.080 ;
        RECT 89.420 27.365 89.870 27.835 ;
        RECT 90.290 26.535 90.810 27.015 ;
        RECT 95.820 27.335 96.340 27.835 ;
        RECT 96.620 26.545 96.890 26.995 ;
        RECT 89.420 23.240 89.870 23.710 ;
        RECT 90.290 22.410 90.810 22.890 ;
        RECT 92.870 20.910 93.455 21.680 ;
        RECT 95.820 23.210 96.340 23.710 ;
        RECT 96.620 22.420 96.890 22.870 ;
        RECT 89.420 18.685 89.870 19.155 ;
        RECT 90.290 17.855 90.810 18.335 ;
        RECT 95.820 18.655 96.340 19.155 ;
        RECT 96.620 17.865 96.890 18.315 ;
      LAYER met2 ;
        RECT 107.250 153.820 107.860 153.850 ;
        RECT 90.020 152.910 107.860 153.820 ;
        RECT 90.020 151.670 100.870 152.910 ;
        RECT 104.270 151.670 107.860 152.910 ;
        RECT 96.530 147.980 99.090 150.790 ;
        RECT 87.690 143.050 88.920 146.890 ;
        RECT 92.815 145.715 93.515 146.635 ;
        RECT 101.685 145.870 102.385 146.640 ;
        RECT 89.390 144.790 96.380 145.360 ;
        RECT 98.820 144.790 105.810 145.360 ;
        RECT 107.250 144.860 107.860 151.670 ;
        RECT 108.175 147.380 109.105 147.400 ;
        RECT 122.670 147.380 124.180 147.460 ;
        RECT 108.150 146.400 124.180 147.380 ;
        RECT 108.175 146.380 109.105 146.400 ;
        RECT 110.640 146.395 124.180 146.400 ;
        RECT 122.670 146.160 124.180 146.395 ;
        RECT 136.890 145.730 137.610 145.850 ;
        RECT 147.470 145.760 148.020 145.930 ;
        RECT 138.550 145.730 141.070 145.740 ;
        RECT 141.690 145.730 148.030 145.760 ;
        RECT 136.890 145.360 148.030 145.730 ;
        RECT 136.890 145.280 137.610 145.360 ;
        RECT 138.550 145.340 141.070 145.360 ;
        RECT 141.690 145.310 148.030 145.360 ;
        RECT 141.730 145.240 148.030 145.310 ;
        RECT 137.170 144.890 137.800 144.920 ;
        RECT 139.220 144.890 140.160 145.190 ;
        RECT 147.470 144.970 148.020 145.240 ;
        RECT 90.230 143.980 96.930 144.550 ;
        RECT 98.270 143.980 104.970 144.550 ;
        RECT 107.250 143.590 108.400 144.860 ;
        RECT 112.650 144.040 113.570 144.460 ;
        RECT 115.220 144.060 116.450 144.410 ;
        RECT 120.100 144.280 121.560 144.760 ;
        RECT 127.150 144.380 129.070 144.810 ;
        RECT 137.170 144.490 140.160 144.890 ;
        RECT 137.170 144.450 137.800 144.490 ;
        RECT 139.220 144.430 140.160 144.490 ;
        RECT 129.760 144.060 130.870 144.420 ;
        RECT 115.220 143.770 130.870 144.060 ;
        RECT 115.220 143.760 124.640 143.770 ;
        RECT 89.450 142.340 105.750 143.160 ;
        RECT 106.030 142.640 109.650 143.300 ;
        RECT 115.220 143.270 116.450 143.760 ;
        RECT 120.630 143.360 124.610 143.370 ;
        RECT 108.550 142.630 109.650 142.640 ;
        RECT 117.010 142.470 129.050 143.360 ;
        RECT 129.760 143.070 130.870 143.770 ;
        RECT 132.270 143.650 147.270 144.290 ;
        RECT 112.650 141.460 113.570 141.880 ;
        RECT 123.170 141.460 126.720 141.470 ;
        RECT 89.390 140.790 96.380 141.360 ;
        RECT 98.820 140.730 105.810 141.300 ;
        RECT 118.010 140.970 119.470 141.450 ;
        RECT 120.150 140.820 126.720 141.460 ;
        RECT 127.200 141.330 132.590 142.220 ;
        RECT 141.770 141.270 142.710 141.340 ;
        RECT 136.940 141.200 137.660 141.270 ;
        RECT 140.630 141.230 142.710 141.270 ;
        RECT 138.640 141.200 142.710 141.230 ;
        RECT 136.930 140.920 142.710 141.200 ;
        RECT 136.930 140.830 138.990 140.920 ;
        RECT 140.630 140.900 142.710 140.920 ;
        RECT 141.770 140.870 142.710 140.900 ;
        RECT 123.170 140.800 126.720 140.820 ;
        RECT 136.940 140.700 137.660 140.830 ;
        RECT 90.230 139.980 96.930 140.550 ;
        RECT 98.270 139.920 104.970 140.490 ;
        RECT 108.590 140.180 109.600 140.640 ;
        RECT 139.480 140.470 140.140 140.590 ;
        RECT 139.480 140.460 142.460 140.470 ;
        RECT 123.380 140.420 130.080 140.430 ;
        RECT 108.130 139.530 114.010 139.980 ;
        RECT 122.010 139.460 130.080 140.420 ;
        RECT 139.480 140.070 142.710 140.460 ;
        RECT 139.480 139.790 140.140 140.070 ;
        RECT 141.740 139.740 142.710 140.070 ;
        RECT 122.010 139.450 123.880 139.460 ;
        RECT 129.450 139.450 130.080 139.460 ;
        RECT 112.640 138.870 113.580 139.300 ;
        RECT 118.080 139.280 119.430 139.400 ;
        RECT 118.080 139.210 128.930 139.280 ;
        RECT 118.080 138.910 129.050 139.210 ;
        RECT 118.080 138.820 119.430 138.910 ;
        RECT 108.590 137.620 109.590 138.080 ;
        RECT 112.650 137.640 117.580 138.510 ;
        RECT 120.130 138.270 121.590 138.750 ;
        RECT 127.120 138.210 129.050 138.910 ;
        RECT 127.150 138.170 129.040 138.210 ;
        RECT 117.000 137.350 125.350 137.380 ;
        RECT 89.390 136.690 96.380 137.260 ;
        RECT 98.820 136.670 105.810 137.240 ;
        RECT 90.230 135.880 96.930 136.450 ;
        RECT 98.270 135.860 104.970 136.430 ;
        RECT 112.650 136.360 113.570 136.730 ;
        RECT 117.000 136.720 129.000 137.350 ;
        RECT 117.000 136.480 121.980 136.720 ;
        RECT 124.020 136.450 129.000 136.720 ;
        RECT 136.900 136.730 137.720 136.820 ;
        RECT 136.900 136.690 138.990 136.730 ;
        RECT 141.710 136.700 142.710 136.800 ;
        RECT 140.650 136.690 142.710 136.700 ;
        RECT 106.920 133.620 108.390 135.090 ;
        RECT 108.620 135.030 109.570 135.460 ;
        RECT 118.030 134.960 119.490 135.440 ;
        RECT 122.110 135.410 122.540 136.420 ;
        RECT 122.760 134.990 123.870 136.320 ;
        RECT 129.810 135.890 134.780 136.470 ;
        RECT 136.900 136.380 142.710 136.690 ;
        RECT 136.900 136.360 138.990 136.380 ;
        RECT 136.900 136.320 137.720 136.360 ;
        RECT 140.650 136.330 142.710 136.380 ;
        RECT 139.460 135.890 140.110 136.050 ;
        RECT 129.810 135.490 140.110 135.890 ;
        RECT 124.990 134.800 126.720 135.350 ;
        RECT 129.810 135.160 137.850 135.490 ;
        RECT 139.460 135.440 140.110 135.490 ;
        RECT 129.820 134.340 130.460 135.160 ;
        RECT 120.170 134.330 130.460 134.340 ;
        RECT 112.640 133.790 113.580 134.160 ;
        RECT 113.950 133.770 130.460 134.330 ;
        RECT 113.950 133.430 121.630 133.770 ;
        RECT 89.390 132.640 96.380 133.210 ;
        RECT 98.820 132.610 105.810 133.180 ;
        RECT 90.230 131.830 96.930 132.400 ;
        RECT 98.270 131.800 104.970 132.370 ;
        RECT 106.460 130.970 108.040 132.010 ;
        RECT 127.490 131.790 132.040 133.420 ;
        RECT 115.230 131.490 132.040 131.790 ;
        RECT 115.230 131.080 132.030 131.490 ;
        RECT 125.890 130.500 127.570 131.080 ;
        RECT 89.390 128.590 96.380 129.160 ;
        RECT 98.820 128.550 105.810 129.120 ;
        RECT 116.760 129.010 118.600 129.090 ;
        RECT 90.230 127.780 96.930 128.350 ;
        RECT 98.270 127.740 104.970 128.310 ;
        RECT 106.900 127.150 113.130 128.390 ;
        RECT 116.760 127.770 121.770 129.010 ;
        RECT 116.850 127.640 121.770 127.770 ;
        RECT 122.740 128.910 123.650 130.220 ;
        RECT 122.740 126.690 125.880 128.910 ;
        RECT 122.770 126.350 125.880 126.690 ;
        RECT 89.390 124.540 96.380 125.110 ;
        RECT 98.820 124.490 105.810 125.060 ;
        RECT 107.120 124.760 111.960 125.100 ;
        RECT 110.810 124.320 112.020 124.340 ;
        RECT 90.230 123.730 96.930 124.300 ;
        RECT 98.270 123.680 104.970 124.250 ;
        RECT 107.160 123.980 112.020 124.320 ;
        RECT 110.810 123.940 112.020 123.980 ;
        RECT 113.820 123.700 115.000 125.200 ;
        RECT 115.210 124.570 120.050 124.910 ;
        RECT 118.910 124.080 120.030 124.090 ;
        RECT 115.190 123.740 120.030 124.080 ;
        RECT 107.210 123.190 112.050 123.530 ;
        RECT 115.310 123.350 116.570 123.360 ;
        RECT 115.160 123.010 120.000 123.350 ;
        RECT 115.310 123.000 116.570 123.010 ;
        RECT 107.180 122.360 112.020 122.700 ;
        RECT 115.200 122.180 120.060 122.520 ;
        RECT 118.910 122.130 120.060 122.180 ;
        RECT 107.290 121.930 108.570 121.950 ;
        RECT 107.230 121.590 112.070 121.930 ;
        RECT 115.320 121.760 116.580 121.770 ;
        RECT 107.290 121.550 108.570 121.590 ;
        RECT 115.200 121.420 120.040 121.760 ;
        RECT 115.320 121.410 116.580 121.420 ;
        RECT 110.800 121.130 112.040 121.140 ;
        RECT 89.390 120.490 96.380 121.060 ;
        RECT 98.820 120.430 105.810 121.000 ;
        RECT 107.200 120.790 112.040 121.130 ;
        RECT 120.790 121.000 121.220 121.370 ;
        RECT 118.910 120.930 121.220 121.000 ;
        RECT 115.160 120.590 121.220 120.930 ;
        RECT 118.910 120.520 121.220 120.590 ;
        RECT 90.230 119.680 96.930 120.250 ;
        RECT 98.270 119.620 104.970 120.190 ;
        RECT 107.150 119.990 111.990 120.330 ;
        RECT 113.260 120.180 113.590 120.200 ;
        RECT 113.260 120.170 116.110 120.180 ;
        RECT 113.260 120.160 116.580 120.170 ;
        RECT 113.260 119.820 120.100 120.160 ;
        RECT 113.260 119.810 116.580 119.820 ;
        RECT 113.260 119.530 113.590 119.810 ;
        RECT 120.790 119.780 121.220 120.520 ;
        RECT 110.790 119.520 113.590 119.530 ;
        RECT 107.100 119.180 113.590 119.520 ;
        RECT 118.920 119.370 120.080 119.400 ;
        RECT 110.790 119.170 113.590 119.180 ;
        RECT 110.860 119.160 113.590 119.170 ;
        RECT 113.260 119.140 113.590 119.160 ;
        RECT 115.250 119.030 120.090 119.370 ;
        RECT 118.920 118.980 120.080 119.030 ;
        RECT 106.030 118.840 106.450 118.980 ;
        RECT 106.030 118.770 108.570 118.840 ;
        RECT 106.030 118.430 111.940 118.770 ;
        RECT 106.030 118.380 108.570 118.430 ;
        RECT 106.030 118.120 106.450 118.380 ;
        RECT 115.270 118.230 120.110 118.570 ;
        RECT 107.080 117.630 111.920 117.970 ;
        RECT 118.920 117.810 120.070 117.850 ;
        RECT 115.230 117.470 120.070 117.810 ;
        RECT 118.920 117.390 120.070 117.470 ;
        RECT 89.390 116.440 96.380 117.010 ;
        RECT 98.820 116.370 105.810 116.940 ;
        RECT 107.110 116.840 111.950 117.180 ;
        RECT 115.210 116.700 120.050 117.040 ;
        RECT 110.800 116.370 111.950 116.380 ;
        RECT 90.230 115.630 96.930 116.200 ;
        RECT 98.270 115.560 104.970 116.130 ;
        RECT 107.110 116.030 111.950 116.370 ;
        RECT 118.920 116.210 120.020 116.250 ;
        RECT 115.140 115.870 120.020 116.210 ;
        RECT 118.920 115.830 120.020 115.870 ;
        RECT 107.160 115.270 112.000 115.610 ;
        RECT 115.150 115.070 119.990 115.410 ;
        RECT 110.800 114.800 111.990 114.810 ;
        RECT 107.150 114.460 111.990 114.800 ;
        RECT 118.920 114.640 120.000 114.680 ;
        RECT 110.800 114.450 111.990 114.460 ;
        RECT 115.150 114.300 120.000 114.640 ;
        RECT 118.920 114.250 120.000 114.300 ;
        RECT 107.130 113.670 111.970 114.010 ;
        RECT 115.320 113.820 116.580 113.830 ;
        RECT 115.170 113.480 120.010 113.820 ;
        RECT 89.390 112.390 96.380 112.960 ;
        RECT 107.110 112.880 111.950 113.220 ;
        RECT 98.820 112.310 105.810 112.880 ;
        RECT 110.800 112.870 111.950 112.880 ;
        RECT 107.300 112.420 108.570 112.430 ;
        RECT 90.230 111.580 96.930 112.150 ;
        RECT 107.100 112.080 111.940 112.420 ;
        RECT 98.270 111.500 104.970 112.070 ;
        RECT 107.300 112.040 108.570 112.080 ;
        RECT 110.810 111.660 111.990 111.710 ;
        RECT 107.110 111.320 111.990 111.660 ;
        RECT 110.810 111.290 111.990 111.320 ;
        RECT 107.300 110.840 108.580 110.850 ;
        RECT 107.110 110.500 111.950 110.840 ;
        RECT 107.300 110.490 108.580 110.500 ;
        RECT 110.790 110.050 111.990 110.060 ;
        RECT 97.465 109.505 106.615 109.895 ;
        RECT 107.100 109.710 111.990 110.050 ;
        RECT 110.790 109.700 111.990 109.710 ;
        RECT 89.390 108.340 96.380 108.910 ;
        RECT 106.225 108.855 106.615 109.505 ;
        RECT 109.635 108.855 110.025 108.885 ;
        RECT 98.820 108.250 105.810 108.820 ;
        RECT 106.225 108.465 110.025 108.855 ;
        RECT 109.635 108.435 110.025 108.465 ;
        RECT 90.230 107.530 96.930 108.100 ;
        RECT 98.270 107.440 104.970 108.010 ;
        RECT 136.890 107.810 137.610 107.930 ;
        RECT 147.470 107.840 148.020 108.010 ;
        RECT 138.550 107.810 141.070 107.820 ;
        RECT 141.690 107.810 148.030 107.840 ;
        RECT 130.120 107.675 130.510 107.705 ;
        RECT 115.960 107.285 130.510 107.675 ;
        RECT 136.890 107.440 148.030 107.810 ;
        RECT 136.890 107.360 137.610 107.440 ;
        RECT 138.550 107.420 141.070 107.440 ;
        RECT 141.690 107.390 148.030 107.440 ;
        RECT 141.730 107.320 148.030 107.390 ;
        RECT 130.120 107.255 130.510 107.285 ;
        RECT 137.170 106.970 137.800 107.000 ;
        RECT 139.220 106.970 140.160 107.270 ;
        RECT 147.470 107.050 148.020 107.320 ;
        RECT 112.650 106.120 113.570 106.540 ;
        RECT 120.100 106.360 121.560 106.840 ;
        RECT 127.150 106.460 129.070 106.890 ;
        RECT 137.170 106.570 140.160 106.970 ;
        RECT 137.170 106.530 137.800 106.570 ;
        RECT 139.220 106.510 140.160 106.570 ;
        RECT 120.630 105.440 124.610 105.450 ;
        RECT 89.390 104.290 96.380 104.860 ;
        RECT 98.820 104.190 105.810 104.760 ;
        RECT 106.030 104.720 109.650 105.380 ;
        RECT 108.550 104.710 109.650 104.720 ;
        RECT 117.010 104.550 129.050 105.440 ;
        RECT 129.760 105.150 130.870 106.500 ;
        RECT 132.270 105.730 147.270 106.370 ;
        RECT 90.230 103.480 96.930 104.050 ;
        RECT 98.270 103.380 104.970 103.950 ;
        RECT 112.650 103.540 113.570 103.960 ;
        RECT 123.170 103.540 126.720 103.550 ;
        RECT 118.010 103.050 119.470 103.530 ;
        RECT 120.150 102.900 126.720 103.540 ;
        RECT 127.200 103.410 132.590 104.300 ;
        RECT 141.770 103.350 142.710 103.420 ;
        RECT 136.940 103.280 137.660 103.350 ;
        RECT 140.630 103.310 142.710 103.350 ;
        RECT 138.640 103.280 142.710 103.310 ;
        RECT 136.930 103.000 142.710 103.280 ;
        RECT 136.930 102.910 138.990 103.000 ;
        RECT 140.630 102.980 142.710 103.000 ;
        RECT 141.770 102.950 142.710 102.980 ;
        RECT 123.170 102.880 126.720 102.900 ;
        RECT 136.940 102.780 137.660 102.910 ;
        RECT 107.100 101.220 107.680 102.580 ;
        RECT 108.590 102.260 109.600 102.720 ;
        RECT 139.480 102.550 140.140 102.670 ;
        RECT 139.480 102.540 142.460 102.550 ;
        RECT 123.380 102.500 130.080 102.510 ;
        RECT 108.130 101.610 114.010 102.060 ;
        RECT 122.010 101.540 130.080 102.500 ;
        RECT 139.480 102.150 142.710 102.540 ;
        RECT 139.480 101.870 140.140 102.150 ;
        RECT 141.740 101.820 142.710 102.150 ;
        RECT 122.010 101.530 123.880 101.540 ;
        RECT 129.450 101.530 130.080 101.540 ;
        RECT 112.640 100.950 113.580 101.380 ;
        RECT 118.080 101.360 119.430 101.480 ;
        RECT 118.080 101.290 128.930 101.360 ;
        RECT 118.080 100.990 129.050 101.290 ;
        RECT 118.080 100.900 119.430 100.990 ;
        RECT 89.390 100.240 96.380 100.810 ;
        RECT 98.820 100.130 105.810 100.700 ;
        RECT 90.230 99.430 96.930 100.000 ;
        RECT 98.270 99.320 104.970 99.890 ;
        RECT 108.590 99.700 109.590 100.160 ;
        RECT 112.650 99.720 117.580 100.590 ;
        RECT 120.130 100.350 121.590 100.830 ;
        RECT 127.120 100.290 129.050 100.990 ;
        RECT 127.150 100.250 129.040 100.290 ;
        RECT 117.000 99.430 125.350 99.460 ;
        RECT 112.650 98.440 113.570 98.810 ;
        RECT 117.000 98.800 129.000 99.430 ;
        RECT 117.000 98.560 121.980 98.800 ;
        RECT 124.020 98.530 129.000 98.800 ;
        RECT 136.900 98.810 137.720 98.900 ;
        RECT 136.900 98.770 138.990 98.810 ;
        RECT 141.710 98.780 142.710 98.880 ;
        RECT 140.650 98.770 142.710 98.780 ;
        RECT 89.390 96.190 96.380 96.760 ;
        RECT 98.820 96.070 105.810 96.640 ;
        RECT 90.230 95.380 96.930 95.950 ;
        RECT 98.270 95.260 104.970 95.830 ;
        RECT 106.920 95.700 108.390 97.170 ;
        RECT 108.620 97.110 109.570 97.540 ;
        RECT 118.030 97.040 119.490 97.520 ;
        RECT 122.110 97.490 122.540 98.500 ;
        RECT 122.760 97.070 123.870 98.400 ;
        RECT 129.810 97.970 134.780 98.550 ;
        RECT 136.900 98.460 142.710 98.770 ;
        RECT 136.900 98.440 138.990 98.460 ;
        RECT 136.900 98.400 137.720 98.440 ;
        RECT 140.650 98.410 142.710 98.460 ;
        RECT 139.460 97.970 140.110 98.130 ;
        RECT 129.810 97.570 140.110 97.970 ;
        RECT 124.990 96.880 126.720 97.430 ;
        RECT 129.810 97.240 137.850 97.570 ;
        RECT 139.460 97.520 140.110 97.570 ;
        RECT 129.820 96.420 130.460 97.240 ;
        RECT 120.170 96.410 130.460 96.420 ;
        RECT 112.640 95.870 113.580 96.240 ;
        RECT 113.950 95.850 130.460 96.410 ;
        RECT 113.950 95.510 121.630 95.850 ;
        RECT 106.460 93.050 108.040 94.090 ;
        RECT 127.490 93.870 132.040 95.500 ;
        RECT 115.230 93.570 132.040 93.870 ;
        RECT 115.230 93.160 132.030 93.570 ;
        RECT 89.390 92.140 96.380 92.710 ;
        RECT 125.890 92.580 127.570 93.160 ;
        RECT 98.820 92.010 105.810 92.580 ;
        RECT 90.230 91.330 96.930 91.900 ;
        RECT 98.270 91.200 104.970 91.770 ;
        RECT 116.760 91.090 118.600 91.170 ;
        RECT 106.900 89.230 113.130 90.470 ;
        RECT 116.760 89.850 121.770 91.090 ;
        RECT 116.850 89.720 121.770 89.850 ;
        RECT 122.740 90.990 123.650 92.300 ;
        RECT 122.740 88.770 125.880 90.990 ;
        RECT 89.390 88.090 96.380 88.660 ;
        RECT 98.820 87.950 105.810 88.520 ;
        RECT 122.770 88.430 125.880 88.770 ;
        RECT 90.230 87.280 96.930 87.850 ;
        RECT 98.270 87.140 104.970 87.710 ;
        RECT 107.120 86.840 111.960 87.180 ;
        RECT 110.810 86.400 112.020 86.420 ;
        RECT 107.160 86.060 112.020 86.400 ;
        RECT 110.810 86.020 112.020 86.060 ;
        RECT 113.820 85.780 115.000 87.280 ;
        RECT 115.210 86.650 120.050 86.990 ;
        RECT 118.910 86.160 120.030 86.170 ;
        RECT 115.190 85.820 120.030 86.160 ;
        RECT 107.210 85.270 112.050 85.610 ;
        RECT 115.310 85.430 116.570 85.440 ;
        RECT 115.160 85.090 120.000 85.430 ;
        RECT 115.310 85.080 116.570 85.090 ;
        RECT 89.390 84.040 96.380 84.610 ;
        RECT 98.820 83.890 105.810 84.460 ;
        RECT 107.180 84.440 112.020 84.780 ;
        RECT 115.200 84.260 120.060 84.600 ;
        RECT 118.910 84.210 120.060 84.260 ;
        RECT 107.290 84.010 108.570 84.030 ;
        RECT 90.230 83.230 96.930 83.800 ;
        RECT 107.230 83.670 112.070 84.010 ;
        RECT 115.320 83.840 116.580 83.850 ;
        RECT 98.270 83.080 104.970 83.650 ;
        RECT 107.290 83.630 108.570 83.670 ;
        RECT 115.200 83.500 120.040 83.840 ;
        RECT 115.320 83.490 116.580 83.500 ;
        RECT 110.800 83.210 112.040 83.220 ;
        RECT 107.200 82.870 112.040 83.210 ;
        RECT 120.790 83.080 121.220 83.450 ;
        RECT 118.910 83.010 121.220 83.080 ;
        RECT 115.160 82.670 121.220 83.010 ;
        RECT 118.910 82.600 121.220 82.670 ;
        RECT 107.150 82.070 111.990 82.410 ;
        RECT 113.260 82.260 113.590 82.280 ;
        RECT 113.260 82.250 116.110 82.260 ;
        RECT 113.260 82.240 116.580 82.250 ;
        RECT 113.260 81.900 120.100 82.240 ;
        RECT 113.260 81.890 116.580 81.900 ;
        RECT 113.260 81.610 113.590 81.890 ;
        RECT 120.790 81.860 121.220 82.600 ;
        RECT 122.440 82.380 124.340 84.310 ;
        RECT 110.790 81.600 113.590 81.610 ;
        RECT 107.100 81.260 113.590 81.600 ;
        RECT 118.920 81.450 120.080 81.480 ;
        RECT 110.790 81.250 113.590 81.260 ;
        RECT 110.860 81.240 113.590 81.250 ;
        RECT 113.260 81.220 113.590 81.240 ;
        RECT 115.250 81.110 120.090 81.450 ;
        RECT 118.920 81.060 120.080 81.110 ;
        RECT 106.030 80.920 106.450 81.060 ;
        RECT 106.030 80.850 108.570 80.920 ;
        RECT 89.390 79.990 96.380 80.560 ;
        RECT 106.030 80.510 111.940 80.850 ;
        RECT 106.030 80.460 108.570 80.510 ;
        RECT 98.820 79.830 105.810 80.400 ;
        RECT 106.030 80.200 106.450 80.460 ;
        RECT 115.270 80.310 120.110 80.650 ;
        RECT 90.230 79.180 96.930 79.750 ;
        RECT 107.080 79.710 111.920 80.050 ;
        RECT 118.920 79.890 120.070 79.930 ;
        RECT 98.270 79.020 104.970 79.590 ;
        RECT 115.230 79.550 120.070 79.890 ;
        RECT 118.920 79.470 120.070 79.550 ;
        RECT 107.110 78.920 111.950 79.260 ;
        RECT 115.210 78.780 120.050 79.120 ;
        RECT 110.800 78.450 111.950 78.460 ;
        RECT 107.110 78.110 111.950 78.450 ;
        RECT 118.920 78.290 120.020 78.330 ;
        RECT 115.140 77.950 120.020 78.290 ;
        RECT 118.920 77.910 120.020 77.950 ;
        RECT 107.160 77.350 112.000 77.690 ;
        RECT 115.150 77.150 119.990 77.490 ;
        RECT 110.800 76.880 111.990 76.890 ;
        RECT 107.150 76.540 111.990 76.880 ;
        RECT 118.920 76.720 120.000 76.760 ;
        RECT 110.800 76.530 111.990 76.540 ;
        RECT 89.390 75.940 96.380 76.510 ;
        RECT 115.150 76.380 120.000 76.720 ;
        RECT 98.820 75.770 105.810 76.340 ;
        RECT 118.920 76.330 120.000 76.380 ;
        RECT 107.130 75.750 111.970 76.090 ;
        RECT 115.320 75.900 116.580 75.910 ;
        RECT 90.230 75.130 96.930 75.700 ;
        RECT 115.170 75.560 120.010 75.900 ;
        RECT 98.270 74.960 104.970 75.530 ;
        RECT 107.110 74.960 111.950 75.300 ;
        RECT 110.800 74.950 111.950 74.960 ;
        RECT 107.300 74.500 108.570 74.510 ;
        RECT 107.100 74.160 111.940 74.500 ;
        RECT 107.300 74.120 108.570 74.160 ;
        RECT 110.810 73.740 111.990 73.790 ;
        RECT 107.110 73.400 111.990 73.740 ;
        RECT 110.810 73.370 111.990 73.400 ;
        RECT 107.300 72.920 108.580 72.930 ;
        RECT 107.110 72.580 111.950 72.920 ;
        RECT 107.300 72.570 108.580 72.580 ;
        RECT 89.390 71.890 96.380 72.460 ;
        RECT 98.820 71.710 105.810 72.280 ;
        RECT 110.790 72.130 111.990 72.140 ;
        RECT 107.100 71.790 111.990 72.130 ;
        RECT 110.790 71.780 111.990 71.790 ;
        RECT 90.230 71.080 96.930 71.650 ;
        RECT 98.270 70.900 104.970 71.470 ;
        RECT 89.390 67.840 96.380 68.410 ;
        RECT 98.820 67.650 105.810 68.220 ;
        RECT 90.230 67.030 96.930 67.600 ;
        RECT 98.270 66.840 104.970 67.410 ;
        RECT 89.390 63.790 96.380 64.360 ;
        RECT 98.820 63.590 105.810 64.160 ;
        RECT 90.230 62.980 96.930 63.550 ;
        RECT 98.270 62.780 104.970 63.350 ;
        RECT 101.685 61.200 102.385 62.070 ;
        RECT 89.390 59.740 96.380 60.310 ;
        RECT 90.230 58.930 96.930 59.500 ;
        RECT 98.820 59.050 105.810 59.620 ;
        RECT 98.270 58.240 104.970 58.810 ;
        RECT 89.390 55.690 96.380 56.260 ;
        RECT 90.230 54.880 96.930 55.450 ;
        RECT 105.810 53.260 107.100 54.540 ;
        RECT 89.390 51.640 96.380 52.210 ;
        RECT 90.230 50.830 96.930 51.400 ;
        RECT 89.390 47.590 96.380 48.160 ;
        RECT 90.230 46.780 96.930 47.350 ;
        RECT 89.390 43.540 96.380 44.110 ;
        RECT 90.230 42.730 96.930 43.300 ;
        RECT 89.390 39.490 96.380 40.060 ;
        RECT 90.230 38.680 96.930 39.250 ;
        RECT 89.390 35.440 96.380 36.010 ;
        RECT 90.230 34.630 96.930 35.200 ;
        RECT 89.390 31.390 96.380 31.960 ;
        RECT 90.230 30.580 96.930 31.150 ;
        RECT 89.390 27.305 96.380 27.875 ;
        RECT 90.230 26.495 96.930 27.065 ;
        RECT 89.390 23.180 96.380 23.750 ;
        RECT 90.230 22.370 96.930 22.940 ;
        RECT 92.815 20.830 93.515 21.790 ;
        RECT 89.390 18.625 96.380 19.195 ;
        RECT 90.230 17.815 96.930 18.385 ;
      LAYER via2 ;
        RECT 96.920 148.310 98.670 150.440 ;
        RECT 87.920 143.230 88.630 146.590 ;
        RECT 92.895 145.815 93.445 146.580 ;
        RECT 101.765 145.960 102.325 146.550 ;
        RECT 108.175 146.425 109.105 147.355 ;
        RECT 122.830 146.410 123.990 147.290 ;
        RECT 107.410 143.760 108.070 144.630 ;
        RECT 112.700 144.090 113.530 144.400 ;
        RECT 115.310 143.440 116.300 144.320 ;
        RECT 120.210 144.310 121.450 144.700 ;
        RECT 127.210 144.410 128.970 144.760 ;
        RECT 108.650 142.800 109.500 143.170 ;
        RECT 117.050 142.550 117.520 143.270 ;
        RECT 124.050 142.530 124.500 143.320 ;
        RECT 129.940 143.320 130.720 144.230 ;
        RECT 112.680 141.520 113.510 141.830 ;
        RECT 127.350 141.470 128.880 142.110 ;
        RECT 118.040 141.050 119.430 141.400 ;
        RECT 120.190 140.890 121.450 141.370 ;
        RECT 125.060 140.910 126.640 141.260 ;
        RECT 108.670 140.240 109.530 140.580 ;
        RECT 122.220 139.510 122.510 140.360 ;
        RECT 112.680 138.930 113.510 139.240 ;
        RECT 118.180 138.860 119.310 139.360 ;
        RECT 108.680 137.700 109.530 138.000 ;
        RECT 112.700 137.770 113.510 138.430 ;
        RECT 117.070 137.700 117.520 138.400 ;
        RECT 120.250 138.300 121.490 138.690 ;
        RECT 127.190 138.420 128.960 138.720 ;
        RECT 112.730 136.400 113.520 136.690 ;
        RECT 117.070 136.530 117.540 137.250 ;
        RECT 124.030 136.500 124.530 137.280 ;
        RECT 122.180 135.460 122.500 136.360 ;
        RECT 108.670 135.080 109.520 135.440 ;
        RECT 118.080 135.060 119.410 135.360 ;
        RECT 106.980 133.780 107.980 134.980 ;
        RECT 123.090 135.120 123.740 135.820 ;
        RECT 125.030 134.910 126.610 135.260 ;
        RECT 112.690 133.800 113.500 134.110 ;
        RECT 114.020 133.530 114.630 134.230 ;
        RECT 120.350 133.670 121.420 134.180 ;
        RECT 125.050 133.900 126.190 134.250 ;
        RECT 107.010 131.060 107.980 131.940 ;
        RECT 115.440 131.200 116.430 131.650 ;
        RECT 127.780 131.520 131.830 133.190 ;
        RECT 107.030 127.320 107.990 128.240 ;
        RECT 120.630 127.790 121.660 128.830 ;
        RECT 125.310 126.790 125.770 128.610 ;
        RECT 107.390 124.790 108.430 125.070 ;
        RECT 110.850 124.000 111.960 124.280 ;
        RECT 113.900 123.860 114.820 125.090 ;
        RECT 115.380 124.580 116.510 124.860 ;
        RECT 118.990 123.750 119.960 124.040 ;
        RECT 107.450 123.200 108.490 123.480 ;
        RECT 115.390 123.040 116.530 123.320 ;
        RECT 110.860 122.370 111.930 122.650 ;
        RECT 119.000 122.170 119.980 122.460 ;
        RECT 107.390 121.600 108.500 121.880 ;
        RECT 115.390 121.450 116.530 121.730 ;
        RECT 110.850 120.830 111.980 121.110 ;
        RECT 118.970 120.620 119.970 120.910 ;
        RECT 107.350 120.030 108.480 120.310 ;
        RECT 115.390 119.840 116.530 120.120 ;
        RECT 110.850 119.200 111.890 119.490 ;
        RECT 118.970 119.030 120.020 119.370 ;
        RECT 107.350 118.430 108.510 118.730 ;
        RECT 115.370 118.260 116.540 118.550 ;
        RECT 110.850 117.630 111.860 117.920 ;
        RECT 118.970 117.460 120.000 117.800 ;
        RECT 107.360 116.850 108.520 117.130 ;
        RECT 115.370 116.710 116.540 117.000 ;
        RECT 110.850 116.050 111.870 116.330 ;
        RECT 119.000 115.890 119.960 116.200 ;
        RECT 107.370 115.290 108.520 115.580 ;
        RECT 115.380 115.090 116.540 115.370 ;
        RECT 110.850 114.490 111.870 114.770 ;
        RECT 118.980 114.310 119.940 114.630 ;
        RECT 107.360 113.680 108.530 113.960 ;
        RECT 115.370 113.510 116.530 113.790 ;
        RECT 110.850 112.890 111.870 113.170 ;
        RECT 107.360 112.090 108.520 112.370 ;
        RECT 110.850 111.350 111.910 111.630 ;
        RECT 107.340 110.530 108.520 110.820 ;
        RECT 110.840 109.740 111.910 110.020 ;
        RECT 116.005 107.285 116.395 107.675 ;
        RECT 112.700 106.170 113.530 106.480 ;
        RECT 120.210 106.390 121.450 106.780 ;
        RECT 127.210 106.490 128.970 106.840 ;
        RECT 108.650 104.880 109.500 105.250 ;
        RECT 117.050 104.630 117.520 105.350 ;
        RECT 124.050 104.610 124.500 105.400 ;
        RECT 129.940 105.400 130.720 106.310 ;
        RECT 112.680 103.600 113.510 103.910 ;
        RECT 127.350 103.550 128.880 104.190 ;
        RECT 118.040 103.130 119.430 103.480 ;
        RECT 120.190 102.970 121.450 103.450 ;
        RECT 125.060 102.990 126.640 103.340 ;
        RECT 107.180 101.310 107.630 102.500 ;
        RECT 108.670 102.320 109.530 102.660 ;
        RECT 122.220 101.590 122.510 102.440 ;
        RECT 112.680 101.010 113.510 101.320 ;
        RECT 118.180 100.940 119.310 101.440 ;
        RECT 108.680 99.780 109.530 100.080 ;
        RECT 112.700 99.850 113.510 100.510 ;
        RECT 117.070 99.780 117.520 100.480 ;
        RECT 120.250 100.380 121.490 100.770 ;
        RECT 127.190 100.500 128.960 100.800 ;
        RECT 112.730 98.480 113.520 98.770 ;
        RECT 117.070 98.610 117.540 99.330 ;
        RECT 124.030 98.580 124.530 99.360 ;
        RECT 122.180 97.540 122.500 98.440 ;
        RECT 108.670 97.160 109.520 97.520 ;
        RECT 118.080 97.140 119.410 97.440 ;
        RECT 106.980 95.860 107.980 97.060 ;
        RECT 123.090 97.200 123.740 97.900 ;
        RECT 125.030 96.990 126.610 97.340 ;
        RECT 112.690 95.880 113.500 96.190 ;
        RECT 114.020 95.610 114.630 96.310 ;
        RECT 120.350 95.750 121.420 96.260 ;
        RECT 125.050 95.980 126.190 96.330 ;
        RECT 107.010 93.140 107.980 94.020 ;
        RECT 115.440 93.280 116.430 93.730 ;
        RECT 127.780 93.600 131.830 95.270 ;
        RECT 107.030 89.400 107.990 90.320 ;
        RECT 120.630 89.870 121.660 90.910 ;
        RECT 125.310 88.870 125.770 90.690 ;
        RECT 107.390 86.870 108.430 87.150 ;
        RECT 110.850 86.080 111.960 86.360 ;
        RECT 113.900 85.940 114.820 87.170 ;
        RECT 115.380 86.660 116.510 86.940 ;
        RECT 118.990 85.830 119.960 86.120 ;
        RECT 107.450 85.280 108.490 85.560 ;
        RECT 115.390 85.120 116.530 85.400 ;
        RECT 110.860 84.450 111.930 84.730 ;
        RECT 119.000 84.250 119.980 84.540 ;
        RECT 107.390 83.680 108.500 83.960 ;
        RECT 115.390 83.530 116.530 83.810 ;
        RECT 110.850 82.910 111.980 83.190 ;
        RECT 118.970 82.700 119.970 82.990 ;
        RECT 107.350 82.110 108.480 82.390 ;
        RECT 115.390 81.920 116.530 82.200 ;
        RECT 122.660 82.590 124.190 84.000 ;
        RECT 110.850 81.280 111.890 81.570 ;
        RECT 118.970 81.110 120.020 81.450 ;
        RECT 107.350 80.510 108.510 80.810 ;
        RECT 115.370 80.340 116.540 80.630 ;
        RECT 110.850 79.710 111.860 80.000 ;
        RECT 118.970 79.540 120.000 79.880 ;
        RECT 107.360 78.930 108.520 79.210 ;
        RECT 115.370 78.790 116.540 79.080 ;
        RECT 110.850 78.130 111.870 78.410 ;
        RECT 119.000 77.970 119.960 78.280 ;
        RECT 107.370 77.370 108.520 77.660 ;
        RECT 115.380 77.170 116.540 77.450 ;
        RECT 110.850 76.570 111.870 76.850 ;
        RECT 118.980 76.390 119.940 76.710 ;
        RECT 107.360 75.760 108.530 76.040 ;
        RECT 115.370 75.590 116.530 75.870 ;
        RECT 110.850 74.970 111.870 75.250 ;
        RECT 107.360 74.170 108.520 74.450 ;
        RECT 110.850 73.430 111.910 73.710 ;
        RECT 107.340 72.610 108.520 72.900 ;
        RECT 110.840 71.820 111.910 72.100 ;
        RECT 101.755 61.250 102.325 62.020 ;
        RECT 105.965 53.400 106.945 54.380 ;
        RECT 92.870 20.910 93.455 21.680 ;
      LAYER met3 ;
        RECT 96.530 150.670 99.090 150.790 ;
        RECT 0.880 148.190 99.090 150.670 ;
        RECT 2.500 148.170 99.090 148.190 ;
        RECT 96.530 147.980 99.090 148.170 ;
        RECT 105.965 147.375 109.130 147.380 ;
        RECT 87.690 146.320 88.920 146.890 ;
        RECT 49.010 143.460 88.920 146.320 ;
        RECT 87.690 143.050 88.920 143.460 ;
        RECT 92.815 20.795 93.510 146.635 ;
        RECT 101.685 61.200 102.385 146.640 ;
        RECT 105.940 146.405 109.130 147.375 ;
        RECT 105.965 146.400 109.130 146.405 ;
        RECT 122.670 146.160 124.180 147.460 ;
        RECT 107.260 144.340 108.180 144.880 ;
        RECT 105.310 143.360 108.180 144.340 ;
        RECT 105.310 143.290 108.050 143.360 ;
        RECT 105.310 142.380 106.990 143.290 ;
        RECT 108.630 143.230 109.550 144.390 ;
        RECT 108.540 142.700 109.600 143.230 ;
        RECT 105.310 102.590 106.270 142.380 ;
        RECT 108.630 140.630 109.550 142.700 ;
        RECT 108.590 140.170 109.610 140.630 ;
        RECT 108.630 138.090 109.550 140.170 ;
        RECT 108.580 137.590 109.620 138.090 ;
        RECT 108.630 135.520 109.550 137.590 ;
        RECT 112.650 135.750 113.570 144.430 ;
        RECT 106.910 127.160 108.070 135.090 ;
        RECT 108.630 133.300 109.560 135.520 ;
        RECT 112.650 133.530 113.580 135.750 ;
        RECT 113.950 125.250 114.740 134.330 ;
        RECT 115.150 131.840 116.560 144.950 ;
        RECT 120.150 143.690 121.540 144.780 ;
        RECT 117.010 136.480 117.580 143.370 ;
        RECT 117.930 140.920 119.540 141.540 ;
        RECT 118.040 140.230 119.440 140.920 ;
        RECT 118.050 135.760 119.420 140.230 ;
        RECT 118.040 135.540 119.420 135.760 ;
        RECT 117.940 134.920 119.530 135.540 ;
        RECT 118.040 134.660 119.420 134.920 ;
        RECT 120.160 133.540 121.530 143.690 ;
        RECT 122.010 135.410 122.540 140.420 ;
        RECT 122.950 135.990 123.470 146.160 ;
        RECT 127.140 143.840 129.060 144.920 ;
        RECT 123.990 136.470 124.560 143.360 ;
        RECT 122.950 134.880 124.080 135.990 ;
        RECT 122.970 134.660 124.080 134.880 ;
        RECT 124.980 134.790 126.730 141.350 ;
        RECT 127.150 138.380 129.060 143.840 ;
        RECT 129.760 143.070 130.870 144.420 ;
        RECT 124.990 132.170 126.260 134.490 ;
        RECT 124.990 131.940 125.910 132.170 ;
        RECT 115.150 125.690 116.600 131.840 ;
        RECT 124.990 130.370 125.900 131.940 ;
        RECT 127.490 131.280 132.080 133.420 ;
        RECT 107.300 110.850 108.570 125.160 ;
        RECT 107.300 110.490 108.580 110.850 ;
        RECT 107.300 109.750 108.570 110.490 ;
        RECT 110.800 110.060 112.070 125.140 ;
        RECT 113.720 123.750 114.900 125.250 ;
        RECT 115.240 123.830 116.600 125.690 ;
        RECT 115.270 123.370 116.580 123.830 ;
        RECT 115.150 111.690 116.580 123.370 ;
        RECT 118.920 113.140 120.180 125.010 ;
        RECT 120.550 123.360 122.090 129.000 ;
        RECT 124.990 126.350 125.880 130.370 ;
        RECT 110.790 109.730 112.070 110.060 ;
        RECT 110.790 109.700 111.990 109.730 ;
        RECT 115.320 109.180 116.580 111.690 ;
        RECT 127.190 109.420 140.590 131.280 ;
        RECT 115.320 108.815 120.090 109.180 ;
        RECT 115.320 108.220 125.830 108.815 ;
        RECT 118.920 108.120 125.830 108.220 ;
        RECT 115.980 107.260 116.420 107.700 ;
        RECT 118.920 107.645 144.035 108.120 ;
        RECT 125.370 107.340 144.030 107.645 ;
        RECT 108.630 105.310 109.550 106.470 ;
        RECT 108.540 104.780 109.600 105.310 ;
        RECT 108.630 102.710 109.550 104.780 ;
        RECT 105.310 101.220 107.760 102.590 ;
        RECT 108.590 102.250 109.610 102.710 ;
        RECT 105.310 98.720 106.270 101.220 ;
        RECT 108.630 100.170 109.550 102.250 ;
        RECT 108.580 99.670 109.620 100.170 ;
        RECT 108.630 97.600 109.550 99.670 ;
        RECT 112.650 97.830 113.570 106.510 ;
        RECT 106.910 89.240 108.070 97.170 ;
        RECT 108.630 95.380 109.560 97.600 ;
        RECT 112.650 95.610 113.580 97.830 ;
        RECT 113.950 87.330 114.740 96.410 ;
        RECT 116.005 93.920 116.395 107.260 ;
        RECT 120.150 105.770 121.540 106.860 ;
        RECT 127.140 105.920 129.060 107.000 ;
        RECT 132.050 106.870 144.030 107.340 ;
        RECT 117.010 98.560 117.580 105.450 ;
        RECT 117.930 103.000 119.540 103.620 ;
        RECT 118.040 102.310 119.440 103.000 ;
        RECT 118.050 97.840 119.420 102.310 ;
        RECT 118.040 97.620 119.420 97.840 ;
        RECT 117.940 97.000 119.530 97.620 ;
        RECT 118.040 96.740 119.420 97.000 ;
        RECT 120.160 95.620 121.530 105.770 ;
        RECT 122.010 97.490 122.540 102.500 ;
        RECT 123.990 98.550 124.560 105.440 ;
        RECT 122.970 97.410 124.080 98.070 ;
        RECT 107.300 72.930 108.570 87.240 ;
        RECT 107.300 72.570 108.580 72.930 ;
        RECT 107.300 71.830 108.570 72.570 ;
        RECT 110.800 72.140 112.070 87.220 ;
        RECT 113.720 85.830 114.900 87.330 ;
        RECT 115.240 85.910 116.600 93.920 ;
        RECT 110.790 71.810 112.070 72.140 ;
        RECT 110.790 71.780 111.990 71.810 ;
        RECT 115.320 66.480 116.580 85.910 ;
        RECT 118.920 75.220 120.180 87.090 ;
        RECT 120.550 85.440 122.090 91.080 ;
        RECT 122.890 84.310 124.300 97.410 ;
        RECT 124.980 96.870 126.730 103.430 ;
        RECT 127.150 100.460 129.060 105.920 ;
        RECT 129.760 105.150 130.870 106.500 ;
        RECT 124.990 94.250 126.260 96.570 ;
        RECT 124.990 94.020 125.910 94.250 ;
        RECT 124.990 92.450 125.900 94.020 ;
        RECT 127.490 93.360 132.080 95.500 ;
        RECT 124.990 88.430 125.880 92.450 ;
        RECT 122.440 82.380 124.340 84.310 ;
        RECT 127.190 71.500 140.590 93.360 ;
        RECT 105.810 53.260 107.100 54.540 ;
        RECT 115.350 8.130 116.550 66.480 ;
        RECT 134.200 11.670 135.430 11.770 ;
        RECT 142.875 11.670 144.030 106.870 ;
        RECT 132.800 10.515 144.030 11.670 ;
        RECT 132.800 10.490 143.220 10.515 ;
        RECT 134.200 10.370 135.430 10.490 ;
        RECT 156.110 8.130 157.380 8.210 ;
        RECT 115.350 6.930 158.390 8.130 ;
        RECT 156.110 6.810 157.380 6.930 ;
      LAYER via3 ;
        RECT 1.210 148.360 2.330 150.490 ;
        RECT 49.200 143.590 50.240 146.090 ;
        RECT 105.970 146.405 106.940 147.375 ;
        RECT 127.740 131.500 131.850 133.280 ;
        RECT 127.330 130.860 140.450 131.180 ;
        RECT 120.780 123.560 121.930 124.440 ;
        RECT 120.780 85.640 121.930 86.520 ;
        RECT 127.740 93.580 131.850 95.360 ;
        RECT 127.330 92.940 140.450 93.260 ;
        RECT 105.940 53.375 106.970 54.405 ;
        RECT 134.420 10.540 135.160 11.530 ;
        RECT 156.340 7.050 157.110 7.980 ;
      LAYER met4 ;
        RECT 3.990 223.220 4.290 224.760 ;
        RECT 7.670 223.220 7.970 224.760 ;
        RECT 11.350 223.220 11.650 224.760 ;
        RECT 15.030 223.220 15.330 224.760 ;
        RECT 18.710 223.220 19.010 224.760 ;
        RECT 22.390 223.220 22.690 224.760 ;
        RECT 26.070 223.220 26.370 224.760 ;
        RECT 29.750 223.220 30.050 224.760 ;
        RECT 33.430 223.220 33.730 224.760 ;
        RECT 37.110 223.220 37.410 224.760 ;
        RECT 40.790 223.220 41.090 224.760 ;
        RECT 44.470 223.220 44.770 224.760 ;
        RECT 48.150 223.220 48.450 224.760 ;
        RECT 51.830 223.220 52.130 224.760 ;
        RECT 55.510 223.220 55.810 224.760 ;
        RECT 59.190 223.220 59.490 224.760 ;
        RECT 62.870 223.220 63.170 224.760 ;
        RECT 66.550 223.220 66.850 224.760 ;
        RECT 70.230 223.220 70.530 224.760 ;
        RECT 73.910 223.220 74.210 224.760 ;
        RECT 77.590 223.220 77.890 224.760 ;
        RECT 81.270 223.220 81.570 224.760 ;
        RECT 84.950 223.220 85.250 224.760 ;
        RECT 88.630 223.220 88.930 224.760 ;
        RECT 2.970 221.620 89.590 223.220 ;
        RECT 49.000 220.760 50.500 221.620 ;
        RECT 105.965 54.410 106.945 147.380 ;
        RECT 127.490 131.460 132.040 133.470 ;
        RECT 127.490 131.260 140.560 131.460 ;
        RECT 127.250 130.800 140.560 131.260 ;
        RECT 127.250 130.780 140.530 130.800 ;
        RECT 127.580 124.640 140.200 129.430 ;
        RECT 124.660 124.620 140.200 124.640 ;
        RECT 120.600 123.400 140.200 124.620 ;
        RECT 124.660 121.850 140.200 123.400 ;
        RECT 127.580 109.810 140.200 121.850 ;
        RECT 127.490 93.540 132.040 95.550 ;
        RECT 127.490 93.340 140.560 93.540 ;
        RECT 127.250 92.880 140.560 93.340 ;
        RECT 127.250 92.860 140.530 92.880 ;
        RECT 127.580 86.720 140.200 91.510 ;
        RECT 124.660 86.700 140.200 86.720 ;
        RECT 120.600 85.480 140.200 86.700 ;
        RECT 124.660 83.930 140.200 85.480 ;
        RECT 127.580 71.890 140.200 83.930 ;
        RECT 105.935 53.370 106.975 54.410 ;
        RECT 134.200 10.370 135.430 11.770 ;
        RECT 134.345 2.495 135.220 10.370 ;
        RECT 156.110 6.810 157.380 8.210 ;
        RECT 134.355 1.000 135.205 2.495 ;
        RECT 156.535 1.000 157.130 6.810 ;
  END
END tt_um_devinatkin_dual_oscillator
END LIBRARY

