VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_rejunity_ay8913
  CLASS BLOCK ;
  FOREIGN tt_um_rejunity_ay8913 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.148600 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.148600 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 13.148600 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1077.790771 ;
    ANTENNADIFFAREA 991.837952 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 9.000 5.000 10.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 22.835 209.135 23.005 209.325 ;
        RECT 31.575 209.135 31.745 209.325 ;
        RECT 32.035 209.135 32.205 209.325 ;
        RECT 36.175 209.135 36.345 209.325 ;
        RECT 38.010 209.185 38.130 209.295 ;
        RECT 39.395 209.135 39.565 209.325 ;
        RECT 39.855 209.135 40.025 209.325 ;
        RECT 45.375 209.135 45.545 209.325 ;
        RECT 48.130 209.185 48.250 209.295 ;
        RECT 49.050 209.185 49.170 209.295 ;
        RECT 50.435 209.135 50.605 209.325 ;
        RECT 50.895 209.135 51.065 209.325 ;
        RECT 56.410 209.185 56.530 209.295 ;
        RECT 57.795 209.135 57.965 209.325 ;
        RECT 58.255 209.135 58.425 209.325 ;
        RECT 61.010 209.185 61.130 209.295 ;
        RECT 62.855 209.135 63.025 209.325 ;
        RECT 63.325 209.180 63.485 209.290 ;
        RECT 64.245 209.135 64.415 209.325 ;
        RECT 65.615 209.135 65.785 209.325 ;
        RECT 67.455 209.135 67.625 209.325 ;
        RECT 73.895 209.135 74.065 209.325 ;
        RECT 74.815 209.135 74.985 209.325 ;
        RECT 79.415 209.135 79.585 209.325 ;
        RECT 79.875 209.135 80.045 209.325 ;
        RECT 82.640 209.135 82.810 209.325 ;
        RECT 83.095 209.135 83.265 209.325 ;
        RECT 86.770 209.185 86.890 209.295 ;
        RECT 90.915 209.135 91.085 209.325 ;
        RECT 91.375 209.135 91.545 209.325 ;
        RECT 93.210 209.185 93.330 209.295 ;
        RECT 93.675 209.135 93.845 209.325 ;
        RECT 96.435 209.135 96.605 209.325 ;
        RECT 96.895 209.135 97.065 209.325 ;
        RECT 99.650 209.185 99.770 209.295 ;
        RECT 100.570 209.185 100.690 209.295 ;
        RECT 101.035 209.135 101.205 209.325 ;
        RECT 102.415 209.135 102.585 209.325 ;
        RECT 104.250 209.185 104.370 209.295 ;
        RECT 104.715 209.135 104.885 209.325 ;
        RECT 106.095 209.135 106.265 209.325 ;
        RECT 107.930 209.185 108.050 209.295 ;
        RECT 109.775 209.135 109.945 209.325 ;
        RECT 110.235 209.135 110.405 209.325 ;
        RECT 111.615 209.135 111.785 209.325 ;
        RECT 113.455 209.135 113.625 209.325 ;
        RECT 118.975 209.135 119.145 209.325 ;
        RECT 119.435 209.135 119.605 209.325 ;
        RECT 124.495 209.135 124.665 209.325 ;
        RECT 124.965 209.180 125.125 209.290 ;
        RECT 127.715 209.135 127.885 209.325 ;
        RECT 128.175 209.135 128.345 209.325 ;
        RECT 131.855 209.135 132.025 209.325 ;
        RECT 138.295 209.135 138.465 209.325 ;
        RECT 139.215 209.135 139.385 209.325 ;
        RECT 141.055 209.135 141.225 209.325 ;
        RECT 146.575 209.135 146.745 209.325 ;
        RECT 150.255 209.135 150.425 209.325 ;
        RECT 152.090 209.185 152.210 209.295 ;
        RECT 153.465 209.135 153.635 209.325 ;
        RECT 153.935 209.135 154.105 209.325 ;
        RECT 156.695 209.135 156.865 209.325 ;
        RECT 22.695 208.325 24.065 209.135 ;
        RECT 24.155 208.455 31.885 209.135 ;
        RECT 24.155 208.225 25.925 208.455 ;
        RECT 27.460 208.235 28.370 208.455 ;
        RECT 31.895 208.325 35.565 209.135 ;
        RECT 35.585 208.265 36.015 209.050 ;
        RECT 36.035 208.325 37.865 209.135 ;
        RECT 38.335 208.355 39.705 209.135 ;
        RECT 39.715 208.325 45.225 209.135 ;
        RECT 45.235 208.325 47.985 209.135 ;
        RECT 48.465 208.265 48.895 209.050 ;
        RECT 49.375 208.355 50.745 209.135 ;
        RECT 50.755 208.325 56.265 209.135 ;
        RECT 56.735 208.355 58.105 209.135 ;
        RECT 58.115 208.325 60.865 209.135 ;
        RECT 61.345 208.265 61.775 209.050 ;
        RECT 61.805 208.225 63.155 209.135 ;
        RECT 64.095 208.355 65.465 209.135 ;
        RECT 65.475 208.325 67.305 209.135 ;
        RECT 67.315 208.225 70.525 209.135 ;
        RECT 70.630 208.455 74.095 209.135 ;
        RECT 70.630 208.225 71.550 208.455 ;
        RECT 74.225 208.265 74.655 209.050 ;
        RECT 74.675 208.355 76.045 209.135 ;
        RECT 76.150 208.455 79.615 209.135 ;
        RECT 79.735 208.455 81.565 209.135 ;
        RECT 76.150 208.225 77.070 208.455 ;
        RECT 80.220 208.225 81.565 208.455 ;
        RECT 81.575 208.225 82.925 209.135 ;
        RECT 82.955 208.325 86.625 209.135 ;
        RECT 87.105 208.265 87.535 209.050 ;
        RECT 87.650 208.455 91.115 209.135 ;
        RECT 91.235 208.455 93.065 209.135 ;
        RECT 93.535 208.455 95.365 209.135 ;
        RECT 87.650 208.225 88.570 208.455 ;
        RECT 91.720 208.225 93.065 208.455 ;
        RECT 94.020 208.225 95.365 208.455 ;
        RECT 95.375 208.355 96.745 209.135 ;
        RECT 96.755 208.325 99.505 209.135 ;
        RECT 99.985 208.265 100.415 209.050 ;
        RECT 100.895 208.355 102.265 209.135 ;
        RECT 102.275 208.325 104.105 209.135 ;
        RECT 104.575 208.355 105.945 209.135 ;
        RECT 105.955 208.325 107.785 209.135 ;
        RECT 108.255 208.455 110.085 209.135 ;
        RECT 110.095 208.355 111.465 209.135 ;
        RECT 111.475 208.325 112.845 209.135 ;
        RECT 112.865 208.265 113.295 209.050 ;
        RECT 113.315 208.325 116.065 209.135 ;
        RECT 116.075 208.225 119.285 209.135 ;
        RECT 119.295 208.455 121.125 209.135 ;
        RECT 121.230 208.455 124.695 209.135 ;
        RECT 121.230 208.225 122.150 208.455 ;
        RECT 125.745 208.265 126.175 209.050 ;
        RECT 126.195 208.455 128.025 209.135 ;
        RECT 128.145 208.455 131.610 209.135 ;
        RECT 131.825 208.455 135.290 209.135 ;
        RECT 126.195 208.225 127.540 208.455 ;
        RECT 130.690 208.225 131.610 208.455 ;
        RECT 134.370 208.225 135.290 208.455 ;
        RECT 135.395 208.225 138.605 209.135 ;
        RECT 138.625 208.265 139.055 209.050 ;
        RECT 139.075 208.455 140.905 209.135 ;
        RECT 139.560 208.225 140.905 208.455 ;
        RECT 140.915 208.325 146.425 209.135 ;
        RECT 146.435 208.325 150.105 209.135 ;
        RECT 150.115 208.325 151.485 209.135 ;
        RECT 151.505 208.265 151.935 209.050 ;
        RECT 152.415 208.355 153.785 209.135 ;
        RECT 153.795 208.325 155.625 209.135 ;
        RECT 155.635 208.325 157.005 209.135 ;
      LAYER nwell ;
        RECT 22.500 205.105 157.200 207.935 ;
      LAYER pwell ;
        RECT 22.695 203.905 24.065 204.715 ;
        RECT 24.075 203.905 27.745 204.715 ;
        RECT 31.270 204.585 32.180 204.805 ;
        RECT 33.715 204.585 35.485 204.815 ;
        RECT 27.755 203.905 35.485 204.585 ;
        RECT 35.585 203.990 36.015 204.775 ;
        RECT 40.010 204.585 40.920 204.805 ;
        RECT 42.455 204.585 43.805 204.815 ;
        RECT 45.675 204.585 46.605 204.815 ;
        RECT 36.495 203.905 43.805 204.585 ;
        RECT 43.855 203.905 46.605 204.585 ;
        RECT 46.615 204.615 47.560 204.815 ;
        RECT 46.615 203.935 49.365 204.615 ;
        RECT 46.615 203.905 47.560 203.935 ;
        RECT 22.835 203.695 23.005 203.905 ;
        RECT 24.215 203.695 24.385 203.905 ;
        RECT 27.895 203.715 28.065 203.905 ;
        RECT 29.735 203.695 29.905 203.885 ;
        RECT 36.170 203.745 36.290 203.855 ;
        RECT 36.635 203.715 36.805 203.905 ;
        RECT 22.695 202.885 24.065 203.695 ;
        RECT 24.075 202.885 29.585 203.695 ;
        RECT 29.595 203.015 37.325 203.695 ;
        RECT 37.560 203.665 37.730 203.885 ;
        RECT 40.770 203.745 40.890 203.855 ;
        RECT 41.230 203.695 41.400 203.885 ;
        RECT 42.615 203.715 42.785 203.885 ;
        RECT 43.995 203.715 44.165 203.905 ;
        RECT 49.050 203.885 49.220 203.935 ;
        RECT 49.375 203.905 50.745 204.685 ;
        RECT 54.270 204.585 55.180 204.805 ;
        RECT 56.715 204.585 58.065 204.815 ;
        RECT 50.755 203.905 58.065 204.585 ;
        RECT 58.115 204.585 59.045 204.815 ;
        RECT 58.115 203.905 60.865 204.585 ;
        RECT 61.345 203.990 61.775 204.775 ;
        RECT 62.755 204.585 64.105 204.815 ;
        RECT 65.640 204.585 66.550 204.805 ;
        RECT 70.575 204.585 71.925 204.815 ;
        RECT 73.460 204.585 74.370 204.805 ;
        RECT 81.410 204.585 82.320 204.805 ;
        RECT 83.855 204.585 85.205 204.815 ;
        RECT 62.755 203.905 70.065 204.585 ;
        RECT 70.575 203.905 77.885 204.585 ;
        RECT 77.895 203.905 85.205 204.585 ;
        RECT 85.275 203.905 86.625 204.815 ;
        RECT 87.105 203.990 87.535 204.775 ;
        RECT 87.555 203.905 88.925 204.715 ;
        RECT 92.450 204.585 93.360 204.805 ;
        RECT 94.895 204.585 96.245 204.815 ;
        RECT 88.935 203.905 96.245 204.585 ;
        RECT 96.305 203.905 97.655 204.815 ;
        RECT 98.595 204.615 99.540 204.815 ;
        RECT 100.875 204.615 101.805 204.815 ;
        RECT 98.595 204.135 101.805 204.615 ;
        RECT 98.595 203.935 101.665 204.135 ;
        RECT 98.595 203.905 99.540 203.935 ;
        RECT 42.620 203.695 42.785 203.715 ;
        RECT 44.915 203.695 45.085 203.885 ;
        RECT 48.130 203.745 48.250 203.855 ;
        RECT 49.050 203.715 49.225 203.885 ;
        RECT 49.515 203.715 49.685 203.905 ;
        RECT 50.895 203.715 51.065 203.905 ;
        RECT 49.075 203.695 49.225 203.715 ;
        RECT 51.355 203.695 51.525 203.885 ;
        RECT 54.120 203.695 54.290 203.885 ;
        RECT 56.420 203.695 56.590 203.885 ;
        RECT 60.555 203.715 60.725 203.905 ;
        RECT 61.945 203.855 62.105 203.860 ;
        RECT 61.010 203.745 61.130 203.855 ;
        RECT 61.930 203.750 62.105 203.855 ;
        RECT 61.930 203.745 62.050 203.750 ;
        RECT 63.315 203.695 63.485 203.885 ;
        RECT 63.775 203.695 63.945 203.885 ;
        RECT 68.375 203.695 68.545 203.885 ;
        RECT 68.835 203.695 69.005 203.885 ;
        RECT 69.755 203.715 69.925 203.905 ;
        RECT 70.215 203.855 70.385 203.885 ;
        RECT 70.210 203.745 70.385 203.855 ;
        RECT 70.215 203.695 70.385 203.745 ;
        RECT 73.445 203.740 73.605 203.850 ;
        RECT 74.815 203.695 74.985 203.885 ;
        RECT 77.575 203.715 77.745 203.905 ;
        RECT 78.035 203.715 78.205 203.905 ;
        RECT 82.180 203.695 82.350 203.885 ;
        RECT 85.390 203.715 85.560 203.905 ;
        RECT 86.770 203.745 86.890 203.855 ;
        RECT 87.695 203.715 87.865 203.905 ;
        RECT 89.075 203.715 89.245 203.905 ;
        RECT 90.000 203.695 90.170 203.885 ;
        RECT 90.450 203.745 90.570 203.855 ;
        RECT 90.910 203.695 91.080 203.885 ;
        RECT 92.295 203.715 92.465 203.885 ;
        RECT 92.300 203.695 92.465 203.715 ;
        RECT 94.595 203.695 94.765 203.885 ;
        RECT 96.905 203.740 97.065 203.850 ;
        RECT 97.355 203.715 97.525 203.905 ;
        RECT 97.815 203.695 97.985 203.885 ;
        RECT 100.575 203.695 100.745 203.885 ;
        RECT 101.495 203.715 101.665 203.935 ;
        RECT 101.815 203.905 104.425 204.815 ;
        RECT 105.075 204.585 106.425 204.815 ;
        RECT 107.960 204.585 108.870 204.805 ;
        RECT 105.075 203.905 112.385 204.585 ;
        RECT 112.865 203.990 113.295 204.775 ;
        RECT 113.315 203.905 116.065 204.715 ;
        RECT 120.050 204.585 120.960 204.805 ;
        RECT 122.495 204.585 123.845 204.815 ;
        RECT 124.380 204.585 125.725 204.815 ;
        RECT 129.710 204.585 130.620 204.805 ;
        RECT 132.155 204.585 133.505 204.815 ;
        RECT 116.535 203.905 123.845 204.585 ;
        RECT 123.895 203.905 125.725 204.585 ;
        RECT 126.195 203.905 133.505 204.585 ;
        RECT 133.555 203.905 136.765 204.815 ;
        RECT 136.785 203.905 138.135 204.815 ;
        RECT 138.625 203.990 139.055 204.775 ;
        RECT 139.075 204.585 140.210 204.815 ;
        RECT 139.075 203.905 142.285 204.585 ;
        RECT 142.315 203.905 143.665 204.815 ;
        RECT 143.685 203.905 145.035 204.815 ;
        RECT 145.055 203.905 150.565 204.715 ;
        RECT 150.575 203.905 154.245 204.715 ;
        RECT 154.255 203.905 155.625 204.715 ;
        RECT 155.635 203.905 157.005 204.715 ;
        RECT 101.960 203.715 102.130 203.905 ;
        RECT 104.710 203.745 104.830 203.855 ;
        RECT 39.690 203.665 40.625 203.695 ;
        RECT 37.560 203.465 40.625 203.665 ;
        RECT 33.110 202.795 34.020 203.015 ;
        RECT 35.555 202.785 37.325 203.015 ;
        RECT 37.415 202.985 40.625 203.465 ;
        RECT 37.415 202.785 38.345 202.985 ;
        RECT 39.675 202.785 40.625 202.985 ;
        RECT 41.115 202.785 42.465 203.695 ;
        RECT 42.620 203.015 44.455 203.695 ;
        RECT 43.525 202.785 44.455 203.015 ;
        RECT 44.875 202.785 47.985 203.695 ;
        RECT 48.465 202.825 48.895 203.610 ;
        RECT 49.075 202.875 51.005 203.695 ;
        RECT 51.215 202.885 53.965 203.695 ;
        RECT 50.055 202.785 51.005 202.875 ;
        RECT 53.975 202.785 56.265 203.695 ;
        RECT 56.275 202.785 61.595 203.695 ;
        RECT 62.265 202.785 63.615 203.695 ;
        RECT 63.745 203.015 67.210 203.695 ;
        RECT 66.290 202.785 67.210 203.015 ;
        RECT 67.325 202.785 68.675 203.695 ;
        RECT 68.695 202.885 70.065 203.695 ;
        RECT 70.075 202.785 73.285 203.695 ;
        RECT 74.225 202.825 74.655 203.610 ;
        RECT 74.675 203.015 81.985 203.695 ;
        RECT 82.035 203.015 86.165 203.695 ;
        RECT 78.190 202.795 79.100 203.015 ;
        RECT 80.635 202.785 81.985 203.015 ;
        RECT 84.775 202.785 86.165 203.015 ;
        RECT 86.175 202.785 90.280 203.695 ;
        RECT 90.795 202.785 92.145 203.695 ;
        RECT 92.300 203.015 94.135 203.695 ;
        RECT 94.455 203.015 96.745 203.695 ;
        RECT 97.675 203.015 99.965 203.695 ;
        RECT 93.205 202.785 94.135 203.015 ;
        RECT 95.825 202.785 96.745 203.015 ;
        RECT 99.045 202.785 99.965 203.015 ;
        RECT 99.985 202.825 100.415 203.610 ;
        RECT 100.435 203.015 103.645 203.695 ;
        RECT 102.510 202.785 103.645 203.015 ;
        RECT 103.655 203.665 104.590 203.695 ;
        RECT 106.550 203.665 106.720 203.885 ;
        RECT 107.010 203.745 107.130 203.855 ;
        RECT 112.075 203.715 112.245 203.905 ;
        RECT 112.530 203.745 112.650 203.855 ;
        RECT 113.455 203.715 113.625 203.905 ;
        RECT 114.375 203.695 114.545 203.885 ;
        RECT 114.835 203.695 115.005 203.885 ;
        RECT 116.675 203.855 116.845 203.905 ;
        RECT 116.210 203.745 116.330 203.855 ;
        RECT 116.670 203.745 116.845 203.855 ;
        RECT 116.675 203.715 116.845 203.745 ;
        RECT 117.135 203.695 117.305 203.885 ;
        RECT 124.035 203.715 124.205 203.905 ;
        RECT 124.495 203.695 124.665 203.885 ;
        RECT 125.870 203.745 125.990 203.855 ;
        RECT 126.335 203.715 126.505 203.905 ;
        RECT 133.235 203.695 133.405 203.885 ;
        RECT 133.700 203.695 133.870 203.885 ;
        RECT 136.455 203.715 136.625 203.905 ;
        RECT 136.915 203.715 137.085 203.905 ;
        RECT 137.375 203.715 137.545 203.885 ;
        RECT 138.290 203.745 138.410 203.855 ;
        RECT 137.385 203.695 137.545 203.715 ;
        RECT 141.520 203.695 141.690 203.885 ;
        RECT 141.975 203.715 142.145 203.905 ;
        RECT 142.430 203.715 142.600 203.905 ;
        RECT 144.735 203.715 144.905 203.905 ;
        RECT 145.195 203.715 145.365 203.905 ;
        RECT 103.655 203.465 106.720 203.665 ;
        RECT 103.655 202.985 106.865 203.465 ;
        RECT 103.655 202.785 104.605 202.985 ;
        RECT 105.935 202.785 106.865 202.985 ;
        RECT 107.375 203.015 114.685 203.695 ;
        RECT 107.375 202.785 108.725 203.015 ;
        RECT 110.260 202.795 111.170 203.015 ;
        RECT 114.695 202.885 116.525 203.695 ;
        RECT 116.995 203.015 124.305 203.695 ;
        RECT 120.510 202.795 121.420 203.015 ;
        RECT 122.955 202.785 124.305 203.015 ;
        RECT 124.355 202.885 125.725 203.695 ;
        RECT 125.745 202.825 126.175 203.610 ;
        RECT 126.235 203.015 133.545 203.695 ;
        RECT 133.555 203.015 137.225 203.695 ;
        RECT 126.235 202.785 127.585 203.015 ;
        RECT 129.120 202.795 130.030 203.015 ;
        RECT 133.555 202.785 134.480 203.015 ;
        RECT 137.385 202.785 141.040 203.695 ;
        RECT 141.375 203.015 145.045 203.695 ;
        RECT 145.055 203.665 146.000 203.695 ;
        RECT 147.490 203.665 147.660 203.885 ;
        RECT 147.955 203.695 148.125 203.885 ;
        RECT 150.715 203.715 150.885 203.905 ;
        RECT 152.095 203.695 152.265 203.885 ;
        RECT 154.395 203.715 154.565 203.905 ;
        RECT 156.695 203.695 156.865 203.905 ;
        RECT 141.375 202.785 142.300 203.015 ;
        RECT 145.055 202.985 147.805 203.665 ;
        RECT 145.055 202.785 146.000 202.985 ;
        RECT 147.815 202.885 151.485 203.695 ;
        RECT 151.505 202.825 151.935 203.610 ;
        RECT 151.955 202.885 155.625 203.695 ;
        RECT 155.635 202.885 157.005 203.695 ;
      LAYER nwell ;
        RECT 22.500 199.665 157.200 202.495 ;
      LAYER pwell ;
        RECT 22.695 198.465 24.065 199.275 ;
        RECT 24.075 198.465 29.585 199.275 ;
        RECT 29.595 198.465 35.105 199.275 ;
        RECT 35.585 198.550 36.015 199.335 ;
        RECT 36.035 198.465 37.865 199.275 ;
        RECT 38.335 198.465 39.685 199.375 ;
        RECT 40.645 198.465 41.995 199.375 ;
        RECT 42.015 198.465 43.365 199.375 ;
        RECT 45.225 199.145 46.145 199.375 ;
        RECT 43.855 198.465 46.145 199.145 ;
        RECT 46.155 198.465 47.525 199.245 ;
        RECT 47.535 198.465 51.205 199.275 ;
        RECT 51.675 198.465 54.885 199.375 ;
        RECT 54.895 198.465 58.105 199.375 ;
        RECT 58.115 198.465 61.325 199.375 ;
        RECT 61.345 198.550 61.775 199.335 ;
        RECT 61.795 198.465 63.165 199.275 ;
        RECT 63.175 198.465 66.385 199.375 ;
        RECT 66.480 198.465 75.585 199.145 ;
        RECT 75.595 198.465 78.345 199.275 ;
        RECT 78.355 198.465 81.565 199.375 ;
        RECT 81.670 199.145 82.590 199.375 ;
        RECT 81.670 198.465 85.135 199.145 ;
        RECT 85.255 198.465 87.085 199.275 ;
        RECT 87.105 198.550 87.535 199.335 ;
        RECT 87.565 199.145 89.525 199.375 ;
        RECT 87.565 198.465 90.015 199.145 ;
        RECT 90.315 198.465 93.985 199.275 ;
        RECT 94.475 198.465 95.825 199.375 ;
        RECT 95.835 198.465 97.205 199.275 ;
        RECT 97.225 198.465 98.575 199.375 ;
        RECT 98.605 198.465 99.955 199.375 ;
        RECT 99.975 198.465 103.645 199.275 ;
        RECT 103.655 199.175 104.585 199.375 ;
        RECT 105.915 199.175 106.865 199.375 ;
        RECT 103.655 198.695 106.865 199.175 ;
        RECT 107.925 199.145 108.855 199.375 ;
        RECT 103.800 198.495 106.865 198.695 ;
        RECT 22.835 198.255 23.005 198.465 ;
        RECT 24.215 198.255 24.385 198.465 ;
        RECT 27.895 198.255 28.065 198.445 ;
        RECT 29.275 198.255 29.445 198.445 ;
        RECT 29.735 198.275 29.905 198.465 ;
        RECT 35.250 198.305 35.370 198.415 ;
        RECT 36.175 198.275 36.345 198.465 ;
        RECT 36.645 198.300 36.805 198.410 ;
        RECT 38.010 198.305 38.130 198.415 ;
        RECT 38.480 198.275 38.650 198.465 ;
        RECT 39.855 198.255 40.025 198.445 ;
        RECT 41.695 198.275 41.865 198.465 ;
        RECT 42.155 198.255 42.325 198.445 ;
        RECT 42.615 198.255 42.785 198.445 ;
        RECT 43.080 198.275 43.250 198.465 ;
        RECT 43.530 198.305 43.650 198.415 ;
        RECT 43.995 198.275 44.165 198.465 ;
        RECT 46.295 198.275 46.465 198.465 ;
        RECT 47.675 198.275 47.845 198.465 ;
        RECT 48.130 198.305 48.250 198.415 ;
        RECT 49.055 198.255 49.225 198.445 ;
        RECT 51.350 198.305 51.470 198.415 ;
        RECT 54.575 198.275 54.745 198.465 ;
        RECT 55.035 198.275 55.205 198.465 ;
        RECT 57.340 198.255 57.510 198.445 ;
        RECT 58.255 198.275 58.425 198.465 ;
        RECT 58.720 198.255 58.890 198.445 ;
        RECT 59.175 198.255 59.345 198.445 ;
        RECT 61.935 198.275 62.105 198.465 ;
        RECT 62.855 198.255 63.025 198.445 ;
        RECT 63.315 198.255 63.485 198.445 ;
        RECT 66.075 198.275 66.245 198.465 ;
        RECT 73.895 198.255 74.065 198.445 ;
        RECT 74.815 198.255 74.985 198.445 ;
        RECT 75.275 198.275 75.445 198.465 ;
        RECT 75.735 198.275 75.905 198.465 ;
        RECT 81.255 198.275 81.425 198.465 ;
        RECT 82.175 198.255 82.345 198.445 ;
        RECT 84.015 198.255 84.185 198.445 ;
        RECT 84.935 198.275 85.105 198.465 ;
        RECT 85.395 198.275 85.565 198.465 ;
        RECT 89.995 198.445 90.015 198.465 ;
        RECT 89.995 198.275 90.165 198.445 ;
        RECT 90.455 198.275 90.625 198.465 ;
        RECT 94.590 198.445 94.760 198.465 ;
        RECT 94.130 198.305 94.250 198.415 ;
        RECT 94.590 198.275 94.765 198.445 ;
        RECT 95.975 198.275 96.145 198.465 ;
        RECT 94.595 198.255 94.765 198.275 ;
        RECT 22.695 197.445 24.065 198.255 ;
        RECT 24.075 197.445 27.745 198.255 ;
        RECT 27.755 197.445 29.125 198.255 ;
        RECT 29.135 197.575 36.445 198.255 ;
        RECT 32.650 197.355 33.560 197.575 ;
        RECT 35.095 197.345 36.445 197.575 ;
        RECT 37.425 197.345 40.155 198.255 ;
        RECT 40.175 197.575 42.465 198.255 ;
        RECT 40.175 197.345 41.095 197.575 ;
        RECT 42.475 197.445 47.985 198.255 ;
        RECT 48.465 197.385 48.895 198.170 ;
        RECT 48.915 197.575 56.225 198.255 ;
        RECT 52.430 197.355 53.340 197.575 ;
        RECT 54.875 197.345 56.225 197.575 ;
        RECT 56.275 197.345 57.625 198.255 ;
        RECT 57.655 197.345 59.005 198.255 ;
        RECT 59.035 197.445 61.785 198.255 ;
        RECT 61.805 197.345 63.155 198.255 ;
        RECT 63.175 197.575 70.485 198.255 ;
        RECT 66.690 197.355 67.600 197.575 ;
        RECT 69.135 197.345 70.485 197.575 ;
        RECT 70.630 197.575 74.095 198.255 ;
        RECT 70.630 197.345 71.550 197.575 ;
        RECT 74.225 197.385 74.655 198.170 ;
        RECT 74.675 197.575 81.985 198.255 ;
        RECT 78.190 197.355 79.100 197.575 ;
        RECT 80.635 197.345 81.985 197.575 ;
        RECT 82.035 197.445 83.865 198.255 ;
        RECT 83.875 197.575 91.185 198.255 ;
        RECT 87.390 197.355 88.300 197.575 ;
        RECT 89.835 197.345 91.185 197.575 ;
        RECT 91.330 197.575 94.795 198.255 ;
        RECT 94.915 198.225 95.860 198.255 ;
        RECT 97.350 198.225 97.520 198.445 ;
        RECT 97.810 198.255 97.980 198.445 ;
        RECT 98.275 198.275 98.445 198.465 ;
        RECT 98.735 198.275 98.905 198.465 ;
        RECT 99.205 198.300 99.365 198.410 ;
        RECT 100.115 198.275 100.285 198.465 ;
        RECT 100.585 198.300 100.745 198.410 ;
        RECT 101.495 198.255 101.665 198.445 ;
        RECT 103.800 198.415 103.970 198.495 ;
        RECT 105.930 198.465 106.865 198.495 ;
        RECT 107.020 198.465 108.855 199.145 ;
        RECT 109.635 198.465 112.845 199.375 ;
        RECT 112.865 198.550 113.295 199.335 ;
        RECT 113.315 198.465 114.685 199.245 ;
        RECT 114.695 198.465 117.905 199.375 ;
        RECT 117.915 198.465 119.745 199.275 ;
        RECT 119.850 199.145 120.770 199.375 ;
        RECT 123.530 199.145 124.450 199.375 ;
        RECT 119.850 198.465 123.315 199.145 ;
        RECT 123.530 198.465 126.995 199.145 ;
        RECT 127.115 198.465 128.485 199.245 ;
        RECT 128.495 198.465 134.005 199.275 ;
        RECT 134.015 198.465 137.685 199.275 ;
        RECT 138.625 198.550 139.055 199.335 ;
        RECT 139.075 199.175 140.005 199.375 ;
        RECT 141.335 199.175 142.285 199.375 ;
        RECT 139.075 198.695 142.285 199.175 ;
        RECT 139.220 198.495 142.285 198.695 ;
        RECT 107.020 198.445 107.185 198.465 ;
        RECT 103.790 198.305 103.970 198.415 ;
        RECT 103.800 198.275 103.970 198.305 ;
        RECT 91.330 197.345 92.250 197.575 ;
        RECT 94.915 197.545 97.665 198.225 ;
        RECT 94.915 197.345 95.860 197.545 ;
        RECT 97.695 197.345 99.045 198.255 ;
        RECT 99.985 197.385 100.415 198.170 ;
        RECT 101.355 197.575 103.645 198.255 ;
        RECT 104.260 198.225 104.430 198.445 ;
        RECT 107.015 198.275 107.185 198.445 ;
        RECT 107.475 198.275 107.645 198.445 ;
        RECT 109.310 198.305 109.430 198.415 ;
        RECT 109.775 198.275 109.945 198.465 ;
        RECT 113.455 198.275 113.625 198.465 ;
        RECT 114.835 198.275 115.005 198.465 ;
        RECT 107.480 198.255 107.645 198.275 ;
        RECT 116.675 198.255 116.845 198.445 ;
        RECT 117.130 198.305 117.250 198.415 ;
        RECT 117.595 198.255 117.765 198.445 ;
        RECT 118.055 198.275 118.225 198.465 ;
        RECT 123.115 198.275 123.285 198.465 ;
        RECT 124.965 198.300 125.125 198.410 ;
        RECT 126.335 198.255 126.505 198.445 ;
        RECT 126.795 198.275 126.965 198.465 ;
        RECT 128.175 198.275 128.345 198.465 ;
        RECT 128.635 198.275 128.805 198.465 ;
        RECT 133.705 198.300 133.865 198.410 ;
        RECT 134.155 198.275 134.325 198.465 ;
        RECT 135.535 198.255 135.705 198.445 ;
        RECT 135.995 198.255 136.165 198.445 ;
        RECT 137.845 198.310 138.005 198.420 ;
        RECT 139.220 198.275 139.390 198.495 ;
        RECT 141.350 198.465 142.285 198.495 ;
        RECT 142.295 199.145 143.225 199.375 ;
        RECT 142.295 198.465 145.045 199.145 ;
        RECT 145.055 198.465 146.425 199.275 ;
        RECT 146.475 199.145 147.825 199.375 ;
        RECT 149.360 199.145 150.270 199.365 ;
        RECT 146.475 198.465 153.785 199.145 ;
        RECT 153.795 198.465 155.625 199.275 ;
        RECT 155.635 198.465 157.005 199.275 ;
        RECT 141.515 198.255 141.685 198.445 ;
        RECT 142.895 198.255 143.065 198.445 ;
        RECT 144.735 198.275 144.905 198.465 ;
        RECT 145.195 198.275 145.365 198.465 ;
        RECT 146.115 198.255 146.285 198.445 ;
        RECT 146.570 198.255 146.740 198.445 ;
        RECT 147.955 198.255 148.125 198.445 ;
        RECT 149.335 198.255 149.505 198.445 ;
        RECT 150.725 198.300 150.885 198.410 ;
        RECT 152.095 198.255 152.265 198.445 ;
        RECT 153.475 198.275 153.645 198.465 ;
        RECT 153.935 198.275 154.105 198.465 ;
        RECT 156.695 198.255 156.865 198.465 ;
        RECT 106.390 198.225 107.325 198.255 ;
        RECT 104.260 198.025 107.325 198.225 ;
        RECT 102.725 197.345 103.645 197.575 ;
        RECT 104.115 197.545 107.325 198.025 ;
        RECT 107.480 197.575 109.315 198.255 ;
        RECT 104.115 197.345 105.045 197.545 ;
        RECT 106.375 197.345 107.325 197.545 ;
        RECT 108.385 197.345 109.315 197.575 ;
        RECT 109.675 197.575 116.985 198.255 ;
        RECT 117.455 197.575 124.765 198.255 ;
        RECT 109.675 197.345 111.025 197.575 ;
        RECT 112.560 197.355 113.470 197.575 ;
        RECT 120.970 197.355 121.880 197.575 ;
        RECT 123.415 197.345 124.765 197.575 ;
        RECT 125.745 197.385 126.175 198.170 ;
        RECT 126.195 197.575 133.505 198.255 ;
        RECT 129.710 197.355 130.620 197.575 ;
        RECT 132.155 197.345 133.505 197.575 ;
        RECT 134.475 197.475 135.845 198.255 ;
        RECT 135.855 197.445 141.365 198.255 ;
        RECT 141.375 197.445 142.745 198.255 ;
        RECT 142.755 197.475 144.125 198.255 ;
        RECT 144.135 197.575 146.425 198.255 ;
        RECT 144.135 197.345 145.055 197.575 ;
        RECT 146.455 197.345 147.805 198.255 ;
        RECT 147.825 197.345 149.175 198.255 ;
        RECT 149.195 197.475 150.565 198.255 ;
        RECT 151.505 197.385 151.935 198.170 ;
        RECT 151.955 197.445 155.625 198.255 ;
        RECT 155.635 197.445 157.005 198.255 ;
      LAYER nwell ;
        RECT 22.500 194.225 157.200 197.055 ;
      LAYER pwell ;
        RECT 22.695 193.025 24.065 193.835 ;
        RECT 24.075 193.025 29.585 193.835 ;
        RECT 29.595 193.025 30.965 193.835 ;
        RECT 30.975 193.025 32.345 193.805 ;
        RECT 32.355 193.025 33.725 193.805 ;
        RECT 33.735 193.025 35.565 193.935 ;
        RECT 35.585 193.110 36.015 193.895 ;
        RECT 36.035 193.025 45.140 193.705 ;
        RECT 45.235 193.025 50.745 193.835 ;
        RECT 50.755 193.025 52.585 193.835 ;
        RECT 53.055 193.025 54.885 193.935 ;
        RECT 58.775 193.845 59.725 193.935 ;
        RECT 54.895 193.025 58.565 193.835 ;
        RECT 58.775 193.025 60.705 193.845 ;
        RECT 61.345 193.110 61.775 193.895 ;
        RECT 62.265 193.025 63.615 193.935 ;
        RECT 64.095 193.025 67.305 193.935 ;
        RECT 70.830 193.705 71.740 193.925 ;
        RECT 73.275 193.705 74.625 193.935 ;
        RECT 67.315 193.025 74.625 193.705 ;
        RECT 74.770 193.705 75.690 193.935 ;
        RECT 74.770 193.025 78.235 193.705 ;
        RECT 78.355 193.025 79.725 193.835 ;
        RECT 79.830 193.705 80.750 193.935 ;
        RECT 79.830 193.025 83.295 193.705 ;
        RECT 83.415 193.025 86.625 193.935 ;
        RECT 87.105 193.110 87.535 193.895 ;
        RECT 87.565 193.025 88.915 193.935 ;
        RECT 88.935 193.025 92.605 193.835 ;
        RECT 93.225 193.025 96.880 193.935 ;
        RECT 97.215 193.705 98.140 193.935 ;
        RECT 97.215 193.025 100.885 193.705 ;
        RECT 102.010 193.025 105.485 193.935 ;
        RECT 109.010 193.705 109.920 193.925 ;
        RECT 111.455 193.705 112.805 193.935 ;
        RECT 105.495 193.025 112.805 193.705 ;
        RECT 112.865 193.110 113.295 193.895 ;
        RECT 113.315 193.025 118.825 193.835 ;
        RECT 128.035 193.735 128.985 193.935 ;
        RECT 130.315 193.735 131.245 193.935 ;
        RECT 118.920 193.025 128.025 193.705 ;
        RECT 128.035 193.255 131.245 193.735 ;
        RECT 134.770 193.705 135.680 193.925 ;
        RECT 137.215 193.705 138.565 193.935 ;
        RECT 128.035 193.055 131.100 193.255 ;
        RECT 128.035 193.025 128.970 193.055 ;
        RECT 22.835 192.815 23.005 193.025 ;
        RECT 24.215 192.815 24.385 193.025 ;
        RECT 29.735 192.815 29.905 193.025 ;
        RECT 31.115 192.815 31.285 193.005 ;
        RECT 32.035 192.835 32.205 193.025 ;
        RECT 33.415 192.835 33.585 193.025 ;
        RECT 33.880 192.835 34.050 193.025 ;
        RECT 36.175 192.835 36.345 193.025 ;
        RECT 40.315 192.815 40.485 193.005 ;
        RECT 42.615 192.835 42.785 193.005 ;
        RECT 42.615 192.815 42.780 192.835 ;
        RECT 44.000 192.815 44.170 193.005 ;
        RECT 44.455 192.815 44.625 193.005 ;
        RECT 45.375 192.835 45.545 193.025 ;
        RECT 46.295 192.815 46.465 193.005 ;
        RECT 47.685 192.860 47.845 192.970 ;
        RECT 49.055 192.815 49.225 193.005 ;
        RECT 50.895 192.835 51.065 193.025 ;
        RECT 52.730 192.865 52.850 192.975 ;
        RECT 53.200 192.835 53.370 193.025 ;
        RECT 55.035 192.835 55.205 193.025 ;
        RECT 60.555 193.005 60.705 193.025 ;
        RECT 56.425 192.860 56.585 192.970 ;
        RECT 57.335 192.815 57.505 193.005 ;
        RECT 60.555 192.835 60.725 193.005 ;
        RECT 61.010 192.865 61.130 192.975 ;
        RECT 61.475 192.815 61.645 193.005 ;
        RECT 61.930 192.865 62.050 192.975 ;
        RECT 63.315 192.835 63.485 193.025 ;
        RECT 63.770 192.865 63.890 192.975 ;
        RECT 64.695 192.815 64.865 193.005 ;
        RECT 66.995 192.835 67.165 193.025 ;
        RECT 67.455 192.835 67.625 193.025 ;
        RECT 71.135 192.815 71.305 193.005 ;
        RECT 72.515 192.815 72.685 193.005 ;
        RECT 72.975 192.815 73.145 193.005 ;
        RECT 74.815 192.815 74.985 193.005 ;
        RECT 78.035 192.835 78.205 193.025 ;
        RECT 78.495 192.835 78.665 193.025 ;
        RECT 82.175 192.815 82.345 193.005 ;
        RECT 83.095 192.835 83.265 193.025 ;
        RECT 84.015 192.815 84.185 193.005 ;
        RECT 86.315 192.835 86.485 193.025 ;
        RECT 86.770 192.865 86.890 192.975 ;
        RECT 87.695 192.835 87.865 193.025 ;
        RECT 89.075 192.835 89.245 193.025 ;
        RECT 93.225 193.005 93.385 193.025 ;
        RECT 91.385 192.860 91.545 192.970 ;
        RECT 92.750 192.865 92.870 192.975 ;
        RECT 93.215 192.835 93.385 193.005 ;
        RECT 95.510 192.815 95.680 193.005 ;
        RECT 22.695 192.005 24.065 192.815 ;
        RECT 24.075 192.005 29.585 192.815 ;
        RECT 29.595 192.005 30.965 192.815 ;
        RECT 30.975 192.135 38.285 192.815 ;
        RECT 34.490 191.915 35.400 192.135 ;
        RECT 36.935 191.905 38.285 192.135 ;
        RECT 38.335 192.135 40.625 192.815 ;
        RECT 40.945 192.135 42.780 192.815 ;
        RECT 38.335 191.905 39.255 192.135 ;
        RECT 40.945 191.905 41.875 192.135 ;
        RECT 42.935 191.905 44.285 192.815 ;
        RECT 44.315 192.005 46.145 192.815 ;
        RECT 46.155 192.035 47.525 192.815 ;
        RECT 48.465 191.945 48.895 192.730 ;
        RECT 48.915 192.135 56.225 192.815 ;
        RECT 52.430 191.915 53.340 192.135 ;
        RECT 54.875 191.905 56.225 192.135 ;
        RECT 57.195 191.905 60.405 192.815 ;
        RECT 61.335 191.905 64.545 192.815 ;
        RECT 64.665 192.135 68.130 192.815 ;
        RECT 67.210 191.905 68.130 192.135 ;
        RECT 68.235 191.905 71.445 192.815 ;
        RECT 71.465 191.905 72.815 192.815 ;
        RECT 72.835 192.005 74.205 192.815 ;
        RECT 74.225 191.945 74.655 192.730 ;
        RECT 74.675 192.135 81.985 192.815 ;
        RECT 78.190 191.915 79.100 192.135 ;
        RECT 80.635 191.905 81.985 192.135 ;
        RECT 82.035 192.005 83.865 192.815 ;
        RECT 83.875 192.135 91.185 192.815 ;
        RECT 92.155 192.135 95.825 192.815 ;
        RECT 95.980 192.785 96.150 193.005 ;
        RECT 97.360 192.835 97.530 193.025 ;
        RECT 99.205 192.860 99.365 192.970 ;
        RECT 100.575 192.815 100.745 193.005 ;
        RECT 101.045 192.870 101.205 192.980 ;
        RECT 102.410 192.865 102.530 192.975 ;
        RECT 102.875 192.815 103.045 193.005 ;
        RECT 105.170 192.835 105.340 193.025 ;
        RECT 105.635 192.835 105.805 193.025 ;
        RECT 108.395 192.815 108.565 193.005 ;
        RECT 109.775 192.815 109.945 193.005 ;
        RECT 110.245 192.860 110.405 192.970 ;
        RECT 113.455 192.835 113.625 193.025 ;
        RECT 118.055 192.815 118.225 193.005 ;
        RECT 121.275 192.815 121.445 193.005 ;
        RECT 121.735 192.815 121.905 193.005 ;
        RECT 125.410 192.865 125.530 192.975 ;
        RECT 127.715 192.835 127.885 193.025 ;
        RECT 129.555 192.815 129.725 193.005 ;
        RECT 130.010 192.815 130.180 193.005 ;
        RECT 130.930 192.835 131.100 193.055 ;
        RECT 131.255 193.025 138.565 193.705 ;
        RECT 138.625 193.110 139.055 193.895 ;
        RECT 139.075 193.025 142.285 193.935 ;
        RECT 143.805 193.705 144.735 193.935 ;
        RECT 142.900 193.025 144.735 193.705 ;
        RECT 145.055 193.735 145.985 193.935 ;
        RECT 147.315 193.735 148.265 193.935 ;
        RECT 145.055 193.255 148.265 193.735 ;
        RECT 145.200 193.055 148.265 193.255 ;
        RECT 131.395 192.975 131.565 193.025 ;
        RECT 131.390 192.865 131.565 192.975 ;
        RECT 131.395 192.835 131.565 192.865 ;
        RECT 98.110 192.785 99.045 192.815 ;
        RECT 95.980 192.585 99.045 192.785 ;
        RECT 87.390 191.915 88.300 192.135 ;
        RECT 89.835 191.905 91.185 192.135 ;
        RECT 94.900 191.905 95.825 192.135 ;
        RECT 95.835 192.105 99.045 192.585 ;
        RECT 95.835 191.905 96.765 192.105 ;
        RECT 98.095 191.905 99.045 192.105 ;
        RECT 99.985 191.945 100.415 192.730 ;
        RECT 100.435 192.005 102.265 192.815 ;
        RECT 102.735 192.135 105.025 192.815 ;
        RECT 104.105 191.905 105.025 192.135 ;
        RECT 105.130 192.135 108.595 192.815 ;
        RECT 105.130 191.905 106.050 192.135 ;
        RECT 108.725 191.905 110.075 192.815 ;
        RECT 111.055 192.135 118.365 192.815 ;
        RECT 111.055 191.905 112.405 192.135 ;
        RECT 113.940 191.915 114.850 192.135 ;
        RECT 118.375 191.905 121.585 192.815 ;
        RECT 121.595 192.005 125.265 192.815 ;
        RECT 125.745 191.945 126.175 192.730 ;
        RECT 126.290 192.135 129.755 192.815 ;
        RECT 126.290 191.905 127.210 192.135 ;
        RECT 129.895 191.905 131.245 192.815 ;
        RECT 131.860 192.785 132.030 193.005 ;
        RECT 135.075 192.815 135.245 193.005 ;
        RECT 136.455 192.815 136.625 193.005 ;
        RECT 139.205 192.835 139.375 193.025 ;
        RECT 142.900 193.005 143.065 193.025 ;
        RECT 140.135 192.815 140.305 193.005 ;
        RECT 142.435 192.975 142.605 193.005 ;
        RECT 142.430 192.865 142.605 192.975 ;
        RECT 142.435 192.815 142.605 192.865 ;
        RECT 142.895 192.815 143.065 193.005 ;
        RECT 145.200 192.835 145.370 193.055 ;
        RECT 147.330 193.025 148.265 193.055 ;
        RECT 148.315 193.705 149.665 193.935 ;
        RECT 151.200 193.705 152.110 193.925 ;
        RECT 148.315 193.025 155.625 193.705 ;
        RECT 155.635 193.025 157.005 193.835 ;
        RECT 147.955 192.815 148.125 193.005 ;
        RECT 149.340 192.815 149.510 193.005 ;
        RECT 149.795 192.815 149.965 193.005 ;
        RECT 152.095 192.815 152.265 193.005 ;
        RECT 155.315 192.835 155.485 193.025 ;
        RECT 156.695 192.815 156.865 193.025 ;
        RECT 133.990 192.785 134.925 192.815 ;
        RECT 131.860 192.585 134.925 192.785 ;
        RECT 131.715 192.105 134.925 192.585 ;
        RECT 131.715 191.905 132.645 192.105 ;
        RECT 133.975 191.905 134.925 192.105 ;
        RECT 134.945 191.905 136.295 192.815 ;
        RECT 136.315 192.005 139.985 192.815 ;
        RECT 139.995 192.005 141.365 192.815 ;
        RECT 141.385 191.905 142.735 192.815 ;
        RECT 142.755 192.135 145.965 192.815 ;
        RECT 144.830 191.905 145.965 192.135 ;
        RECT 145.975 192.135 148.265 192.815 ;
        RECT 145.975 191.905 146.895 192.135 ;
        RECT 148.275 191.905 149.625 192.815 ;
        RECT 149.655 192.005 151.485 192.815 ;
        RECT 151.505 191.945 151.935 192.730 ;
        RECT 151.955 192.005 155.625 192.815 ;
        RECT 155.635 192.005 157.005 192.815 ;
      LAYER nwell ;
        RECT 22.500 188.785 157.200 191.615 ;
      LAYER pwell ;
        RECT 22.695 187.585 24.065 188.395 ;
        RECT 24.075 187.585 29.585 188.395 ;
        RECT 29.595 187.585 30.965 188.395 ;
        RECT 32.025 188.265 32.955 188.495 ;
        RECT 31.120 187.585 32.955 188.265 ;
        RECT 33.275 187.585 35.105 188.395 ;
        RECT 35.585 187.670 36.015 188.455 ;
        RECT 36.035 187.585 41.545 188.395 ;
        RECT 41.555 187.585 43.385 188.395 ;
        RECT 43.395 188.295 44.325 188.495 ;
        RECT 45.655 188.295 46.605 188.495 ;
        RECT 43.395 187.815 46.605 188.295 ;
        RECT 43.540 187.615 46.605 187.815 ;
        RECT 22.835 187.375 23.005 187.585 ;
        RECT 24.215 187.535 24.385 187.585 ;
        RECT 24.210 187.425 24.385 187.535 ;
        RECT 24.215 187.395 24.385 187.425 ;
        RECT 24.675 187.375 24.845 187.565 ;
        RECT 29.735 187.395 29.905 187.585 ;
        RECT 31.120 187.565 31.285 187.585 ;
        RECT 31.115 187.395 31.285 187.565 ;
        RECT 33.415 187.395 33.585 187.585 ;
        RECT 22.695 186.565 24.065 187.375 ;
        RECT 24.535 186.695 31.845 187.375 ;
        RECT 28.050 186.475 28.960 186.695 ;
        RECT 30.495 186.465 31.845 186.695 ;
        RECT 31.895 187.345 32.830 187.375 ;
        RECT 34.790 187.345 34.960 187.565 ;
        RECT 35.255 187.535 35.425 187.565 ;
        RECT 35.250 187.425 35.425 187.535 ;
        RECT 35.255 187.395 35.425 187.425 ;
        RECT 36.175 187.395 36.345 187.585 ;
        RECT 37.550 187.425 37.670 187.535 ;
        RECT 31.895 187.145 34.960 187.345 ;
        RECT 35.260 187.375 35.425 187.395 ;
        RECT 38.935 187.375 39.105 187.565 ;
        RECT 39.395 187.375 39.565 187.565 ;
        RECT 41.695 187.395 41.865 187.585 ;
        RECT 43.075 187.375 43.245 187.565 ;
        RECT 43.540 187.395 43.710 187.615 ;
        RECT 45.670 187.585 46.605 187.615 ;
        RECT 46.615 188.265 47.535 188.495 ;
        RECT 49.965 188.265 50.895 188.495 ;
        RECT 46.615 187.585 48.905 188.265 ;
        RECT 49.060 187.585 50.895 188.265 ;
        RECT 51.215 187.585 53.045 188.395 ;
        RECT 53.685 187.585 57.185 188.495 ;
        RECT 57.195 188.295 58.140 188.495 ;
        RECT 59.475 188.295 60.405 188.495 ;
        RECT 57.195 187.815 60.405 188.295 ;
        RECT 57.195 187.615 60.265 187.815 ;
        RECT 61.345 187.670 61.775 188.455 ;
        RECT 61.995 188.405 62.945 188.495 ;
        RECT 57.195 187.585 58.140 187.615 ;
        RECT 44.455 187.395 44.625 187.565 ;
        RECT 44.475 187.375 44.625 187.395 ;
        RECT 47.675 187.375 47.845 187.565 ;
        RECT 48.130 187.425 48.250 187.535 ;
        RECT 48.595 187.395 48.765 187.585 ;
        RECT 49.060 187.565 49.225 187.585 ;
        RECT 49.055 187.375 49.225 187.565 ;
        RECT 50.435 187.395 50.605 187.565 ;
        RECT 51.355 187.395 51.525 187.585 ;
        RECT 53.685 187.565 53.820 187.585 ;
        RECT 52.735 187.395 52.905 187.565 ;
        RECT 53.190 187.425 53.310 187.535 ;
        RECT 53.650 187.395 53.820 187.565 ;
        RECT 50.455 187.375 50.605 187.395 ;
        RECT 52.735 187.375 52.935 187.395 ;
        RECT 31.895 186.665 35.105 187.145 ;
        RECT 35.260 186.695 37.095 187.375 ;
        RECT 31.895 186.465 32.845 186.665 ;
        RECT 34.175 186.465 35.105 186.665 ;
        RECT 36.165 186.465 37.095 186.695 ;
        RECT 37.875 186.595 39.245 187.375 ;
        RECT 39.255 186.565 42.925 187.375 ;
        RECT 42.935 186.565 44.305 187.375 ;
        RECT 44.475 186.555 46.405 187.375 ;
        RECT 45.455 186.465 46.405 186.555 ;
        RECT 46.625 186.465 47.975 187.375 ;
        RECT 48.465 186.505 48.895 187.290 ;
        RECT 48.915 186.565 50.285 187.375 ;
        RECT 50.455 186.555 52.385 187.375 ;
        RECT 52.735 186.695 56.265 187.375 ;
        RECT 56.420 187.345 56.590 187.565 ;
        RECT 59.185 187.420 59.345 187.530 ;
        RECT 60.095 187.395 60.265 187.615 ;
        RECT 61.995 187.585 63.925 188.405 ;
        RECT 64.595 188.265 65.945 188.495 ;
        RECT 67.480 188.265 68.390 188.485 ;
        RECT 64.595 187.585 71.905 188.265 ;
        RECT 71.915 187.585 74.665 188.395 ;
        RECT 74.675 187.585 77.885 188.495 ;
        RECT 77.895 187.585 87.000 188.265 ;
        RECT 87.105 187.670 87.535 188.455 ;
        RECT 87.650 188.265 88.570 188.495 ;
        RECT 87.650 187.585 91.115 188.265 ;
        RECT 91.235 187.585 94.905 188.395 ;
        RECT 97.450 188.265 98.585 188.495 ;
        RECT 95.375 187.585 98.585 188.265 ;
        RECT 98.595 188.265 99.525 188.495 ;
        RECT 98.595 187.585 101.345 188.265 ;
        RECT 101.355 187.585 105.025 188.395 ;
        RECT 105.055 187.585 106.405 188.495 ;
        RECT 107.465 188.265 108.395 188.495 ;
        RECT 110.085 188.265 111.005 188.495 ;
        RECT 106.560 187.585 108.395 188.265 ;
        RECT 108.715 187.585 111.005 188.265 ;
        RECT 111.025 187.585 112.375 188.495 ;
        RECT 112.865 187.670 113.295 188.455 ;
        RECT 113.315 187.585 114.665 188.495 ;
        RECT 114.695 187.585 116.065 188.365 ;
        RECT 116.075 187.585 117.445 188.395 ;
        RECT 120.970 188.265 121.880 188.485 ;
        RECT 123.415 188.265 124.765 188.495 ;
        RECT 117.455 187.585 124.765 188.265 ;
        RECT 125.755 187.585 127.105 188.495 ;
        RECT 128.485 188.265 129.405 188.495 ;
        RECT 127.115 187.585 129.405 188.265 ;
        RECT 129.415 188.265 130.335 188.495 ;
        RECT 132.765 188.265 133.695 188.495 ;
        RECT 129.415 187.585 131.705 188.265 ;
        RECT 131.860 187.585 133.695 188.265 ;
        RECT 134.015 187.585 135.845 188.395 ;
        RECT 137.660 188.295 138.605 188.495 ;
        RECT 135.855 187.615 138.605 188.295 ;
        RECT 138.625 187.670 139.055 188.455 ;
        RECT 63.775 187.565 63.925 187.585 ;
        RECT 60.565 187.430 60.725 187.540 ;
        RECT 62.855 187.375 63.025 187.565 ;
        RECT 63.775 187.395 63.945 187.565 ;
        RECT 64.230 187.425 64.350 187.535 ;
        RECT 66.075 187.375 66.245 187.565 ;
        RECT 69.755 187.375 69.925 187.565 ;
        RECT 71.595 187.395 71.765 187.585 ;
        RECT 72.055 187.395 72.225 187.585 ;
        RECT 73.435 187.375 73.605 187.565 ;
        RECT 73.890 187.425 74.010 187.535 ;
        RECT 74.815 187.375 74.985 187.565 ;
        RECT 77.575 187.395 77.745 187.585 ;
        RECT 78.035 187.395 78.205 187.585 ;
        RECT 78.955 187.375 79.125 187.565 ;
        RECT 82.635 187.375 82.805 187.565 ;
        RECT 85.855 187.375 86.025 187.565 ;
        RECT 86.310 187.425 86.430 187.535 ;
        RECT 58.080 187.345 59.025 187.375 ;
        RECT 51.435 186.465 52.385 186.555 ;
        RECT 53.440 186.465 56.265 186.695 ;
        RECT 56.275 186.665 59.025 187.345 ;
        RECT 58.080 186.465 59.025 186.665 ;
        RECT 59.955 186.465 63.165 187.375 ;
        RECT 63.175 186.465 66.385 187.375 ;
        RECT 66.490 186.695 69.955 187.375 ;
        RECT 70.170 186.695 73.635 187.375 ;
        RECT 66.490 186.465 67.410 186.695 ;
        RECT 70.170 186.465 71.090 186.695 ;
        RECT 74.225 186.505 74.655 187.290 ;
        RECT 74.675 186.565 76.045 187.375 ;
        RECT 76.055 186.465 79.265 187.375 ;
        RECT 79.370 186.695 82.835 187.375 ;
        RECT 79.370 186.465 80.290 186.695 ;
        RECT 82.955 186.465 86.165 187.375 ;
        RECT 86.780 187.345 86.950 187.565 ;
        RECT 90.915 187.395 91.085 187.585 ;
        RECT 91.375 187.395 91.545 187.585 ;
        RECT 88.440 187.345 89.385 187.375 ;
        RECT 86.635 186.665 89.385 187.345 ;
        RECT 88.440 186.465 89.385 186.665 ;
        RECT 89.395 187.345 90.340 187.375 ;
        RECT 91.830 187.345 92.000 187.565 ;
        RECT 92.295 187.375 92.465 187.565 ;
        RECT 95.050 187.425 95.170 187.535 ;
        RECT 95.515 187.395 95.685 187.585 ;
        RECT 95.970 187.425 96.090 187.535 ;
        RECT 96.425 187.375 96.595 187.565 ;
        RECT 99.650 187.425 99.770 187.535 ;
        RECT 100.585 187.420 100.745 187.530 ;
        RECT 101.035 187.395 101.205 187.585 ;
        RECT 101.495 187.375 101.665 187.585 ;
        RECT 104.250 187.425 104.370 187.535 ;
        RECT 104.715 187.375 104.885 187.565 ;
        RECT 105.170 187.395 105.340 187.585 ;
        RECT 106.560 187.565 106.725 187.585 ;
        RECT 106.555 187.535 106.725 187.565 ;
        RECT 106.550 187.425 106.725 187.535 ;
        RECT 106.555 187.395 106.725 187.425 ;
        RECT 107.935 187.375 108.105 187.565 ;
        RECT 108.390 187.425 108.510 187.535 ;
        RECT 108.855 187.375 109.025 187.585 ;
        RECT 111.155 187.395 111.325 187.585 ;
        RECT 112.530 187.425 112.650 187.535 ;
        RECT 114.380 187.395 114.550 187.585 ;
        RECT 114.835 187.395 115.005 187.585 ;
        RECT 116.215 187.395 116.385 187.585 ;
        RECT 117.595 187.395 117.765 187.585 ;
        RECT 118.975 187.375 119.145 187.565 ;
        RECT 119.435 187.375 119.605 187.565 ;
        RECT 123.110 187.425 123.230 187.535 ;
        RECT 124.495 187.375 124.665 187.565 ;
        RECT 124.965 187.420 125.125 187.540 ;
        RECT 126.790 187.395 126.960 187.585 ;
        RECT 127.255 187.395 127.425 187.585 ;
        RECT 128.175 187.375 128.345 187.565 ;
        RECT 128.640 187.375 128.810 187.565 ;
        RECT 130.475 187.375 130.645 187.565 ;
        RECT 131.395 187.395 131.565 187.585 ;
        RECT 131.860 187.565 132.025 187.585 ;
        RECT 131.855 187.395 132.030 187.565 ;
        RECT 134.155 187.395 134.325 187.585 ;
        RECT 134.625 187.420 134.785 187.530 ;
        RECT 136.000 187.395 136.170 187.615 ;
        RECT 137.660 187.585 138.605 187.615 ;
        RECT 139.075 187.585 144.585 188.395 ;
        RECT 144.595 187.585 146.425 188.395 ;
        RECT 146.435 187.585 155.540 188.265 ;
        RECT 155.635 187.585 157.005 188.395 ;
        RECT 89.395 186.665 92.145 187.345 ;
        RECT 89.395 186.465 90.340 186.665 ;
        RECT 92.155 186.565 95.825 187.375 ;
        RECT 96.295 186.465 99.505 187.375 ;
        RECT 99.985 186.505 100.415 187.290 ;
        RECT 101.355 186.695 104.105 187.375 ;
        RECT 104.575 186.695 106.405 187.375 ;
        RECT 103.175 186.465 104.105 186.695 ;
        RECT 105.060 186.465 106.405 186.695 ;
        RECT 106.885 186.465 108.235 187.375 ;
        RECT 108.715 186.695 111.005 187.375 ;
        RECT 110.085 186.465 111.005 186.695 ;
        RECT 111.975 186.695 119.285 187.375 ;
        RECT 111.975 186.465 113.325 186.695 ;
        RECT 114.860 186.475 115.770 186.695 ;
        RECT 119.295 186.565 122.965 187.375 ;
        RECT 123.435 186.595 124.805 187.375 ;
        RECT 125.745 186.505 126.175 187.290 ;
        RECT 126.195 186.695 128.485 187.375 ;
        RECT 126.195 186.465 127.115 186.695 ;
        RECT 128.495 186.465 130.325 187.375 ;
        RECT 130.335 186.565 131.705 187.375 ;
        RECT 131.860 187.345 132.030 187.395 ;
        RECT 138.295 187.375 138.465 187.565 ;
        RECT 138.755 187.375 138.925 187.565 ;
        RECT 139.215 187.395 139.385 187.585 ;
        RECT 144.735 187.565 144.905 187.585 ;
        RECT 141.975 187.375 142.145 187.565 ;
        RECT 144.735 187.395 144.910 187.565 ;
        RECT 146.575 187.395 146.745 187.585 ;
        RECT 133.520 187.345 134.465 187.375 ;
        RECT 131.715 186.665 134.465 187.345 ;
        RECT 133.520 186.465 134.465 186.665 ;
        RECT 135.395 186.695 138.605 187.375 ;
        RECT 135.395 186.465 136.530 186.695 ;
        RECT 138.615 186.465 141.825 187.375 ;
        RECT 141.835 186.565 144.585 187.375 ;
        RECT 144.740 187.345 144.910 187.395 ;
        RECT 149.795 187.375 149.965 187.565 ;
        RECT 151.175 187.375 151.345 187.565 ;
        RECT 152.095 187.375 152.265 187.565 ;
        RECT 156.695 187.375 156.865 187.585 ;
        RECT 146.870 187.345 147.805 187.375 ;
        RECT 144.740 187.145 147.805 187.345 ;
        RECT 144.595 186.665 147.805 187.145 ;
        RECT 144.595 186.465 145.525 186.665 ;
        RECT 146.855 186.465 147.805 186.665 ;
        RECT 147.815 186.695 150.105 187.375 ;
        RECT 147.815 186.465 148.735 186.695 ;
        RECT 150.115 186.595 151.485 187.375 ;
        RECT 151.505 186.505 151.935 187.290 ;
        RECT 151.955 186.565 155.625 187.375 ;
        RECT 155.635 186.565 157.005 187.375 ;
      LAYER nwell ;
        RECT 22.500 183.345 157.200 186.175 ;
      LAYER pwell ;
        RECT 32.115 182.965 33.065 183.055 ;
        RECT 22.695 182.145 24.065 182.955 ;
        RECT 24.075 182.145 26.825 182.955 ;
        RECT 26.835 182.145 28.205 182.925 ;
        RECT 28.215 182.145 30.965 182.955 ;
        RECT 31.135 182.145 33.065 182.965 ;
        RECT 34.645 182.825 35.565 183.055 ;
        RECT 33.275 182.145 35.565 182.825 ;
        RECT 35.585 182.230 36.015 183.015 ;
        RECT 39.550 182.825 40.460 183.045 ;
        RECT 41.995 182.825 43.345 183.055 ;
        RECT 36.035 182.145 43.345 182.825 ;
        RECT 43.395 182.145 44.765 182.955 ;
        RECT 48.290 182.825 49.200 183.045 ;
        RECT 50.735 182.825 52.085 183.055 ;
        RECT 44.775 182.145 52.085 182.825 ;
        RECT 52.230 182.825 53.150 183.055 ;
        RECT 52.230 182.145 55.695 182.825 ;
        RECT 55.815 182.145 59.025 183.055 ;
        RECT 59.045 182.145 60.395 183.055 ;
        RECT 61.345 182.230 61.775 183.015 ;
        RECT 61.805 182.145 63.155 183.055 ;
        RECT 66.690 182.825 67.600 183.045 ;
        RECT 69.135 182.825 70.485 183.055 ;
        RECT 74.050 182.825 74.960 183.045 ;
        RECT 76.495 182.825 77.845 183.055 ;
        RECT 81.410 182.825 82.320 183.045 ;
        RECT 83.855 182.825 85.205 183.055 ;
        RECT 63.175 182.145 70.485 182.825 ;
        RECT 70.535 182.145 77.845 182.825 ;
        RECT 77.895 182.145 85.205 182.825 ;
        RECT 85.735 182.145 87.085 183.055 ;
        RECT 87.105 182.230 87.535 183.015 ;
        RECT 87.650 182.825 88.570 183.055 ;
        RECT 87.650 182.145 91.115 182.825 ;
        RECT 91.695 182.145 94.905 183.055 ;
        RECT 95.875 182.825 97.225 183.055 ;
        RECT 98.760 182.825 99.670 183.045 ;
        RECT 95.875 182.145 103.185 182.825 ;
        RECT 103.195 182.145 108.705 182.955 ;
        RECT 110.225 182.825 111.155 183.055 ;
        RECT 109.320 182.145 111.155 182.825 ;
        RECT 111.485 182.145 112.835 183.055 ;
        RECT 112.865 182.230 113.295 183.015 ;
        RECT 113.315 182.145 114.685 182.925 ;
        RECT 114.695 182.145 120.205 182.955 ;
        RECT 124.650 182.825 125.560 183.045 ;
        RECT 127.095 182.825 128.445 183.055 ;
        RECT 121.135 182.145 128.445 182.825 ;
        RECT 128.505 182.145 131.235 183.055 ;
        RECT 133.520 182.855 134.465 183.055 ;
        RECT 136.740 182.855 137.685 183.055 ;
        RECT 131.715 182.175 134.465 182.855 ;
        RECT 134.935 182.175 137.685 182.855 ;
        RECT 138.625 182.230 139.055 183.015 ;
        RECT 22.835 181.935 23.005 182.145 ;
        RECT 24.215 181.955 24.385 182.145 ;
        RECT 26.055 181.935 26.225 182.125 ;
        RECT 26.515 181.935 26.685 182.125 ;
        RECT 27.895 181.955 28.065 182.145 ;
        RECT 28.355 181.955 28.525 182.145 ;
        RECT 31.135 182.125 31.285 182.145 ;
        RECT 30.205 181.980 30.365 182.090 ;
        RECT 31.115 181.955 31.285 182.125 ;
        RECT 31.120 181.935 31.285 181.955 ;
        RECT 33.415 181.935 33.585 182.145 ;
        RECT 36.175 182.125 36.345 182.145 ;
        RECT 36.175 181.955 36.350 182.125 ;
        RECT 22.695 181.125 24.065 181.935 ;
        RECT 24.995 181.155 26.365 181.935 ;
        RECT 26.375 181.125 30.045 181.935 ;
        RECT 31.120 181.255 32.955 181.935 ;
        RECT 32.025 181.025 32.955 181.255 ;
        RECT 33.275 181.125 36.025 181.935 ;
        RECT 36.180 181.905 36.350 181.955 ;
        RECT 39.395 181.935 39.565 182.125 ;
        RECT 42.150 181.985 42.270 182.095 ;
        RECT 43.535 181.955 43.705 182.145 ;
        RECT 44.915 181.955 45.085 182.145 ;
        RECT 45.830 181.935 46.000 182.125 ;
        RECT 46.295 181.935 46.465 182.125 ;
        RECT 48.130 181.985 48.250 182.095 ;
        RECT 49.055 181.935 49.225 182.125 ;
        RECT 52.735 181.935 52.905 182.125 ;
        RECT 55.035 181.935 55.205 182.125 ;
        RECT 55.495 181.935 55.665 182.145 ;
        RECT 58.715 181.955 58.885 182.145 ;
        RECT 59.170 181.985 59.290 182.095 ;
        RECT 59.635 181.935 59.805 182.125 ;
        RECT 60.095 181.955 60.265 182.145 ;
        RECT 60.565 181.990 60.725 182.100 ;
        RECT 62.855 181.955 63.025 182.145 ;
        RECT 63.315 181.955 63.485 182.145 ;
        RECT 70.215 181.935 70.385 182.125 ;
        RECT 70.675 181.935 70.845 182.145 ;
        RECT 74.815 181.935 74.985 182.125 ;
        RECT 78.035 181.955 78.205 182.145 ;
        RECT 85.850 182.125 86.020 182.145 ;
        RECT 78.490 181.985 78.610 182.095 ;
        RECT 81.715 181.935 81.885 182.125 ;
        RECT 82.175 181.935 82.345 182.125 ;
        RECT 85.390 181.985 85.510 182.095 ;
        RECT 85.850 181.955 86.030 182.125 ;
        RECT 38.310 181.905 39.245 181.935 ;
        RECT 36.180 181.705 39.245 181.905 ;
        RECT 36.035 181.225 39.245 181.705 ;
        RECT 36.035 181.025 36.965 181.225 ;
        RECT 38.295 181.025 39.245 181.225 ;
        RECT 39.255 181.125 42.005 181.935 ;
        RECT 42.670 181.025 46.145 181.935 ;
        RECT 46.155 181.125 47.985 181.935 ;
        RECT 48.465 181.065 48.895 181.850 ;
        RECT 48.915 181.125 52.585 181.935 ;
        RECT 52.595 181.125 53.965 181.935 ;
        RECT 53.985 181.025 55.335 181.935 ;
        RECT 55.355 181.125 59.025 181.935 ;
        RECT 59.495 181.255 66.805 181.935 ;
        RECT 63.010 181.035 63.920 181.255 ;
        RECT 65.455 181.025 66.805 181.255 ;
        RECT 66.950 181.255 70.415 181.935 ;
        RECT 66.950 181.025 67.870 181.255 ;
        RECT 70.535 181.125 74.205 181.935 ;
        RECT 74.225 181.065 74.655 181.850 ;
        RECT 74.675 181.125 78.345 181.935 ;
        RECT 78.815 181.025 82.025 181.935 ;
        RECT 82.035 181.125 85.705 181.935 ;
        RECT 85.860 181.905 86.030 181.955 ;
        RECT 88.615 181.935 88.785 182.125 ;
        RECT 90.915 181.955 91.085 182.145 ;
        RECT 91.370 181.985 91.490 182.095 ;
        RECT 91.835 181.955 92.005 182.145 ;
        RECT 87.520 181.905 88.465 181.935 ;
        RECT 85.715 181.225 88.465 181.905 ;
        RECT 88.475 181.255 91.685 181.935 ;
        RECT 92.760 181.905 92.930 182.125 ;
        RECT 95.065 181.990 95.225 182.100 ;
        RECT 95.985 181.980 96.145 182.090 ;
        RECT 96.895 181.935 97.065 182.125 ;
        RECT 99.205 181.980 99.365 182.090 ;
        RECT 100.575 181.935 100.745 182.125 ;
        RECT 102.875 181.955 103.045 182.145 ;
        RECT 103.335 182.125 103.505 182.145 ;
        RECT 109.320 182.125 109.485 182.145 ;
        RECT 103.335 181.955 103.510 182.125 ;
        RECT 103.340 181.935 103.510 181.955 ;
        RECT 104.715 181.935 104.885 182.125 ;
        RECT 108.395 181.935 108.565 182.125 ;
        RECT 108.850 181.985 108.970 182.095 ;
        RECT 109.315 181.955 109.485 182.125 ;
        RECT 109.775 181.955 109.945 182.125 ;
        RECT 109.925 181.935 109.945 181.955 ;
        RECT 112.535 181.935 112.705 182.145 ;
        RECT 113.455 181.955 113.625 182.145 ;
        RECT 114.835 181.955 115.005 182.145 ;
        RECT 116.215 181.935 116.385 182.125 ;
        RECT 116.675 181.935 116.845 182.125 ;
        RECT 120.365 181.990 120.525 182.100 ;
        RECT 121.275 181.955 121.445 182.145 ;
        RECT 121.735 181.935 121.905 182.125 ;
        RECT 124.955 181.935 125.125 182.125 ;
        RECT 125.410 181.985 125.530 182.095 ;
        RECT 128.635 181.955 128.805 182.145 ;
        RECT 129.555 181.935 129.725 182.125 ;
        RECT 130.015 181.935 130.185 182.125 ;
        RECT 131.390 181.985 131.510 182.095 ;
        RECT 131.860 181.955 132.030 182.175 ;
        RECT 133.520 182.145 134.465 182.175 ;
        RECT 132.775 181.935 132.945 182.125 ;
        RECT 134.610 181.985 134.730 182.095 ;
        RECT 135.080 181.955 135.250 182.175 ;
        RECT 136.740 182.145 137.685 182.175 ;
        RECT 139.095 182.145 140.445 183.055 ;
        RECT 140.915 182.825 142.260 183.055 ;
        RECT 143.065 182.825 143.995 183.055 ;
        RECT 145.055 182.855 145.985 183.055 ;
        RECT 147.315 182.855 148.265 183.055 ;
        RECT 140.915 182.145 142.745 182.825 ;
        RECT 143.065 182.145 144.900 182.825 ;
        RECT 145.055 182.375 148.265 182.855 ;
        RECT 139.210 182.125 139.380 182.145 ;
        RECT 135.535 181.935 135.705 182.125 ;
        RECT 137.845 181.990 138.005 182.100 ;
        RECT 139.210 181.955 139.385 182.125 ;
        RECT 140.590 181.985 140.710 182.095 ;
        RECT 139.215 181.935 139.385 181.955 ;
        RECT 141.975 181.935 142.145 182.125 ;
        RECT 142.435 181.955 142.605 182.145 ;
        RECT 144.735 182.125 144.900 182.145 ;
        RECT 145.200 182.175 148.265 182.375 ;
        RECT 143.810 181.985 143.930 182.095 ;
        RECT 144.735 181.955 144.905 182.125 ;
        RECT 145.200 181.955 145.370 182.175 ;
        RECT 147.330 182.145 148.265 182.175 ;
        RECT 148.315 182.825 149.665 183.055 ;
        RECT 151.200 182.825 152.110 183.045 ;
        RECT 148.315 182.145 155.625 182.825 ;
        RECT 155.635 182.145 157.005 182.955 ;
        RECT 151.175 181.935 151.345 182.125 ;
        RECT 152.095 181.955 152.265 182.125 ;
        RECT 152.100 181.935 152.265 181.955 ;
        RECT 155.315 181.935 155.485 182.145 ;
        RECT 156.695 181.935 156.865 182.145 ;
        RECT 94.890 181.905 95.825 181.935 ;
        RECT 92.760 181.705 95.825 181.905 ;
        RECT 87.520 181.025 88.465 181.225 ;
        RECT 90.550 181.025 91.685 181.255 ;
        RECT 92.615 181.225 95.825 181.705 ;
        RECT 96.755 181.255 99.045 181.935 ;
        RECT 92.615 181.025 93.545 181.225 ;
        RECT 94.875 181.025 95.825 181.225 ;
        RECT 98.125 181.025 99.045 181.255 ;
        RECT 99.985 181.065 100.415 181.850 ;
        RECT 100.435 181.125 103.185 181.935 ;
        RECT 103.195 181.025 104.545 181.935 ;
        RECT 104.575 181.125 108.245 181.935 ;
        RECT 108.255 181.125 109.625 181.935 ;
        RECT 109.925 181.255 112.375 181.935 ;
        RECT 110.415 181.025 112.375 181.255 ;
        RECT 112.395 181.125 115.145 181.935 ;
        RECT 115.165 181.025 116.515 181.935 ;
        RECT 116.535 181.125 118.365 181.935 ;
        RECT 118.470 181.255 121.935 181.935 ;
        RECT 118.470 181.025 119.390 181.255 ;
        RECT 122.055 181.025 125.265 181.935 ;
        RECT 125.745 181.065 126.175 181.850 ;
        RECT 126.290 181.255 129.755 181.935 ;
        RECT 126.290 181.025 127.210 181.255 ;
        RECT 129.875 181.125 132.625 181.935 ;
        RECT 132.635 181.255 135.385 181.935 ;
        RECT 134.455 181.025 135.385 181.255 ;
        RECT 135.395 181.125 139.065 181.935 ;
        RECT 139.075 181.255 141.825 181.935 ;
        RECT 140.895 181.025 141.825 181.255 ;
        RECT 141.835 181.125 143.665 181.935 ;
        RECT 144.175 181.255 151.485 181.935 ;
        RECT 144.175 181.025 145.525 181.255 ;
        RECT 147.060 181.035 147.970 181.255 ;
        RECT 151.505 181.065 151.935 181.850 ;
        RECT 152.100 181.255 153.935 181.935 ;
        RECT 153.005 181.025 153.935 181.255 ;
        RECT 154.255 181.155 155.625 181.935 ;
        RECT 155.635 181.125 157.005 181.935 ;
      LAYER nwell ;
        RECT 22.500 177.905 157.200 180.735 ;
      LAYER pwell ;
        RECT 22.695 176.705 24.065 177.515 ;
        RECT 27.590 177.385 28.500 177.605 ;
        RECT 30.035 177.385 31.385 177.615 ;
        RECT 24.075 176.705 31.385 177.385 ;
        RECT 31.435 177.415 32.385 177.615 ;
        RECT 33.715 177.415 34.645 177.615 ;
        RECT 31.435 176.935 34.645 177.415 ;
        RECT 31.435 176.735 34.500 176.935 ;
        RECT 35.585 176.790 36.015 177.575 ;
        RECT 36.035 177.385 36.955 177.615 ;
        RECT 31.435 176.705 32.370 176.735 ;
        RECT 22.835 176.495 23.005 176.705 ;
        RECT 24.215 176.515 24.385 176.705 ;
        RECT 26.055 176.495 26.225 176.685 ;
        RECT 26.515 176.495 26.685 176.685 ;
        RECT 28.355 176.515 28.525 176.685 ;
        RECT 28.375 176.495 28.525 176.515 ;
        RECT 22.695 175.685 24.065 176.495 ;
        RECT 24.995 175.715 26.365 176.495 ;
        RECT 26.375 175.685 28.205 176.495 ;
        RECT 28.375 175.675 30.305 176.495 ;
        RECT 30.660 176.465 30.830 176.685 ;
        RECT 34.330 176.515 34.500 176.735 ;
        RECT 36.035 176.705 38.325 177.385 ;
        RECT 38.335 176.705 42.005 177.515 ;
        RECT 44.550 177.385 45.685 177.615 ;
        RECT 42.475 176.705 45.685 177.385 ;
        RECT 45.695 177.385 46.830 177.615 ;
        RECT 45.695 176.705 48.905 177.385 ;
        RECT 48.925 176.705 50.275 177.615 ;
        RECT 53.960 177.385 54.885 177.615 ;
        RECT 56.700 177.415 57.645 177.615 ;
        RECT 51.215 176.705 54.885 177.385 ;
        RECT 54.895 176.735 57.645 177.415 ;
        RECT 34.805 176.550 34.965 176.660 ;
        RECT 35.715 176.515 35.885 176.685 ;
        RECT 35.715 176.495 35.880 176.515 ;
        RECT 36.175 176.495 36.345 176.685 ;
        RECT 38.015 176.515 38.185 176.705 ;
        RECT 38.475 176.515 38.645 176.705 ;
        RECT 42.150 176.545 42.270 176.655 ;
        RECT 42.615 176.515 42.785 176.705 ;
        RECT 43.545 176.540 43.705 176.650 ;
        RECT 44.455 176.495 44.625 176.685 ;
        RECT 45.835 176.495 46.005 176.685 ;
        RECT 48.595 176.515 48.765 176.705 ;
        RECT 49.055 176.515 49.225 176.705 ;
        RECT 49.975 176.495 50.145 176.685 ;
        RECT 50.445 176.550 50.605 176.660 ;
        RECT 54.570 176.515 54.740 176.705 ;
        RECT 55.040 176.515 55.210 176.735 ;
        RECT 56.700 176.705 57.645 176.735 ;
        RECT 57.655 176.705 59.005 177.615 ;
        RECT 59.035 176.705 60.865 177.515 ;
        RECT 61.345 176.790 61.775 177.575 ;
        RECT 61.835 177.385 63.185 177.615 ;
        RECT 64.720 177.385 65.630 177.605 ;
        RECT 61.835 176.705 69.145 177.385 ;
        RECT 69.155 176.705 72.365 177.615 ;
        RECT 75.030 177.385 75.950 177.615 ;
        RECT 72.485 176.705 75.950 177.385 ;
        RECT 76.055 176.705 77.885 177.515 ;
        RECT 81.870 177.385 82.780 177.605 ;
        RECT 84.315 177.385 85.665 177.615 ;
        RECT 78.355 176.705 85.665 177.385 ;
        RECT 85.715 176.705 87.085 177.515 ;
        RECT 87.105 176.790 87.535 177.575 ;
        RECT 87.555 176.705 89.385 177.515 ;
        RECT 91.200 177.415 92.145 177.615 ;
        RECT 89.395 176.735 92.145 177.415 ;
        RECT 93.665 177.385 94.595 177.615 ;
        RECT 56.875 176.515 57.045 176.685 ;
        RECT 56.875 176.495 57.035 176.515 ;
        RECT 57.340 176.495 57.510 176.685 ;
        RECT 58.720 176.515 58.890 176.705 ;
        RECT 59.175 176.515 59.345 176.705 ;
        RECT 61.010 176.545 61.130 176.655 ;
        RECT 61.940 176.495 62.110 176.685 ;
        RECT 62.405 176.540 62.565 176.650 ;
        RECT 66.075 176.495 66.245 176.685 ;
        RECT 66.530 176.545 66.650 176.655 ;
        RECT 68.835 176.515 69.005 176.705 ;
        RECT 72.055 176.515 72.225 176.705 ;
        RECT 72.515 176.515 72.685 176.705 ;
        RECT 73.895 176.495 74.065 176.685 ;
        RECT 76.195 176.515 76.365 176.705 ;
        RECT 78.035 176.655 78.205 176.685 ;
        RECT 78.030 176.545 78.205 176.655 ;
        RECT 78.035 176.495 78.205 176.545 ;
        RECT 78.495 176.515 78.665 176.705 ;
        RECT 81.255 176.495 81.425 176.685 ;
        RECT 81.725 176.540 81.885 176.650 ;
        RECT 83.555 176.495 83.725 176.685 ;
        RECT 84.940 176.495 85.110 176.685 ;
        RECT 85.855 176.515 86.025 176.705 ;
        RECT 87.695 176.515 87.865 176.705 ;
        RECT 32.790 176.465 33.725 176.495 ;
        RECT 30.660 176.265 33.725 176.465 ;
        RECT 29.355 175.585 30.305 175.675 ;
        RECT 30.515 175.785 33.725 176.265 ;
        RECT 30.515 175.585 31.445 175.785 ;
        RECT 32.775 175.585 33.725 175.785 ;
        RECT 34.045 175.815 35.880 176.495 ;
        RECT 36.035 175.815 43.345 176.495 ;
        RECT 34.045 175.585 34.975 175.815 ;
        RECT 39.550 175.595 40.460 175.815 ;
        RECT 41.995 175.585 43.345 175.815 ;
        RECT 44.325 175.585 45.675 176.495 ;
        RECT 45.695 175.815 48.435 176.495 ;
        RECT 48.465 175.625 48.895 176.410 ;
        RECT 49.835 175.585 53.045 176.495 ;
        RECT 53.380 175.585 57.035 176.495 ;
        RECT 57.195 175.815 60.865 176.495 ;
        RECT 57.195 175.585 58.120 175.815 ;
        RECT 60.875 175.585 62.225 176.495 ;
        RECT 63.175 175.585 66.385 176.495 ;
        RECT 66.895 175.815 74.205 176.495 ;
        RECT 66.895 175.585 68.245 175.815 ;
        RECT 69.780 175.595 70.690 175.815 ;
        RECT 74.225 175.625 74.655 176.410 ;
        RECT 74.770 175.815 78.235 176.495 ;
        RECT 74.770 175.585 75.690 175.815 ;
        RECT 78.355 175.585 81.565 176.495 ;
        RECT 82.505 175.585 83.855 176.495 ;
        RECT 83.875 175.585 85.225 176.495 ;
        RECT 85.255 176.465 86.190 176.495 ;
        RECT 88.150 176.465 88.320 176.685 ;
        RECT 88.615 176.495 88.785 176.685 ;
        RECT 89.540 176.515 89.710 176.735 ;
        RECT 91.200 176.705 92.145 176.735 ;
        RECT 92.760 176.705 94.595 177.385 ;
        RECT 94.915 177.385 95.835 177.615 ;
        RECT 94.915 176.705 97.205 177.385 ;
        RECT 97.215 176.705 98.585 177.485 ;
        RECT 99.055 176.705 101.805 177.615 ;
        RECT 101.995 176.935 104.330 177.615 ;
        RECT 107.325 177.385 108.245 177.615 ;
        RECT 101.995 176.705 103.845 176.935 ;
        RECT 104.660 176.705 108.245 177.385 ;
        RECT 108.255 176.705 111.925 177.515 ;
        RECT 112.865 176.790 113.295 177.575 ;
        RECT 116.830 177.385 117.740 177.605 ;
        RECT 119.275 177.385 120.625 177.615 ;
        RECT 124.190 177.385 125.100 177.605 ;
        RECT 126.635 177.385 127.985 177.615 ;
        RECT 129.855 177.385 130.785 177.615 ;
        RECT 113.315 176.705 120.625 177.385 ;
        RECT 120.675 176.705 127.985 177.385 ;
        RECT 128.035 176.705 130.785 177.385 ;
        RECT 130.795 176.705 132.625 177.515 ;
        RECT 133.095 176.705 137.225 177.615 ;
        RECT 137.245 176.705 138.595 177.615 ;
        RECT 138.625 176.790 139.055 177.575 ;
        RECT 139.075 176.705 141.825 177.615 ;
        RECT 141.835 177.385 142.755 177.615 ;
        RECT 141.835 176.705 144.125 177.385 ;
        RECT 144.330 176.705 147.805 177.615 ;
        RECT 151.330 177.385 152.240 177.605 ;
        RECT 153.775 177.385 155.125 177.615 ;
        RECT 147.815 176.705 155.125 177.385 ;
        RECT 155.635 176.705 157.005 177.515 ;
        RECT 92.760 176.685 92.925 176.705 ;
        RECT 90.915 176.495 91.085 176.685 ;
        RECT 92.290 176.545 92.410 176.655 ;
        RECT 92.755 176.515 92.925 176.685 ;
        RECT 96.895 176.515 97.065 176.705 ;
        RECT 97.355 176.495 97.525 176.705 ;
        RECT 97.815 176.495 97.985 176.685 ;
        RECT 98.730 176.545 98.850 176.655 ;
        RECT 99.195 176.515 99.365 176.705 ;
        RECT 101.995 176.685 102.125 176.705 ;
        RECT 101.955 176.495 102.125 176.685 ;
        RECT 102.410 176.545 102.530 176.655 ;
        RECT 105.635 176.495 105.805 176.685 ;
        RECT 106.100 176.495 106.270 176.685 ;
        RECT 107.930 176.515 108.100 176.705 ;
        RECT 108.395 176.515 108.565 176.705 ;
        RECT 109.770 176.545 109.890 176.655 ;
        RECT 110.240 176.495 110.410 176.685 ;
        RECT 112.085 176.550 112.245 176.660 ;
        RECT 113.455 176.515 113.625 176.705 ;
        RECT 113.910 176.545 114.030 176.655 ;
        RECT 116.675 176.495 116.845 176.685 ;
        RECT 117.135 176.495 117.305 176.685 ;
        RECT 118.515 176.495 118.685 176.685 ;
        RECT 120.815 176.515 120.985 176.705 ;
        RECT 128.175 176.515 128.345 176.705 ;
        RECT 129.555 176.495 129.725 176.685 ;
        RECT 85.255 176.265 88.320 176.465 ;
        RECT 85.255 175.785 88.465 176.265 ;
        RECT 88.475 175.815 90.765 176.495 ;
        RECT 90.775 175.815 93.525 176.495 ;
        RECT 85.255 175.585 86.205 175.785 ;
        RECT 87.535 175.585 88.465 175.785 ;
        RECT 89.845 175.585 90.765 175.815 ;
        RECT 92.595 175.585 93.525 175.815 ;
        RECT 93.535 175.585 97.665 176.495 ;
        RECT 97.685 175.585 99.035 176.495 ;
        RECT 99.985 175.625 100.415 176.410 ;
        RECT 100.435 175.585 102.250 176.495 ;
        RECT 102.735 175.585 105.945 176.495 ;
        RECT 105.955 175.585 109.430 176.495 ;
        RECT 110.095 175.815 113.765 176.495 ;
        RECT 114.235 175.815 116.985 176.495 ;
        RECT 110.095 175.585 111.020 175.815 ;
        RECT 114.235 175.585 115.165 175.815 ;
        RECT 116.995 175.685 118.365 176.495 ;
        RECT 118.375 175.815 125.685 176.495 ;
        RECT 121.890 175.595 122.800 175.815 ;
        RECT 124.335 175.585 125.685 175.815 ;
        RECT 125.745 175.625 126.175 176.410 ;
        RECT 126.290 175.815 129.755 176.495 ;
        RECT 130.020 176.465 130.190 176.685 ;
        RECT 130.935 176.515 131.105 176.705 ;
        RECT 132.780 176.655 132.950 176.685 ;
        RECT 132.770 176.545 132.950 176.655 ;
        RECT 131.680 176.465 132.625 176.495 ;
        RECT 132.780 176.465 132.950 176.545 ;
        RECT 136.915 176.515 137.085 176.705 ;
        RECT 137.375 176.515 137.545 176.705 ;
        RECT 137.835 176.495 138.005 176.685 ;
        RECT 138.290 176.545 138.410 176.655 ;
        RECT 139.215 176.515 139.385 176.705 ;
        RECT 140.135 176.495 140.305 176.685 ;
        RECT 140.595 176.495 140.765 176.685 ;
        RECT 143.355 176.495 143.525 176.685 ;
        RECT 143.815 176.515 143.985 176.705 ;
        RECT 144.735 176.495 144.905 176.685 ;
        RECT 147.490 176.515 147.660 176.705 ;
        RECT 147.955 176.495 148.125 176.705 ;
        RECT 148.415 176.495 148.585 176.685 ;
        RECT 149.790 176.495 149.960 176.685 ;
        RECT 155.315 176.655 155.485 176.685 ;
        RECT 151.170 176.545 151.290 176.655 ;
        RECT 155.310 176.545 155.485 176.655 ;
        RECT 155.315 176.495 155.485 176.545 ;
        RECT 156.695 176.495 156.865 176.705 ;
        RECT 134.440 176.465 135.385 176.495 ;
        RECT 126.290 175.585 127.210 175.815 ;
        RECT 129.875 175.785 132.625 176.465 ;
        RECT 132.635 175.785 135.385 176.465 ;
        RECT 131.680 175.585 132.625 175.785 ;
        RECT 134.440 175.585 135.385 175.785 ;
        RECT 135.405 175.585 138.135 176.495 ;
        RECT 138.615 175.585 140.430 176.495 ;
        RECT 140.455 175.685 142.285 176.495 ;
        RECT 142.305 175.585 143.655 176.495 ;
        RECT 144.595 175.815 146.885 176.495 ;
        RECT 145.965 175.585 146.885 175.815 ;
        RECT 146.905 175.585 148.255 176.495 ;
        RECT 148.275 175.685 149.645 176.495 ;
        RECT 149.675 175.585 151.025 176.495 ;
        RECT 151.505 175.625 151.935 176.410 ;
        RECT 152.050 175.815 155.515 176.495 ;
        RECT 152.050 175.585 152.970 175.815 ;
        RECT 155.635 175.685 157.005 176.495 ;
      LAYER nwell ;
        RECT 22.500 172.465 157.200 175.295 ;
      LAYER pwell ;
        RECT 22.695 171.265 24.065 172.075 ;
        RECT 27.590 171.945 28.500 172.165 ;
        RECT 30.035 171.945 31.385 172.175 ;
        RECT 24.075 171.265 31.385 171.945 ;
        RECT 31.435 171.265 33.265 172.075 ;
        RECT 34.325 171.945 35.255 172.175 ;
        RECT 33.420 171.265 35.255 171.945 ;
        RECT 35.585 171.350 36.015 172.135 ;
        RECT 36.495 171.265 37.865 172.045 ;
        RECT 37.875 171.265 41.545 172.075 ;
        RECT 42.475 171.945 43.610 172.175 ;
        RECT 42.475 171.265 45.685 171.945 ;
        RECT 45.695 171.265 48.445 172.175 ;
        RECT 48.455 171.265 53.965 172.075 ;
        RECT 53.975 171.265 55.345 172.075 ;
        RECT 55.355 171.945 56.490 172.175 ;
        RECT 55.355 171.265 58.565 171.945 ;
        RECT 58.585 171.265 59.935 172.175 ;
        RECT 59.965 171.265 61.315 172.175 ;
        RECT 61.345 171.350 61.775 172.135 ;
        RECT 62.255 171.265 65.465 172.175 ;
        RECT 65.570 171.945 66.490 172.175 ;
        RECT 73.130 171.945 74.040 172.165 ;
        RECT 75.575 171.945 76.925 172.175 ;
        RECT 80.490 171.945 81.400 172.165 ;
        RECT 82.935 171.945 84.285 172.175 ;
        RECT 65.570 171.265 69.035 171.945 ;
        RECT 69.615 171.265 76.925 171.945 ;
        RECT 76.975 171.265 84.285 171.945 ;
        RECT 84.335 171.265 85.705 172.045 ;
        RECT 85.715 171.265 87.085 172.075 ;
        RECT 87.105 171.350 87.535 172.135 ;
        RECT 87.650 171.945 88.570 172.175 ;
        RECT 87.650 171.265 91.115 171.945 ;
        RECT 91.255 171.265 92.605 172.175 ;
        RECT 95.340 171.975 96.285 172.175 ;
        RECT 93.535 171.295 96.285 171.975 ;
        RECT 22.835 171.055 23.005 171.265 ;
        RECT 24.215 171.055 24.385 171.265 ;
        RECT 29.735 171.055 29.905 171.245 ;
        RECT 31.115 171.075 31.285 171.245 ;
        RECT 31.575 171.075 31.745 171.265 ;
        RECT 33.420 171.245 33.585 171.265 ;
        RECT 33.415 171.075 33.590 171.245 ;
        RECT 36.170 171.105 36.290 171.215 ;
        RECT 36.635 171.075 36.805 171.265 ;
        RECT 38.015 171.075 38.185 171.265 ;
        RECT 31.135 171.055 31.285 171.075 ;
        RECT 22.695 170.245 24.065 171.055 ;
        RECT 24.075 170.245 29.585 171.055 ;
        RECT 29.595 170.245 30.965 171.055 ;
        RECT 31.135 170.235 33.065 171.055 ;
        RECT 33.420 171.025 33.590 171.075 ;
        RECT 38.475 171.055 38.645 171.245 ;
        RECT 39.855 171.055 40.025 171.245 ;
        RECT 40.315 171.055 40.485 171.245 ;
        RECT 41.705 171.110 41.865 171.220 ;
        RECT 42.150 171.105 42.270 171.215 ;
        RECT 42.615 171.055 42.785 171.245 ;
        RECT 45.375 171.075 45.545 171.265 ;
        RECT 45.840 171.245 46.010 171.265 ;
        RECT 45.835 171.075 46.010 171.245 ;
        RECT 48.595 171.075 48.765 171.265 ;
        RECT 54.115 171.245 54.285 171.265 ;
        RECT 45.835 171.055 46.005 171.075 ;
        RECT 35.550 171.025 36.485 171.055 ;
        RECT 33.420 170.825 36.485 171.025 ;
        RECT 32.115 170.145 33.065 170.235 ;
        RECT 33.275 170.345 36.485 170.825 ;
        RECT 33.275 170.145 34.205 170.345 ;
        RECT 35.535 170.145 36.485 170.345 ;
        RECT 36.495 170.375 38.785 171.055 ;
        RECT 36.495 170.145 37.415 170.375 ;
        RECT 38.795 170.275 40.165 171.055 ;
        RECT 40.175 170.245 42.005 171.055 ;
        RECT 42.475 170.375 45.685 171.055 ;
        RECT 44.550 170.145 45.685 170.375 ;
        RECT 45.695 170.245 48.445 171.055 ;
        RECT 49.060 171.025 49.230 171.245 ;
        RECT 51.815 171.055 51.985 171.245 ;
        RECT 53.650 171.105 53.770 171.215 ;
        RECT 54.115 171.075 54.290 171.245 ;
        RECT 54.120 171.055 54.290 171.075 ;
        RECT 57.335 171.055 57.505 171.245 ;
        RECT 57.795 171.055 57.965 171.245 ;
        RECT 58.255 171.075 58.425 171.265 ;
        RECT 58.715 171.075 58.885 171.265 ;
        RECT 61.015 171.075 61.185 171.265 ;
        RECT 61.930 171.105 62.050 171.215 ;
        RECT 62.395 171.075 62.565 171.265 ;
        RECT 67.455 171.055 67.625 171.245 ;
        RECT 67.910 171.105 68.030 171.215 ;
        RECT 68.835 171.075 69.005 171.265 ;
        RECT 69.290 171.105 69.410 171.215 ;
        RECT 69.755 171.075 69.925 171.265 ;
        RECT 70.210 171.055 70.380 171.245 ;
        RECT 70.675 171.055 70.845 171.245 ;
        RECT 73.890 171.105 74.010 171.215 ;
        RECT 74.815 171.055 74.985 171.245 ;
        RECT 77.115 171.075 77.285 171.265 ;
        RECT 78.955 171.055 79.125 171.245 ;
        RECT 82.175 171.055 82.345 171.245 ;
        RECT 85.395 171.075 85.565 171.265 ;
        RECT 85.855 171.055 86.025 171.265 ;
        RECT 86.315 171.055 86.485 171.245 ;
        RECT 89.995 171.055 90.165 171.245 ;
        RECT 90.915 171.075 91.085 171.265 ;
        RECT 50.720 171.025 51.665 171.055 ;
        RECT 48.465 170.185 48.895 170.970 ;
        RECT 48.915 170.345 51.665 171.025 ;
        RECT 50.720 170.145 51.665 170.345 ;
        RECT 51.675 170.245 53.505 171.055 ;
        RECT 53.975 170.145 55.805 171.055 ;
        RECT 55.815 170.145 57.630 171.055 ;
        RECT 57.655 170.245 60.405 171.055 ;
        RECT 60.455 170.375 67.765 171.055 ;
        RECT 60.455 170.145 61.805 170.375 ;
        RECT 63.340 170.155 64.250 170.375 ;
        RECT 68.315 170.145 70.525 171.055 ;
        RECT 70.535 170.145 73.745 171.055 ;
        RECT 74.225 170.185 74.655 170.970 ;
        RECT 74.675 170.245 76.045 171.055 ;
        RECT 76.055 170.145 79.265 171.055 ;
        RECT 79.275 170.145 82.485 171.055 ;
        RECT 82.590 170.375 86.055 171.055 ;
        RECT 82.590 170.145 83.510 170.375 ;
        RECT 86.175 170.245 89.845 171.055 ;
        RECT 89.855 170.245 91.225 171.055 ;
        RECT 91.380 171.025 91.550 171.245 ;
        RECT 92.290 171.075 92.460 171.265 ;
        RECT 92.765 171.110 92.925 171.220 ;
        RECT 93.680 171.075 93.850 171.295 ;
        RECT 95.340 171.265 96.285 171.295 ;
        RECT 96.305 171.265 99.035 172.175 ;
        RECT 99.055 171.265 104.565 172.075 ;
        RECT 104.575 171.265 110.085 172.075 ;
        RECT 110.095 171.265 112.845 172.075 ;
        RECT 112.865 171.350 113.295 172.135 ;
        RECT 113.315 171.265 115.130 172.175 ;
        RECT 115.155 171.265 118.825 172.075 ;
        RECT 119.755 171.265 122.965 172.175 ;
        RECT 122.975 171.265 128.485 172.075 ;
        RECT 128.955 171.265 130.305 172.175 ;
        RECT 130.335 171.265 132.165 172.075 ;
        RECT 132.270 171.945 133.190 172.175 ;
        RECT 132.270 171.265 135.735 171.945 ;
        RECT 135.855 171.265 138.605 172.075 ;
        RECT 138.625 171.350 139.055 172.135 ;
        RECT 139.075 171.265 142.745 172.075 ;
        RECT 142.935 171.495 145.270 172.175 ;
        RECT 142.935 171.265 144.785 171.495 ;
        RECT 145.515 171.265 148.265 172.075 ;
        RECT 151.790 171.945 152.700 172.165 ;
        RECT 154.235 171.945 155.585 172.175 ;
        RECT 148.275 171.265 155.585 171.945 ;
        RECT 155.635 171.265 157.005 172.075 ;
        RECT 94.135 171.055 94.305 171.245 ;
        RECT 96.895 171.055 97.065 171.245 ;
        RECT 98.735 171.075 98.905 171.265 ;
        RECT 99.195 171.075 99.365 171.265 ;
        RECT 99.650 171.105 99.770 171.215 ;
        RECT 104.715 171.075 104.885 171.265 ;
        RECT 107.475 171.055 107.645 171.245 ;
        RECT 107.935 171.055 108.105 171.245 ;
        RECT 109.775 171.055 109.945 171.245 ;
        RECT 110.235 171.075 110.405 171.265 ;
        RECT 114.835 171.075 115.005 171.265 ;
        RECT 115.295 171.075 115.465 171.265 ;
        RECT 118.985 171.110 119.145 171.220 ;
        RECT 120.355 171.055 120.525 171.245 ;
        RECT 122.655 171.075 122.825 171.265 ;
        RECT 123.115 171.245 123.285 171.265 ;
        RECT 123.110 171.075 123.285 171.245 ;
        RECT 123.110 171.055 123.280 171.075 ;
        RECT 123.575 171.055 123.745 171.245 ;
        RECT 125.410 171.105 125.530 171.215 ;
        RECT 126.335 171.055 126.505 171.245 ;
        RECT 128.630 171.105 128.750 171.215 ;
        RECT 129.555 171.055 129.725 171.245 ;
        RECT 130.020 171.075 130.190 171.265 ;
        RECT 130.475 171.075 130.645 171.265 ;
        RECT 135.535 171.075 135.705 171.265 ;
        RECT 135.995 171.075 136.165 171.265 ;
        RECT 136.915 171.055 137.085 171.245 ;
        RECT 138.300 171.055 138.470 171.245 ;
        RECT 139.215 171.075 139.385 171.265 ;
        RECT 142.935 171.245 143.065 171.265 ;
        RECT 139.675 171.055 139.845 171.245 ;
        RECT 142.895 171.055 143.065 171.245 ;
        RECT 144.280 171.055 144.450 171.245 ;
        RECT 145.655 171.075 145.825 171.265 ;
        RECT 148.415 171.075 148.585 171.265 ;
        RECT 149.795 171.055 149.965 171.245 ;
        RECT 151.175 171.055 151.345 171.245 ;
        RECT 152.095 171.075 152.265 171.245 ;
        RECT 152.100 171.055 152.265 171.075 ;
        RECT 154.395 171.055 154.565 171.245 ;
        RECT 156.695 171.055 156.865 171.265 ;
        RECT 93.040 171.025 93.985 171.055 ;
        RECT 91.235 170.345 93.985 171.025 ;
        RECT 93.995 170.375 96.745 171.055 ;
        RECT 93.040 170.145 93.985 170.345 ;
        RECT 95.815 170.145 96.745 170.375 ;
        RECT 96.755 170.245 99.505 171.055 ;
        RECT 99.985 170.185 100.415 170.970 ;
        RECT 100.475 170.375 107.785 171.055 ;
        RECT 100.475 170.145 101.825 170.375 ;
        RECT 103.360 170.155 104.270 170.375 ;
        RECT 107.795 170.245 109.625 171.055 ;
        RECT 109.635 170.375 116.945 171.055 ;
        RECT 113.150 170.155 114.060 170.375 ;
        RECT 115.595 170.145 116.945 170.375 ;
        RECT 117.090 170.375 120.555 171.055 ;
        RECT 117.090 170.145 118.010 170.375 ;
        RECT 120.815 170.145 123.425 171.055 ;
        RECT 123.435 170.245 125.265 171.055 ;
        RECT 125.745 170.185 126.175 170.970 ;
        RECT 126.295 170.145 129.405 171.055 ;
        RECT 129.415 170.375 136.725 171.055 ;
        RECT 132.930 170.155 133.840 170.375 ;
        RECT 135.375 170.145 136.725 170.375 ;
        RECT 136.775 170.245 138.145 171.055 ;
        RECT 138.155 170.145 139.505 171.055 ;
        RECT 139.535 170.145 142.745 171.055 ;
        RECT 142.755 170.245 144.125 171.055 ;
        RECT 144.135 170.375 147.720 171.055 ;
        RECT 147.815 170.375 150.105 171.055 ;
        RECT 144.135 170.145 145.055 170.375 ;
        RECT 147.815 170.145 148.735 170.375 ;
        RECT 150.125 170.145 151.475 171.055 ;
        RECT 151.505 170.185 151.935 170.970 ;
        RECT 152.100 170.375 153.935 171.055 ;
        RECT 153.005 170.145 153.935 170.375 ;
        RECT 154.265 170.145 155.615 171.055 ;
        RECT 155.635 170.245 157.005 171.055 ;
      LAYER nwell ;
        RECT 22.500 167.025 157.200 169.855 ;
      LAYER pwell ;
        RECT 22.695 165.825 24.065 166.635 ;
        RECT 27.590 166.505 28.500 166.725 ;
        RECT 30.035 166.505 31.385 166.735 ;
        RECT 24.075 165.825 31.385 166.505 ;
        RECT 31.435 166.535 32.385 166.735 ;
        RECT 33.715 166.535 34.645 166.735 ;
        RECT 31.435 166.055 34.645 166.535 ;
        RECT 31.435 165.855 34.500 166.055 ;
        RECT 35.585 165.910 36.015 166.695 ;
        RECT 40.470 166.505 41.380 166.725 ;
        RECT 42.915 166.505 44.265 166.735 ;
        RECT 31.435 165.825 32.370 165.855 ;
        RECT 22.835 165.615 23.005 165.825 ;
        RECT 24.215 165.615 24.385 165.825 ;
        RECT 34.330 165.805 34.500 165.855 ;
        RECT 36.955 165.825 44.265 166.505 ;
        RECT 44.315 165.825 47.235 166.735 ;
        RECT 47.535 165.825 48.905 166.635 ;
        RECT 51.655 166.505 52.585 166.735 ;
        RECT 48.915 165.825 52.585 166.505 ;
        RECT 52.595 166.535 53.540 166.735 ;
        RECT 52.595 165.855 55.345 166.535 ;
        RECT 55.435 166.055 58.495 166.735 ;
        RECT 52.595 165.825 53.540 165.855 ;
        RECT 26.975 165.615 27.145 165.805 ;
        RECT 27.435 165.615 27.605 165.805 ;
        RECT 31.125 165.660 31.285 165.770 ;
        RECT 33.875 165.635 34.045 165.805 ;
        RECT 34.330 165.635 34.505 165.805 ;
        RECT 34.805 165.670 34.965 165.780 ;
        RECT 36.185 165.670 36.345 165.780 ;
        RECT 37.095 165.775 37.265 165.825 ;
        RECT 44.460 165.805 44.630 165.825 ;
        RECT 37.090 165.665 37.265 165.775 ;
        RECT 37.095 165.635 37.265 165.665 ;
        RECT 33.875 165.615 34.040 165.635 ;
        RECT 34.335 165.615 34.505 165.635 ;
        RECT 22.695 164.805 24.065 165.615 ;
        RECT 24.075 164.805 25.905 165.615 ;
        RECT 25.915 164.835 27.285 165.615 ;
        RECT 27.295 164.805 30.965 165.615 ;
        RECT 32.205 164.935 34.040 165.615 ;
        RECT 32.205 164.705 33.135 164.935 ;
        RECT 34.195 164.805 36.945 165.615 ;
        RECT 37.560 165.585 37.730 165.805 ;
        RECT 40.775 165.615 40.945 165.805 ;
        RECT 44.455 165.635 44.630 165.805 ;
        RECT 44.455 165.615 44.625 165.635 ;
        RECT 45.835 165.615 46.005 165.805 ;
        RECT 47.675 165.635 47.845 165.825 ;
        RECT 49.055 165.805 49.225 165.825 ;
        RECT 49.055 165.635 49.230 165.805 ;
        RECT 39.690 165.585 40.625 165.615 ;
        RECT 37.560 165.385 40.625 165.585 ;
        RECT 37.415 164.905 40.625 165.385 ;
        RECT 37.415 164.705 38.345 164.905 ;
        RECT 39.675 164.705 40.625 164.905 ;
        RECT 40.635 164.805 44.305 165.615 ;
        RECT 44.315 164.805 45.685 165.615 ;
        RECT 45.695 164.935 48.445 165.615 ;
        RECT 49.060 165.585 49.230 165.635 ;
        RECT 53.195 165.615 53.365 165.805 ;
        RECT 53.665 165.660 53.825 165.770 ;
        RECT 54.570 165.615 54.740 165.805 ;
        RECT 55.030 165.635 55.200 165.855 ;
        RECT 55.435 165.825 58.425 166.055 ;
        RECT 58.575 165.825 61.325 166.635 ;
        RECT 61.345 165.910 61.775 166.695 ;
        RECT 61.795 165.825 64.545 166.635 ;
        RECT 65.015 165.825 68.225 166.735 ;
        RECT 68.330 166.505 69.250 166.735 ;
        RECT 68.330 165.825 71.795 166.505 ;
        RECT 71.915 165.825 73.745 166.635 ;
        RECT 73.840 165.825 82.945 166.505 ;
        RECT 83.035 165.825 85.245 166.735 ;
        RECT 85.255 165.825 87.085 166.635 ;
        RECT 87.105 165.910 87.535 166.695 ;
        RECT 88.925 166.505 89.845 166.735 ;
        RECT 87.555 165.825 89.845 166.505 ;
        RECT 89.855 165.825 91.685 166.735 ;
        RECT 91.695 165.825 97.205 166.635 ;
        RECT 97.215 165.825 100.885 166.635 ;
        RECT 100.895 165.825 102.265 166.635 ;
        RECT 104.930 166.505 105.850 166.735 ;
        RECT 102.385 165.825 105.850 166.505 ;
        RECT 105.955 165.825 109.165 166.735 ;
        RECT 109.175 165.825 112.385 166.735 ;
        RECT 112.865 165.910 113.295 166.695 ;
        RECT 113.325 165.825 114.675 166.735 ;
        RECT 115.155 165.825 118.365 166.735 ;
        RECT 122.350 166.505 123.260 166.725 ;
        RECT 124.795 166.505 126.145 166.735 ;
        RECT 118.835 165.825 126.145 166.505 ;
        RECT 126.195 165.825 129.405 166.735 ;
        RECT 132.930 166.505 133.840 166.725 ;
        RECT 135.375 166.505 136.725 166.735 ;
        RECT 129.415 165.825 136.725 166.505 ;
        RECT 136.775 165.825 138.605 166.635 ;
        RECT 138.625 165.910 139.055 166.695 ;
        RECT 139.170 166.505 140.090 166.735 ;
        RECT 139.170 165.825 142.635 166.505 ;
        RECT 142.950 165.825 146.425 166.735 ;
        RECT 146.895 165.825 148.265 166.605 ;
        RECT 148.315 166.505 149.665 166.735 ;
        RECT 151.200 166.505 152.110 166.725 ;
        RECT 148.315 165.825 155.625 166.505 ;
        RECT 155.635 165.825 157.005 166.635 ;
        RECT 58.255 165.635 58.425 165.825 ;
        RECT 58.715 165.635 58.885 165.825 ;
        RECT 59.635 165.635 59.805 165.805 ;
        RECT 59.635 165.615 59.785 165.635 ;
        RECT 60.095 165.615 60.265 165.805 ;
        RECT 61.935 165.635 62.105 165.825 ;
        RECT 62.850 165.665 62.970 165.775 ;
        RECT 63.315 165.615 63.485 165.805 ;
        RECT 64.690 165.665 64.810 165.775 ;
        RECT 65.160 165.635 65.330 165.825 ;
        RECT 71.595 165.635 71.765 165.825 ;
        RECT 72.055 165.635 72.225 165.825 ;
        RECT 73.895 165.615 74.065 165.805 ;
        RECT 74.815 165.615 74.985 165.805 ;
        RECT 76.650 165.665 76.770 165.775 ;
        RECT 77.115 165.615 77.285 165.805 ;
        RECT 82.635 165.635 82.805 165.825 ;
        RECT 84.485 165.660 84.645 165.770 ;
        RECT 84.930 165.635 85.100 165.825 ;
        RECT 85.395 165.635 85.565 165.825 ;
        RECT 87.695 165.635 87.865 165.825 ;
        RECT 91.370 165.635 91.540 165.825 ;
        RECT 91.835 165.635 92.005 165.825 ;
        RECT 92.295 165.615 92.465 165.805 ;
        RECT 97.355 165.635 97.525 165.825 ;
        RECT 99.655 165.615 99.825 165.805 ;
        RECT 101.035 165.635 101.205 165.825 ;
        RECT 102.415 165.635 102.585 165.825 ;
        RECT 102.875 165.615 103.045 165.805 ;
        RECT 104.260 165.615 104.430 165.805 ;
        RECT 104.720 165.615 104.890 165.805 ;
        RECT 106.095 165.615 106.265 165.805 ;
        RECT 107.930 165.665 108.050 165.775 ;
        RECT 108.855 165.635 109.025 165.825 ;
        RECT 111.155 165.615 111.325 165.805 ;
        RECT 111.615 165.615 111.785 165.805 ;
        RECT 112.075 165.635 112.245 165.825 ;
        RECT 112.530 165.665 112.650 165.775 ;
        RECT 114.375 165.635 114.545 165.825 ;
        RECT 114.830 165.665 114.950 165.775 ;
        RECT 116.215 165.615 116.385 165.805 ;
        RECT 118.050 165.635 118.220 165.825 ;
        RECT 118.510 165.615 118.680 165.805 ;
        RECT 118.975 165.775 119.145 165.825 ;
        RECT 118.970 165.665 119.145 165.775 ;
        RECT 118.975 165.635 119.145 165.665 ;
        RECT 122.195 165.615 122.365 165.805 ;
        RECT 122.655 165.615 122.825 165.805 ;
        RECT 125.410 165.665 125.530 165.775 ;
        RECT 126.335 165.635 126.505 165.825 ;
        RECT 129.555 165.615 129.725 165.825 ;
        RECT 130.015 165.615 130.185 165.805 ;
        RECT 134.615 165.615 134.785 165.805 ;
        RECT 136.915 165.635 137.085 165.825 ;
        RECT 138.295 165.615 138.465 165.805 ;
        RECT 138.755 165.615 138.925 165.805 ;
        RECT 142.435 165.635 142.605 165.825 ;
        RECT 144.275 165.615 144.445 165.805 ;
        RECT 146.110 165.635 146.280 165.825 ;
        RECT 146.570 165.665 146.690 165.775 ;
        RECT 147.035 165.635 147.205 165.825 ;
        RECT 147.955 165.615 148.125 165.805 ;
        RECT 148.415 165.635 148.585 165.805 ;
        RECT 151.170 165.665 151.290 165.775 ;
        RECT 148.565 165.615 148.585 165.635 ;
        RECT 152.095 165.615 152.265 165.805 ;
        RECT 155.315 165.615 155.485 165.825 ;
        RECT 156.695 165.615 156.865 165.825 ;
        RECT 50.720 165.585 51.665 165.615 ;
        RECT 47.515 164.705 48.445 164.935 ;
        RECT 48.465 164.745 48.895 165.530 ;
        RECT 48.915 164.905 51.665 165.585 ;
        RECT 50.720 164.705 51.665 164.905 ;
        RECT 51.675 164.705 53.490 165.615 ;
        RECT 54.445 164.705 57.645 165.615 ;
        RECT 57.855 164.795 59.785 165.615 ;
        RECT 59.955 164.805 62.705 165.615 ;
        RECT 63.175 164.935 70.485 165.615 ;
        RECT 57.855 164.705 58.805 164.795 ;
        RECT 66.690 164.715 67.600 164.935 ;
        RECT 69.135 164.705 70.485 164.935 ;
        RECT 70.630 164.935 74.095 165.615 ;
        RECT 70.630 164.705 71.550 164.935 ;
        RECT 74.225 164.745 74.655 165.530 ;
        RECT 74.675 164.805 76.505 165.615 ;
        RECT 76.975 164.935 84.285 165.615 ;
        RECT 80.490 164.715 81.400 164.935 ;
        RECT 82.935 164.705 84.285 164.935 ;
        RECT 85.295 164.935 92.605 165.615 ;
        RECT 92.655 164.935 99.965 165.615 ;
        RECT 85.295 164.705 86.645 164.935 ;
        RECT 88.180 164.715 89.090 164.935 ;
        RECT 92.655 164.705 94.005 164.935 ;
        RECT 95.540 164.715 96.450 164.935 ;
        RECT 99.985 164.745 100.415 165.530 ;
        RECT 100.435 164.705 103.185 165.615 ;
        RECT 103.195 164.705 104.545 165.615 ;
        RECT 104.575 164.705 105.925 165.615 ;
        RECT 105.955 164.805 107.785 165.615 ;
        RECT 108.255 164.705 111.465 165.615 ;
        RECT 111.475 164.805 112.845 165.615 ;
        RECT 112.950 164.935 116.415 165.615 ;
        RECT 112.950 164.705 113.870 164.935 ;
        RECT 116.615 164.705 118.825 165.615 ;
        RECT 119.295 164.705 122.505 165.615 ;
        RECT 122.515 164.805 125.265 165.615 ;
        RECT 125.745 164.745 126.175 165.530 ;
        RECT 126.290 164.935 129.755 165.615 ;
        RECT 126.290 164.705 127.210 164.935 ;
        RECT 129.875 164.805 131.245 165.615 ;
        RECT 131.350 164.935 134.815 165.615 ;
        RECT 135.030 164.935 138.495 165.615 ;
        RECT 131.350 164.705 132.270 164.935 ;
        RECT 135.030 164.705 135.950 164.935 ;
        RECT 138.615 164.805 142.285 165.615 ;
        RECT 143.225 164.705 144.575 165.615 ;
        RECT 144.690 164.935 148.155 165.615 ;
        RECT 148.565 164.935 151.015 165.615 ;
        RECT 144.690 164.705 145.610 164.935 ;
        RECT 149.055 164.705 151.015 164.935 ;
        RECT 151.505 164.745 151.935 165.530 ;
        RECT 151.955 164.935 154.245 165.615 ;
        RECT 153.325 164.705 154.245 164.935 ;
        RECT 154.255 164.835 155.625 165.615 ;
        RECT 155.635 164.805 157.005 165.615 ;
      LAYER nwell ;
        RECT 22.500 161.585 157.200 164.415 ;
      LAYER pwell ;
        RECT 22.695 160.385 24.065 161.195 ;
        RECT 24.995 160.385 26.810 161.295 ;
        RECT 26.835 160.385 28.665 161.295 ;
        RECT 28.770 161.065 29.690 161.295 ;
        RECT 28.770 160.385 32.235 161.065 ;
        RECT 32.355 160.385 33.725 161.165 ;
        RECT 33.735 160.385 35.565 161.195 ;
        RECT 35.585 160.470 36.015 161.255 ;
        RECT 36.505 160.385 39.235 161.295 ;
        RECT 40.590 161.095 41.545 161.295 ;
        RECT 39.265 160.415 41.545 161.095 ;
        RECT 22.835 160.175 23.005 160.385 ;
        RECT 24.225 160.220 24.385 160.340 ;
        RECT 26.515 160.195 26.685 160.385 ;
        RECT 26.980 160.195 27.150 160.385 ;
        RECT 28.355 160.175 28.525 160.365 ;
        RECT 32.035 160.195 32.205 160.385 ;
        RECT 32.495 160.195 32.665 160.385 ;
        RECT 33.875 160.195 34.045 160.385 ;
        RECT 36.170 160.225 36.290 160.335 ;
        RECT 36.635 160.195 36.805 160.385 ;
        RECT 37.555 160.175 37.725 160.365 ;
        RECT 38.015 160.175 38.185 160.365 ;
        RECT 39.390 160.195 39.560 160.415 ;
        RECT 40.590 160.385 41.545 160.415 ;
        RECT 41.555 160.385 44.305 161.195 ;
        RECT 44.315 160.385 46.145 161.295 ;
        RECT 46.155 160.385 51.665 161.195 ;
        RECT 51.675 160.385 54.425 161.195 ;
        RECT 54.445 160.385 57.175 161.295 ;
        RECT 57.195 161.095 58.140 161.295 ;
        RECT 57.195 160.415 59.945 161.095 ;
        RECT 57.195 160.385 58.140 160.415 ;
        RECT 41.695 160.195 41.865 160.385 ;
        RECT 45.375 160.175 45.545 160.365 ;
        RECT 45.830 160.195 46.000 160.385 ;
        RECT 46.295 160.195 46.465 160.385 ;
        RECT 48.130 160.225 48.250 160.335 ;
        RECT 49.055 160.175 49.225 160.365 ;
        RECT 51.815 160.195 51.985 160.385 ;
        RECT 52.730 160.225 52.850 160.335 ;
        RECT 53.195 160.175 53.365 160.365 ;
        RECT 54.575 160.195 54.745 160.385 ;
        RECT 55.955 160.175 56.125 160.365 ;
        RECT 59.630 160.195 59.800 160.415 ;
        RECT 59.955 160.385 61.325 161.195 ;
        RECT 61.345 160.470 61.775 161.255 ;
        RECT 61.795 160.385 63.625 161.195 ;
        RECT 63.635 160.385 66.845 161.295 ;
        RECT 66.855 160.385 69.605 161.195 ;
        RECT 70.115 161.065 71.465 161.295 ;
        RECT 73.000 161.065 73.910 161.285 ;
        RECT 70.115 160.385 77.425 161.065 ;
        RECT 77.435 160.385 79.265 161.195 ;
        RECT 79.735 160.385 82.945 161.295 ;
        RECT 82.955 160.385 86.625 161.195 ;
        RECT 87.105 160.470 87.535 161.255 ;
        RECT 88.025 160.385 90.755 161.295 ;
        RECT 90.775 160.385 92.145 161.165 ;
        RECT 92.155 160.385 93.985 161.195 ;
        RECT 96.650 161.065 97.570 161.295 ;
        RECT 94.105 160.385 97.570 161.065 ;
        RECT 97.775 160.385 100.885 161.295 ;
        RECT 100.895 160.385 102.725 161.195 ;
        RECT 103.235 161.065 104.585 161.295 ;
        RECT 106.120 161.065 107.030 161.285 ;
        RECT 103.235 160.385 110.545 161.065 ;
        RECT 110.555 160.385 112.385 161.195 ;
        RECT 112.865 160.470 113.295 161.255 ;
        RECT 113.315 160.385 115.145 161.195 ;
        RECT 115.615 160.385 118.365 161.295 ;
        RECT 118.395 160.385 119.745 161.295 ;
        RECT 119.755 160.385 125.265 161.195 ;
        RECT 125.735 160.385 128.945 161.295 ;
        RECT 132.470 161.065 133.380 161.285 ;
        RECT 134.915 161.065 136.265 161.295 ;
        RECT 128.955 160.385 136.265 161.065 ;
        RECT 137.245 160.385 138.595 161.295 ;
        RECT 138.625 160.470 139.055 161.255 ;
        RECT 141.820 161.065 142.745 161.295 ;
        RECT 144.575 161.065 145.505 161.295 ;
        RECT 139.075 160.385 142.745 161.065 ;
        RECT 142.755 160.385 145.505 161.065 ;
        RECT 146.435 160.385 155.540 161.065 ;
        RECT 155.635 160.385 157.005 161.195 ;
        RECT 60.095 160.195 60.265 160.385 ;
        RECT 61.935 160.195 62.105 160.385 ;
        RECT 66.535 160.175 66.705 160.385 ;
        RECT 66.995 160.195 67.165 160.385 ;
        RECT 69.750 160.225 69.870 160.335 ;
        RECT 73.895 160.175 74.065 160.365 ;
        RECT 74.815 160.175 74.985 160.365 ;
        RECT 76.655 160.175 76.825 160.365 ;
        RECT 77.115 160.195 77.285 160.385 ;
        RECT 77.575 160.195 77.745 160.385 ;
        RECT 79.410 160.225 79.530 160.335 ;
        RECT 79.880 160.195 80.050 160.385 ;
        RECT 80.335 160.195 80.505 160.365 ;
        RECT 83.095 160.195 83.265 160.385 ;
        RECT 80.355 160.175 80.505 160.195 ;
        RECT 83.555 160.175 83.725 160.365 ;
        RECT 84.015 160.175 84.185 160.365 ;
        RECT 86.770 160.225 86.890 160.335 ;
        RECT 22.695 159.365 24.065 160.175 ;
        RECT 25.090 159.495 28.555 160.175 ;
        RECT 28.760 159.495 37.865 160.175 ;
        RECT 37.875 159.495 45.185 160.175 ;
        RECT 25.090 159.265 26.010 159.495 ;
        RECT 41.390 159.275 42.300 159.495 ;
        RECT 43.835 159.265 45.185 159.495 ;
        RECT 45.245 159.265 47.975 160.175 ;
        RECT 48.465 159.305 48.895 160.090 ;
        RECT 48.915 159.365 52.585 160.175 ;
        RECT 53.055 159.495 55.805 160.175 ;
        RECT 55.815 159.495 59.485 160.175 ;
        RECT 54.875 159.265 55.805 159.495 ;
        RECT 58.555 159.265 59.485 159.495 ;
        RECT 59.535 159.495 66.845 160.175 ;
        RECT 66.895 159.495 74.205 160.175 ;
        RECT 59.535 159.265 60.885 159.495 ;
        RECT 62.420 159.275 63.330 159.495 ;
        RECT 66.895 159.265 68.245 159.495 ;
        RECT 69.780 159.275 70.690 159.495 ;
        RECT 74.225 159.305 74.655 160.090 ;
        RECT 74.675 159.495 76.505 160.175 ;
        RECT 75.160 159.265 76.505 159.495 ;
        RECT 76.515 159.365 80.185 160.175 ;
        RECT 80.355 159.355 82.285 160.175 ;
        RECT 82.495 159.395 83.865 160.175 ;
        RECT 83.875 159.365 86.625 160.175 ;
        RECT 87.235 160.145 87.405 160.365 ;
        RECT 87.690 160.225 87.810 160.335 ;
        RECT 88.155 160.195 88.325 160.385 ;
        RECT 90.455 160.175 90.625 160.365 ;
        RECT 91.835 160.195 92.005 160.385 ;
        RECT 92.295 160.195 92.465 160.385 ;
        RECT 93.215 160.175 93.385 160.365 ;
        RECT 94.135 160.195 94.305 160.385 ;
        RECT 94.595 160.195 94.765 160.365 ;
        RECT 94.615 160.175 94.765 160.195 ;
        RECT 96.895 160.175 97.065 160.365 ;
        RECT 97.815 160.195 97.985 160.385 ;
        RECT 98.275 160.175 98.445 160.365 ;
        RECT 101.035 160.195 101.205 160.385 ;
        RECT 102.870 160.225 102.990 160.335 ;
        RECT 109.315 160.175 109.485 160.365 ;
        RECT 109.775 160.175 109.945 160.365 ;
        RECT 110.235 160.195 110.405 160.385 ;
        RECT 110.695 160.195 110.865 160.385 ;
        RECT 112.530 160.225 112.650 160.335 ;
        RECT 113.455 160.195 113.625 160.385 ;
        RECT 115.290 160.225 115.410 160.335 ;
        RECT 118.055 160.175 118.225 160.385 ;
        RECT 118.515 160.175 118.685 160.365 ;
        RECT 119.430 160.195 119.600 160.385 ;
        RECT 119.895 160.195 120.065 160.385 ;
        RECT 122.195 160.175 122.365 160.365 ;
        RECT 123.575 160.175 123.745 160.365 ;
        RECT 124.965 160.220 125.125 160.330 ;
        RECT 125.410 160.225 125.530 160.335 ;
        RECT 125.875 160.195 126.045 160.385 ;
        RECT 126.335 160.175 126.505 160.365 ;
        RECT 129.095 160.195 129.265 160.385 ;
        RECT 129.555 160.175 129.725 160.365 ;
        RECT 136.465 160.230 136.625 160.340 ;
        RECT 136.915 160.175 137.085 160.365 ;
        RECT 137.375 160.195 137.545 160.385 ;
        RECT 141.055 160.175 141.225 160.365 ;
        RECT 141.515 160.175 141.685 160.365 ;
        RECT 142.430 160.195 142.600 160.385 ;
        RECT 142.895 160.195 143.065 160.385 ;
        RECT 145.665 160.230 145.825 160.340 ;
        RECT 146.575 160.195 146.745 160.385 ;
        RECT 151.175 160.175 151.345 160.365 ;
        RECT 153.935 160.195 154.105 160.365 ;
        RECT 153.935 160.175 154.100 160.195 ;
        RECT 154.390 160.175 154.560 160.365 ;
        RECT 156.695 160.175 156.865 160.385 ;
        RECT 89.360 160.145 90.305 160.175 ;
        RECT 87.235 159.945 90.305 160.145 ;
        RECT 87.095 159.465 90.305 159.945 ;
        RECT 90.315 159.495 93.055 160.175 ;
        RECT 81.335 159.265 82.285 159.355 ;
        RECT 87.095 159.265 88.025 159.465 ;
        RECT 89.360 159.265 90.305 159.465 ;
        RECT 93.075 159.365 94.445 160.175 ;
        RECT 94.615 159.355 96.545 160.175 ;
        RECT 96.755 159.395 98.125 160.175 ;
        RECT 98.135 159.365 99.965 160.175 ;
        RECT 95.595 159.265 96.545 159.355 ;
        RECT 99.985 159.305 100.415 160.090 ;
        RECT 100.520 159.495 109.625 160.175 ;
        RECT 109.635 159.495 116.945 160.175 ;
        RECT 113.150 159.275 114.060 159.495 ;
        RECT 115.595 159.265 116.945 159.495 ;
        RECT 116.995 159.395 118.365 160.175 ;
        RECT 118.375 159.365 122.045 160.175 ;
        RECT 122.055 159.365 123.425 160.175 ;
        RECT 123.435 159.395 124.805 160.175 ;
        RECT 125.745 159.305 126.175 160.090 ;
        RECT 126.195 159.265 129.405 160.175 ;
        RECT 129.415 159.495 136.725 160.175 ;
        RECT 132.930 159.275 133.840 159.495 ;
        RECT 135.375 159.265 136.725 159.495 ;
        RECT 136.775 159.365 139.525 160.175 ;
        RECT 139.535 159.265 141.350 160.175 ;
        RECT 141.375 159.365 144.125 160.175 ;
        RECT 144.175 159.495 151.485 160.175 ;
        RECT 144.175 159.265 145.525 159.495 ;
        RECT 147.060 159.275 147.970 159.495 ;
        RECT 151.505 159.305 151.935 160.090 ;
        RECT 152.265 159.495 154.100 160.175 ;
        RECT 152.265 159.265 153.195 159.495 ;
        RECT 154.275 159.265 155.625 160.175 ;
        RECT 155.635 159.365 157.005 160.175 ;
      LAYER nwell ;
        RECT 22.500 156.145 157.200 158.975 ;
      LAYER pwell ;
        RECT 22.695 154.945 24.065 155.755 ;
        RECT 27.590 155.625 28.500 155.845 ;
        RECT 30.035 155.625 31.385 155.855 ;
        RECT 24.075 154.945 31.385 155.625 ;
        RECT 32.355 155.655 33.285 155.855 ;
        RECT 34.615 155.655 35.565 155.855 ;
        RECT 32.355 155.175 35.565 155.655 ;
        RECT 32.500 154.975 35.565 155.175 ;
        RECT 35.585 155.030 36.015 155.815 ;
        RECT 37.405 155.625 38.325 155.855 ;
        RECT 41.850 155.625 42.760 155.845 ;
        RECT 44.295 155.625 45.645 155.855 ;
        RECT 22.835 154.735 23.005 154.945 ;
        RECT 24.215 154.735 24.385 154.945 ;
        RECT 26.975 154.735 27.145 154.925 ;
        RECT 27.435 154.735 27.605 154.925 ;
        RECT 31.585 154.790 31.745 154.900 ;
        RECT 32.500 154.755 32.670 154.975 ;
        RECT 34.630 154.945 35.565 154.975 ;
        RECT 36.035 154.945 38.325 155.625 ;
        RECT 38.335 154.945 45.645 155.625 ;
        RECT 46.175 154.945 47.525 155.855 ;
        RECT 51.050 155.625 51.960 155.845 ;
        RECT 53.495 155.625 55.265 155.855 ;
        RECT 47.535 154.945 55.265 155.625 ;
        RECT 55.355 154.945 56.725 155.755 ;
        RECT 56.735 155.655 57.680 155.855 ;
        RECT 56.735 154.975 59.485 155.655 ;
        RECT 56.735 154.945 57.680 154.975 ;
        RECT 32.955 154.735 33.125 154.925 ;
        RECT 36.175 154.755 36.345 154.945 ;
        RECT 38.475 154.755 38.645 154.945 ;
        RECT 40.315 154.735 40.485 154.925 ;
        RECT 42.615 154.735 42.785 154.925 ;
        RECT 43.085 154.780 43.245 154.890 ;
        RECT 43.995 154.735 44.165 154.925 ;
        RECT 45.830 154.785 45.950 154.895 ;
        RECT 46.290 154.755 46.460 154.945 ;
        RECT 47.215 154.735 47.385 154.925 ;
        RECT 47.675 154.755 47.845 154.945 ;
        RECT 49.050 154.785 49.170 154.895 ;
        RECT 49.515 154.735 49.685 154.925 ;
        RECT 52.735 154.735 52.905 154.925 ;
        RECT 55.495 154.755 55.665 154.945 ;
        RECT 57.795 154.735 57.965 154.925 ;
        RECT 59.170 154.755 59.340 154.975 ;
        RECT 59.495 154.945 61.325 155.755 ;
        RECT 61.345 155.030 61.775 155.815 ;
        RECT 64.450 155.625 65.370 155.855 ;
        RECT 61.905 154.945 65.370 155.625 ;
        RECT 65.475 154.945 66.845 155.755 ;
        RECT 69.510 155.625 70.430 155.855 ;
        RECT 74.970 155.625 75.880 155.845 ;
        RECT 77.415 155.625 78.765 155.855 ;
        RECT 82.330 155.625 83.240 155.845 ;
        RECT 84.775 155.625 86.125 155.855 ;
        RECT 66.965 154.945 70.430 155.625 ;
        RECT 71.455 154.945 78.765 155.625 ;
        RECT 78.815 154.945 86.125 155.625 ;
        RECT 87.105 155.030 87.535 155.815 ;
        RECT 88.040 155.625 91.650 155.855 ;
        RECT 93.065 155.625 93.985 155.855 ;
        RECT 87.555 154.945 91.650 155.625 ;
        RECT 91.695 154.945 93.985 155.625 ;
        RECT 94.035 155.625 95.385 155.855 ;
        RECT 96.920 155.625 97.830 155.845 ;
        RECT 94.035 154.945 101.345 155.625 ;
        RECT 101.355 154.945 104.105 155.755 ;
        RECT 106.770 155.625 107.690 155.855 ;
        RECT 104.225 154.945 107.690 155.625 ;
        RECT 107.795 154.945 111.005 155.855 ;
        RECT 111.015 154.945 112.845 155.755 ;
        RECT 112.865 155.030 113.295 155.815 ;
        RECT 117.750 155.625 118.660 155.845 ;
        RECT 120.195 155.625 121.545 155.855 ;
        RECT 114.235 154.945 121.545 155.625 ;
        RECT 121.795 155.765 122.745 155.855 ;
        RECT 121.795 154.945 123.725 155.765 ;
        RECT 124.395 155.625 125.745 155.855 ;
        RECT 127.280 155.625 128.190 155.845 ;
        RECT 124.395 154.945 131.705 155.625 ;
        RECT 131.715 154.945 137.225 155.755 ;
        RECT 137.235 154.945 138.605 155.725 ;
        RECT 138.625 155.030 139.055 155.815 ;
        RECT 139.075 154.945 144.585 155.755 ;
        RECT 144.595 154.945 148.265 155.755 ;
        RECT 151.790 155.625 152.700 155.845 ;
        RECT 154.235 155.625 155.585 155.855 ;
        RECT 148.275 154.945 155.585 155.625 ;
        RECT 155.635 154.945 157.005 155.755 ;
        RECT 59.635 154.755 59.805 154.945 ;
        RECT 22.695 153.925 24.065 154.735 ;
        RECT 24.075 153.925 25.905 154.735 ;
        RECT 25.915 153.955 27.285 154.735 ;
        RECT 27.295 153.925 32.805 154.735 ;
        RECT 32.815 153.925 38.325 154.735 ;
        RECT 39.255 153.955 40.625 154.735 ;
        RECT 40.635 154.055 42.925 154.735 ;
        RECT 40.635 153.825 41.555 154.055 ;
        RECT 43.955 153.825 47.065 154.735 ;
        RECT 47.075 153.925 48.445 154.735 ;
        RECT 48.465 153.865 48.895 154.650 ;
        RECT 49.475 153.825 52.585 154.735 ;
        RECT 52.595 153.925 54.425 154.735 ;
        RECT 54.530 154.055 57.995 154.735 ;
        RECT 58.115 154.705 59.060 154.735 ;
        RECT 60.550 154.705 60.720 154.925 ;
        RECT 61.015 154.735 61.185 154.925 ;
        RECT 61.935 154.755 62.105 154.945 ;
        RECT 62.850 154.785 62.970 154.895 ;
        RECT 63.315 154.735 63.485 154.925 ;
        RECT 65.615 154.755 65.785 154.945 ;
        RECT 66.995 154.755 67.165 154.945 ;
        RECT 69.295 154.735 69.465 154.925 ;
        RECT 69.755 154.735 69.925 154.925 ;
        RECT 70.685 154.790 70.845 154.900 ;
        RECT 71.595 154.755 71.765 154.945 ;
        RECT 73.895 154.735 74.065 154.925 ;
        RECT 74.810 154.785 74.930 154.895 ;
        RECT 78.035 154.735 78.205 154.925 ;
        RECT 78.955 154.755 79.125 154.945 ;
        RECT 81.715 154.735 81.885 154.925 ;
        RECT 82.185 154.780 82.345 154.890 ;
        RECT 83.370 154.735 83.540 154.925 ;
        RECT 86.325 154.790 86.485 154.900 ;
        RECT 87.230 154.785 87.350 154.895 ;
        RECT 87.700 154.755 87.870 154.945 ;
        RECT 91.835 154.755 92.005 154.945 ;
        RECT 94.590 154.735 94.760 154.925 ;
        RECT 95.065 154.780 95.225 154.890 ;
        RECT 96.250 154.735 96.420 154.925 ;
        RECT 101.035 154.755 101.205 154.945 ;
        RECT 101.495 154.735 101.665 154.945 ;
        RECT 101.955 154.735 102.125 154.925 ;
        RECT 104.255 154.755 104.425 154.945 ;
        RECT 104.715 154.735 104.885 154.925 ;
        RECT 106.095 154.735 106.265 154.925 ;
        RECT 107.935 154.755 108.105 154.945 ;
        RECT 111.155 154.755 111.325 154.945 ;
        RECT 113.455 154.735 113.625 154.925 ;
        RECT 114.375 154.755 114.545 154.945 ;
        RECT 123.575 154.925 123.725 154.945 ;
        RECT 118.700 154.735 118.870 154.925 ;
        RECT 121.275 154.755 121.445 154.925 ;
        RECT 121.275 154.735 121.425 154.755 ;
        RECT 122.655 154.735 122.825 154.925 ;
        RECT 123.110 154.785 123.230 154.895 ;
        RECT 123.575 154.755 123.745 154.925 ;
        RECT 124.030 154.785 124.150 154.895 ;
        RECT 123.595 154.735 123.745 154.755 ;
        RECT 126.610 154.735 126.780 154.925 ;
        RECT 130.470 154.785 130.590 154.895 ;
        RECT 130.935 154.735 131.105 154.925 ;
        RECT 131.395 154.755 131.565 154.945 ;
        RECT 131.855 154.755 132.025 154.945 ;
        RECT 132.315 154.735 132.485 154.925 ;
        RECT 134.150 154.785 134.270 154.895 ;
        RECT 134.615 154.735 134.785 154.925 ;
        RECT 138.295 154.755 138.465 154.945 ;
        RECT 139.215 154.755 139.385 154.945 ;
        RECT 143.815 154.735 143.985 154.925 ;
        RECT 144.735 154.755 144.905 154.945 ;
        RECT 148.415 154.755 148.585 154.945 ;
        RECT 149.335 154.735 149.505 154.925 ;
        RECT 151.170 154.785 151.290 154.895 ;
        RECT 155.315 154.735 155.485 154.925 ;
        RECT 156.695 154.735 156.865 154.945 ;
        RECT 54.530 153.825 55.450 154.055 ;
        RECT 58.115 154.025 60.865 154.705 ;
        RECT 58.115 153.825 59.060 154.025 ;
        RECT 60.875 153.925 62.705 154.735 ;
        RECT 63.175 153.825 66.385 154.735 ;
        RECT 66.395 153.825 69.605 154.735 ;
        RECT 69.615 154.055 72.365 154.735 ;
        RECT 71.435 153.825 72.365 154.055 ;
        RECT 72.375 154.055 74.205 154.735 ;
        RECT 72.375 153.825 73.720 154.055 ;
        RECT 74.225 153.865 74.655 154.650 ;
        RECT 75.135 153.825 78.345 154.735 ;
        RECT 78.450 154.055 81.915 154.735 ;
        RECT 82.955 154.055 86.855 154.735 ;
        RECT 78.450 153.825 79.370 154.055 ;
        RECT 82.955 153.825 83.885 154.055 ;
        RECT 87.795 153.825 94.905 154.735 ;
        RECT 95.835 154.055 99.735 154.735 ;
        RECT 95.835 153.825 96.765 154.055 ;
        RECT 99.985 153.865 100.415 154.650 ;
        RECT 100.435 153.955 101.805 154.735 ;
        RECT 101.815 153.925 104.565 154.735 ;
        RECT 104.575 153.955 105.945 154.735 ;
        RECT 105.955 154.055 113.265 154.735 ;
        RECT 109.470 153.835 110.380 154.055 ;
        RECT 111.915 153.825 113.265 154.055 ;
        RECT 113.315 153.925 115.145 154.735 ;
        RECT 115.385 154.055 119.285 154.735 ;
        RECT 118.355 153.825 119.285 154.055 ;
        RECT 119.495 153.915 121.425 154.735 ;
        RECT 121.595 153.955 122.965 154.735 ;
        RECT 123.595 153.915 125.525 154.735 ;
        RECT 119.495 153.825 120.445 153.915 ;
        RECT 124.575 153.825 125.525 153.915 ;
        RECT 125.745 153.865 126.175 154.650 ;
        RECT 126.195 154.055 130.095 154.735 ;
        RECT 126.195 153.825 127.125 154.055 ;
        RECT 130.805 153.825 132.155 154.735 ;
        RECT 132.175 153.925 134.005 154.735 ;
        RECT 134.475 154.055 143.580 154.735 ;
        RECT 143.675 153.925 149.185 154.735 ;
        RECT 149.195 153.925 151.025 154.735 ;
        RECT 151.505 153.865 151.935 154.650 ;
        RECT 152.050 154.055 155.515 154.735 ;
        RECT 152.050 153.825 152.970 154.055 ;
        RECT 155.635 153.925 157.005 154.735 ;
      LAYER nwell ;
        RECT 22.500 150.705 157.200 153.535 ;
      LAYER pwell ;
        RECT 22.695 149.505 24.065 150.315 ;
        RECT 27.590 150.185 28.500 150.405 ;
        RECT 30.035 150.185 31.385 150.415 ;
        RECT 24.075 149.505 31.385 150.185 ;
        RECT 31.435 149.505 32.805 150.315 ;
        RECT 32.835 149.505 34.185 150.415 ;
        RECT 34.195 149.505 35.565 150.315 ;
        RECT 35.585 149.590 36.015 150.375 ;
        RECT 36.035 149.505 37.405 150.315 ;
        RECT 37.900 150.185 39.245 150.415 ;
        RECT 37.415 149.505 39.245 150.185 ;
        RECT 39.395 149.505 42.005 150.415 ;
        RECT 42.015 150.185 42.935 150.415 ;
        RECT 45.790 150.185 46.710 150.415 ;
        RECT 42.015 149.505 45.600 150.185 ;
        RECT 45.790 149.505 49.255 150.185 ;
        RECT 49.375 149.505 58.480 150.185 ;
        RECT 58.575 149.505 61.325 150.315 ;
        RECT 61.345 149.590 61.775 150.375 ;
        RECT 61.795 149.505 64.715 150.415 ;
        RECT 66.385 150.185 67.305 150.415 ;
        RECT 65.015 149.505 67.305 150.185 ;
        RECT 67.775 149.505 70.985 150.415 ;
        RECT 70.995 150.185 73.820 150.415 ;
        RECT 78.250 150.185 79.170 150.415 ;
        RECT 70.995 149.505 74.525 150.185 ;
        RECT 75.705 149.505 79.170 150.185 ;
        RECT 79.275 149.505 82.485 150.415 ;
        RECT 82.495 149.505 85.245 150.415 ;
        RECT 85.255 149.505 87.085 150.315 ;
        RECT 87.105 149.590 87.535 150.375 ;
        RECT 87.635 149.505 89.845 150.415 ;
        RECT 90.315 150.215 91.265 150.415 ;
        RECT 92.595 150.215 93.525 150.415 ;
        RECT 90.315 149.735 93.525 150.215 ;
        RECT 93.545 149.735 96.745 150.415 ;
        RECT 97.895 150.325 98.845 150.415 ;
        RECT 90.315 149.535 93.380 149.735 ;
        RECT 90.315 149.505 91.250 149.535 ;
        RECT 22.835 149.295 23.005 149.505 ;
        RECT 24.215 149.315 24.385 149.505 ;
        RECT 25.135 149.295 25.305 149.485 ;
        RECT 27.895 149.295 28.065 149.485 ;
        RECT 31.575 149.315 31.745 149.505 ;
        RECT 31.575 149.295 31.725 149.315 ;
        RECT 32.035 149.295 32.205 149.485 ;
        RECT 33.870 149.315 34.040 149.505 ;
        RECT 34.335 149.315 34.505 149.505 ;
        RECT 36.175 149.315 36.345 149.505 ;
        RECT 37.555 149.315 37.725 149.505 ;
        RECT 39.390 149.345 39.510 149.455 ;
        RECT 39.855 149.295 40.025 149.485 ;
        RECT 41.690 149.315 41.860 149.505 ;
        RECT 42.160 149.315 42.330 149.505 ;
        RECT 48.140 149.295 48.310 149.485 ;
        RECT 49.055 149.295 49.225 149.505 ;
        RECT 49.515 149.315 49.685 149.505 ;
        RECT 50.895 149.295 51.065 149.485 ;
        RECT 58.265 149.340 58.425 149.450 ;
        RECT 58.715 149.315 58.885 149.505 ;
        RECT 61.940 149.485 62.110 149.505 ;
        RECT 61.935 149.315 62.110 149.485 ;
        RECT 61.935 149.295 62.105 149.315 ;
        RECT 62.400 149.295 62.570 149.485 ;
        RECT 65.155 149.315 65.325 149.505 ;
        RECT 67.450 149.345 67.570 149.455 ;
        RECT 67.915 149.315 68.085 149.505 ;
        RECT 74.325 149.485 74.525 149.505 ;
        RECT 71.135 149.295 71.305 149.485 ;
        RECT 72.515 149.295 72.685 149.485 ;
        RECT 72.975 149.295 73.145 149.485 ;
        RECT 74.355 149.315 74.525 149.485 ;
        RECT 74.825 149.455 74.985 149.460 ;
        RECT 74.810 149.350 74.985 149.455 ;
        RECT 74.810 149.345 74.930 149.350 ;
        RECT 75.735 149.315 75.905 149.505 ;
        RECT 79.415 149.315 79.585 149.505 ;
        RECT 82.175 149.295 82.345 149.485 ;
        RECT 82.635 149.295 82.805 149.505 ;
        RECT 84.015 149.295 84.185 149.485 ;
        RECT 85.395 149.315 85.565 149.505 ;
        RECT 87.705 149.340 87.865 149.450 ;
        RECT 88.615 149.315 88.785 149.485 ;
        RECT 89.530 149.315 89.700 149.505 ;
        RECT 89.990 149.345 90.110 149.455 ;
        RECT 88.635 149.295 88.785 149.315 ;
        RECT 91.190 149.295 91.360 149.485 ;
        RECT 93.210 149.315 93.380 149.535 ;
        RECT 93.545 149.505 96.600 149.735 ;
        RECT 95.055 149.295 95.225 149.485 ;
        RECT 96.430 149.315 96.600 149.505 ;
        RECT 96.915 149.505 98.845 150.325 ;
        RECT 102.570 150.185 103.480 150.405 ;
        RECT 105.015 150.185 106.365 150.415 ;
        RECT 99.055 149.505 106.365 150.185 ;
        RECT 106.415 150.185 107.345 150.415 ;
        RECT 110.755 150.325 111.705 150.415 ;
        RECT 106.415 149.505 110.315 150.185 ;
        RECT 110.755 149.505 112.685 150.325 ;
        RECT 112.865 149.590 113.295 150.375 ;
        RECT 122.975 150.185 123.905 150.415 ;
        RECT 113.775 149.505 122.880 150.185 ;
        RECT 122.975 149.505 126.875 150.185 ;
        RECT 127.115 149.505 129.865 150.315 ;
        RECT 130.335 149.505 133.085 150.415 ;
        RECT 133.565 149.505 134.915 150.415 ;
        RECT 134.945 149.505 136.295 150.415 ;
        RECT 137.685 150.185 138.605 150.415 ;
        RECT 136.315 149.505 138.605 150.185 ;
        RECT 138.625 149.590 139.055 150.375 ;
        RECT 139.085 149.505 141.815 150.415 ;
        RECT 142.395 149.505 145.505 150.415 ;
        RECT 145.535 149.505 146.885 150.415 ;
        RECT 146.935 150.185 148.285 150.415 ;
        RECT 149.820 150.185 150.730 150.405 ;
        RECT 146.935 149.505 154.245 150.185 ;
        RECT 154.255 149.505 155.625 150.315 ;
        RECT 155.635 149.505 157.005 150.315 ;
        RECT 96.915 149.485 97.065 149.505 ;
        RECT 96.895 149.315 97.065 149.485 ;
        RECT 98.735 149.295 98.905 149.485 ;
        RECT 99.195 149.315 99.365 149.505 ;
        RECT 100.850 149.295 101.020 149.485 ;
        RECT 104.710 149.345 104.830 149.455 ;
        RECT 105.175 149.295 105.345 149.485 ;
        RECT 106.555 149.295 106.725 149.485 ;
        RECT 106.830 149.315 107.000 149.505 ;
        RECT 112.535 149.485 112.685 149.505 ;
        RECT 112.535 149.315 112.705 149.485 ;
        RECT 113.450 149.345 113.570 149.455 ;
        RECT 113.915 149.315 114.085 149.505 ;
        RECT 114.835 149.295 115.005 149.485 ;
        RECT 123.115 149.295 123.285 149.485 ;
        RECT 123.390 149.315 123.560 149.505 ;
        RECT 125.415 149.315 125.585 149.485 ;
        RECT 125.415 149.295 125.565 149.315 ;
        RECT 126.335 149.295 126.505 149.485 ;
        RECT 127.255 149.315 127.425 149.505 ;
        RECT 129.090 149.345 129.210 149.455 ;
        RECT 130.010 149.345 130.130 149.455 ;
        RECT 130.475 149.315 130.645 149.505 ;
        RECT 132.770 149.295 132.940 149.485 ;
        RECT 133.235 149.455 133.405 149.485 ;
        RECT 133.230 149.345 133.405 149.455 ;
        RECT 133.235 149.295 133.405 149.345 ;
        RECT 134.615 149.295 134.785 149.505 ;
        RECT 135.995 149.315 136.165 149.505 ;
        RECT 136.455 149.315 136.625 149.505 ;
        RECT 139.215 149.315 139.385 149.505 ;
        RECT 141.975 149.455 142.145 149.485 ;
        RECT 141.970 149.345 142.145 149.455 ;
        RECT 141.975 149.295 142.145 149.345 ;
        RECT 142.435 149.315 142.605 149.505 ;
        RECT 22.695 148.485 24.065 149.295 ;
        RECT 24.995 148.615 27.745 149.295 ;
        RECT 26.815 148.385 27.745 148.615 ;
        RECT 27.755 148.485 29.585 149.295 ;
        RECT 29.795 148.475 31.725 149.295 ;
        RECT 31.895 148.615 39.205 149.295 ;
        RECT 39.715 148.615 47.025 149.295 ;
        RECT 29.795 148.385 30.745 148.475 ;
        RECT 35.410 148.395 36.320 148.615 ;
        RECT 37.855 148.385 39.205 148.615 ;
        RECT 43.230 148.395 44.140 148.615 ;
        RECT 45.675 148.385 47.025 148.615 ;
        RECT 47.075 148.385 48.425 149.295 ;
        RECT 48.465 148.425 48.895 149.210 ;
        RECT 48.915 148.485 50.745 149.295 ;
        RECT 50.755 148.615 58.065 149.295 ;
        RECT 54.270 148.395 55.180 148.615 ;
        RECT 56.715 148.385 58.065 148.615 ;
        RECT 59.035 148.615 62.245 149.295 ;
        RECT 59.035 148.385 60.170 148.615 ;
        RECT 62.255 148.385 64.085 149.295 ;
        RECT 64.135 148.615 71.445 149.295 ;
        RECT 64.135 148.385 65.485 148.615 ;
        RECT 67.020 148.395 67.930 148.615 ;
        RECT 71.455 148.515 72.825 149.295 ;
        RECT 72.835 148.485 74.205 149.295 ;
        RECT 74.225 148.425 74.655 149.210 ;
        RECT 75.175 148.615 82.485 149.295 ;
        RECT 75.175 148.385 76.525 148.615 ;
        RECT 78.060 148.395 78.970 148.615 ;
        RECT 82.505 148.385 83.855 149.295 ;
        RECT 83.875 148.485 87.545 149.295 ;
        RECT 88.635 148.475 90.565 149.295 ;
        RECT 89.615 148.385 90.565 148.475 ;
        RECT 90.775 148.615 94.675 149.295 ;
        RECT 90.775 148.385 91.705 148.615 ;
        RECT 94.915 148.485 98.585 149.295 ;
        RECT 98.595 148.485 99.965 149.295 ;
        RECT 99.985 148.425 100.415 149.210 ;
        RECT 100.435 148.615 104.335 149.295 ;
        RECT 100.435 148.385 101.365 148.615 ;
        RECT 105.035 148.515 106.405 149.295 ;
        RECT 106.415 148.615 113.725 149.295 ;
        RECT 114.695 148.615 122.005 149.295 ;
        RECT 109.930 148.395 110.840 148.615 ;
        RECT 112.375 148.385 113.725 148.615 ;
        RECT 118.210 148.395 119.120 148.615 ;
        RECT 120.655 148.385 122.005 148.615 ;
        RECT 122.055 148.515 123.425 149.295 ;
        RECT 123.635 148.475 125.565 149.295 ;
        RECT 123.635 148.385 124.585 148.475 ;
        RECT 125.745 148.425 126.175 149.210 ;
        RECT 126.195 148.485 128.945 149.295 ;
        RECT 129.610 148.385 133.085 149.295 ;
        RECT 133.095 148.485 134.465 149.295 ;
        RECT 134.475 148.615 141.785 149.295 ;
        RECT 141.835 148.615 145.045 149.295 ;
        RECT 145.200 149.265 145.370 149.485 ;
        RECT 145.650 149.315 145.820 149.505 ;
        RECT 148.415 149.295 148.585 149.485 ;
        RECT 149.795 149.295 149.965 149.485 ;
        RECT 152.095 149.295 152.265 149.485 ;
        RECT 153.935 149.315 154.105 149.505 ;
        RECT 154.395 149.315 154.565 149.505 ;
        RECT 156.695 149.295 156.865 149.505 ;
        RECT 147.330 149.265 148.265 149.295 ;
        RECT 145.200 149.065 148.265 149.265 ;
        RECT 137.990 148.395 138.900 148.615 ;
        RECT 140.435 148.385 141.785 148.615 ;
        RECT 143.910 148.385 145.045 148.615 ;
        RECT 145.055 148.585 148.265 149.065 ;
        RECT 145.055 148.385 145.985 148.585 ;
        RECT 147.315 148.385 148.265 148.585 ;
        RECT 148.275 148.515 149.645 149.295 ;
        RECT 149.655 148.485 151.485 149.295 ;
        RECT 151.505 148.425 151.935 149.210 ;
        RECT 151.955 148.485 155.625 149.295 ;
        RECT 155.635 148.485 157.005 149.295 ;
      LAYER nwell ;
        RECT 22.500 145.265 157.200 148.095 ;
      LAYER pwell ;
        RECT 22.695 144.065 24.065 144.875 ;
        RECT 24.075 144.065 26.825 144.875 ;
        RECT 27.615 144.745 29.575 144.975 ;
        RECT 27.125 144.065 29.575 144.745 ;
        RECT 29.595 144.065 33.265 144.875 ;
        RECT 33.275 144.065 35.105 144.975 ;
        RECT 35.585 144.150 36.015 144.935 ;
        RECT 37.050 144.745 37.970 144.975 ;
        RECT 37.050 144.065 40.515 144.745 ;
        RECT 40.635 144.065 44.305 144.875 ;
        RECT 44.315 144.065 51.005 144.975 ;
        RECT 52.155 144.065 53.505 144.975 ;
        RECT 53.515 144.065 55.345 144.875 ;
        RECT 55.355 144.775 56.305 144.975 ;
        RECT 57.635 144.775 58.565 144.975 ;
        RECT 55.355 144.295 58.565 144.775 ;
        RECT 55.355 144.095 58.420 144.295 ;
        RECT 55.355 144.065 56.290 144.095 ;
        RECT 22.835 143.855 23.005 144.065 ;
        RECT 24.215 143.855 24.385 144.065 ;
        RECT 27.125 144.045 27.145 144.065 ;
        RECT 26.975 143.875 27.145 144.045 ;
        RECT 29.735 143.875 29.905 144.065 ;
        RECT 34.790 144.045 34.960 144.065 ;
        RECT 34.790 143.875 34.965 144.045 ;
        RECT 35.250 144.010 35.370 144.015 ;
        RECT 35.250 143.905 35.425 144.010 ;
        RECT 36.185 143.910 36.345 144.020 ;
        RECT 35.265 143.900 35.425 143.905 ;
        RECT 34.795 143.855 34.965 143.875 ;
        RECT 38.930 143.855 39.100 144.045 ;
        RECT 22.695 143.045 24.065 143.855 ;
        RECT 24.075 143.175 31.385 143.855 ;
        RECT 27.590 142.955 28.500 143.175 ;
        RECT 30.035 142.945 31.385 143.175 ;
        RECT 31.530 143.175 34.995 143.855 ;
        RECT 31.530 142.945 32.450 143.175 ;
        RECT 36.325 142.945 39.245 143.855 ;
        RECT 39.400 143.825 39.570 144.045 ;
        RECT 40.315 143.875 40.485 144.065 ;
        RECT 40.775 143.875 40.945 144.065 ;
        RECT 43.075 143.855 43.245 144.045 ;
        RECT 43.535 143.855 43.705 144.045 ;
        RECT 44.455 143.875 44.625 144.065 ;
        RECT 44.915 143.875 45.085 144.045 ;
        RECT 44.935 143.855 45.085 143.875 ;
        RECT 48.135 143.855 48.305 144.045 ;
        RECT 49.055 143.855 49.225 144.045 ;
        RECT 51.365 143.910 51.525 144.020 ;
        RECT 51.815 143.855 51.985 144.045 ;
        RECT 52.270 143.875 52.440 144.065 ;
        RECT 53.655 143.875 53.825 144.065 ;
        RECT 58.250 143.875 58.420 144.095 ;
        RECT 58.575 144.065 61.325 144.875 ;
        RECT 61.345 144.150 61.775 144.935 ;
        RECT 61.795 144.065 63.625 144.875 ;
        RECT 63.635 144.745 66.460 144.975 ;
        RECT 67.410 144.745 68.330 144.975 ;
        RECT 72.010 144.745 72.930 144.975 ;
        RECT 63.635 144.065 67.165 144.745 ;
        RECT 67.410 144.065 70.875 144.745 ;
        RECT 72.010 144.065 75.475 144.745 ;
        RECT 75.595 144.065 84.700 144.745 ;
        RECT 84.795 144.065 86.625 144.875 ;
        RECT 87.105 144.150 87.535 144.935 ;
        RECT 91.990 144.745 92.900 144.965 ;
        RECT 94.435 144.745 95.785 144.975 ;
        RECT 96.885 144.745 97.815 144.975 ;
        RECT 98.620 144.745 99.965 144.975 ;
        RECT 88.475 144.065 95.785 144.745 ;
        RECT 95.980 144.065 97.815 144.745 ;
        RECT 98.135 144.065 99.965 144.745 ;
        RECT 99.975 144.065 103.645 144.875 ;
        RECT 103.655 144.065 107.545 144.975 ;
        RECT 108.715 144.745 109.645 144.975 ;
        RECT 108.715 144.065 112.615 144.745 ;
        RECT 112.865 144.150 113.295 144.935 ;
        RECT 113.315 144.065 115.145 144.875 ;
        RECT 118.355 144.745 119.285 144.975 ;
        RECT 115.385 144.065 119.285 144.745 ;
        RECT 119.295 144.065 121.125 144.875 ;
        RECT 125.110 144.745 126.020 144.965 ;
        RECT 127.555 144.745 128.905 144.975 ;
        RECT 121.595 144.065 128.905 144.745 ;
        RECT 129.875 144.065 133.085 144.975 ;
        RECT 133.095 144.065 136.305 144.975 ;
        RECT 137.650 144.775 138.605 144.975 ;
        RECT 136.325 144.095 138.605 144.775 ;
        RECT 138.625 144.150 139.055 144.935 ;
        RECT 58.715 143.875 58.885 144.065 ;
        RECT 59.175 143.855 59.345 144.045 ;
        RECT 61.475 143.855 61.645 144.045 ;
        RECT 61.935 143.875 62.105 144.065 ;
        RECT 66.965 144.045 67.165 144.065 ;
        RECT 64.235 143.855 64.405 144.045 ;
        RECT 64.695 143.855 64.865 144.045 ;
        RECT 66.995 143.875 67.165 144.045 ;
        RECT 67.910 143.905 68.030 144.015 ;
        RECT 68.375 143.875 68.545 144.045 ;
        RECT 70.675 143.875 70.845 144.065 ;
        RECT 71.145 143.910 71.305 144.020 ;
        RECT 68.385 143.855 68.545 143.875 ;
        RECT 72.515 143.855 72.685 144.045 ;
        RECT 74.825 143.900 74.985 144.010 ;
        RECT 75.275 143.875 75.445 144.065 ;
        RECT 75.735 143.855 75.905 144.065 ;
        RECT 84.935 143.875 85.105 144.065 ;
        RECT 86.315 143.855 86.485 144.045 ;
        RECT 86.775 144.015 86.945 144.045 ;
        RECT 86.770 143.905 86.945 144.015 ;
        RECT 87.705 143.910 87.865 144.020 ;
        RECT 86.775 143.855 86.945 143.905 ;
        RECT 88.615 143.875 88.785 144.065 ;
        RECT 95.980 144.045 96.145 144.065 ;
        RECT 91.830 143.855 92.000 144.045 ;
        RECT 93.220 143.855 93.390 144.045 ;
        RECT 93.670 143.905 93.790 144.015 ;
        RECT 95.975 143.875 96.145 144.045 ;
        RECT 41.060 143.825 42.005 143.855 ;
        RECT 39.255 143.145 42.005 143.825 ;
        RECT 41.060 142.945 42.005 143.145 ;
        RECT 42.015 143.075 43.385 143.855 ;
        RECT 43.395 143.045 44.765 143.855 ;
        RECT 44.935 143.035 46.865 143.855 ;
        RECT 47.075 143.075 48.445 143.855 ;
        RECT 45.915 142.945 46.865 143.035 ;
        RECT 48.465 142.985 48.895 143.770 ;
        RECT 48.915 143.045 51.665 143.855 ;
        RECT 51.675 143.175 58.985 143.855 ;
        RECT 55.190 142.955 56.100 143.175 ;
        RECT 57.635 142.945 58.985 143.175 ;
        RECT 59.035 143.045 60.405 143.855 ;
        RECT 60.425 142.945 61.775 143.855 ;
        RECT 61.805 142.945 64.535 143.855 ;
        RECT 64.555 142.945 67.765 143.855 ;
        RECT 68.385 142.945 72.040 143.855 ;
        RECT 72.375 143.045 74.205 143.855 ;
        RECT 74.225 142.985 74.655 143.770 ;
        RECT 75.705 143.175 79.170 143.855 ;
        RECT 78.250 142.945 79.170 143.175 ;
        RECT 79.315 143.175 86.625 143.855 ;
        RECT 79.315 142.945 80.665 143.175 ;
        RECT 82.200 142.955 83.110 143.175 ;
        RECT 86.635 142.945 89.845 143.855 ;
        RECT 89.870 143.175 92.145 143.855 ;
        RECT 89.870 142.945 91.240 143.175 ;
        RECT 92.155 142.945 93.505 143.855 ;
        RECT 93.995 143.825 94.940 143.855 ;
        RECT 96.430 143.825 96.600 144.045 ;
        RECT 96.900 143.825 97.070 144.045 ;
        RECT 98.275 143.875 98.445 144.065 ;
        RECT 100.115 143.875 100.285 144.065 ;
        RECT 100.575 143.855 100.745 144.045 ;
        RECT 103.800 143.875 103.970 144.065 ;
        RECT 104.710 143.855 104.880 144.045 ;
        RECT 105.175 143.855 105.345 144.045 ;
        RECT 107.945 143.910 108.105 144.020 ;
        RECT 108.855 143.855 109.025 144.045 ;
        RECT 109.130 143.875 109.300 144.065 ;
        RECT 109.315 143.855 109.485 144.045 ;
        RECT 111.150 143.905 111.270 144.015 ;
        RECT 113.455 143.875 113.625 144.065 ;
        RECT 113.455 143.855 113.605 143.875 ;
        RECT 113.915 143.855 114.085 144.045 ;
        RECT 115.295 143.855 115.465 144.045 ;
        RECT 116.675 143.855 116.845 144.045 ;
        RECT 118.700 143.875 118.870 144.065 ;
        RECT 119.435 143.875 119.605 144.065 ;
        RECT 119.895 143.875 120.065 144.045 ;
        RECT 119.895 143.855 120.045 143.875 ;
        RECT 120.355 143.855 120.525 144.045 ;
        RECT 121.270 143.905 121.390 144.015 ;
        RECT 121.735 143.875 121.905 144.065 ;
        RECT 126.335 143.875 126.505 144.045 ;
        RECT 126.355 143.855 126.505 143.875 ;
        RECT 128.635 143.855 128.805 144.045 ;
        RECT 129.105 143.910 129.265 144.020 ;
        RECT 130.015 143.875 130.185 144.065 ;
        RECT 130.470 143.905 130.590 144.015 ;
        RECT 130.935 143.855 131.105 144.045 ;
        RECT 133.235 143.875 133.405 144.065 ;
        RECT 136.450 144.045 136.620 144.095 ;
        RECT 137.650 144.065 138.605 144.095 ;
        RECT 139.085 144.065 140.435 144.975 ;
        RECT 140.475 144.065 141.825 144.975 ;
        RECT 141.845 144.065 143.195 144.975 ;
        RECT 143.215 144.065 146.885 144.875 ;
        RECT 146.895 144.065 148.265 144.875 ;
        RECT 151.790 144.745 152.700 144.965 ;
        RECT 154.235 144.745 155.585 144.975 ;
        RECT 148.275 144.065 155.585 144.745 ;
        RECT 155.635 144.065 157.005 144.875 ;
        RECT 134.165 143.900 134.325 144.010 ;
        RECT 135.995 143.855 136.165 144.045 ;
        RECT 136.450 143.875 136.625 144.045 ;
        RECT 139.210 143.905 139.330 144.015 ;
        RECT 140.135 143.875 140.305 144.065 ;
        RECT 140.590 144.045 140.760 144.065 ;
        RECT 140.590 143.875 140.770 144.045 ;
        RECT 136.455 143.855 136.625 143.875 ;
        RECT 140.600 143.855 140.770 143.875 ;
        RECT 141.055 143.855 141.225 144.045 ;
        RECT 142.895 143.875 143.065 144.065 ;
        RECT 143.355 144.015 143.525 144.065 ;
        RECT 143.350 143.905 143.525 144.015 ;
        RECT 143.355 143.875 143.525 143.905 ;
        RECT 143.815 143.875 143.985 144.045 ;
        RECT 143.820 143.855 143.985 143.875 ;
        RECT 146.115 143.855 146.285 144.045 ;
        RECT 147.035 143.875 147.205 144.065 ;
        RECT 148.415 143.855 148.585 144.065 ;
        RECT 149.795 143.855 149.965 144.045 ;
        RECT 152.095 143.855 152.265 144.045 ;
        RECT 156.695 143.855 156.865 144.065 ;
        RECT 99.030 143.825 99.965 143.855 ;
        RECT 93.995 143.145 96.745 143.825 ;
        RECT 96.900 143.625 99.965 143.825 ;
        RECT 96.755 143.145 99.965 143.625 ;
        RECT 93.995 142.945 94.940 143.145 ;
        RECT 96.755 142.945 97.685 143.145 ;
        RECT 99.015 142.945 99.965 143.145 ;
        RECT 99.985 142.985 100.415 143.770 ;
        RECT 100.435 143.045 101.805 143.855 ;
        RECT 102.815 143.625 105.020 143.855 ;
        RECT 101.875 142.945 105.020 143.625 ;
        RECT 105.035 143.175 107.775 143.855 ;
        RECT 107.795 143.075 109.165 143.855 ;
        RECT 109.175 143.045 111.005 143.855 ;
        RECT 111.675 143.035 113.605 143.855 ;
        RECT 113.775 143.045 115.145 143.855 ;
        RECT 115.155 143.075 116.525 143.855 ;
        RECT 116.535 143.045 117.905 143.855 ;
        RECT 118.115 143.035 120.045 143.855 ;
        RECT 120.215 143.045 125.725 143.855 ;
        RECT 111.675 142.945 112.625 143.035 ;
        RECT 118.115 142.945 119.065 143.035 ;
        RECT 125.745 142.985 126.175 143.770 ;
        RECT 126.355 143.035 128.285 143.855 ;
        RECT 128.495 143.045 130.325 143.855 ;
        RECT 127.335 142.945 128.285 143.035 ;
        RECT 130.795 142.945 134.005 143.855 ;
        RECT 134.945 142.945 136.295 143.855 ;
        RECT 136.315 143.045 139.065 143.855 ;
        RECT 139.535 142.945 140.885 143.855 ;
        RECT 140.915 143.175 143.205 143.855 ;
        RECT 143.820 143.175 145.655 143.855 ;
        RECT 145.975 143.175 148.265 143.855 ;
        RECT 142.285 142.945 143.205 143.175 ;
        RECT 144.725 142.945 145.655 143.175 ;
        RECT 147.345 142.945 148.265 143.175 ;
        RECT 148.275 143.075 149.645 143.855 ;
        RECT 149.655 143.045 151.485 143.855 ;
        RECT 151.505 142.985 151.935 143.770 ;
        RECT 151.955 143.045 155.625 143.855 ;
        RECT 155.635 143.045 157.005 143.855 ;
      LAYER nwell ;
        RECT 22.500 139.825 157.200 142.655 ;
      LAYER pwell ;
        RECT 22.695 138.625 24.065 139.435 ;
        RECT 24.075 138.625 26.825 139.435 ;
        RECT 26.835 138.625 29.585 139.535 ;
        RECT 29.595 138.625 32.345 139.435 ;
        RECT 32.815 139.305 33.735 139.535 ;
        RECT 32.815 138.625 35.105 139.305 ;
        RECT 35.585 138.710 36.015 139.495 ;
        RECT 36.130 139.305 37.050 139.535 ;
        RECT 39.715 139.335 40.645 139.535 ;
        RECT 41.975 139.335 42.925 139.535 ;
        RECT 36.130 138.625 39.595 139.305 ;
        RECT 39.715 138.855 42.925 139.335 ;
        RECT 46.450 139.305 47.360 139.525 ;
        RECT 48.895 139.305 50.245 139.535 ;
        RECT 52.100 139.335 53.045 139.535 ;
        RECT 39.860 138.655 42.925 138.855 ;
        RECT 22.835 138.415 23.005 138.625 ;
        RECT 24.215 138.435 24.385 138.625 ;
        RECT 25.135 138.415 25.305 138.605 ;
        RECT 26.975 138.435 27.145 138.625 ;
        RECT 29.735 138.435 29.905 138.625 ;
        RECT 32.495 138.575 32.665 138.605 ;
        RECT 32.490 138.465 32.665 138.575 ;
        RECT 32.495 138.415 32.665 138.465 ;
        RECT 34.795 138.435 34.965 138.625 ;
        RECT 35.250 138.570 35.370 138.575 ;
        RECT 35.250 138.465 35.425 138.570 ;
        RECT 35.265 138.460 35.425 138.465 ;
        RECT 39.395 138.435 39.565 138.625 ;
        RECT 39.860 138.435 40.030 138.655 ;
        RECT 41.990 138.625 42.925 138.655 ;
        RECT 42.935 138.625 50.245 139.305 ;
        RECT 50.295 138.655 53.045 139.335 ;
        RECT 43.075 138.415 43.245 138.625 ;
        RECT 43.535 138.415 43.705 138.605 ;
        RECT 47.215 138.415 47.385 138.605 ;
        RECT 49.055 138.415 49.225 138.605 ;
        RECT 50.440 138.435 50.610 138.655 ;
        RECT 52.100 138.625 53.045 138.655 ;
        RECT 53.975 138.625 55.345 139.405 ;
        RECT 55.355 138.625 58.105 139.435 ;
        RECT 59.355 139.305 61.315 139.535 ;
        RECT 58.865 138.625 61.315 139.305 ;
        RECT 61.345 138.710 61.775 139.495 ;
        RECT 65.310 139.305 66.220 139.525 ;
        RECT 67.755 139.305 69.105 139.535 ;
        RECT 61.795 138.625 69.105 139.305 ;
        RECT 69.480 138.625 73.135 139.535 ;
        RECT 73.305 138.625 74.655 139.535 ;
        RECT 74.685 138.625 76.035 139.535 ;
        RECT 78.710 139.305 79.630 139.535 ;
        RECT 76.165 138.625 79.630 139.305 ;
        RECT 79.775 139.305 81.125 139.535 ;
        RECT 82.660 139.305 83.570 139.525 ;
        RECT 79.775 138.625 87.085 139.305 ;
        RECT 87.105 138.710 87.535 139.495 ;
        RECT 87.570 139.305 88.940 139.535 ;
        RECT 87.570 138.625 89.845 139.305 ;
        RECT 89.855 138.625 91.225 139.405 ;
        RECT 91.780 138.625 100.885 139.305 ;
        RECT 100.975 138.625 103.185 139.535 ;
        RECT 103.195 138.625 105.405 139.535 ;
        RECT 105.980 139.305 107.325 139.535 ;
        RECT 105.495 138.625 107.325 139.305 ;
        RECT 107.335 139.305 108.265 139.535 ;
        RECT 107.335 138.625 111.235 139.305 ;
        RECT 111.475 138.625 112.845 139.435 ;
        RECT 112.865 138.710 113.295 139.495 ;
        RECT 117.750 139.305 118.660 139.525 ;
        RECT 120.195 139.305 121.545 139.535 ;
        RECT 125.570 139.305 126.480 139.525 ;
        RECT 128.015 139.305 129.365 139.535 ;
        RECT 114.235 138.625 121.545 139.305 ;
        RECT 122.055 138.625 129.365 139.305 ;
        RECT 129.415 138.625 131.245 139.435 ;
        RECT 131.730 138.625 135.385 139.535 ;
        RECT 135.595 139.445 136.545 139.535 ;
        RECT 135.595 138.625 137.525 139.445 ;
        RECT 138.625 138.710 139.055 139.495 ;
        RECT 139.085 138.625 140.435 139.535 ;
        RECT 140.455 139.305 141.590 139.535 ;
        RECT 144.725 139.305 145.655 139.535 ;
        RECT 140.455 138.625 143.665 139.305 ;
        RECT 143.820 138.625 145.655 139.305 ;
        RECT 145.975 138.625 147.325 139.535 ;
        RECT 150.870 139.305 151.780 139.525 ;
        RECT 153.315 139.305 154.665 139.535 ;
        RECT 147.355 138.625 154.665 139.305 ;
        RECT 155.635 138.625 157.005 139.435 ;
        RECT 52.730 138.465 52.850 138.575 ;
        RECT 53.205 138.470 53.365 138.580 ;
        RECT 54.115 138.415 54.285 138.605 ;
        RECT 54.580 138.415 54.750 138.605 ;
        RECT 55.035 138.435 55.205 138.625 ;
        RECT 55.495 138.435 55.665 138.625 ;
        RECT 58.865 138.605 58.885 138.625 ;
        RECT 57.790 138.465 57.910 138.575 ;
        RECT 58.250 138.415 58.420 138.605 ;
        RECT 58.715 138.435 58.885 138.605 ;
        RECT 59.635 138.435 59.805 138.605 ;
        RECT 59.640 138.415 59.805 138.435 ;
        RECT 61.935 138.415 62.105 138.625 ;
        RECT 72.975 138.605 73.135 138.625 ;
        RECT 65.615 138.415 65.785 138.605 ;
        RECT 67.915 138.415 68.085 138.605 ;
        RECT 69.755 138.415 69.925 138.605 ;
        RECT 72.975 138.415 73.145 138.605 ;
        RECT 74.355 138.435 74.525 138.625 ;
        RECT 75.735 138.435 75.905 138.625 ;
        RECT 76.195 138.435 76.365 138.625 ;
        RECT 81.715 138.415 81.885 138.605 ;
        RECT 82.175 138.415 82.345 138.605 ;
        RECT 84.930 138.465 85.050 138.575 ;
        RECT 85.395 138.415 85.565 138.605 ;
        RECT 86.775 138.435 86.945 138.625 ;
        RECT 87.235 138.415 87.405 138.605 ;
        RECT 89.075 138.415 89.245 138.605 ;
        RECT 89.530 138.435 89.700 138.625 ;
        RECT 90.915 138.435 91.085 138.625 ;
        RECT 91.370 138.465 91.490 138.575 ;
        RECT 98.275 138.435 98.445 138.605 ;
        RECT 98.275 138.415 98.425 138.435 ;
        RECT 98.735 138.415 98.905 138.605 ;
        RECT 100.575 138.415 100.745 138.625 ;
        RECT 102.870 138.435 103.040 138.625 ;
        RECT 103.340 138.435 103.510 138.625 ;
        RECT 103.795 138.415 103.965 138.605 ;
        RECT 104.265 138.460 104.425 138.570 ;
        RECT 105.175 138.415 105.345 138.605 ;
        RECT 105.635 138.435 105.805 138.625 ;
        RECT 107.750 138.435 107.920 138.625 ;
        RECT 111.615 138.435 111.785 138.625 ;
        RECT 113.465 138.470 113.625 138.580 ;
        RECT 114.375 138.435 114.545 138.625 ;
        RECT 114.830 138.465 114.950 138.575 ;
        RECT 114.375 138.415 114.525 138.435 ;
        RECT 115.570 138.415 115.740 138.605 ;
        RECT 119.435 138.415 119.605 138.605 ;
        RECT 122.195 138.575 122.365 138.625 ;
        RECT 121.730 138.465 121.850 138.575 ;
        RECT 122.190 138.465 122.365 138.575 ;
        RECT 122.195 138.435 122.365 138.465 ;
        RECT 123.575 138.415 123.745 138.605 ;
        RECT 124.035 138.415 124.205 138.605 ;
        RECT 126.610 138.415 126.780 138.605 ;
        RECT 129.555 138.435 129.725 138.625 ;
        RECT 130.485 138.460 130.645 138.570 ;
        RECT 131.390 138.465 131.510 138.575 ;
        RECT 22.695 137.605 24.065 138.415 ;
        RECT 24.995 137.735 32.305 138.415 ;
        RECT 28.510 137.515 29.420 137.735 ;
        RECT 30.955 137.505 32.305 137.735 ;
        RECT 32.355 137.505 35.105 138.415 ;
        RECT 36.075 137.735 43.385 138.415 ;
        RECT 36.075 137.505 37.425 137.735 ;
        RECT 38.960 137.515 39.870 137.735 ;
        RECT 43.395 137.605 47.065 138.415 ;
        RECT 47.075 137.605 48.445 138.415 ;
        RECT 48.465 137.545 48.895 138.330 ;
        RECT 48.915 137.605 52.585 138.415 ;
        RECT 53.055 137.635 54.425 138.415 ;
        RECT 54.440 138.185 56.645 138.415 ;
        RECT 54.440 137.505 57.585 138.185 ;
        RECT 58.135 137.505 59.485 138.415 ;
        RECT 59.640 137.735 61.475 138.415 ;
        RECT 61.905 137.735 65.370 138.415 ;
        RECT 65.475 137.735 67.765 138.415 ;
        RECT 60.545 137.505 61.475 137.735 ;
        RECT 64.450 137.505 65.370 137.735 ;
        RECT 66.845 137.505 67.765 137.735 ;
        RECT 67.775 137.605 69.605 138.415 ;
        RECT 69.615 137.505 72.825 138.415 ;
        RECT 72.835 137.605 74.205 138.415 ;
        RECT 74.225 137.545 74.655 138.330 ;
        RECT 74.715 137.735 82.025 138.415 ;
        RECT 74.715 137.505 76.065 137.735 ;
        RECT 77.600 137.515 78.510 137.735 ;
        RECT 82.035 137.605 84.785 138.415 ;
        RECT 85.255 137.735 87.085 138.415 ;
        RECT 85.740 137.505 87.085 137.735 ;
        RECT 87.095 137.605 88.925 138.415 ;
        RECT 88.935 137.735 96.245 138.415 ;
        RECT 92.450 137.515 93.360 137.735 ;
        RECT 94.895 137.505 96.245 137.735 ;
        RECT 96.495 137.595 98.425 138.415 ;
        RECT 98.595 137.605 99.965 138.415 ;
        RECT 96.495 137.505 97.445 137.595 ;
        RECT 99.985 137.545 100.415 138.330 ;
        RECT 100.435 137.735 102.265 138.415 ;
        RECT 100.920 137.505 102.265 137.735 ;
        RECT 102.275 137.735 104.105 138.415 ;
        RECT 105.035 137.735 112.345 138.415 ;
        RECT 102.275 137.505 103.620 137.735 ;
        RECT 108.550 137.515 109.460 137.735 ;
        RECT 110.995 137.505 112.345 137.735 ;
        RECT 112.595 137.595 114.525 138.415 ;
        RECT 115.155 137.735 119.055 138.415 ;
        RECT 112.595 137.505 113.545 137.595 ;
        RECT 115.155 137.505 116.085 137.735 ;
        RECT 119.295 137.605 122.045 138.415 ;
        RECT 122.515 137.635 123.885 138.415 ;
        RECT 123.895 137.605 125.725 138.415 ;
        RECT 125.745 137.545 126.175 138.330 ;
        RECT 126.195 137.735 130.095 138.415 ;
        RECT 131.255 138.385 132.205 138.415 ;
        RECT 134.610 138.385 134.780 138.605 ;
        RECT 135.070 138.385 135.240 138.625 ;
        RECT 137.375 138.605 137.525 138.625 ;
        RECT 140.135 138.605 140.305 138.625 ;
        RECT 137.375 138.415 137.545 138.605 ;
        RECT 137.845 138.470 138.005 138.580 ;
        RECT 140.130 138.435 140.305 138.605 ;
        RECT 140.130 138.415 140.300 138.435 ;
        RECT 136.270 138.385 137.225 138.415 ;
        RECT 126.195 137.505 127.125 137.735 ;
        RECT 131.255 137.705 134.925 138.385 ;
        RECT 134.945 137.705 137.225 138.385 ;
        RECT 131.255 137.505 132.205 137.705 ;
        RECT 136.270 137.505 137.225 137.705 ;
        RECT 137.235 137.605 139.985 138.415 ;
        RECT 140.015 137.505 141.365 138.415 ;
        RECT 141.520 138.385 141.690 138.605 ;
        RECT 143.355 138.435 143.525 138.625 ;
        RECT 143.820 138.605 143.985 138.625 ;
        RECT 143.815 138.435 143.985 138.605 ;
        RECT 145.655 138.415 145.825 138.605 ;
        RECT 146.110 138.465 146.230 138.575 ;
        RECT 146.575 138.415 146.745 138.605 ;
        RECT 147.040 138.435 147.210 138.625 ;
        RECT 147.495 138.435 147.665 138.625 ;
        RECT 147.955 138.415 148.125 138.605 ;
        RECT 149.335 138.415 149.505 138.605 ;
        RECT 151.170 138.465 151.290 138.575 ;
        RECT 152.095 138.415 152.265 138.605 ;
        RECT 154.865 138.470 155.025 138.580 ;
        RECT 156.695 138.415 156.865 138.625 ;
        RECT 143.650 138.385 144.585 138.415 ;
        RECT 141.520 138.185 144.585 138.385 ;
        RECT 141.375 137.705 144.585 138.185 ;
        RECT 141.375 137.505 142.305 137.705 ;
        RECT 143.635 137.505 144.585 137.705 ;
        RECT 144.605 137.505 145.955 138.415 ;
        RECT 146.435 137.635 147.805 138.415 ;
        RECT 147.815 137.635 149.185 138.415 ;
        RECT 149.195 137.605 151.025 138.415 ;
        RECT 151.505 137.545 151.935 138.330 ;
        RECT 151.955 137.605 155.625 138.415 ;
        RECT 155.635 137.605 157.005 138.415 ;
      LAYER nwell ;
        RECT 22.500 134.385 157.200 137.215 ;
      LAYER pwell ;
        RECT 22.695 133.185 24.065 133.995 ;
        RECT 24.075 133.185 27.745 133.995 ;
        RECT 28.675 133.185 32.150 134.095 ;
        RECT 33.135 133.865 35.095 134.095 ;
        RECT 32.645 133.185 35.095 133.865 ;
        RECT 35.585 133.270 36.015 134.055 ;
        RECT 36.345 133.865 37.275 134.095 ;
        RECT 36.345 133.185 38.180 133.865 ;
        RECT 38.335 133.185 42.005 133.995 ;
        RECT 45.990 133.865 46.900 134.085 ;
        RECT 48.435 133.865 49.785 134.095 ;
        RECT 53.350 133.865 54.260 134.085 ;
        RECT 55.795 133.865 57.145 134.095 ;
        RECT 42.475 133.185 49.785 133.865 ;
        RECT 49.835 133.185 57.145 133.865 ;
        RECT 57.290 133.865 58.210 134.095 ;
        RECT 57.290 133.185 60.755 133.865 ;
        RECT 61.345 133.270 61.775 134.055 ;
        RECT 61.880 133.185 70.985 133.865 ;
        RECT 70.995 133.185 72.365 133.995 ;
        RECT 72.515 133.185 75.125 134.095 ;
        RECT 75.135 133.185 78.345 134.095 ;
        RECT 78.355 133.185 79.725 133.995 ;
        RECT 79.735 133.185 82.475 133.865 ;
        RECT 82.495 133.185 86.165 133.995 ;
        RECT 87.105 133.270 87.535 134.055 ;
        RECT 87.555 133.185 91.225 133.995 ;
        RECT 91.235 133.185 92.605 133.965 ;
        RECT 93.075 133.865 94.005 134.095 ;
        RECT 93.075 133.185 96.975 133.865 ;
        RECT 97.215 133.185 100.325 134.095 ;
        RECT 100.530 133.865 101.450 134.095 ;
        RECT 110.755 134.005 111.705 134.095 ;
        RECT 100.530 133.185 103.995 133.865 ;
        RECT 104.115 133.185 106.865 133.995 ;
        RECT 107.335 133.185 108.705 133.965 ;
        RECT 108.715 133.185 110.545 133.995 ;
        RECT 110.755 133.185 112.685 134.005 ;
        RECT 112.865 133.270 113.295 134.055 ;
        RECT 123.000 133.865 124.345 134.095 ;
        RECT 113.315 133.185 122.420 133.865 ;
        RECT 122.515 133.185 124.345 133.865 ;
        RECT 124.355 133.185 125.705 134.095 ;
        RECT 125.735 133.185 131.245 133.995 ;
        RECT 131.255 133.185 136.765 133.995 ;
        RECT 136.775 133.185 138.605 133.995 ;
        RECT 138.625 133.270 139.055 134.055 ;
        RECT 139.995 133.185 141.825 133.865 ;
        RECT 141.835 133.185 145.505 133.995 ;
        RECT 145.515 133.185 146.885 133.995 ;
        RECT 146.935 133.865 148.285 134.095 ;
        RECT 149.820 133.865 150.730 134.085 ;
        RECT 146.935 133.185 154.245 133.865 ;
        RECT 154.255 133.185 155.625 133.995 ;
        RECT 155.635 133.185 157.005 133.995 ;
        RECT 22.835 132.975 23.005 133.185 ;
        RECT 24.215 133.135 24.385 133.185 ;
        RECT 28.820 133.165 28.990 133.185 ;
        RECT 32.645 133.165 32.665 133.185 ;
        RECT 38.015 133.165 38.180 133.185 ;
        RECT 24.210 133.025 24.385 133.135 ;
        RECT 24.215 132.995 24.385 133.025 ;
        RECT 24.680 132.975 24.850 133.165 ;
        RECT 27.905 133.030 28.065 133.140 ;
        RECT 28.350 133.025 28.470 133.135 ;
        RECT 28.815 132.995 28.990 133.165 ;
        RECT 32.495 132.995 32.665 133.165 ;
        RECT 35.250 133.025 35.370 133.135 ;
        RECT 28.815 132.975 28.985 132.995 ;
        RECT 35.715 132.975 35.885 133.165 ;
        RECT 36.175 132.975 36.345 133.165 ;
        RECT 38.015 132.995 38.185 133.165 ;
        RECT 38.475 132.995 38.645 133.185 ;
        RECT 42.150 133.025 42.270 133.135 ;
        RECT 42.615 132.995 42.785 133.185 ;
        RECT 46.755 132.975 46.925 133.165 ;
        RECT 48.135 132.975 48.305 133.165 ;
        RECT 49.055 132.975 49.225 133.165 ;
        RECT 49.975 132.995 50.145 133.185 ;
        RECT 51.815 132.995 51.985 133.165 ;
        RECT 51.835 132.975 51.985 132.995 ;
        RECT 54.120 132.975 54.290 133.165 ;
        RECT 58.265 133.020 58.425 133.130 ;
        RECT 59.175 132.975 59.345 133.165 ;
        RECT 60.555 132.995 60.725 133.185 ;
        RECT 61.010 133.025 61.130 133.135 ;
        RECT 64.695 132.975 64.865 133.165 ;
        RECT 70.675 132.995 70.845 133.185 ;
        RECT 71.135 132.995 71.305 133.185 ;
        RECT 74.810 133.165 74.980 133.185 ;
        RECT 72.055 132.975 72.225 133.165 ;
        RECT 73.435 132.975 73.605 133.165 ;
        RECT 73.890 133.025 74.010 133.135 ;
        RECT 74.810 132.995 74.985 133.165 ;
        RECT 78.035 132.995 78.205 133.185 ;
        RECT 78.495 132.995 78.665 133.185 ;
        RECT 79.875 132.995 80.045 133.185 ;
        RECT 74.815 132.975 74.985 132.995 ;
        RECT 82.175 132.975 82.345 133.165 ;
        RECT 82.635 132.995 82.805 133.185 ;
        RECT 86.325 133.030 86.485 133.140 ;
        RECT 87.695 132.995 87.865 133.185 ;
        RECT 89.810 132.975 89.980 133.165 ;
        RECT 92.295 132.995 92.465 133.185 ;
        RECT 92.750 133.025 92.870 133.135 ;
        RECT 93.490 132.995 93.660 133.185 ;
        RECT 93.670 133.025 93.790 133.135 ;
        RECT 94.410 132.975 94.580 133.165 ;
        RECT 98.270 133.025 98.390 133.135 ;
        RECT 98.730 132.975 98.900 133.165 ;
        RECT 100.115 132.995 100.285 133.185 ;
        RECT 103.795 132.995 103.965 133.185 ;
        RECT 104.255 132.995 104.425 133.185 ;
        RECT 107.010 133.025 107.130 133.135 ;
        RECT 107.475 132.975 107.645 133.185 ;
        RECT 107.935 132.975 108.105 133.165 ;
        RECT 108.855 132.995 109.025 133.185 ;
        RECT 112.535 133.165 112.685 133.185 ;
        RECT 112.535 132.995 112.705 133.165 ;
        RECT 113.455 132.995 113.625 133.185 ;
        RECT 122.195 132.975 122.365 133.165 ;
        RECT 122.655 133.135 122.825 133.185 ;
        RECT 122.650 133.025 122.825 133.135 ;
        RECT 122.655 132.995 122.825 133.025 ;
        RECT 123.115 132.975 123.285 133.165 ;
        RECT 125.420 132.995 125.590 133.185 ;
        RECT 125.875 132.995 126.045 133.185 ;
        RECT 126.335 132.975 126.505 133.165 ;
        RECT 130.010 133.025 130.130 133.135 ;
        RECT 130.470 132.975 130.640 133.165 ;
        RECT 131.395 132.995 131.565 133.185 ;
        RECT 135.070 132.975 135.240 133.165 ;
        RECT 136.915 132.995 137.085 133.185 ;
        RECT 137.835 132.975 138.005 133.165 ;
        RECT 138.295 132.995 138.465 133.165 ;
        RECT 139.225 133.030 139.385 133.140 ;
        RECT 140.135 132.995 140.305 133.185 ;
        RECT 138.315 132.975 138.465 132.995 ;
        RECT 140.595 132.975 140.765 133.165 ;
        RECT 141.975 132.995 142.145 133.185 ;
        RECT 141.980 132.975 142.145 132.995 ;
        RECT 144.275 132.975 144.445 133.165 ;
        RECT 145.655 132.995 145.825 133.185 ;
        RECT 147.035 132.975 147.205 133.165 ;
        RECT 148.415 132.975 148.585 133.165 ;
        RECT 151.170 133.025 151.290 133.135 ;
        RECT 152.095 132.975 152.265 133.165 ;
        RECT 153.935 132.995 154.105 133.185 ;
        RECT 154.395 132.995 154.565 133.185 ;
        RECT 156.695 132.975 156.865 133.185 ;
        RECT 22.695 132.165 24.065 132.975 ;
        RECT 24.535 132.065 28.010 132.975 ;
        RECT 28.785 132.295 32.250 132.975 ;
        RECT 31.330 132.065 32.250 132.295 ;
        RECT 32.450 132.295 35.915 132.975 ;
        RECT 36.035 132.295 43.345 132.975 ;
        RECT 32.450 132.065 33.370 132.295 ;
        RECT 39.550 132.075 40.460 132.295 ;
        RECT 41.995 132.065 43.345 132.295 ;
        RECT 43.490 132.295 46.955 132.975 ;
        RECT 43.490 132.065 44.410 132.295 ;
        RECT 47.085 132.065 48.435 132.975 ;
        RECT 48.465 132.105 48.895 132.890 ;
        RECT 48.915 132.295 51.655 132.975 ;
        RECT 51.835 132.155 53.765 132.975 ;
        RECT 52.815 132.065 53.765 132.155 ;
        RECT 53.975 132.065 57.865 132.975 ;
        RECT 59.035 132.295 61.325 132.975 ;
        RECT 60.405 132.065 61.325 132.295 ;
        RECT 61.430 132.295 64.895 132.975 ;
        RECT 65.055 132.295 72.365 132.975 ;
        RECT 61.430 132.065 62.350 132.295 ;
        RECT 65.055 132.065 66.405 132.295 ;
        RECT 67.940 132.075 68.850 132.295 ;
        RECT 72.375 132.195 73.745 132.975 ;
        RECT 74.225 132.105 74.655 132.890 ;
        RECT 74.675 132.295 81.985 132.975 ;
        RECT 82.035 132.295 89.345 132.975 ;
        RECT 78.190 132.075 79.100 132.295 ;
        RECT 80.635 132.065 81.985 132.295 ;
        RECT 85.550 132.075 86.460 132.295 ;
        RECT 87.995 132.065 89.345 132.295 ;
        RECT 89.395 132.295 93.295 132.975 ;
        RECT 93.995 132.295 97.895 132.975 ;
        RECT 89.395 132.065 90.325 132.295 ;
        RECT 93.995 132.065 94.925 132.295 ;
        RECT 98.615 132.065 99.965 132.975 ;
        RECT 99.985 132.105 100.415 132.890 ;
        RECT 100.475 132.295 107.785 132.975 ;
        RECT 107.795 132.295 115.105 132.975 ;
        RECT 100.475 132.065 101.825 132.295 ;
        RECT 103.360 132.075 104.270 132.295 ;
        RECT 111.310 132.075 112.220 132.295 ;
        RECT 113.755 132.065 115.105 132.295 ;
        RECT 115.195 132.065 122.475 132.975 ;
        RECT 122.975 132.295 125.715 132.975 ;
        RECT 125.745 132.105 126.175 132.890 ;
        RECT 126.305 132.295 129.770 132.975 ;
        RECT 128.850 132.065 129.770 132.295 ;
        RECT 130.355 132.065 131.705 132.975 ;
        RECT 131.715 132.295 135.385 132.975 ;
        RECT 134.460 132.065 135.385 132.295 ;
        RECT 135.425 132.065 138.145 132.975 ;
        RECT 138.315 132.155 140.245 132.975 ;
        RECT 140.455 132.165 141.825 132.975 ;
        RECT 141.980 132.295 143.815 132.975 ;
        RECT 139.295 132.065 140.245 132.155 ;
        RECT 142.885 132.065 143.815 132.295 ;
        RECT 144.135 132.165 146.885 132.975 ;
        RECT 146.895 132.195 148.265 132.975 ;
        RECT 148.275 132.165 151.025 132.975 ;
        RECT 151.505 132.105 151.935 132.890 ;
        RECT 151.955 132.165 155.625 132.975 ;
        RECT 155.635 132.165 157.005 132.975 ;
      LAYER nwell ;
        RECT 22.500 128.945 157.200 131.775 ;
      LAYER pwell ;
        RECT 22.695 127.745 24.065 128.555 ;
        RECT 24.630 128.425 25.550 128.655 ;
        RECT 31.730 128.425 32.640 128.645 ;
        RECT 34.175 128.425 35.525 128.655 ;
        RECT 24.630 127.745 28.095 128.425 ;
        RECT 28.215 127.745 35.525 128.425 ;
        RECT 35.585 127.830 36.015 128.615 ;
        RECT 36.230 127.745 39.705 128.655 ;
        RECT 49.390 128.425 50.760 128.655 ;
        RECT 40.175 127.745 49.280 128.425 ;
        RECT 49.390 127.745 51.665 128.425 ;
        RECT 51.675 127.745 53.965 128.655 ;
        RECT 57.490 128.425 58.400 128.645 ;
        RECT 59.935 128.425 61.285 128.655 ;
        RECT 53.975 127.745 61.285 128.425 ;
        RECT 61.345 127.830 61.775 128.615 ;
        RECT 62.265 127.745 64.995 128.655 ;
        RECT 68.530 128.425 69.440 128.645 ;
        RECT 70.975 128.425 72.325 128.655 ;
        RECT 65.015 127.745 72.325 128.425 ;
        RECT 72.470 128.425 73.390 128.655 ;
        RECT 72.470 127.745 75.935 128.425 ;
        RECT 76.055 127.745 77.885 128.555 ;
        RECT 78.360 127.975 81.505 128.655 ;
        RECT 85.935 128.565 86.885 128.655 ;
        RECT 78.360 127.745 80.565 127.975 ;
        RECT 81.575 127.745 83.405 128.555 ;
        RECT 83.415 127.745 84.785 128.525 ;
        RECT 84.955 127.745 86.885 128.565 ;
        RECT 87.105 127.830 87.535 128.615 ;
        RECT 92.375 128.565 93.325 128.655 ;
        RECT 87.555 127.745 90.295 128.425 ;
        RECT 91.395 127.745 93.325 128.565 ;
        RECT 93.575 127.745 100.855 128.655 ;
        RECT 100.895 127.745 106.405 128.555 ;
        RECT 106.415 127.745 107.785 128.555 ;
        RECT 107.795 128.425 108.725 128.655 ;
        RECT 107.795 127.745 111.695 128.425 ;
        RECT 112.865 127.830 113.295 128.615 ;
        RECT 113.315 127.745 115.145 128.555 ;
        RECT 117.955 128.425 119.305 128.655 ;
        RECT 120.840 128.425 121.750 128.645 ;
        RECT 115.165 127.745 117.905 128.425 ;
        RECT 117.955 127.745 125.265 128.425 ;
        RECT 126.195 127.745 129.305 128.655 ;
        RECT 129.415 127.745 131.245 128.555 ;
        RECT 131.350 128.425 132.270 128.655 ;
        RECT 134.935 128.455 135.880 128.655 ;
        RECT 131.350 127.745 134.815 128.425 ;
        RECT 134.935 127.775 137.685 128.455 ;
        RECT 138.625 127.830 139.055 128.615 ;
        RECT 134.935 127.745 135.880 127.775 ;
        RECT 22.835 127.535 23.005 127.745 ;
        RECT 24.215 127.695 24.385 127.725 ;
        RECT 24.210 127.585 24.385 127.695 ;
        RECT 24.215 127.535 24.385 127.585 ;
        RECT 27.895 127.555 28.065 127.745 ;
        RECT 28.355 127.555 28.525 127.745 ;
        RECT 31.575 127.535 31.745 127.725 ;
        RECT 36.170 127.535 36.340 127.725 ;
        RECT 36.635 127.535 36.805 127.725 ;
        RECT 39.390 127.555 39.560 127.745 ;
        RECT 39.850 127.585 39.970 127.695 ;
        RECT 40.315 127.555 40.485 127.745 ;
        RECT 43.535 127.535 43.705 127.725 ;
        RECT 44.005 127.580 44.165 127.690 ;
        RECT 44.915 127.535 45.085 127.725 ;
        RECT 49.050 127.585 49.170 127.695 ;
        RECT 51.350 127.555 51.520 127.745 ;
        RECT 51.815 127.555 51.985 127.745 ;
        RECT 52.735 127.535 52.905 127.725 ;
        RECT 53.190 127.585 53.310 127.695 ;
        RECT 53.655 127.535 53.825 127.725 ;
        RECT 54.115 127.555 54.285 127.745 ;
        RECT 61.010 127.585 61.130 127.695 ;
        RECT 61.475 127.535 61.645 127.725 ;
        RECT 61.930 127.585 62.050 127.695 ;
        RECT 62.395 127.555 62.565 127.745 ;
        RECT 65.155 127.555 65.325 127.745 ;
        RECT 66.075 127.535 66.245 127.725 ;
        RECT 66.530 127.585 66.650 127.695 ;
        RECT 66.995 127.535 67.165 127.725 ;
        RECT 71.595 127.535 71.765 127.725 ;
        RECT 72.055 127.535 72.225 127.725 ;
        RECT 73.445 127.580 73.605 127.690 ;
        RECT 74.815 127.535 74.985 127.725 ;
        RECT 75.735 127.555 75.905 127.745 ;
        RECT 76.195 127.555 76.365 127.745 ;
        RECT 78.030 127.585 78.150 127.695 ;
        RECT 78.500 127.555 78.670 127.745 ;
        RECT 81.715 127.555 81.885 127.745 ;
        RECT 82.820 127.535 82.990 127.725 ;
        RECT 83.555 127.535 83.725 127.725 ;
        RECT 84.475 127.555 84.645 127.745 ;
        RECT 84.955 127.725 85.105 127.745 ;
        RECT 84.935 127.555 85.105 127.725 ;
        RECT 87.245 127.580 87.405 127.690 ;
        RECT 87.695 127.555 87.865 127.745 ;
        RECT 91.395 127.725 91.545 127.745 ;
        RECT 88.155 127.535 88.325 127.725 ;
        RECT 89.535 127.535 89.705 127.725 ;
        RECT 90.465 127.590 90.625 127.700 ;
        RECT 91.375 127.555 91.545 127.725 ;
        RECT 96.895 127.535 97.065 127.725 ;
        RECT 99.650 127.585 99.770 127.695 ;
        RECT 100.575 127.535 100.745 127.745 ;
        RECT 101.035 127.555 101.205 127.745 ;
        RECT 104.255 127.555 104.425 127.725 ;
        RECT 104.255 127.535 104.405 127.555 ;
        RECT 104.715 127.535 104.885 127.725 ;
        RECT 106.555 127.555 106.725 127.745 ;
        RECT 108.210 127.555 108.380 127.745 ;
        RECT 112.085 127.590 112.245 127.700 ;
        RECT 113.455 127.555 113.625 127.745 ;
        RECT 117.595 127.725 117.765 127.745 ;
        RECT 114.375 127.535 114.545 127.725 ;
        RECT 114.835 127.535 115.005 127.725 ;
        RECT 117.595 127.555 117.770 127.725 ;
        RECT 117.600 127.535 117.770 127.555 ;
        RECT 119.435 127.535 119.605 127.725 ;
        RECT 122.195 127.555 122.365 127.725 ;
        RECT 122.290 127.535 122.365 127.555 ;
        RECT 124.495 127.535 124.665 127.725 ;
        RECT 124.955 127.555 125.125 127.745 ;
        RECT 125.425 127.590 125.585 127.700 ;
        RECT 129.095 127.535 129.265 127.745 ;
        RECT 129.555 127.535 129.725 127.745 ;
        RECT 132.315 127.535 132.485 127.725 ;
        RECT 134.615 127.555 134.785 127.745 ;
        RECT 137.370 127.725 137.540 127.775 ;
        RECT 139.085 127.745 140.435 128.655 ;
        RECT 140.455 127.745 141.805 128.655 ;
        RECT 141.855 127.745 143.205 128.655 ;
        RECT 144.585 128.425 145.505 128.655 ;
        RECT 146.565 128.425 147.495 128.655 ;
        RECT 143.215 127.745 145.505 128.425 ;
        RECT 145.660 127.745 147.495 128.425 ;
        RECT 147.855 128.425 149.205 128.655 ;
        RECT 150.740 128.425 151.650 128.645 ;
        RECT 147.855 127.745 155.165 128.425 ;
        RECT 155.635 127.745 157.005 128.555 ;
        RECT 135.995 127.535 136.165 127.725 ;
        RECT 137.370 127.555 137.545 127.725 ;
        RECT 137.845 127.590 138.005 127.700 ;
        RECT 140.135 127.555 140.305 127.745 ;
        RECT 141.050 127.585 141.170 127.695 ;
        RECT 141.520 127.555 141.690 127.745 ;
        RECT 141.970 127.555 142.140 127.745 ;
        RECT 143.355 127.555 143.525 127.745 ;
        RECT 145.660 127.725 145.825 127.745 ;
        RECT 137.375 127.535 137.545 127.555 ;
        RECT 144.275 127.535 144.445 127.725 ;
        RECT 22.695 126.725 24.065 127.535 ;
        RECT 24.075 126.855 31.385 127.535 ;
        RECT 27.590 126.635 28.500 126.855 ;
        RECT 30.035 126.625 31.385 126.855 ;
        RECT 31.435 126.725 32.805 127.535 ;
        RECT 33.010 126.625 36.485 127.535 ;
        RECT 36.605 126.855 40.070 127.535 ;
        RECT 39.150 126.625 40.070 126.855 ;
        RECT 40.270 126.855 43.735 127.535 ;
        RECT 44.885 126.855 48.350 127.535 ;
        RECT 40.270 126.625 41.190 126.855 ;
        RECT 47.430 126.625 48.350 126.855 ;
        RECT 48.465 126.665 48.895 127.450 ;
        RECT 49.470 126.855 52.935 127.535 ;
        RECT 53.515 126.855 60.825 127.535 ;
        RECT 49.470 126.625 50.390 126.855 ;
        RECT 57.030 126.635 57.940 126.855 ;
        RECT 59.475 126.625 60.825 126.855 ;
        RECT 61.345 126.625 64.075 127.535 ;
        RECT 64.095 126.855 66.385 127.535 ;
        RECT 64.095 126.625 65.015 126.855 ;
        RECT 66.865 126.625 69.595 127.535 ;
        RECT 69.615 126.855 71.905 127.535 ;
        RECT 69.615 126.625 70.535 126.855 ;
        RECT 71.925 126.625 73.275 127.535 ;
        RECT 74.225 126.665 74.655 127.450 ;
        RECT 74.785 126.855 78.250 127.535 ;
        RECT 79.505 126.855 83.405 127.535 ;
        RECT 77.330 126.625 78.250 126.855 ;
        RECT 82.475 126.625 83.405 126.855 ;
        RECT 83.415 126.725 87.085 127.535 ;
        RECT 88.015 126.755 89.385 127.535 ;
        RECT 89.395 126.855 96.705 127.535 ;
        RECT 92.910 126.635 93.820 126.855 ;
        RECT 95.355 126.625 96.705 126.855 ;
        RECT 96.755 126.725 99.505 127.535 ;
        RECT 99.985 126.665 100.415 127.450 ;
        RECT 100.435 126.725 102.265 127.535 ;
        RECT 102.475 126.715 104.405 127.535 ;
        RECT 104.575 126.725 107.325 127.535 ;
        RECT 102.475 126.625 103.425 126.715 ;
        RECT 107.375 126.625 114.655 127.535 ;
        RECT 114.695 126.725 117.445 127.535 ;
        RECT 117.455 126.625 119.285 127.535 ;
        RECT 119.295 126.855 122.035 127.535 ;
        RECT 122.290 126.855 124.125 127.535 ;
        RECT 122.775 126.625 124.125 126.855 ;
        RECT 124.355 126.725 125.725 127.535 ;
        RECT 125.745 126.665 126.175 127.450 ;
        RECT 126.195 126.625 129.405 127.535 ;
        RECT 129.415 126.855 132.155 127.535 ;
        RECT 132.175 126.625 135.845 127.535 ;
        RECT 135.865 126.625 137.215 127.535 ;
        RECT 137.235 126.725 140.905 127.535 ;
        RECT 141.375 126.855 144.585 127.535 ;
        RECT 144.740 127.505 144.910 127.725 ;
        RECT 145.655 127.555 145.825 127.725 ;
        RECT 147.955 127.535 148.125 127.725 ;
        RECT 150.255 127.535 150.425 127.725 ;
        RECT 153.015 127.535 153.185 127.725 ;
        RECT 153.475 127.535 153.645 127.725 ;
        RECT 154.855 127.555 155.025 127.745 ;
        RECT 155.310 127.585 155.430 127.695 ;
        RECT 156.695 127.535 156.865 127.745 ;
        RECT 146.870 127.505 147.805 127.535 ;
        RECT 144.740 127.305 147.805 127.505 ;
        RECT 141.375 126.625 142.510 126.855 ;
        RECT 144.595 126.825 147.805 127.305 ;
        RECT 147.815 126.855 150.105 127.535 ;
        RECT 144.595 126.625 145.525 126.825 ;
        RECT 146.855 126.625 147.805 126.825 ;
        RECT 149.185 126.625 150.105 126.855 ;
        RECT 150.115 126.755 151.485 127.535 ;
        RECT 151.505 126.665 151.935 127.450 ;
        RECT 151.955 126.755 153.325 127.535 ;
        RECT 153.335 126.725 155.165 127.535 ;
        RECT 155.635 126.725 157.005 127.535 ;
      LAYER nwell ;
        RECT 22.500 123.505 157.200 126.335 ;
      LAYER pwell ;
        RECT 22.695 122.305 24.065 123.115 ;
        RECT 26.045 122.985 26.975 123.215 ;
        RECT 29.950 122.985 30.870 123.215 ;
        RECT 25.140 122.305 26.975 122.985 ;
        RECT 27.405 122.305 30.870 122.985 ;
        RECT 31.070 122.985 31.990 123.215 ;
        RECT 31.070 122.305 34.535 122.985 ;
        RECT 35.585 122.390 36.015 123.175 ;
        RECT 36.075 122.985 37.425 123.215 ;
        RECT 38.960 122.985 39.870 123.205 ;
        RECT 43.895 122.985 45.245 123.215 ;
        RECT 46.780 122.985 47.690 123.205 ;
        RECT 52.265 122.985 53.195 123.215 ;
        RECT 36.075 122.305 43.385 122.985 ;
        RECT 43.895 122.305 51.205 122.985 ;
        RECT 51.360 122.305 53.195 122.985 ;
        RECT 53.515 122.305 55.330 123.215 ;
        RECT 55.355 122.305 57.185 123.215 ;
        RECT 57.195 122.305 60.865 123.115 ;
        RECT 61.345 122.390 61.775 123.175 ;
        RECT 61.795 122.305 64.545 123.115 ;
        RECT 65.015 122.305 74.120 122.985 ;
        RECT 74.215 122.305 76.045 123.115 ;
        RECT 79.570 122.985 80.480 123.205 ;
        RECT 82.015 122.985 83.365 123.215 ;
        RECT 76.055 122.305 83.365 122.985 ;
        RECT 83.615 123.125 84.565 123.215 ;
        RECT 83.615 122.305 85.545 123.125 ;
        RECT 85.715 122.305 87.085 123.115 ;
        RECT 87.105 122.390 87.535 123.175 ;
        RECT 88.695 123.125 89.645 123.215 ;
        RECT 94.215 123.125 95.165 123.215 ;
        RECT 87.715 122.305 89.645 123.125 ;
        RECT 89.855 122.305 91.685 123.115 ;
        RECT 91.695 122.305 93.065 123.085 ;
        RECT 93.235 122.305 95.165 123.125 ;
        RECT 95.375 122.305 97.205 123.115 ;
        RECT 97.215 122.305 98.585 123.085 ;
        RECT 102.110 122.985 103.020 123.205 ;
        RECT 104.555 122.985 105.905 123.215 ;
        RECT 98.595 122.305 105.905 122.985 ;
        RECT 105.955 122.305 107.325 123.085 ;
        RECT 107.335 122.985 108.265 123.215 ;
        RECT 107.335 122.305 111.235 122.985 ;
        RECT 111.475 122.305 112.845 123.115 ;
        RECT 112.865 122.390 113.295 123.175 ;
        RECT 113.315 122.305 116.985 123.115 ;
        RECT 130.630 122.985 131.540 123.205 ;
        RECT 133.075 122.985 134.425 123.215 ;
        RECT 117.915 122.305 127.020 122.985 ;
        RECT 127.115 122.305 134.425 122.985 ;
        RECT 134.570 122.985 135.490 123.215 ;
        RECT 134.570 122.305 138.035 122.985 ;
        RECT 138.625 122.390 139.055 123.175 ;
        RECT 139.075 122.985 139.995 123.215 ;
        RECT 142.755 123.015 143.700 123.215 ;
        RECT 145.035 123.015 145.965 123.215 ;
        RECT 139.075 122.305 142.660 122.985 ;
        RECT 142.755 122.535 145.965 123.015 ;
        RECT 142.755 122.335 145.825 122.535 ;
        RECT 142.755 122.305 143.700 122.335 ;
        RECT 22.835 122.095 23.005 122.305 ;
        RECT 25.140 122.285 25.305 122.305 ;
        RECT 24.225 122.150 24.385 122.260 ;
        RECT 25.135 122.115 25.305 122.285 ;
        RECT 27.435 122.115 27.605 122.305 ;
        RECT 31.115 122.095 31.285 122.285 ;
        RECT 34.335 122.115 34.505 122.305 ;
        RECT 34.790 122.260 34.960 122.285 ;
        RECT 34.790 122.150 34.965 122.260 ;
        RECT 34.790 122.095 34.960 122.150 ;
        RECT 36.635 122.095 36.805 122.285 ;
        RECT 22.695 121.285 24.065 122.095 ;
        RECT 24.115 121.415 31.425 122.095 ;
        RECT 24.115 121.185 25.465 121.415 ;
        RECT 27.000 121.195 27.910 121.415 ;
        RECT 31.630 121.185 35.105 122.095 ;
        RECT 35.115 121.415 36.945 122.095 ;
        RECT 37.100 122.065 37.270 122.285 ;
        RECT 39.855 122.095 40.025 122.285 ;
        RECT 43.075 122.115 43.245 122.305 ;
        RECT 43.530 122.145 43.650 122.255 ;
        RECT 46.480 122.095 46.650 122.285 ;
        RECT 47.215 122.095 47.385 122.285 ;
        RECT 49.050 122.145 49.170 122.255 ;
        RECT 49.515 122.095 49.685 122.285 ;
        RECT 50.895 122.115 51.065 122.305 ;
        RECT 51.360 122.285 51.525 122.305 ;
        RECT 51.355 122.115 51.525 122.285 ;
        RECT 55.035 122.115 55.205 122.305 ;
        RECT 55.500 122.115 55.670 122.305 ;
        RECT 57.335 122.115 57.505 122.305 ;
        RECT 60.095 122.095 60.265 122.285 ;
        RECT 60.555 122.095 60.725 122.285 ;
        RECT 61.010 122.145 61.130 122.255 ;
        RECT 61.935 122.115 62.105 122.305 ;
        RECT 63.775 122.095 63.945 122.285 ;
        RECT 64.690 122.145 64.810 122.255 ;
        RECT 65.155 122.115 65.325 122.305 ;
        RECT 66.530 122.145 66.650 122.255 ;
        RECT 73.895 122.095 74.065 122.285 ;
        RECT 74.355 122.115 74.525 122.305 ;
        RECT 76.195 122.115 76.365 122.305 ;
        RECT 85.395 122.285 85.545 122.305 ;
        RECT 78.035 122.095 78.205 122.285 ;
        RECT 78.495 122.095 78.665 122.285 ;
        RECT 82.175 122.095 82.345 122.285 ;
        RECT 82.635 122.095 82.805 122.285 ;
        RECT 85.395 122.115 85.565 122.285 ;
        RECT 85.855 122.115 86.025 122.305 ;
        RECT 87.715 122.285 87.865 122.305 ;
        RECT 87.695 122.115 87.865 122.285 ;
        RECT 89.995 122.095 90.165 122.305 ;
        RECT 92.755 122.115 92.925 122.305 ;
        RECT 93.235 122.285 93.385 122.305 ;
        RECT 93.215 122.115 93.385 122.285 ;
        RECT 95.515 122.115 95.685 122.305 ;
        RECT 97.355 122.115 97.525 122.305 ;
        RECT 97.815 122.095 97.985 122.285 ;
        RECT 98.735 122.115 98.905 122.305 ;
        RECT 99.650 122.145 99.770 122.255 ;
        RECT 100.850 122.095 101.020 122.285 ;
        RECT 104.710 122.145 104.830 122.255 ;
        RECT 105.175 122.095 105.345 122.285 ;
        RECT 107.015 122.115 107.185 122.305 ;
        RECT 107.750 122.115 107.920 122.305 ;
        RECT 111.615 122.115 111.785 122.305 ;
        RECT 112.535 122.095 112.705 122.285 ;
        RECT 113.455 122.115 113.625 122.305 ;
        RECT 117.145 122.150 117.305 122.260 ;
        RECT 118.055 122.115 118.225 122.305 ;
        RECT 120.815 122.095 120.985 122.285 ;
        RECT 121.285 122.140 121.445 122.250 ;
        RECT 124.955 122.095 125.125 122.285 ;
        RECT 125.410 122.145 125.530 122.255 ;
        RECT 126.335 122.095 126.505 122.285 ;
        RECT 127.255 122.115 127.425 122.305 ;
        RECT 133.700 122.095 133.870 122.285 ;
        RECT 136.905 122.095 137.075 122.285 ;
        RECT 137.835 122.115 138.005 122.305 ;
        RECT 138.290 122.145 138.410 122.255 ;
        RECT 139.220 122.115 139.390 122.305 ;
        RECT 140.140 122.095 140.310 122.285 ;
        RECT 143.355 122.115 143.525 122.285 ;
        RECT 143.810 122.145 143.930 122.255 ;
        RECT 145.655 122.115 145.825 122.335 ;
        RECT 145.985 122.305 147.335 123.215 ;
        RECT 147.855 122.985 149.205 123.215 ;
        RECT 150.740 122.985 151.650 123.205 ;
        RECT 147.855 122.305 155.165 122.985 ;
        RECT 155.635 122.305 157.005 123.115 ;
        RECT 146.115 122.115 146.285 122.305 ;
        RECT 147.490 122.145 147.610 122.255 ;
        RECT 143.355 122.095 143.505 122.115 ;
        RECT 151.175 122.095 151.345 122.285 ;
        RECT 152.095 122.095 152.265 122.285 ;
        RECT 154.855 122.115 155.025 122.305 ;
        RECT 155.310 122.145 155.430 122.255 ;
        RECT 156.695 122.095 156.865 122.305 ;
        RECT 38.760 122.065 39.705 122.095 ;
        RECT 36.955 121.385 39.705 122.065 ;
        RECT 38.760 121.185 39.705 121.385 ;
        RECT 39.795 121.185 42.795 122.095 ;
        RECT 43.165 121.415 47.065 122.095 ;
        RECT 46.135 121.185 47.065 121.415 ;
        RECT 47.075 121.285 48.445 122.095 ;
        RECT 48.465 121.225 48.895 122.010 ;
        RECT 49.375 121.415 56.685 122.095 ;
        RECT 52.890 121.195 53.800 121.415 ;
        RECT 55.335 121.185 56.685 121.415 ;
        RECT 56.830 121.415 60.295 122.095 ;
        RECT 56.830 121.185 57.750 121.415 ;
        RECT 60.515 121.185 63.625 122.095 ;
        RECT 63.635 121.285 66.385 122.095 ;
        RECT 66.895 121.415 74.205 122.095 ;
        RECT 66.895 121.185 68.245 121.415 ;
        RECT 69.780 121.195 70.690 121.415 ;
        RECT 74.225 121.225 74.655 122.010 ;
        RECT 74.770 121.415 78.235 122.095 ;
        RECT 74.770 121.185 75.690 121.415 ;
        RECT 78.365 121.185 81.095 122.095 ;
        RECT 81.115 121.315 82.485 122.095 ;
        RECT 82.495 121.415 89.805 122.095 ;
        RECT 89.855 121.415 97.585 122.095 ;
        RECT 86.010 121.195 86.920 121.415 ;
        RECT 88.455 121.185 89.805 121.415 ;
        RECT 93.370 121.195 94.280 121.415 ;
        RECT 95.815 121.185 97.585 121.415 ;
        RECT 97.675 121.285 99.505 122.095 ;
        RECT 99.985 121.225 100.415 122.010 ;
        RECT 100.435 121.415 104.335 122.095 ;
        RECT 105.035 121.415 112.345 122.095 ;
        RECT 100.435 121.185 101.365 121.415 ;
        RECT 108.550 121.195 109.460 121.415 ;
        RECT 110.995 121.185 112.345 121.415 ;
        RECT 112.395 121.285 113.765 122.095 ;
        RECT 113.815 121.415 121.125 122.095 ;
        RECT 113.815 121.185 115.165 121.415 ;
        RECT 116.700 121.195 117.610 121.415 ;
        RECT 122.055 121.185 125.265 122.095 ;
        RECT 125.745 121.225 126.175 122.010 ;
        RECT 126.195 121.415 133.505 122.095 ;
        RECT 129.710 121.195 130.620 121.415 ;
        RECT 132.155 121.185 133.505 121.415 ;
        RECT 133.555 121.185 136.475 122.095 ;
        RECT 136.775 121.185 139.985 122.095 ;
        RECT 139.995 121.185 141.345 122.095 ;
        RECT 141.575 121.275 143.505 122.095 ;
        RECT 144.175 121.415 151.485 122.095 ;
        RECT 141.575 121.185 142.525 121.275 ;
        RECT 144.175 121.185 145.525 121.415 ;
        RECT 147.060 121.195 147.970 121.415 ;
        RECT 151.505 121.225 151.935 122.010 ;
        RECT 151.955 121.285 155.625 122.095 ;
        RECT 155.635 121.285 157.005 122.095 ;
      LAYER nwell ;
        RECT 22.500 118.065 157.200 120.895 ;
      LAYER pwell ;
        RECT 22.695 116.865 24.065 117.675 ;
        RECT 24.075 116.865 25.905 117.675 ;
        RECT 26.965 117.545 27.895 117.775 ;
        RECT 26.060 116.865 27.895 117.545 ;
        RECT 28.255 117.545 29.605 117.775 ;
        RECT 31.140 117.545 32.050 117.765 ;
        RECT 28.255 116.865 35.565 117.545 ;
        RECT 35.585 116.950 36.015 117.735 ;
        RECT 36.130 117.545 37.050 117.775 ;
        RECT 36.130 116.865 39.595 117.545 ;
        RECT 39.715 116.865 43.190 117.775 ;
        RECT 43.490 117.545 44.410 117.775 ;
        RECT 43.490 116.865 46.955 117.545 ;
        RECT 48.190 116.865 51.665 117.775 ;
        RECT 54.330 117.545 55.250 117.775 ;
        RECT 51.785 116.865 55.250 117.545 ;
        RECT 55.665 117.545 56.595 117.775 ;
        RECT 57.655 117.575 58.600 117.775 ;
        RECT 55.665 116.865 57.500 117.545 ;
        RECT 57.655 116.895 60.405 117.575 ;
        RECT 61.345 116.950 61.775 117.735 ;
        RECT 57.655 116.865 58.600 116.895 ;
        RECT 22.835 116.655 23.005 116.865 ;
        RECT 24.215 116.675 24.385 116.865 ;
        RECT 26.060 116.845 26.225 116.865 ;
        RECT 25.135 116.675 25.305 116.845 ;
        RECT 26.055 116.675 26.225 116.845 ;
        RECT 25.140 116.655 25.305 116.675 ;
        RECT 30.650 116.655 30.820 116.845 ;
        RECT 31.115 116.655 31.285 116.845 ;
        RECT 22.695 115.845 24.065 116.655 ;
        RECT 25.140 115.975 26.975 116.655 ;
        RECT 26.045 115.745 26.975 115.975 ;
        RECT 27.490 115.745 30.965 116.655 ;
        RECT 31.085 115.975 34.550 116.655 ;
        RECT 34.800 116.625 34.970 116.845 ;
        RECT 35.255 116.675 35.425 116.865 ;
        RECT 37.555 116.655 37.725 116.845 ;
        RECT 39.395 116.675 39.565 116.865 ;
        RECT 39.860 116.675 40.030 116.865 ;
        RECT 46.755 116.675 46.925 116.865 ;
        RECT 47.225 116.710 47.385 116.820 ;
        RECT 48.130 116.655 48.300 116.845 ;
        RECT 49.055 116.655 49.225 116.845 ;
        RECT 51.350 116.675 51.520 116.865 ;
        RECT 51.815 116.675 51.985 116.865 ;
        RECT 57.335 116.845 57.500 116.865 ;
        RECT 57.335 116.675 57.505 116.845 ;
        RECT 57.795 116.655 57.965 116.845 ;
        RECT 58.255 116.655 58.425 116.845 ;
        RECT 59.635 116.655 59.805 116.845 ;
        RECT 60.090 116.675 60.260 116.895 ;
        RECT 61.795 116.865 65.465 117.675 ;
        RECT 65.935 117.545 66.865 117.775 ;
        RECT 65.935 116.865 69.835 117.545 ;
        RECT 70.085 116.865 71.435 117.775 ;
        RECT 71.455 116.865 76.965 117.675 ;
        RECT 78.805 117.545 79.725 117.775 ;
        RECT 81.775 117.685 82.725 117.775 ;
        RECT 77.435 116.865 79.725 117.545 ;
        RECT 79.735 116.865 81.105 117.645 ;
        RECT 81.775 116.865 83.705 117.685 ;
        RECT 83.875 116.865 85.245 117.645 ;
        RECT 85.255 116.865 87.085 117.675 ;
        RECT 87.105 116.950 87.535 117.735 ;
        RECT 87.555 117.545 88.485 117.775 ;
        RECT 92.615 117.545 93.545 117.775 ;
        RECT 87.555 116.865 91.455 117.545 ;
        RECT 92.615 116.865 96.515 117.545 ;
        RECT 96.755 116.865 98.585 117.675 ;
        RECT 99.055 117.545 99.985 117.775 ;
        RECT 110.755 117.685 111.705 117.775 ;
        RECT 99.055 116.865 102.955 117.545 ;
        RECT 103.195 116.865 108.705 117.675 ;
        RECT 108.715 116.865 110.545 117.675 ;
        RECT 110.755 116.865 112.685 117.685 ;
        RECT 112.865 116.950 113.295 117.735 ;
        RECT 113.315 116.865 115.925 117.775 ;
        RECT 118.730 117.545 119.650 117.775 ;
        RECT 116.185 116.865 119.650 117.545 ;
        RECT 119.765 116.865 122.495 117.775 ;
        RECT 122.515 116.865 123.885 117.645 ;
        RECT 124.355 116.865 127.565 117.775 ;
        RECT 127.575 116.865 128.945 117.675 ;
        RECT 129.050 117.545 129.970 117.775 ;
        RECT 129.050 116.865 132.515 117.545 ;
        RECT 132.635 116.865 135.845 117.775 ;
        RECT 136.165 117.545 137.095 117.775 ;
        RECT 136.165 116.865 138.000 117.545 ;
        RECT 138.625 116.950 139.055 117.735 ;
        RECT 139.075 116.865 140.425 117.775 ;
        RECT 140.455 117.575 141.385 117.775 ;
        RECT 142.715 117.575 143.665 117.775 ;
        RECT 140.455 117.095 143.665 117.575 ;
        RECT 140.600 116.895 143.665 117.095 ;
        RECT 60.565 116.710 60.725 116.820 ;
        RECT 61.475 116.655 61.645 116.845 ;
        RECT 61.935 116.675 62.105 116.865 ;
        RECT 64.690 116.705 64.810 116.815 ;
        RECT 36.460 116.625 37.405 116.655 ;
        RECT 33.630 115.745 34.550 115.975 ;
        RECT 34.655 115.945 37.405 116.625 ;
        RECT 37.415 115.975 44.725 116.655 ;
        RECT 36.460 115.745 37.405 115.945 ;
        RECT 40.930 115.755 41.840 115.975 ;
        RECT 43.375 115.745 44.725 115.975 ;
        RECT 44.970 115.745 48.445 116.655 ;
        RECT 48.465 115.785 48.895 116.570 ;
        RECT 48.915 115.845 50.745 116.655 ;
        RECT 50.795 115.975 58.105 116.655 ;
        RECT 50.795 115.745 52.145 115.975 ;
        RECT 53.680 115.755 54.590 115.975 ;
        RECT 58.125 115.745 59.475 116.655 ;
        RECT 59.495 115.845 61.325 116.655 ;
        RECT 61.335 115.745 64.545 116.655 ;
        RECT 65.155 116.625 65.325 116.845 ;
        RECT 65.610 116.705 65.730 116.815 ;
        RECT 66.350 116.675 66.520 116.865 ;
        RECT 68.370 116.705 68.490 116.815 ;
        RECT 71.135 116.675 71.305 116.865 ;
        RECT 71.595 116.675 71.765 116.865 ;
        RECT 72.240 116.655 72.410 116.845 ;
        RECT 73.895 116.655 74.065 116.845 ;
        RECT 74.810 116.705 74.930 116.815 ;
        RECT 75.275 116.655 75.445 116.845 ;
        RECT 77.110 116.705 77.230 116.815 ;
        RECT 77.575 116.675 77.745 116.865 ;
        RECT 80.795 116.675 80.965 116.865 ;
        RECT 83.555 116.845 83.705 116.865 ;
        RECT 81.250 116.705 81.370 116.815 ;
        RECT 82.645 116.700 82.805 116.810 ;
        RECT 83.555 116.655 83.725 116.845 ;
        RECT 84.935 116.675 85.105 116.865 ;
        RECT 85.395 116.675 85.565 116.865 ;
        RECT 87.970 116.675 88.140 116.865 ;
        RECT 91.845 116.710 92.005 116.820 ;
        RECT 92.760 116.655 92.930 116.845 ;
        RECT 93.030 116.675 93.200 116.865 ;
        RECT 94.135 116.655 94.305 116.845 ;
        RECT 95.970 116.705 96.090 116.815 ;
        RECT 96.435 116.655 96.605 116.845 ;
        RECT 96.895 116.675 97.065 116.865 ;
        RECT 97.815 116.675 97.985 116.845 ;
        RECT 98.730 116.705 98.850 116.815 ;
        RECT 99.470 116.675 99.640 116.865 ;
        RECT 103.335 116.675 103.505 116.865 ;
        RECT 97.835 116.655 97.985 116.675 ;
        RECT 107.475 116.655 107.645 116.845 ;
        RECT 107.930 116.705 108.050 116.815 ;
        RECT 108.395 116.655 108.565 116.845 ;
        RECT 108.855 116.675 109.025 116.865 ;
        RECT 112.535 116.845 112.685 116.865 ;
        RECT 112.535 116.675 112.705 116.845 ;
        RECT 113.460 116.675 113.630 116.865 ;
        RECT 116.030 116.655 116.200 116.845 ;
        RECT 116.215 116.675 116.385 116.865 ;
        RECT 119.895 116.675 120.065 116.865 ;
        RECT 123.300 116.655 123.470 116.845 ;
        RECT 123.575 116.675 123.745 116.865 ;
        RECT 124.035 116.815 124.205 116.845 ;
        RECT 124.030 116.705 124.205 116.815 ;
        RECT 124.035 116.655 124.205 116.705 ;
        RECT 124.495 116.675 124.665 116.865 ;
        RECT 126.335 116.655 126.505 116.845 ;
        RECT 127.715 116.675 127.885 116.865 ;
        RECT 132.315 116.675 132.485 116.865 ;
        RECT 133.695 116.655 133.865 116.845 ;
        RECT 135.535 116.675 135.705 116.865 ;
        RECT 137.835 116.845 138.000 116.865 ;
        RECT 137.375 116.675 137.545 116.845 ;
        RECT 137.835 116.675 138.005 116.845 ;
        RECT 138.290 116.705 138.410 116.815 ;
        RECT 140.140 116.675 140.310 116.865 ;
        RECT 140.600 116.675 140.770 116.895 ;
        RECT 142.730 116.865 143.665 116.895 ;
        RECT 143.770 117.545 144.690 117.775 ;
        RECT 147.395 117.545 148.745 117.775 ;
        RECT 150.280 117.545 151.190 117.765 ;
        RECT 143.770 116.865 147.235 117.545 ;
        RECT 147.395 116.865 154.705 117.545 ;
        RECT 155.635 116.865 157.005 117.675 ;
        RECT 137.525 116.655 137.545 116.675 ;
        RECT 143.355 116.655 143.525 116.845 ;
        RECT 143.810 116.705 143.930 116.815 ;
        RECT 144.275 116.655 144.445 116.845 ;
        RECT 147.035 116.675 147.205 116.865 ;
        RECT 152.095 116.655 152.265 116.845 ;
        RECT 153.475 116.655 153.645 116.845 ;
        RECT 154.395 116.675 154.565 116.865 ;
        RECT 154.865 116.710 155.025 116.820 ;
        RECT 155.310 116.705 155.430 116.815 ;
        RECT 156.695 116.655 156.865 116.865 ;
        RECT 67.280 116.625 68.225 116.655 ;
        RECT 65.155 116.425 68.225 116.625 ;
        RECT 65.015 115.945 68.225 116.425 ;
        RECT 68.925 115.975 72.825 116.655 ;
        RECT 65.015 115.745 65.945 115.945 ;
        RECT 67.280 115.745 68.225 115.945 ;
        RECT 71.895 115.745 72.825 115.975 ;
        RECT 72.835 115.875 74.205 116.655 ;
        RECT 74.225 115.785 74.655 116.570 ;
        RECT 75.135 115.975 82.445 116.655 ;
        RECT 83.415 115.975 92.520 116.655 ;
        RECT 78.650 115.755 79.560 115.975 ;
        RECT 81.095 115.745 82.445 115.975 ;
        RECT 92.615 115.745 93.965 116.655 ;
        RECT 93.995 115.845 95.825 116.655 ;
        RECT 96.295 115.875 97.665 116.655 ;
        RECT 97.835 115.835 99.765 116.655 ;
        RECT 98.815 115.745 99.765 115.835 ;
        RECT 99.985 115.785 100.415 116.570 ;
        RECT 100.475 115.975 107.785 116.655 ;
        RECT 108.255 115.975 115.565 116.655 ;
        RECT 100.475 115.745 101.825 115.975 ;
        RECT 103.360 115.755 104.270 115.975 ;
        RECT 111.770 115.755 112.680 115.975 ;
        RECT 114.215 115.745 115.565 115.975 ;
        RECT 115.615 115.975 119.515 116.655 ;
        RECT 119.985 115.975 123.885 116.655 ;
        RECT 115.615 115.745 116.545 115.975 ;
        RECT 122.955 115.745 123.885 115.975 ;
        RECT 123.895 115.845 125.725 116.655 ;
        RECT 125.745 115.785 126.175 116.570 ;
        RECT 126.195 115.975 133.505 116.655 ;
        RECT 133.665 115.975 137.130 116.655 ;
        RECT 137.525 115.975 139.975 116.655 ;
        RECT 129.710 115.755 130.620 115.975 ;
        RECT 132.155 115.745 133.505 115.975 ;
        RECT 136.210 115.745 137.130 115.975 ;
        RECT 138.015 115.745 139.975 115.975 ;
        RECT 140.090 115.975 143.555 116.655 ;
        RECT 144.135 115.975 151.445 116.655 ;
        RECT 140.090 115.745 141.010 115.975 ;
        RECT 147.650 115.755 148.560 115.975 ;
        RECT 150.095 115.745 151.445 115.975 ;
        RECT 151.505 115.785 151.935 116.570 ;
        RECT 151.955 115.875 153.325 116.655 ;
        RECT 153.335 115.845 155.165 116.655 ;
        RECT 155.635 115.845 157.005 116.655 ;
      LAYER nwell ;
        RECT 22.500 112.625 157.200 115.455 ;
      LAYER pwell ;
        RECT 22.695 111.425 24.065 112.235 ;
        RECT 25.305 112.105 26.235 112.335 ;
        RECT 25.305 111.425 27.140 112.105 ;
        RECT 27.295 111.425 30.770 112.335 ;
        RECT 31.070 112.105 31.990 112.335 ;
        RECT 31.070 111.425 34.535 112.105 ;
        RECT 35.585 111.510 36.015 112.295 ;
        RECT 36.035 111.425 37.405 112.235 ;
        RECT 37.510 112.105 38.430 112.335 ;
        RECT 41.095 112.105 42.440 112.335 ;
        RECT 45.590 112.105 46.510 112.335 ;
        RECT 50.130 112.105 51.040 112.325 ;
        RECT 52.575 112.105 53.925 112.335 ;
        RECT 57.490 112.105 58.400 112.325 ;
        RECT 59.935 112.105 61.285 112.335 ;
        RECT 37.510 111.425 40.975 112.105 ;
        RECT 41.095 111.425 42.925 112.105 ;
        RECT 43.045 111.425 46.510 112.105 ;
        RECT 46.615 111.425 53.925 112.105 ;
        RECT 53.975 111.425 61.285 112.105 ;
        RECT 61.345 111.510 61.775 112.295 ;
        RECT 61.795 111.425 65.270 112.335 ;
        RECT 65.570 112.105 66.490 112.335 ;
        RECT 73.130 112.105 74.040 112.325 ;
        RECT 75.575 112.105 76.925 112.335 ;
        RECT 65.570 111.425 69.035 112.105 ;
        RECT 69.615 111.425 76.925 112.105 ;
        RECT 76.975 111.425 78.345 112.205 ;
        RECT 81.555 112.105 82.485 112.335 ;
        RECT 78.585 111.425 82.485 112.105 ;
        RECT 82.495 112.105 83.425 112.335 ;
        RECT 82.495 111.425 86.395 112.105 ;
        RECT 87.105 111.510 87.535 112.295 ;
        RECT 91.990 112.105 92.900 112.325 ;
        RECT 94.435 112.105 95.785 112.335 ;
        RECT 88.475 111.425 95.785 112.105 ;
        RECT 95.835 112.105 96.765 112.335 ;
        RECT 95.835 111.425 99.735 112.105 ;
        RECT 99.975 111.425 103.645 112.235 ;
        RECT 103.655 111.425 105.025 112.235 ;
        RECT 105.035 112.105 105.965 112.335 ;
        RECT 105.035 111.425 108.935 112.105 ;
        RECT 109.635 111.425 111.005 112.205 ;
        RECT 111.015 111.425 112.845 112.235 ;
        RECT 112.865 111.510 113.295 112.295 ;
        RECT 114.455 112.245 115.405 112.335 ;
        RECT 113.475 111.425 115.405 112.245 ;
        RECT 115.695 112.105 117.465 112.335 ;
        RECT 119.000 112.105 119.910 112.325 ;
        RECT 115.695 111.425 123.425 112.105 ;
        RECT 123.435 111.425 125.265 112.235 ;
        RECT 128.790 112.105 129.700 112.325 ;
        RECT 131.235 112.105 132.585 112.335 ;
        RECT 125.275 111.425 132.585 112.105 ;
        RECT 133.095 111.425 136.305 112.335 ;
        RECT 136.515 112.245 137.465 112.335 ;
        RECT 136.515 111.425 138.445 112.245 ;
        RECT 138.625 111.510 139.055 112.295 ;
        RECT 139.095 111.425 140.445 112.335 ;
        RECT 140.650 111.425 144.125 112.335 ;
        RECT 144.445 112.105 145.375 112.335 ;
        RECT 144.445 111.425 146.280 112.105 ;
        RECT 146.435 111.425 155.540 112.105 ;
        RECT 155.635 111.425 157.005 112.235 ;
        RECT 22.835 111.215 23.005 111.425 ;
        RECT 26.975 111.405 27.140 111.425 ;
        RECT 24.215 111.215 24.385 111.405 ;
        RECT 26.975 111.235 27.145 111.405 ;
        RECT 27.440 111.235 27.610 111.425 ;
        RECT 32.955 111.215 33.125 111.405 ;
        RECT 33.415 111.215 33.585 111.405 ;
        RECT 34.335 111.235 34.505 111.425 ;
        RECT 34.805 111.270 34.965 111.380 ;
        RECT 36.175 111.235 36.345 111.425 ;
        RECT 40.775 111.235 40.945 111.425 ;
        RECT 42.615 111.235 42.785 111.425 ;
        RECT 43.075 111.405 43.245 111.425 ;
        RECT 43.075 111.235 43.250 111.405 ;
        RECT 40.780 111.215 40.945 111.235 ;
        RECT 43.080 111.215 43.250 111.235 ;
        RECT 46.755 111.215 46.925 111.425 ;
        RECT 49.050 111.265 49.170 111.375 ;
        RECT 52.735 111.215 52.905 111.405 ;
        RECT 22.695 110.405 24.065 111.215 ;
        RECT 24.075 110.535 31.385 111.215 ;
        RECT 27.590 110.315 28.500 110.535 ;
        RECT 30.035 110.305 31.385 110.535 ;
        RECT 31.435 110.535 33.265 111.215 ;
        RECT 33.275 110.535 40.585 111.215 ;
        RECT 40.780 110.535 42.615 111.215 ;
        RECT 31.435 110.305 32.780 110.535 ;
        RECT 36.790 110.315 37.700 110.535 ;
        RECT 39.235 110.305 40.585 110.535 ;
        RECT 41.685 110.305 42.615 110.535 ;
        RECT 42.935 110.305 46.410 111.215 ;
        RECT 46.615 110.405 48.445 111.215 ;
        RECT 48.465 110.345 48.895 111.130 ;
        RECT 49.470 110.535 52.935 111.215 ;
        RECT 53.200 111.185 53.370 111.405 ;
        RECT 54.115 111.235 54.285 111.425 ;
        RECT 61.940 111.405 62.110 111.425 ;
        RECT 57.795 111.235 57.965 111.405 ;
        RECT 58.250 111.265 58.370 111.375 ;
        RECT 61.935 111.235 62.110 111.405 ;
        RECT 57.795 111.215 57.960 111.235 ;
        RECT 61.935 111.215 62.105 111.235 ;
        RECT 54.860 111.185 55.805 111.215 ;
        RECT 49.470 110.305 50.390 110.535 ;
        RECT 53.055 110.505 55.805 111.185 ;
        RECT 54.860 110.305 55.805 110.505 ;
        RECT 56.125 110.535 57.960 111.215 ;
        RECT 58.670 110.535 62.135 111.215 ;
        RECT 62.400 111.185 62.570 111.405 ;
        RECT 65.155 111.215 65.325 111.405 ;
        RECT 66.535 111.215 66.705 111.405 ;
        RECT 68.835 111.235 69.005 111.425 ;
        RECT 69.290 111.265 69.410 111.375 ;
        RECT 69.755 111.235 69.925 111.425 ;
        RECT 71.135 111.215 71.305 111.405 ;
        RECT 71.595 111.215 71.765 111.405 ;
        RECT 74.825 111.260 74.985 111.370 ;
        RECT 75.740 111.215 75.910 111.405 ;
        RECT 77.115 111.235 77.285 111.425 ;
        RECT 78.505 111.260 78.665 111.370 ;
        RECT 79.415 111.215 79.585 111.405 ;
        RECT 81.900 111.235 82.070 111.425 ;
        RECT 82.910 111.235 83.080 111.425 ;
        RECT 86.770 111.265 86.890 111.375 ;
        RECT 87.705 111.270 87.865 111.380 ;
        RECT 88.615 111.235 88.785 111.425 ;
        RECT 89.075 111.235 89.245 111.405 ;
        RECT 89.545 111.260 89.705 111.370 ;
        RECT 89.075 111.215 89.225 111.235 ;
        RECT 91.375 111.215 91.545 111.405 ;
        RECT 92.750 111.215 92.920 111.405 ;
        RECT 93.215 111.235 93.385 111.405 ;
        RECT 93.235 111.215 93.385 111.235 ;
        RECT 95.515 111.215 95.685 111.405 ;
        RECT 96.250 111.235 96.420 111.425 ;
        RECT 99.205 111.260 99.365 111.370 ;
        RECT 100.115 111.235 100.285 111.425 ;
        RECT 100.575 111.215 100.745 111.405 ;
        RECT 102.415 111.215 102.585 111.405 ;
        RECT 103.795 111.215 103.965 111.425 ;
        RECT 105.450 111.235 105.620 111.425 ;
        RECT 109.310 111.265 109.430 111.375 ;
        RECT 110.695 111.235 110.865 111.425 ;
        RECT 111.155 111.235 111.325 111.425 ;
        RECT 113.475 111.405 113.625 111.425 ;
        RECT 112.995 111.235 113.165 111.405 ;
        RECT 112.995 111.215 113.145 111.235 ;
        RECT 113.455 111.215 113.625 111.405 ;
        RECT 117.135 111.235 117.305 111.405 ;
        RECT 117.155 111.215 117.305 111.235 ;
        RECT 119.435 111.215 119.605 111.405 ;
        RECT 123.115 111.235 123.285 111.425 ;
        RECT 123.575 111.235 123.745 111.425 ;
        RECT 124.965 111.260 125.125 111.370 ;
        RECT 125.415 111.235 125.585 111.425 ;
        RECT 126.335 111.215 126.505 111.405 ;
        RECT 131.855 111.215 132.025 111.405 ;
        RECT 132.770 111.265 132.890 111.375 ;
        RECT 133.235 111.235 133.405 111.425 ;
        RECT 138.295 111.405 138.445 111.425 ;
        RECT 134.615 111.215 134.785 111.405 ;
        RECT 135.075 111.215 135.245 111.405 ;
        RECT 137.835 111.215 138.005 111.405 ;
        RECT 138.295 111.215 138.465 111.405 ;
        RECT 139.210 111.235 139.380 111.425 ;
        RECT 143.810 111.235 143.980 111.425 ;
        RECT 146.115 111.405 146.280 111.425 ;
        RECT 145.655 111.215 145.825 111.405 ;
        RECT 146.115 111.235 146.285 111.405 ;
        RECT 146.575 111.235 146.745 111.425 ;
        RECT 149.335 111.215 149.505 111.405 ;
        RECT 150.725 111.260 150.885 111.370 ;
        RECT 152.095 111.215 152.265 111.405 ;
        RECT 156.695 111.215 156.865 111.425 ;
        RECT 64.060 111.185 65.005 111.215 ;
        RECT 56.125 110.305 57.055 110.535 ;
        RECT 58.670 110.305 59.590 110.535 ;
        RECT 62.255 110.505 65.005 111.185 ;
        RECT 64.060 110.305 65.005 110.505 ;
        RECT 65.025 110.305 66.375 111.215 ;
        RECT 66.495 110.305 69.605 111.215 ;
        RECT 69.615 110.305 71.430 111.215 ;
        RECT 71.455 110.405 74.205 111.215 ;
        RECT 74.225 110.345 74.655 111.130 ;
        RECT 75.595 110.305 78.205 111.215 ;
        RECT 79.275 110.535 87.005 111.215 ;
        RECT 82.790 110.315 83.700 110.535 ;
        RECT 85.235 110.305 87.005 110.535 ;
        RECT 87.295 110.395 89.225 111.215 ;
        RECT 90.315 110.435 91.685 111.215 ;
        RECT 87.295 110.305 88.245 110.395 ;
        RECT 91.715 110.305 93.065 111.215 ;
        RECT 93.235 110.395 95.165 111.215 ;
        RECT 95.375 110.405 99.045 111.215 ;
        RECT 94.215 110.305 95.165 110.395 ;
        RECT 99.985 110.345 100.415 111.130 ;
        RECT 100.435 110.405 102.265 111.215 ;
        RECT 102.275 110.435 103.645 111.215 ;
        RECT 103.655 110.535 110.965 111.215 ;
        RECT 107.170 110.315 108.080 110.535 ;
        RECT 109.615 110.305 110.965 110.535 ;
        RECT 111.215 110.395 113.145 111.215 ;
        RECT 113.315 110.405 116.985 111.215 ;
        RECT 117.155 110.395 119.085 111.215 ;
        RECT 119.295 110.405 124.805 111.215 ;
        RECT 111.215 110.305 112.165 110.395 ;
        RECT 118.135 110.305 119.085 110.395 ;
        RECT 125.745 110.345 126.175 111.130 ;
        RECT 126.195 110.405 131.705 111.215 ;
        RECT 131.715 110.405 133.085 111.215 ;
        RECT 133.095 110.305 134.910 111.215 ;
        RECT 134.935 110.405 136.765 111.215 ;
        RECT 136.785 110.305 138.135 111.215 ;
        RECT 138.155 110.535 145.465 111.215 ;
        RECT 145.625 110.535 149.090 111.215 ;
        RECT 141.670 110.315 142.580 110.535 ;
        RECT 144.115 110.305 145.465 110.535 ;
        RECT 148.170 110.305 149.090 110.535 ;
        RECT 149.205 110.305 150.555 111.215 ;
        RECT 151.505 110.345 151.935 111.130 ;
        RECT 151.955 110.405 155.625 111.215 ;
        RECT 155.635 110.405 157.005 111.215 ;
      LAYER nwell ;
        RECT 22.500 107.185 157.200 110.015 ;
      LAYER pwell ;
        RECT 22.695 105.985 24.065 106.795 ;
        RECT 26.045 106.665 26.975 106.895 ;
        RECT 25.140 105.985 26.975 106.665 ;
        RECT 27.390 106.665 28.310 106.895 ;
        RECT 31.990 106.665 32.910 106.895 ;
        RECT 27.390 105.985 30.855 106.665 ;
        RECT 31.990 105.985 35.455 106.665 ;
        RECT 35.585 106.070 36.015 106.855 ;
        RECT 37.150 105.985 40.625 106.895 ;
        RECT 43.290 106.665 44.210 106.895 ;
        RECT 40.745 105.985 44.210 106.665 ;
        RECT 44.315 105.985 47.790 106.895 ;
        RECT 50.650 106.665 51.570 106.895 ;
        RECT 48.105 105.985 51.570 106.665 ;
        RECT 51.675 105.985 55.150 106.895 ;
        RECT 55.665 106.665 56.595 106.895 ;
        RECT 58.705 106.665 59.635 106.895 ;
        RECT 55.665 105.985 57.500 106.665 ;
        RECT 22.835 105.775 23.005 105.985 ;
        RECT 25.140 105.965 25.305 105.985 ;
        RECT 24.215 105.775 24.385 105.965 ;
        RECT 25.135 105.795 25.305 105.965 ;
        RECT 29.270 105.775 29.440 105.965 ;
        RECT 29.745 105.820 29.905 105.930 ;
        RECT 30.655 105.775 30.825 105.985 ;
        RECT 31.125 105.830 31.285 105.940 ;
        RECT 35.255 105.795 35.425 105.985 ;
        RECT 36.185 105.830 36.345 105.940 ;
        RECT 38.015 105.775 38.185 105.965 ;
        RECT 40.310 105.795 40.480 105.985 ;
        RECT 40.775 105.795 40.945 105.985 ;
        RECT 44.460 105.795 44.630 105.985 ;
        RECT 47.215 105.775 47.385 105.965 ;
        RECT 48.135 105.795 48.305 105.985 ;
        RECT 22.695 104.965 24.065 105.775 ;
        RECT 24.075 104.965 25.905 105.775 ;
        RECT 26.110 104.865 29.585 105.775 ;
        RECT 30.515 105.095 37.825 105.775 ;
        RECT 37.875 105.095 46.980 105.775 ;
        RECT 34.030 104.875 34.940 105.095 ;
        RECT 36.475 104.865 37.825 105.095 ;
        RECT 47.075 104.965 48.445 105.775 ;
        RECT 49.060 105.745 49.230 105.965 ;
        RECT 51.820 105.935 51.990 105.985 ;
        RECT 57.335 105.965 57.500 105.985 ;
        RECT 57.800 105.985 59.635 106.665 ;
        RECT 59.955 105.985 61.325 106.765 ;
        RECT 61.345 106.070 61.775 106.855 ;
        RECT 61.795 105.985 65.465 106.795 ;
        RECT 65.935 105.985 67.765 106.895 ;
        RECT 67.870 106.665 68.790 106.895 ;
        RECT 74.110 106.665 75.030 106.895 ;
        RECT 67.870 105.985 71.335 106.665 ;
        RECT 71.565 105.985 75.030 106.665 ;
        RECT 75.135 105.985 78.805 106.795 ;
        RECT 79.275 105.985 82.945 106.895 ;
        RECT 82.955 105.985 85.705 106.795 ;
        RECT 85.735 105.985 87.085 106.895 ;
        RECT 87.105 106.070 87.535 106.855 ;
        RECT 96.035 106.805 96.985 106.895 ;
        RECT 87.555 105.985 93.065 106.795 ;
        RECT 93.535 105.985 94.905 106.765 ;
        RECT 96.035 105.985 97.965 106.805 ;
        RECT 98.135 105.985 99.965 106.795 ;
        RECT 99.975 105.985 101.345 106.765 ;
        RECT 101.355 105.985 106.865 106.795 ;
        RECT 106.875 105.985 112.385 106.795 ;
        RECT 112.865 106.070 113.295 106.855 ;
        RECT 113.315 105.985 114.665 106.895 ;
        RECT 114.715 105.985 116.065 106.895 ;
        RECT 118.595 106.805 119.545 106.895 ;
        RECT 116.075 105.985 117.445 106.795 ;
        RECT 117.615 105.985 119.545 106.805 ;
        RECT 119.755 105.985 121.585 106.795 ;
        RECT 121.595 105.985 125.070 106.895 ;
        RECT 125.370 106.665 126.290 106.895 ;
        RECT 128.965 106.665 130.925 106.895 ;
        RECT 125.370 105.985 128.835 106.665 ;
        RECT 128.965 105.985 131.415 106.665 ;
        RECT 131.715 105.985 137.225 106.795 ;
        RECT 137.235 105.985 138.605 106.795 ;
        RECT 138.625 106.070 139.055 106.855 ;
        RECT 139.075 105.985 142.745 106.795 ;
        RECT 142.755 105.985 144.125 106.795 ;
        RECT 144.135 105.985 145.485 106.895 ;
        RECT 145.515 105.985 151.025 106.795 ;
        RECT 151.035 105.985 154.705 106.795 ;
        RECT 155.635 105.985 157.005 106.795 ;
        RECT 57.800 105.965 57.965 105.985 ;
        RECT 51.810 105.825 51.990 105.935 ;
        RECT 51.820 105.795 51.990 105.825 ;
        RECT 55.495 105.775 55.665 105.965 ;
        RECT 55.955 105.775 56.125 105.965 ;
        RECT 57.335 105.795 57.505 105.965 ;
        RECT 57.795 105.795 57.965 105.965 ;
        RECT 61.015 105.795 61.185 105.985 ;
        RECT 61.935 105.795 62.105 105.985 ;
        RECT 65.615 105.935 65.785 105.965 ;
        RECT 65.610 105.825 65.785 105.935 ;
        RECT 65.615 105.795 65.785 105.825 ;
        RECT 66.085 105.820 66.245 105.930 ;
        RECT 67.450 105.795 67.620 105.985 ;
        RECT 71.135 105.795 71.305 105.985 ;
        RECT 71.595 105.795 71.765 105.985 ;
        RECT 65.615 105.775 65.780 105.795 ;
        RECT 73.895 105.775 74.065 105.965 ;
        RECT 74.815 105.775 74.985 105.965 ;
        RECT 75.275 105.795 75.445 105.985 ;
        RECT 78.950 105.825 79.070 105.935 ;
        RECT 79.420 105.795 79.590 105.985 ;
        RECT 83.095 105.965 83.265 105.985 ;
        RECT 80.795 105.775 80.965 105.965 ;
        RECT 82.630 105.825 82.750 105.935 ;
        RECT 83.095 105.795 83.270 105.965 ;
        RECT 86.770 105.795 86.940 105.985 ;
        RECT 87.695 105.965 87.865 105.985 ;
        RECT 87.690 105.795 87.865 105.965 ;
        RECT 88.150 105.825 88.270 105.935 ;
        RECT 83.100 105.775 83.270 105.795 ;
        RECT 87.690 105.775 87.860 105.795 ;
        RECT 88.620 105.775 88.790 105.965 ;
        RECT 92.295 105.775 92.465 105.965 ;
        RECT 93.210 105.825 93.330 105.935 ;
        RECT 94.595 105.795 94.765 105.985 ;
        RECT 97.815 105.965 97.965 105.985 ;
        RECT 95.065 105.830 95.225 105.940 ;
        RECT 97.815 105.795 97.985 105.965 ;
        RECT 98.275 105.795 98.445 105.985 ;
        RECT 99.650 105.825 99.770 105.935 ;
        RECT 100.115 105.795 100.285 105.985 ;
        RECT 100.850 105.775 101.020 105.965 ;
        RECT 101.495 105.795 101.665 105.985 ;
        RECT 104.715 105.775 104.885 105.965 ;
        RECT 106.550 105.825 106.670 105.935 ;
        RECT 107.015 105.795 107.185 105.985 ;
        RECT 107.290 105.775 107.460 105.965 ;
        RECT 111.160 105.775 111.330 105.965 ;
        RECT 112.530 105.825 112.650 105.935 ;
        RECT 113.460 105.795 113.630 105.985 ;
        RECT 114.830 105.825 114.950 105.935 ;
        RECT 115.750 105.795 115.920 105.985 ;
        RECT 116.215 105.775 116.385 105.985 ;
        RECT 117.615 105.965 117.765 105.985 ;
        RECT 116.950 105.775 117.120 105.965 ;
        RECT 117.595 105.795 117.765 105.965 ;
        RECT 119.895 105.795 120.065 105.985 ;
        RECT 120.815 105.775 120.985 105.965 ;
        RECT 121.740 105.795 121.910 105.985 ;
        RECT 122.655 105.775 122.825 105.965 ;
        RECT 128.635 105.795 128.805 105.985 ;
        RECT 131.395 105.965 131.415 105.985 ;
        RECT 131.395 105.795 131.565 105.965 ;
        RECT 131.855 105.795 132.025 105.985 ;
        RECT 133.235 105.775 133.405 105.965 ;
        RECT 133.695 105.775 133.865 105.965 ;
        RECT 137.375 105.795 137.545 105.985 ;
        RECT 139.215 105.775 139.385 105.985 ;
        RECT 142.895 105.935 143.065 105.985 ;
        RECT 142.890 105.825 143.065 105.935 ;
        RECT 142.895 105.795 143.065 105.825 ;
        RECT 143.355 105.775 143.525 105.965 ;
        RECT 144.735 105.775 144.905 105.965 ;
        RECT 145.200 105.795 145.370 105.985 ;
        RECT 145.655 105.795 145.825 105.985 ;
        RECT 150.255 105.775 150.425 105.965 ;
        RECT 151.175 105.795 151.345 105.985 ;
        RECT 152.095 105.775 152.265 105.965 ;
        RECT 154.865 105.830 155.025 105.940 ;
        RECT 156.695 105.775 156.865 105.985 ;
        RECT 50.720 105.745 51.665 105.775 ;
        RECT 48.465 104.905 48.895 105.690 ;
        RECT 48.915 105.065 51.665 105.745 ;
        RECT 50.720 104.865 51.665 105.065 ;
        RECT 52.230 105.095 55.695 105.775 ;
        RECT 55.815 105.095 63.545 105.775 ;
        RECT 52.230 104.865 53.150 105.095 ;
        RECT 59.330 104.875 60.240 105.095 ;
        RECT 61.775 104.865 63.545 105.095 ;
        RECT 63.945 105.095 65.780 105.775 ;
        RECT 66.895 105.095 74.205 105.775 ;
        RECT 63.945 104.865 64.875 105.095 ;
        RECT 66.895 104.865 68.245 105.095 ;
        RECT 69.780 104.875 70.690 105.095 ;
        RECT 74.225 104.905 74.655 105.690 ;
        RECT 74.675 104.865 80.515 105.775 ;
        RECT 80.655 104.965 82.485 105.775 ;
        RECT 82.955 104.865 86.625 105.775 ;
        RECT 86.655 104.865 88.005 105.775 ;
        RECT 88.475 104.865 92.145 105.775 ;
        RECT 92.155 105.095 99.465 105.775 ;
        RECT 95.670 104.875 96.580 105.095 ;
        RECT 98.115 104.865 99.465 105.095 ;
        RECT 99.985 104.905 100.415 105.690 ;
        RECT 100.435 105.095 104.335 105.775 ;
        RECT 100.435 104.865 101.365 105.095 ;
        RECT 104.575 104.965 106.405 105.775 ;
        RECT 106.875 105.095 110.775 105.775 ;
        RECT 106.875 104.865 107.805 105.095 ;
        RECT 111.015 104.865 114.685 105.775 ;
        RECT 115.155 104.995 116.525 105.775 ;
        RECT 116.535 105.095 120.435 105.775 ;
        RECT 116.535 104.865 117.465 105.095 ;
        RECT 120.675 104.965 122.505 105.775 ;
        RECT 122.555 104.865 125.725 105.775 ;
        RECT 125.745 104.905 126.175 105.690 ;
        RECT 126.235 105.095 133.545 105.775 ;
        RECT 126.235 104.865 127.585 105.095 ;
        RECT 129.120 104.875 130.030 105.095 ;
        RECT 133.555 104.965 139.065 105.775 ;
        RECT 139.075 104.965 142.745 105.775 ;
        RECT 143.215 104.995 144.585 105.775 ;
        RECT 144.595 104.965 150.105 105.775 ;
        RECT 150.115 104.965 151.485 105.775 ;
        RECT 151.505 104.905 151.935 105.690 ;
        RECT 151.955 104.965 155.625 105.775 ;
        RECT 155.635 104.965 157.005 105.775 ;
      LAYER nwell ;
        RECT 22.500 101.745 157.200 104.575 ;
      LAYER pwell ;
        RECT 22.695 100.545 24.065 101.355 ;
        RECT 24.115 101.225 25.465 101.455 ;
        RECT 27.000 101.225 27.910 101.445 ;
        RECT 24.115 100.545 31.425 101.225 ;
        RECT 32.090 100.545 35.565 101.455 ;
        RECT 35.585 100.630 36.015 101.415 ;
        RECT 37.545 101.225 38.475 101.455 ;
        RECT 36.640 100.545 38.475 101.225 ;
        RECT 38.890 101.225 39.810 101.455 ;
        RECT 45.990 101.225 46.900 101.445 ;
        RECT 48.435 101.225 49.785 101.455 ;
        RECT 53.350 101.225 54.260 101.445 ;
        RECT 55.795 101.225 57.145 101.455 ;
        RECT 38.890 100.545 42.355 101.225 ;
        RECT 42.475 100.545 49.785 101.225 ;
        RECT 49.835 100.545 57.145 101.225 ;
        RECT 58.115 101.255 59.045 101.455 ;
        RECT 60.375 101.255 61.325 101.455 ;
        RECT 58.115 100.775 61.325 101.255 ;
        RECT 58.260 100.575 61.325 100.775 ;
        RECT 61.345 100.630 61.775 101.415 ;
        RECT 22.835 100.335 23.005 100.545 ;
        RECT 24.215 100.335 24.385 100.525 ;
        RECT 29.275 100.335 29.445 100.525 ;
        RECT 31.115 100.355 31.285 100.545 ;
        RECT 31.570 100.385 31.690 100.495 ;
        RECT 32.950 100.335 33.120 100.525 ;
        RECT 35.250 100.355 35.420 100.545 ;
        RECT 36.640 100.525 36.805 100.545 ;
        RECT 35.715 100.335 35.885 100.525 ;
        RECT 36.170 100.490 36.290 100.495 ;
        RECT 36.170 100.385 36.345 100.490 ;
        RECT 36.185 100.380 36.345 100.385 ;
        RECT 36.635 100.355 36.805 100.525 ;
        RECT 38.935 100.355 39.105 100.525 ;
        RECT 38.935 100.335 39.100 100.355 ;
        RECT 39.395 100.335 39.565 100.525 ;
        RECT 42.155 100.355 42.325 100.545 ;
        RECT 42.615 100.355 42.785 100.545 ;
        RECT 46.755 100.335 46.925 100.525 ;
        RECT 49.055 100.335 49.225 100.525 ;
        RECT 49.975 100.355 50.145 100.545 ;
        RECT 54.575 100.335 54.745 100.525 ;
        RECT 57.335 100.355 57.505 100.525 ;
        RECT 58.260 100.355 58.430 100.575 ;
        RECT 60.390 100.545 61.325 100.575 ;
        RECT 61.795 100.545 63.165 101.355 ;
        RECT 63.465 100.545 66.385 101.455 ;
        RECT 66.395 101.225 67.530 101.455 ;
        RECT 69.615 101.225 70.535 101.455 ;
        RECT 66.395 100.545 69.605 101.225 ;
        RECT 69.615 100.545 71.905 101.225 ;
        RECT 71.915 100.545 73.745 101.355 ;
        RECT 73.755 100.545 79.595 101.455 ;
        RECT 79.735 100.545 81.565 101.355 ;
        RECT 82.055 100.545 83.405 101.455 ;
        RECT 83.415 100.545 85.245 101.355 ;
        RECT 85.715 100.545 87.065 101.455 ;
        RECT 87.105 100.630 87.535 101.415 ;
        RECT 87.555 100.545 88.925 101.355 ;
        RECT 88.935 100.545 92.605 101.455 ;
        RECT 92.615 100.545 94.445 101.355 ;
        RECT 94.455 101.225 95.385 101.455 ;
        RECT 99.095 101.225 100.445 101.455 ;
        RECT 101.980 101.225 102.890 101.445 ;
        RECT 109.375 101.365 110.325 101.455 ;
        RECT 94.455 100.545 98.355 101.225 ;
        RECT 99.095 100.545 106.405 101.225 ;
        RECT 106.875 100.545 108.245 101.325 ;
        RECT 109.375 100.545 111.305 101.365 ;
        RECT 111.475 100.545 112.845 101.355 ;
        RECT 112.865 100.630 113.295 101.415 ;
        RECT 113.315 100.545 114.685 101.355 ;
        RECT 118.210 101.225 119.120 101.445 ;
        RECT 120.655 101.225 122.005 101.455 ;
        RECT 114.695 100.545 122.005 101.225 ;
        RECT 122.985 100.545 125.715 101.455 ;
        RECT 126.195 100.545 128.945 101.455 ;
        RECT 128.955 100.545 132.625 101.355 ;
        RECT 132.735 100.545 135.845 101.455 ;
        RECT 135.855 100.545 138.605 101.355 ;
        RECT 138.625 100.630 139.055 101.415 ;
        RECT 139.175 100.545 142.285 101.455 ;
        RECT 142.795 101.225 144.145 101.455 ;
        RECT 145.680 101.225 146.590 101.445 ;
        RECT 142.795 100.545 150.105 101.225 ;
        RECT 150.115 100.545 155.625 101.355 ;
        RECT 155.635 100.545 157.005 101.355 ;
        RECT 57.485 100.335 57.505 100.355 ;
        RECT 60.095 100.335 60.265 100.525 ;
        RECT 61.935 100.355 62.105 100.545 ;
        RECT 64.695 100.355 64.865 100.525 ;
        RECT 64.695 100.335 64.845 100.355 ;
        RECT 22.695 99.525 24.065 100.335 ;
        RECT 24.075 99.525 25.905 100.335 ;
        RECT 26.010 99.655 29.475 100.335 ;
        RECT 26.010 99.425 26.930 99.655 ;
        RECT 29.790 99.425 33.265 100.335 ;
        RECT 33.285 99.425 36.015 100.335 ;
        RECT 37.265 99.655 39.100 100.335 ;
        RECT 39.255 99.655 46.565 100.335 ;
        RECT 37.265 99.425 38.195 99.655 ;
        RECT 42.770 99.435 43.680 99.655 ;
        RECT 45.215 99.425 46.565 99.655 ;
        RECT 46.615 99.525 48.445 100.335 ;
        RECT 48.465 99.465 48.895 100.250 ;
        RECT 48.915 99.525 54.425 100.335 ;
        RECT 54.435 99.525 57.185 100.335 ;
        RECT 57.485 99.655 59.935 100.335 ;
        RECT 57.975 99.425 59.935 99.655 ;
        RECT 59.955 99.425 62.705 100.335 ;
        RECT 62.915 99.515 64.845 100.335 ;
        RECT 65.160 100.305 65.330 100.525 ;
        RECT 66.070 100.355 66.240 100.545 ;
        RECT 68.375 100.335 68.545 100.525 ;
        RECT 69.295 100.355 69.465 100.545 ;
        RECT 71.595 100.355 71.765 100.545 ;
        RECT 72.055 100.355 72.225 100.545 ;
        RECT 73.895 100.495 74.065 100.545 ;
        RECT 73.890 100.385 74.065 100.495 ;
        RECT 73.895 100.355 74.065 100.385 ;
        RECT 74.815 100.335 74.985 100.525 ;
        RECT 79.875 100.355 80.045 100.545 ;
        RECT 81.710 100.385 81.830 100.495 ;
        RECT 83.090 100.355 83.260 100.545 ;
        RECT 83.555 100.355 83.725 100.545 ;
        RECT 85.390 100.385 85.510 100.495 ;
        RECT 85.860 100.355 86.030 100.545 ;
        RECT 87.695 100.355 87.865 100.545 ;
        RECT 88.150 100.335 88.320 100.525 ;
        RECT 88.620 100.335 88.790 100.525 ;
        RECT 89.080 100.355 89.250 100.545 ;
        RECT 92.305 100.380 92.465 100.490 ;
        RECT 92.755 100.355 92.925 100.545 ;
        RECT 94.130 100.335 94.300 100.525 ;
        RECT 94.870 100.355 95.040 100.545 ;
        RECT 95.510 100.335 95.680 100.525 ;
        RECT 95.975 100.335 96.145 100.525 ;
        RECT 98.730 100.385 98.850 100.495 ;
        RECT 99.650 100.385 99.770 100.495 ;
        RECT 100.570 100.385 100.690 100.495 ;
        RECT 101.035 100.355 101.205 100.525 ;
        RECT 101.055 100.335 101.205 100.355 ;
        RECT 103.335 100.335 103.505 100.525 ;
        RECT 105.170 100.385 105.290 100.495 ;
        RECT 105.635 100.335 105.805 100.525 ;
        RECT 106.095 100.355 106.265 100.545 ;
        RECT 106.550 100.385 106.670 100.495 ;
        RECT 107.935 100.355 108.105 100.545 ;
        RECT 111.155 100.525 111.305 100.545 ;
        RECT 108.405 100.390 108.565 100.500 ;
        RECT 111.155 100.355 111.325 100.525 ;
        RECT 111.615 100.355 111.785 100.545 ;
        RECT 113.455 100.355 113.625 100.545 ;
        RECT 114.835 100.355 115.005 100.545 ;
        RECT 116.210 100.335 116.380 100.525 ;
        RECT 116.680 100.335 116.850 100.525 ;
        RECT 121.270 100.335 121.440 100.525 ;
        RECT 121.735 100.335 121.905 100.525 ;
        RECT 122.205 100.390 122.365 100.500 ;
        RECT 123.115 100.355 123.285 100.545 ;
        RECT 125.410 100.385 125.530 100.495 ;
        RECT 125.870 100.385 125.990 100.495 ;
        RECT 126.335 100.335 126.505 100.525 ;
        RECT 128.635 100.355 128.805 100.545 ;
        RECT 129.095 100.355 129.265 100.545 ;
        RECT 131.850 100.385 131.970 100.495 ;
        RECT 132.315 100.335 132.485 100.525 ;
        RECT 132.775 100.355 132.945 100.545 ;
        RECT 135.540 100.335 135.710 100.525 ;
        RECT 135.995 100.355 136.165 100.545 ;
        RECT 139.215 100.335 139.385 100.545 ;
        RECT 141.975 100.355 142.145 100.525 ;
        RECT 142.430 100.385 142.550 100.495 ;
        RECT 141.995 100.335 142.145 100.355 ;
        RECT 144.275 100.335 144.445 100.525 ;
        RECT 149.795 100.335 149.965 100.545 ;
        RECT 150.255 100.355 150.425 100.545 ;
        RECT 152.095 100.335 152.265 100.525 ;
        RECT 156.695 100.335 156.865 100.545 ;
        RECT 67.290 100.305 68.225 100.335 ;
        RECT 65.160 100.105 68.225 100.305 ;
        RECT 65.015 99.625 68.225 100.105 ;
        RECT 62.915 99.425 63.865 99.515 ;
        RECT 65.015 99.425 65.945 99.625 ;
        RECT 67.275 99.425 68.225 99.625 ;
        RECT 68.235 99.525 73.745 100.335 ;
        RECT 74.225 99.465 74.655 100.250 ;
        RECT 74.730 99.425 84.750 100.335 ;
        RECT 84.795 99.425 88.465 100.335 ;
        RECT 88.475 99.425 92.145 100.335 ;
        RECT 93.095 99.425 94.445 100.335 ;
        RECT 94.475 99.425 95.825 100.335 ;
        RECT 95.835 99.525 99.505 100.335 ;
        RECT 99.985 99.465 100.415 100.250 ;
        RECT 101.055 99.515 102.985 100.335 ;
        RECT 103.195 99.525 105.025 100.335 ;
        RECT 105.495 99.655 112.805 100.335 ;
        RECT 102.035 99.425 102.985 99.515 ;
        RECT 109.010 99.435 109.920 99.655 ;
        RECT 111.455 99.425 112.805 99.655 ;
        RECT 112.855 99.425 116.525 100.335 ;
        RECT 116.535 99.425 120.205 100.335 ;
        RECT 120.235 99.425 121.585 100.335 ;
        RECT 121.595 99.525 125.265 100.335 ;
        RECT 125.745 99.465 126.175 100.250 ;
        RECT 126.195 99.525 131.705 100.335 ;
        RECT 132.255 99.425 135.255 100.335 ;
        RECT 135.395 99.425 138.870 100.335 ;
        RECT 139.075 99.525 141.825 100.335 ;
        RECT 141.995 99.515 143.925 100.335 ;
        RECT 144.135 99.525 149.645 100.335 ;
        RECT 149.655 99.525 151.485 100.335 ;
        RECT 142.975 99.425 143.925 99.515 ;
        RECT 151.505 99.465 151.935 100.250 ;
        RECT 151.955 99.525 155.625 100.335 ;
        RECT 155.635 99.525 157.005 100.335 ;
      LAYER nwell ;
        RECT 22.500 96.305 157.200 99.135 ;
      LAYER pwell ;
        RECT 22.695 95.105 24.065 95.915 ;
        RECT 24.855 95.785 26.815 96.015 ;
        RECT 24.365 95.105 26.815 95.785 ;
        RECT 26.835 95.105 30.005 96.015 ;
        RECT 30.055 95.105 32.805 96.015 ;
        RECT 33.125 95.785 34.055 96.015 ;
        RECT 33.125 95.105 34.960 95.785 ;
        RECT 35.585 95.190 36.015 95.975 ;
        RECT 39.550 95.785 40.460 96.005 ;
        RECT 41.995 95.785 43.345 96.015 ;
        RECT 36.035 95.105 43.345 95.785 ;
        RECT 43.395 95.105 46.145 95.915 ;
        RECT 49.670 95.785 50.580 96.005 ;
        RECT 52.115 95.785 53.465 96.015 ;
        RECT 57.030 95.785 57.940 96.005 ;
        RECT 59.475 95.785 61.245 96.015 ;
        RECT 46.155 95.105 53.465 95.785 ;
        RECT 53.515 95.105 61.245 95.785 ;
        RECT 61.345 95.190 61.775 95.975 ;
        RECT 61.795 95.105 65.465 95.915 ;
        RECT 69.450 95.785 70.360 96.005 ;
        RECT 71.895 95.785 73.245 96.015 ;
        RECT 65.935 95.105 73.245 95.785 ;
        RECT 73.295 95.105 79.135 96.015 ;
        RECT 79.275 95.105 82.025 95.915 ;
        RECT 82.085 95.105 86.555 96.015 ;
        RECT 87.105 95.190 87.535 95.975 ;
        RECT 87.555 95.105 90.305 95.915 ;
        RECT 90.315 95.105 97.665 96.015 ;
        RECT 97.675 95.105 100.425 95.915 ;
        RECT 100.895 95.105 102.265 95.885 ;
        RECT 102.275 95.105 105.945 95.915 ;
        RECT 106.875 95.105 108.245 95.885 ;
        RECT 108.255 95.105 111.005 95.915 ;
        RECT 111.475 95.105 112.825 96.015 ;
        RECT 112.865 95.190 113.295 95.975 ;
        RECT 123.755 95.785 125.715 96.015 ;
        RECT 113.400 95.105 122.505 95.785 ;
        RECT 123.265 95.105 125.715 95.785 ;
        RECT 126.655 95.815 127.600 96.015 ;
        RECT 126.655 95.135 129.405 95.815 ;
        RECT 126.655 95.105 127.600 95.135 ;
        RECT 22.835 94.895 23.005 95.105 ;
        RECT 24.365 95.085 24.385 95.105 ;
        RECT 24.215 94.895 24.385 95.085 ;
        RECT 29.735 94.895 29.905 95.105 ;
        RECT 30.195 94.915 30.365 95.105 ;
        RECT 34.795 95.085 34.960 95.105 ;
        RECT 33.870 94.895 34.040 95.085 ;
        RECT 34.335 94.895 34.505 95.085 ;
        RECT 34.795 94.915 34.965 95.085 ;
        RECT 35.250 94.945 35.370 95.055 ;
        RECT 36.175 94.915 36.345 95.105 ;
        RECT 38.015 94.915 38.185 95.085 ;
        RECT 38.470 94.945 38.590 95.055 ;
        RECT 40.775 94.915 40.945 95.085 ;
        RECT 38.015 94.895 38.180 94.915 ;
        RECT 40.775 94.895 40.940 94.915 ;
        RECT 41.235 94.895 41.405 95.085 ;
        RECT 43.535 94.915 43.705 95.105 ;
        RECT 45.380 94.895 45.550 95.085 ;
        RECT 46.295 94.915 46.465 95.105 ;
        RECT 47.675 94.915 47.845 95.085 ;
        RECT 48.130 94.945 48.250 95.055 ;
        RECT 47.675 94.895 47.825 94.915 ;
        RECT 49.055 94.895 49.225 95.085 ;
        RECT 52.735 94.895 52.905 95.085 ;
        RECT 53.655 94.915 53.825 95.105 ;
        RECT 55.035 94.915 55.205 95.085 ;
        RECT 55.035 94.895 55.185 94.915 ;
        RECT 55.495 94.895 55.665 95.085 ;
        RECT 61.015 94.895 61.185 95.085 ;
        RECT 61.935 94.915 62.105 95.105 ;
        RECT 65.610 94.945 65.730 95.055 ;
        RECT 66.075 94.915 66.245 95.105 ;
        RECT 66.545 94.940 66.705 95.050 ;
        RECT 68.375 94.895 68.545 95.085 ;
        RECT 68.835 94.895 69.005 95.085 ;
        RECT 73.435 94.915 73.605 95.105 ;
        RECT 74.815 94.895 74.985 95.085 ;
        RECT 77.575 94.915 77.745 95.085 ;
        RECT 79.415 94.915 79.585 95.105 ;
        RECT 77.725 94.895 77.745 94.915 ;
        RECT 80.325 94.895 80.495 95.085 ;
        RECT 82.155 94.915 82.325 95.105 ;
        RECT 83.555 94.895 83.725 95.085 ;
        RECT 86.770 94.945 86.890 95.055 ;
        RECT 87.695 94.915 87.865 95.105 ;
        RECT 89.070 94.945 89.190 95.055 ;
        RECT 89.540 94.895 89.710 95.085 ;
        RECT 93.215 94.895 93.385 95.085 ;
        RECT 96.435 94.895 96.605 95.085 ;
        RECT 97.350 94.915 97.520 95.105 ;
        RECT 97.815 94.915 97.985 95.105 ;
        RECT 99.650 94.945 99.770 95.055 ;
        RECT 100.570 94.945 100.690 95.055 ;
        RECT 101.035 94.915 101.205 95.105 ;
        RECT 102.415 94.915 102.585 95.105 ;
        RECT 106.105 94.950 106.265 95.060 ;
        RECT 107.015 94.915 107.185 95.105 ;
        RECT 107.475 94.895 107.645 95.085 ;
        RECT 108.395 94.915 108.565 95.105 ;
        RECT 111.150 94.945 111.270 95.055 ;
        RECT 111.620 94.915 111.790 95.105 ;
        RECT 114.835 94.895 115.005 95.085 ;
        RECT 118.065 94.895 118.235 95.085 ;
        RECT 118.515 94.895 118.685 95.085 ;
        RECT 122.195 94.915 122.365 95.105 ;
        RECT 123.265 95.085 123.285 95.105 ;
        RECT 129.090 95.085 129.260 95.135 ;
        RECT 129.415 95.105 131.245 96.015 ;
        RECT 131.255 95.105 134.005 95.915 ;
        RECT 134.490 95.105 136.305 96.015 ;
        RECT 137.255 95.105 138.605 96.015 ;
        RECT 138.625 95.190 139.055 95.975 ;
        RECT 139.075 95.105 140.905 96.015 ;
        RECT 140.915 95.105 142.265 96.015 ;
        RECT 142.295 95.105 143.665 95.915 ;
        RECT 145.495 95.785 146.425 96.015 ;
        RECT 148.035 95.925 148.985 96.015 ;
        RECT 143.675 95.105 146.425 95.785 ;
        RECT 147.055 95.105 148.985 95.925 ;
        RECT 149.195 95.105 154.705 95.915 ;
        RECT 155.635 95.105 157.005 95.915 ;
        RECT 122.650 94.945 122.770 95.055 ;
        RECT 123.115 94.915 123.285 95.085 ;
        RECT 125.885 94.950 126.045 95.060 ;
        RECT 126.335 94.895 126.505 95.085 ;
        RECT 129.090 94.915 129.270 95.085 ;
        RECT 129.100 94.895 129.270 94.915 ;
        RECT 130.470 94.895 130.640 95.085 ;
        RECT 130.930 94.915 131.100 95.105 ;
        RECT 131.395 94.915 131.565 95.105 ;
        RECT 131.865 94.940 132.025 95.050 ;
        RECT 132.775 94.895 132.945 95.085 ;
        RECT 134.150 94.945 134.270 95.055 ;
        RECT 134.615 94.915 134.785 95.105 ;
        RECT 137.370 95.085 137.540 95.105 ;
        RECT 135.990 94.895 136.160 95.085 ;
        RECT 136.465 94.940 136.625 95.060 ;
        RECT 137.370 94.915 137.545 95.085 ;
        RECT 139.220 94.915 139.390 95.105 ;
        RECT 139.670 94.945 139.790 95.055 ;
        RECT 137.380 94.895 137.545 94.915 ;
        RECT 141.050 94.895 141.220 95.085 ;
        RECT 141.515 94.895 141.685 95.085 ;
        RECT 141.980 94.915 142.150 95.105 ;
        RECT 142.435 94.915 142.605 95.105 ;
        RECT 143.815 94.915 143.985 95.105 ;
        RECT 147.055 95.085 147.205 95.105 ;
        RECT 146.570 94.945 146.690 95.055 ;
        RECT 147.035 94.915 147.205 95.085 ;
        RECT 149.335 94.915 149.505 95.105 ;
        RECT 151.175 94.895 151.345 95.085 ;
        RECT 153.015 94.895 153.185 95.085 ;
        RECT 153.475 94.895 153.645 95.085 ;
        RECT 154.865 94.950 155.025 95.060 ;
        RECT 155.310 94.945 155.430 95.055 ;
        RECT 156.695 94.895 156.865 95.105 ;
        RECT 22.695 94.085 24.065 94.895 ;
        RECT 24.075 94.085 29.585 94.895 ;
        RECT 29.595 94.085 32.345 94.895 ;
        RECT 32.355 93.985 34.185 94.895 ;
        RECT 34.210 93.985 36.025 94.895 ;
        RECT 36.345 94.215 38.180 94.895 ;
        RECT 39.105 94.215 40.940 94.895 ;
        RECT 36.345 93.985 37.275 94.215 ;
        RECT 39.105 93.985 40.035 94.215 ;
        RECT 41.195 93.985 44.305 94.895 ;
        RECT 44.315 93.985 45.665 94.895 ;
        RECT 45.895 94.075 47.825 94.895 ;
        RECT 45.895 93.985 46.845 94.075 ;
        RECT 48.465 94.025 48.895 94.810 ;
        RECT 48.915 94.085 51.665 94.895 ;
        RECT 51.675 94.115 53.045 94.895 ;
        RECT 53.255 94.075 55.185 94.895 ;
        RECT 55.355 94.085 60.865 94.895 ;
        RECT 60.875 94.085 66.385 94.895 ;
        RECT 67.315 94.115 68.685 94.895 ;
        RECT 68.695 94.085 74.205 94.895 ;
        RECT 53.255 93.985 54.205 94.075 ;
        RECT 74.225 94.025 74.655 94.810 ;
        RECT 74.675 94.085 77.425 94.895 ;
        RECT 77.725 94.215 80.175 94.895 ;
        RECT 78.215 93.985 80.175 94.215 ;
        RECT 80.195 93.985 83.405 94.895 ;
        RECT 83.415 94.085 88.925 94.895 ;
        RECT 89.395 93.985 93.065 94.895 ;
        RECT 93.175 93.985 96.285 94.895 ;
        RECT 96.395 93.985 99.505 94.895 ;
        RECT 99.985 94.025 100.415 94.810 ;
        RECT 100.475 94.215 107.785 94.895 ;
        RECT 107.835 94.215 115.145 94.895 ;
        RECT 100.475 93.985 101.825 94.215 ;
        RECT 103.360 93.995 104.270 94.215 ;
        RECT 107.835 93.985 109.185 94.215 ;
        RECT 110.720 93.995 111.630 94.215 ;
        RECT 115.155 93.985 118.365 94.895 ;
        RECT 118.375 94.215 125.685 94.895 ;
        RECT 121.890 93.995 122.800 94.215 ;
        RECT 124.335 93.985 125.685 94.215 ;
        RECT 125.745 94.025 126.175 94.810 ;
        RECT 126.195 93.985 128.945 94.895 ;
        RECT 128.955 93.985 130.305 94.895 ;
        RECT 130.355 93.985 131.705 94.895 ;
        RECT 132.650 93.985 134.465 94.895 ;
        RECT 134.475 93.985 136.305 94.895 ;
        RECT 137.380 94.215 139.215 94.895 ;
        RECT 138.285 93.985 139.215 94.215 ;
        RECT 140.015 93.985 141.365 94.895 ;
        RECT 141.375 93.985 144.125 94.895 ;
        RECT 144.175 94.215 151.485 94.895 ;
        RECT 144.175 93.985 145.525 94.215 ;
        RECT 147.060 93.995 147.970 94.215 ;
        RECT 151.505 94.025 151.935 94.810 ;
        RECT 151.955 94.115 153.325 94.895 ;
        RECT 153.335 94.085 155.165 94.895 ;
        RECT 155.635 94.085 157.005 94.895 ;
      LAYER nwell ;
        RECT 22.500 90.865 157.200 93.695 ;
      LAYER pwell ;
        RECT 22.695 89.665 24.065 90.475 ;
        RECT 24.075 89.665 26.825 90.475 ;
        RECT 27.615 90.345 29.575 90.575 ;
        RECT 27.125 89.665 29.575 90.345 ;
        RECT 29.605 89.665 32.805 90.575 ;
        RECT 32.815 89.665 35.565 90.475 ;
        RECT 35.585 89.750 36.015 90.535 ;
        RECT 36.115 89.665 39.115 90.575 ;
        RECT 40.175 89.665 42.005 90.575 ;
        RECT 42.015 89.665 43.365 90.575 ;
        RECT 43.395 89.665 46.145 90.475 ;
        RECT 46.155 89.665 47.525 90.445 ;
        RECT 47.535 89.665 51.205 90.475 ;
        RECT 51.215 89.665 52.585 90.475 ;
        RECT 52.595 89.665 55.705 90.575 ;
        RECT 55.815 89.665 61.325 90.475 ;
        RECT 61.345 89.750 61.775 90.535 ;
        RECT 62.455 90.485 63.405 90.575 ;
        RECT 62.455 89.665 64.385 90.485 ;
        RECT 64.555 89.665 68.225 90.475 ;
        RECT 69.155 89.665 72.630 90.575 ;
        RECT 72.835 89.665 74.665 90.475 ;
        RECT 75.175 90.345 76.525 90.575 ;
        RECT 78.060 90.345 78.970 90.565 ;
        RECT 75.175 89.665 82.485 90.345 ;
        RECT 82.495 89.665 85.245 90.575 ;
        RECT 85.255 89.665 87.085 90.475 ;
        RECT 87.105 89.750 87.535 90.535 ;
        RECT 100.655 90.485 101.605 90.575 ;
        RECT 107.095 90.485 108.045 90.575 ;
        RECT 87.555 89.665 93.065 90.475 ;
        RECT 93.075 89.665 98.585 90.475 ;
        RECT 99.675 89.665 101.605 90.485 ;
        RECT 101.815 89.665 105.485 90.475 ;
        RECT 106.115 89.665 108.045 90.485 ;
        RECT 108.255 89.665 111.925 90.475 ;
        RECT 112.865 89.750 113.295 90.535 ;
        RECT 113.315 89.665 114.685 90.475 ;
        RECT 114.765 89.665 119.235 90.575 ;
        RECT 119.295 89.665 124.805 90.475 ;
        RECT 124.815 89.665 127.565 90.475 ;
        RECT 129.415 89.665 131.245 90.475 ;
        RECT 134.770 90.345 135.680 90.565 ;
        RECT 137.215 90.345 138.565 90.575 ;
        RECT 131.255 89.665 138.565 90.345 ;
        RECT 138.625 89.750 139.055 90.535 ;
        RECT 139.075 89.665 142.745 90.475 ;
        RECT 142.755 89.665 144.125 90.475 ;
        RECT 144.235 89.665 147.345 90.575 ;
        RECT 147.355 89.665 148.705 90.575 ;
        RECT 148.735 89.665 154.245 90.475 ;
        RECT 154.255 89.665 155.625 90.475 ;
        RECT 155.635 89.665 157.005 90.475 ;
        RECT 22.835 89.455 23.005 89.665 ;
        RECT 24.215 89.455 24.385 89.665 ;
        RECT 27.125 89.645 27.145 89.665 ;
        RECT 26.975 89.475 27.145 89.645 ;
        RECT 29.730 89.475 29.900 89.665 ;
        RECT 32.955 89.475 33.125 89.665 ;
        RECT 22.695 88.645 24.065 89.455 ;
        RECT 24.075 88.775 31.385 89.455 ;
        RECT 27.590 88.555 28.500 88.775 ;
        RECT 30.035 88.545 31.385 88.775 ;
        RECT 31.435 89.425 32.380 89.455 ;
        RECT 33.870 89.425 34.040 89.645 ;
        RECT 34.335 89.455 34.505 89.645 ;
        RECT 36.175 89.475 36.345 89.665 ;
        RECT 37.095 89.455 37.265 89.645 ;
        RECT 37.560 89.455 37.730 89.645 ;
        RECT 39.405 89.510 39.565 89.620 ;
        RECT 40.320 89.475 40.490 89.665 ;
        RECT 43.080 89.475 43.250 89.665 ;
        RECT 43.535 89.475 43.705 89.665 ;
        RECT 46.295 89.475 46.465 89.665 ;
        RECT 47.675 89.475 47.845 89.665 ;
        RECT 48.135 89.455 48.305 89.645 ;
        RECT 49.055 89.455 49.225 89.645 ;
        RECT 51.355 89.475 51.525 89.665 ;
        RECT 51.810 89.455 51.980 89.645 ;
        RECT 52.275 89.455 52.445 89.645 ;
        RECT 55.495 89.475 55.665 89.665 ;
        RECT 55.955 89.475 56.125 89.665 ;
        RECT 64.235 89.645 64.385 89.665 ;
        RECT 57.335 89.455 57.505 89.645 ;
        RECT 57.790 89.505 57.910 89.615 ;
        RECT 58.255 89.455 58.425 89.645 ;
        RECT 61.930 89.505 62.050 89.615 ;
        RECT 64.235 89.475 64.405 89.645 ;
        RECT 64.695 89.475 64.865 89.665 ;
        RECT 66.535 89.455 66.705 89.645 ;
        RECT 66.995 89.455 67.165 89.645 ;
        RECT 68.385 89.510 68.545 89.620 ;
        RECT 69.300 89.475 69.470 89.665 ;
        RECT 72.055 89.455 72.225 89.645 ;
        RECT 72.515 89.455 72.685 89.645 ;
        RECT 72.975 89.475 73.145 89.665 ;
        RECT 74.815 89.615 74.985 89.645 ;
        RECT 74.810 89.505 74.985 89.615 ;
        RECT 74.815 89.455 74.985 89.505 ;
        RECT 77.580 89.455 77.750 89.645 ;
        RECT 79.410 89.455 79.580 89.645 ;
        RECT 31.435 88.745 34.185 89.425 ;
        RECT 31.435 88.545 32.380 88.745 ;
        RECT 34.195 88.645 35.565 89.455 ;
        RECT 35.575 88.545 37.390 89.455 ;
        RECT 37.415 88.545 40.890 89.455 ;
        RECT 41.135 88.775 48.445 89.455 ;
        RECT 41.135 88.545 42.485 88.775 ;
        RECT 44.020 88.555 44.930 88.775 ;
        RECT 48.465 88.585 48.895 89.370 ;
        RECT 48.915 88.645 50.745 89.455 ;
        RECT 50.775 88.545 52.125 89.455 ;
        RECT 52.135 88.775 54.885 89.455 ;
        RECT 53.955 88.545 54.885 88.775 ;
        RECT 54.895 88.545 57.645 89.455 ;
        RECT 58.115 88.675 59.485 89.455 ;
        RECT 59.535 88.775 66.845 89.455 ;
        RECT 59.535 88.545 60.885 88.775 ;
        RECT 62.420 88.555 63.330 88.775 ;
        RECT 66.855 88.645 69.605 89.455 ;
        RECT 69.625 88.545 72.355 89.455 ;
        RECT 72.375 88.645 74.205 89.455 ;
        RECT 74.225 88.585 74.655 89.370 ;
        RECT 74.675 88.645 76.505 89.455 ;
        RECT 76.515 88.545 77.865 89.455 ;
        RECT 77.895 88.545 79.725 89.455 ;
        RECT 79.880 89.425 80.050 89.645 ;
        RECT 82.175 89.475 82.345 89.665 ;
        RECT 82.635 89.615 82.805 89.665 ;
        RECT 82.630 89.505 82.805 89.615 ;
        RECT 82.635 89.475 82.805 89.505 ;
        RECT 84.475 89.455 84.645 89.645 ;
        RECT 84.935 89.455 85.105 89.645 ;
        RECT 85.395 89.475 85.565 89.665 ;
        RECT 87.695 89.475 87.865 89.665 ;
        RECT 92.295 89.455 92.465 89.645 ;
        RECT 93.215 89.475 93.385 89.665 ;
        RECT 99.675 89.645 99.825 89.665 ;
        RECT 96.890 89.455 97.060 89.645 ;
        RECT 97.355 89.455 97.525 89.645 ;
        RECT 98.745 89.510 98.905 89.620 ;
        RECT 99.655 89.475 99.825 89.645 ;
        RECT 100.575 89.455 100.745 89.645 ;
        RECT 101.955 89.475 102.125 89.665 ;
        RECT 106.115 89.645 106.265 89.665 ;
        RECT 102.410 89.505 102.530 89.615 ;
        RECT 103.800 89.455 103.970 89.645 ;
        RECT 104.255 89.455 104.425 89.645 ;
        RECT 105.630 89.505 105.750 89.615 ;
        RECT 106.095 89.475 106.265 89.645 ;
        RECT 108.395 89.475 108.565 89.665 ;
        RECT 109.775 89.455 109.945 89.645 ;
        RECT 112.085 89.510 112.245 89.620 ;
        RECT 112.535 89.455 112.705 89.645 ;
        RECT 113.455 89.475 113.625 89.665 ;
        RECT 118.995 89.645 119.165 89.665 ;
        RECT 114.375 89.475 114.545 89.645 ;
        RECT 114.395 89.455 114.545 89.475 ;
        RECT 116.675 89.455 116.845 89.645 ;
        RECT 118.065 89.500 118.225 89.610 ;
        RECT 118.975 89.475 119.165 89.645 ;
        RECT 119.435 89.475 119.605 89.665 ;
        RECT 120.355 89.455 120.525 89.645 ;
        RECT 124.955 89.475 125.125 89.665 ;
        RECT 125.415 89.455 125.585 89.645 ;
        RECT 126.340 89.455 126.510 89.645 ;
        RECT 127.710 89.505 127.830 89.615 ;
        RECT 128.180 89.455 128.350 89.645 ;
        RECT 129.095 89.475 129.265 89.645 ;
        RECT 129.555 89.475 129.725 89.665 ;
        RECT 131.395 89.475 131.565 89.665 ;
        RECT 133.695 89.455 133.865 89.645 ;
        RECT 139.215 89.615 139.385 89.665 ;
        RECT 139.210 89.505 139.385 89.615 ;
        RECT 139.215 89.475 139.385 89.505 ;
        RECT 139.675 89.475 139.845 89.645 ;
        RECT 139.695 89.455 139.845 89.475 ;
        RECT 141.975 89.455 142.145 89.645 ;
        RECT 142.895 89.475 143.065 89.665 ;
        RECT 143.355 89.455 143.525 89.645 ;
        RECT 144.275 89.475 144.445 89.665 ;
        RECT 148.420 89.645 148.590 89.665 ;
        RECT 148.875 89.645 149.045 89.665 ;
        RECT 147.030 89.505 147.150 89.615 ;
        RECT 148.410 89.475 148.590 89.645 ;
        RECT 148.870 89.475 149.045 89.645 ;
        RECT 148.410 89.455 148.580 89.475 ;
        RECT 148.870 89.455 149.040 89.475 ;
        RECT 150.255 89.455 150.425 89.645 ;
        RECT 152.095 89.455 152.265 89.645 ;
        RECT 154.395 89.475 154.565 89.665 ;
        RECT 156.695 89.455 156.865 89.665 ;
        RECT 81.540 89.425 82.485 89.455 ;
        RECT 79.735 88.745 82.485 89.425 ;
        RECT 81.540 88.545 82.485 88.745 ;
        RECT 82.955 88.545 84.770 89.455 ;
        RECT 84.795 88.775 92.105 89.455 ;
        RECT 88.310 88.555 89.220 88.775 ;
        RECT 90.755 88.545 92.105 88.775 ;
        RECT 92.235 88.545 95.235 89.455 ;
        RECT 95.375 88.545 97.205 89.455 ;
        RECT 97.215 88.645 99.965 89.455 ;
        RECT 99.985 88.585 100.415 89.370 ;
        RECT 100.435 88.645 102.265 89.455 ;
        RECT 102.735 88.545 104.085 89.455 ;
        RECT 104.115 88.645 109.625 89.455 ;
        RECT 109.635 88.775 112.385 89.455 ;
        RECT 111.455 88.545 112.385 88.775 ;
        RECT 112.395 88.645 114.225 89.455 ;
        RECT 114.395 88.635 116.325 89.455 ;
        RECT 116.535 88.675 117.905 89.455 ;
        RECT 120.215 88.645 122.965 89.455 ;
        RECT 115.375 88.545 116.325 88.635 ;
        RECT 122.975 88.545 125.725 89.455 ;
        RECT 125.745 88.585 126.175 89.370 ;
        RECT 126.195 88.545 127.545 89.455 ;
        RECT 128.035 88.775 133.545 89.455 ;
        RECT 132.155 88.545 133.545 88.775 ;
        RECT 133.555 88.645 139.065 89.455 ;
        RECT 139.695 88.635 141.625 89.455 ;
        RECT 141.835 88.675 143.205 89.455 ;
        RECT 143.215 88.645 146.885 89.455 ;
        RECT 140.675 88.545 141.625 88.635 ;
        RECT 147.375 88.545 148.725 89.455 ;
        RECT 148.755 88.545 150.105 89.455 ;
        RECT 150.115 88.645 151.485 89.455 ;
        RECT 151.505 88.585 151.935 89.370 ;
        RECT 151.955 88.645 155.625 89.455 ;
        RECT 155.635 88.645 157.005 89.455 ;
      LAYER nwell ;
        RECT 22.500 85.425 157.200 88.255 ;
      LAYER pwell ;
        RECT 22.695 84.225 24.065 85.035 ;
        RECT 24.075 84.225 26.825 85.035 ;
        RECT 26.835 84.225 29.585 85.135 ;
        RECT 29.615 84.225 30.965 85.135 ;
        RECT 30.995 84.225 32.345 85.135 ;
        RECT 35.585 84.310 36.015 85.095 ;
        RECT 37.055 84.225 40.165 85.135 ;
        RECT 40.175 84.225 42.925 85.035 ;
        RECT 44.315 84.225 47.985 85.035 ;
        RECT 49.375 84.225 52.125 85.035 ;
        RECT 52.615 84.225 53.965 85.135 ;
        RECT 53.975 84.225 55.805 85.035 ;
        RECT 55.815 84.225 58.565 85.135 ;
        RECT 60.395 84.905 61.325 85.135 ;
        RECT 58.575 84.225 61.325 84.905 ;
        RECT 61.345 84.310 61.775 85.095 ;
        RECT 61.895 84.225 65.005 85.135 ;
        RECT 65.015 84.225 68.685 85.035 ;
        RECT 68.780 84.225 77.885 84.905 ;
        RECT 77.895 84.225 80.645 85.135 ;
        RECT 80.675 84.225 82.025 85.135 ;
        RECT 82.035 84.225 85.705 85.035 ;
        RECT 85.715 84.225 87.085 85.035 ;
        RECT 87.105 84.310 87.535 85.095 ;
        RECT 87.555 84.225 89.385 85.135 ;
        RECT 90.335 84.225 91.685 85.135 ;
        RECT 91.695 84.225 93.510 85.135 ;
        RECT 93.535 84.225 97.010 85.135 ;
        RECT 98.265 84.905 99.195 85.135 ;
        RECT 97.360 84.225 99.195 84.905 ;
        RECT 99.975 84.225 102.725 85.135 ;
        RECT 102.835 84.225 105.945 85.135 ;
        RECT 105.955 84.905 106.885 85.135 ;
        RECT 105.955 84.225 108.705 84.905 ;
        RECT 109.735 84.225 112.845 85.135 ;
        RECT 112.865 84.310 113.295 85.095 ;
        RECT 114.275 84.905 115.625 85.135 ;
        RECT 117.160 84.905 118.070 85.125 ;
        RECT 125.715 84.905 127.105 85.135 ;
        RECT 131.235 84.905 132.625 85.135 ;
        RECT 136.755 84.905 138.145 85.135 ;
        RECT 114.275 84.225 121.585 84.905 ;
        RECT 121.595 84.225 127.105 84.905 ;
        RECT 127.115 84.225 132.625 84.905 ;
        RECT 132.635 84.225 138.145 84.905 ;
        RECT 138.625 84.310 139.055 85.095 ;
        RECT 144.430 84.905 145.340 85.125 ;
        RECT 146.875 84.905 148.225 85.135 ;
        RECT 140.915 84.225 148.225 84.905 ;
        RECT 149.195 84.225 152.305 85.135 ;
        RECT 152.415 84.905 153.345 85.135 ;
        RECT 152.415 84.225 155.165 84.905 ;
        RECT 155.635 84.225 157.005 85.035 ;
        RECT 22.835 84.015 23.005 84.225 ;
        RECT 24.215 84.015 24.385 84.225 ;
        RECT 26.050 84.065 26.170 84.175 ;
        RECT 26.975 84.035 27.145 84.225 ;
        RECT 30.650 84.205 30.820 84.225 ;
        RECT 27.435 84.035 27.605 84.205 ;
        RECT 27.895 84.015 28.065 84.205 ;
        RECT 30.650 84.035 30.825 84.205 ;
        RECT 31.110 84.035 31.280 84.225 ;
        RECT 32.505 84.070 32.665 84.180 ;
        RECT 30.655 84.015 30.825 84.035 ;
        RECT 33.420 84.015 33.590 84.205 ;
        RECT 34.335 84.035 34.505 84.205 ;
        RECT 34.805 84.070 34.965 84.180 ;
        RECT 36.185 84.070 36.345 84.180 ;
        RECT 37.095 84.035 37.265 84.225 ;
        RECT 38.935 84.015 39.105 84.205 ;
        RECT 40.315 84.035 40.485 84.225 ;
        RECT 43.075 84.035 43.245 84.205 ;
        RECT 44.455 84.035 44.625 84.225 ;
        RECT 47.670 84.015 47.840 84.205 ;
        RECT 48.135 84.175 48.305 84.205 ;
        RECT 48.130 84.065 48.305 84.175 ;
        RECT 48.135 84.035 48.305 84.065 ;
        RECT 49.060 84.015 49.230 84.205 ;
        RECT 49.515 84.035 49.685 84.225 ;
        RECT 52.270 84.065 52.390 84.175 ;
        RECT 52.730 84.035 52.900 84.225 ;
        RECT 54.115 84.035 54.285 84.225 ;
        RECT 55.495 84.035 55.665 84.205 ;
        RECT 55.955 84.015 56.125 84.225 ;
        RECT 58.715 84.035 58.885 84.225 ;
        RECT 59.630 84.015 59.800 84.205 ;
        RECT 61.020 84.015 61.190 84.205 ;
        RECT 61.475 84.015 61.645 84.205 ;
        RECT 61.935 84.035 62.105 84.225 ;
        RECT 65.155 84.175 65.325 84.225 ;
        RECT 65.150 84.065 65.325 84.175 ;
        RECT 65.155 84.035 65.325 84.065 ;
        RECT 72.515 84.015 72.685 84.205 ;
        RECT 72.975 84.015 73.145 84.205 ;
        RECT 74.815 84.015 74.985 84.205 ;
        RECT 77.575 84.035 77.745 84.225 ;
        RECT 78.035 84.035 78.205 84.205 ;
        RECT 79.415 84.015 79.585 84.205 ;
        RECT 80.335 84.035 80.505 84.225 ;
        RECT 81.710 84.035 81.880 84.225 ;
        RECT 82.175 84.035 82.345 84.225 ;
        RECT 83.555 84.015 83.725 84.205 ;
        RECT 84.025 84.060 84.185 84.170 ;
        RECT 84.940 84.015 85.110 84.205 ;
        RECT 85.855 84.035 86.025 84.225 ;
        RECT 89.070 84.035 89.240 84.225 ;
        RECT 89.545 84.070 89.705 84.180 ;
        RECT 90.450 84.035 90.620 84.225 ;
        RECT 91.835 84.035 92.005 84.205 ;
        RECT 92.295 84.015 92.465 84.205 ;
        RECT 93.215 84.035 93.385 84.225 ;
        RECT 93.680 84.035 93.850 84.225 ;
        RECT 97.360 84.205 97.525 84.225 ;
        RECT 94.130 84.065 94.250 84.175 ;
        RECT 94.590 84.015 94.760 84.205 ;
        RECT 95.975 84.015 96.145 84.205 ;
        RECT 97.355 84.035 97.525 84.205 ;
        RECT 97.810 84.065 97.930 84.175 ;
        RECT 99.195 84.035 99.365 84.205 ;
        RECT 99.650 84.065 99.770 84.175 ;
        RECT 100.115 84.035 100.285 84.225 ;
        RECT 100.575 84.015 100.745 84.205 ;
        RECT 102.410 84.065 102.530 84.175 ;
        RECT 102.875 84.035 103.045 84.225 ;
        RECT 103.790 84.015 103.960 84.205 ;
        RECT 104.255 84.015 104.425 84.205 ;
        RECT 107.935 84.015 108.105 84.205 ;
        RECT 108.395 84.035 108.565 84.225 ;
        RECT 108.865 84.070 109.025 84.180 ;
        RECT 109.775 84.035 109.945 84.225 ;
        RECT 111.610 84.015 111.780 84.205 ;
        RECT 113.000 84.015 113.170 84.205 ;
        RECT 113.455 84.015 113.625 84.205 ;
        RECT 118.975 84.015 119.145 84.205 ;
        RECT 121.275 84.035 121.445 84.225 ;
        RECT 121.740 84.035 121.910 84.225 ;
        RECT 122.655 84.015 122.825 84.205 ;
        RECT 124.035 84.035 124.205 84.205 ;
        RECT 125.410 84.065 125.530 84.175 ;
        RECT 126.335 84.015 126.505 84.205 ;
        RECT 127.260 84.035 127.430 84.225 ;
        RECT 131.865 84.060 132.025 84.170 ;
        RECT 132.780 84.035 132.950 84.225 ;
        RECT 133.695 84.035 133.865 84.205 ;
        RECT 135.075 84.015 135.245 84.205 ;
        RECT 135.530 84.065 135.650 84.175 ;
        RECT 135.995 84.015 136.165 84.205 ;
        RECT 137.380 84.015 137.550 84.205 ;
        RECT 138.290 84.065 138.410 84.175 ;
        RECT 140.135 84.035 140.305 84.205 ;
        RECT 140.590 84.065 140.710 84.175 ;
        RECT 141.055 84.035 141.225 84.225 ;
        RECT 143.815 84.035 143.985 84.205 ;
        RECT 144.275 84.015 144.445 84.205 ;
        RECT 147.035 84.015 147.205 84.205 ;
        RECT 148.425 84.070 148.585 84.180 ;
        RECT 149.795 84.015 149.965 84.205 ;
        RECT 152.095 84.015 152.265 84.225 ;
        RECT 154.855 84.035 155.025 84.225 ;
        RECT 155.310 84.065 155.430 84.175 ;
        RECT 156.695 84.015 156.865 84.225 ;
        RECT 22.695 83.205 24.065 84.015 ;
        RECT 24.075 83.205 25.905 84.015 ;
        RECT 27.755 83.205 30.505 84.015 ;
        RECT 30.515 83.105 33.265 84.015 ;
        RECT 33.275 83.335 38.785 84.015 ;
        RECT 37.395 83.105 38.785 83.335 ;
        RECT 38.795 83.205 42.465 84.015 ;
        RECT 42.475 83.335 47.985 84.015 ;
        RECT 42.475 83.105 43.865 83.335 ;
        RECT 48.465 83.145 48.895 83.930 ;
        RECT 48.915 83.335 54.425 84.015 ;
        RECT 53.035 83.105 54.425 83.335 ;
        RECT 55.815 83.205 58.565 84.015 ;
        RECT 58.595 83.105 59.945 84.015 ;
        RECT 59.955 83.105 61.305 84.015 ;
        RECT 61.335 83.205 65.005 84.015 ;
        RECT 65.515 83.335 72.825 84.015 ;
        RECT 65.515 83.105 66.865 83.335 ;
        RECT 68.400 83.115 69.310 83.335 ;
        RECT 72.835 83.205 74.205 84.015 ;
        RECT 74.225 83.145 74.655 83.930 ;
        RECT 74.715 83.105 77.885 84.015 ;
        RECT 79.275 83.205 81.105 84.015 ;
        RECT 81.115 83.105 83.865 84.015 ;
        RECT 84.795 83.335 90.305 84.015 ;
        RECT 88.915 83.105 90.305 83.335 ;
        RECT 92.155 83.205 93.985 84.015 ;
        RECT 94.475 83.105 95.825 84.015 ;
        RECT 95.835 83.205 97.665 84.015 ;
        RECT 99.985 83.145 100.415 83.930 ;
        RECT 100.435 83.205 102.265 84.015 ;
        RECT 102.755 83.105 104.105 84.015 ;
        RECT 104.115 83.205 107.785 84.015 ;
        RECT 107.795 83.105 110.545 84.015 ;
        RECT 110.575 83.105 111.925 84.015 ;
        RECT 111.935 83.105 113.285 84.015 ;
        RECT 113.315 83.205 118.825 84.015 ;
        RECT 118.835 83.205 122.505 84.015 ;
        RECT 122.515 83.205 123.885 84.015 ;
        RECT 125.745 83.145 126.175 83.930 ;
        RECT 126.195 83.205 131.705 84.015 ;
        RECT 134.015 83.235 135.385 84.015 ;
        RECT 135.855 83.235 137.225 84.015 ;
        RECT 137.235 83.335 142.745 84.015 ;
        RECT 141.355 83.105 142.745 83.335 ;
        RECT 144.135 83.205 146.885 84.015 ;
        RECT 146.895 83.105 149.645 84.015 ;
        RECT 149.655 83.205 151.485 84.015 ;
        RECT 151.505 83.145 151.935 83.930 ;
        RECT 151.955 83.205 155.625 84.015 ;
        RECT 155.635 83.205 157.005 84.015 ;
      LAYER nwell ;
        RECT 22.500 79.985 157.200 82.815 ;
      LAYER pwell ;
        RECT 22.695 78.785 24.065 79.595 ;
        RECT 30.035 79.465 31.425 79.695 ;
        RECT 25.915 78.785 31.425 79.465 ;
        RECT 31.435 78.785 33.265 79.595 ;
        RECT 33.275 78.785 34.625 79.695 ;
        RECT 35.585 78.870 36.015 79.655 ;
        RECT 36.035 78.785 41.545 79.595 ;
        RECT 41.555 78.785 44.305 79.595 ;
        RECT 44.315 78.785 45.685 79.565 ;
        RECT 45.695 78.785 48.445 79.595 ;
        RECT 48.455 78.785 49.825 79.565 ;
        RECT 49.835 78.785 51.665 79.595 ;
        RECT 51.675 78.785 53.045 79.565 ;
        RECT 57.175 79.465 58.565 79.695 ;
        RECT 53.055 78.785 58.565 79.465 ;
        RECT 58.575 78.785 61.325 79.595 ;
        RECT 61.345 78.870 61.775 79.655 ;
        RECT 62.255 78.785 64.085 79.695 ;
        RECT 64.095 78.785 69.605 79.595 ;
        RECT 70.855 79.465 72.815 79.695 ;
        RECT 70.365 78.785 72.815 79.465 ;
        RECT 74.215 78.785 76.045 79.595 ;
        RECT 76.055 79.465 77.445 79.695 ;
        RECT 76.055 78.785 81.565 79.465 ;
        RECT 82.515 78.785 83.865 79.695 ;
        RECT 87.105 78.870 87.535 79.655 ;
        RECT 87.555 78.785 90.305 79.595 ;
        RECT 94.895 79.465 96.285 79.695 ;
        RECT 90.775 78.785 96.285 79.465 ;
        RECT 96.295 78.785 97.665 79.565 ;
        RECT 101.795 79.465 103.185 79.695 ;
        RECT 97.675 78.785 103.185 79.465 ;
        RECT 103.195 78.785 108.705 79.595 ;
        RECT 108.715 78.785 112.385 79.595 ;
        RECT 112.865 78.870 113.295 79.655 ;
        RECT 113.315 78.785 116.985 79.595 ;
        RECT 118.965 79.465 119.895 79.695 ;
        RECT 118.060 78.785 119.895 79.465 ;
        RECT 120.525 79.465 121.455 79.695 ;
        RECT 120.525 78.785 122.360 79.465 ;
        RECT 122.515 78.785 123.865 79.695 ;
        RECT 123.915 78.785 125.265 79.695 ;
        RECT 127.555 79.465 128.485 79.695 ;
        RECT 129.635 79.605 130.585 79.695 ;
        RECT 125.735 78.785 128.485 79.465 ;
        RECT 128.655 78.785 130.585 79.605 ;
        RECT 130.805 78.785 132.155 79.695 ;
        RECT 132.175 78.785 133.545 79.595 ;
        RECT 134.890 79.495 135.845 79.695 ;
        RECT 133.565 78.815 135.845 79.495 ;
        RECT 22.835 78.575 23.005 78.785 ;
        RECT 24.215 78.735 24.385 78.765 ;
        RECT 24.210 78.625 24.385 78.735 ;
        RECT 24.215 78.575 24.385 78.625 ;
        RECT 24.675 78.595 24.845 78.765 ;
        RECT 26.060 78.575 26.230 78.785 ;
        RECT 31.575 78.575 31.745 78.785 ;
        RECT 33.420 78.735 33.590 78.785 ;
        RECT 33.410 78.625 33.590 78.735 ;
        RECT 34.805 78.630 34.965 78.740 ;
        RECT 33.420 78.595 33.590 78.625 ;
        RECT 35.715 78.595 35.885 78.765 ;
        RECT 36.175 78.595 36.345 78.785 ;
        RECT 35.715 78.575 35.880 78.595 ;
        RECT 37.090 78.575 37.260 78.765 ;
        RECT 37.560 78.575 37.730 78.765 ;
        RECT 38.935 78.575 39.105 78.765 ;
        RECT 40.775 78.575 40.945 78.765 ;
        RECT 41.695 78.595 41.865 78.785 ;
        RECT 43.535 78.595 43.705 78.765 ;
        RECT 44.455 78.595 44.625 78.785 ;
        RECT 45.835 78.765 46.005 78.785 ;
        RECT 45.835 78.595 46.015 78.765 ;
        RECT 43.555 78.575 43.705 78.595 ;
        RECT 45.845 78.575 46.015 78.595 ;
        RECT 47.215 78.575 47.385 78.765 ;
        RECT 48.595 78.595 48.765 78.785 ;
        RECT 49.975 78.595 50.145 78.785 ;
        RECT 22.695 77.765 24.065 78.575 ;
        RECT 24.075 77.765 25.905 78.575 ;
        RECT 25.915 77.895 31.425 78.575 ;
        RECT 30.035 77.665 31.425 77.895 ;
        RECT 31.435 77.765 33.265 78.575 ;
        RECT 34.045 77.895 35.880 78.575 ;
        RECT 34.045 77.665 34.975 77.895 ;
        RECT 36.055 77.665 37.405 78.575 ;
        RECT 37.415 77.665 38.765 78.575 ;
        RECT 38.795 77.765 40.625 78.575 ;
        RECT 40.635 77.895 43.385 78.575 ;
        RECT 42.455 77.665 43.385 77.895 ;
        RECT 43.555 77.755 45.485 78.575 ;
        RECT 45.695 77.795 47.065 78.575 ;
        RECT 47.075 77.765 48.445 78.575 ;
        RECT 48.915 78.545 49.870 78.575 ;
        RECT 50.900 78.545 51.070 78.765 ;
        RECT 51.355 78.575 51.525 78.765 ;
        RECT 51.815 78.595 51.985 78.785 ;
        RECT 53.200 78.595 53.370 78.785 ;
        RECT 55.030 78.625 55.150 78.735 ;
        RECT 56.415 78.595 56.585 78.765 ;
        RECT 56.870 78.625 56.990 78.735 ;
        RECT 58.250 78.575 58.420 78.765 ;
        RECT 58.715 78.595 58.885 78.785 ;
        RECT 58.735 78.575 58.885 78.595 ;
        RECT 61.015 78.575 61.185 78.765 ;
        RECT 61.930 78.625 62.050 78.735 ;
        RECT 62.400 78.595 62.570 78.785 ;
        RECT 64.235 78.595 64.405 78.785 ;
        RECT 70.365 78.765 70.385 78.785 ;
        RECT 64.695 78.575 64.865 78.765 ;
        RECT 66.995 78.575 67.165 78.765 ;
        RECT 68.370 78.625 68.490 78.735 ;
        RECT 69.750 78.625 69.870 78.735 ;
        RECT 70.215 78.595 70.385 78.765 ;
        RECT 72.975 78.595 73.145 78.765 ;
        RECT 73.890 78.575 74.060 78.765 ;
        RECT 74.355 78.595 74.525 78.785 ;
        RECT 81.250 78.765 81.420 78.785 ;
        RECT 83.550 78.765 83.720 78.785 ;
        RECT 76.655 78.595 76.825 78.765 ;
        RECT 77.110 78.625 77.230 78.735 ;
        RECT 79.415 78.595 79.585 78.765 ;
        RECT 76.655 78.575 76.820 78.595 ;
        RECT 79.415 78.575 79.580 78.595 ;
        RECT 80.790 78.575 80.960 78.765 ;
        RECT 81.250 78.595 81.430 78.765 ;
        RECT 81.725 78.630 81.885 78.740 ;
        RECT 82.645 78.620 82.805 78.730 ;
        RECT 83.550 78.595 83.725 78.765 ;
        RECT 84.025 78.630 84.185 78.740 ;
        RECT 85.855 78.595 86.025 78.765 ;
        RECT 86.315 78.595 86.485 78.765 ;
        RECT 87.695 78.595 87.865 78.785 ;
        RECT 90.920 78.765 91.090 78.785 ;
        RECT 81.260 78.575 81.430 78.595 ;
        RECT 83.555 78.575 83.725 78.595 ;
        RECT 86.335 78.575 86.485 78.595 ;
        RECT 88.625 78.575 88.795 78.765 ;
        RECT 90.005 78.620 90.165 78.730 ;
        RECT 90.450 78.625 90.570 78.735 ;
        RECT 90.915 78.595 91.090 78.765 ;
        RECT 90.915 78.575 91.085 78.595 ;
        RECT 92.295 78.575 92.465 78.765 ;
        RECT 44.535 77.665 45.485 77.755 ;
        RECT 48.465 77.705 48.895 78.490 ;
        RECT 48.915 77.865 51.195 78.545 ;
        RECT 48.915 77.665 49.870 77.865 ;
        RECT 51.215 77.765 54.885 78.575 ;
        RECT 57.215 77.665 58.565 78.575 ;
        RECT 58.735 77.755 60.665 78.575 ;
        RECT 59.715 77.665 60.665 77.755 ;
        RECT 60.955 77.665 64.405 78.575 ;
        RECT 64.555 77.895 66.845 78.575 ;
        RECT 65.925 77.665 66.845 77.895 ;
        RECT 66.855 77.795 68.225 78.575 ;
        RECT 68.695 77.895 74.205 78.575 ;
        RECT 68.695 77.665 70.085 77.895 ;
        RECT 74.225 77.705 74.655 78.490 ;
        RECT 74.985 77.895 76.820 78.575 ;
        RECT 77.745 77.895 79.580 78.575 ;
        RECT 74.985 77.665 75.915 77.895 ;
        RECT 77.745 77.665 78.675 77.895 ;
        RECT 79.755 77.665 81.105 78.575 ;
        RECT 81.115 77.665 82.465 78.575 ;
        RECT 83.415 77.895 86.165 78.575 ;
        RECT 85.235 77.665 86.165 77.895 ;
        RECT 86.335 77.755 88.265 78.575 ;
        RECT 88.475 77.795 89.845 78.575 ;
        RECT 90.775 77.795 92.145 78.575 ;
        RECT 92.155 77.765 93.525 78.575 ;
        RECT 93.670 78.545 93.840 78.765 ;
        RECT 95.975 78.575 96.145 78.765 ;
        RECT 96.435 78.595 96.605 78.785 ;
        RECT 97.820 78.595 97.990 78.785 ;
        RECT 98.735 78.595 98.905 78.765 ;
        RECT 100.585 78.620 100.745 78.730 ;
        RECT 101.500 78.575 101.670 78.765 ;
        RECT 103.335 78.595 103.505 78.785 ;
        RECT 107.010 78.625 107.130 78.735 ;
        RECT 108.855 78.595 109.025 78.785 ;
        RECT 110.695 78.575 110.865 78.765 ;
        RECT 112.530 78.625 112.650 78.735 ;
        RECT 113.455 78.595 113.625 78.785 ;
        RECT 118.060 78.765 118.225 78.785 ;
        RECT 122.195 78.765 122.360 78.785 ;
        RECT 117.145 78.630 117.305 78.740 ;
        RECT 118.055 78.575 118.225 78.765 ;
        RECT 118.525 78.620 118.685 78.730 ;
        RECT 119.435 78.575 119.605 78.765 ;
        RECT 120.815 78.575 120.985 78.765 ;
        RECT 122.195 78.595 122.365 78.765 ;
        RECT 122.660 78.595 122.830 78.785 ;
        RECT 124.495 78.575 124.665 78.765 ;
        RECT 124.950 78.595 125.120 78.785 ;
        RECT 125.410 78.625 125.530 78.735 ;
        RECT 125.875 78.595 126.045 78.785 ;
        RECT 128.655 78.765 128.805 78.785 ;
        RECT 126.335 78.575 126.505 78.765 ;
        RECT 128.635 78.575 128.805 78.765 ;
        RECT 130.025 78.575 130.195 78.765 ;
        RECT 130.935 78.595 131.105 78.785 ;
        RECT 131.395 78.575 131.565 78.765 ;
        RECT 132.315 78.595 132.485 78.785 ;
        RECT 132.775 78.575 132.945 78.765 ;
        RECT 133.690 78.595 133.860 78.815 ;
        RECT 134.890 78.785 135.845 78.815 ;
        RECT 135.855 78.785 138.605 79.595 ;
        RECT 138.625 78.870 139.055 79.655 ;
        RECT 139.075 78.785 140.445 79.595 ;
        RECT 153.290 79.495 154.245 79.695 ;
        RECT 142.755 78.785 151.860 79.465 ;
        RECT 151.965 78.815 154.245 79.495 ;
        RECT 134.610 78.625 134.730 78.735 ;
        RECT 94.870 78.545 95.825 78.575 ;
        RECT 93.545 77.865 95.825 78.545 ;
        RECT 87.315 77.665 88.265 77.755 ;
        RECT 94.870 77.665 95.825 77.865 ;
        RECT 95.835 77.765 98.585 78.575 ;
        RECT 99.985 77.705 100.415 78.490 ;
        RECT 101.355 77.895 106.865 78.575 ;
        RECT 105.475 77.665 106.865 77.895 ;
        RECT 107.475 77.665 110.925 78.575 ;
        RECT 111.055 77.895 118.365 78.575 ;
        RECT 111.055 77.665 112.405 77.895 ;
        RECT 113.940 77.675 114.850 77.895 ;
        RECT 119.305 77.665 120.655 78.575 ;
        RECT 120.675 77.765 124.345 78.575 ;
        RECT 124.355 77.765 125.725 78.575 ;
        RECT 125.745 77.705 126.175 78.490 ;
        RECT 126.195 77.895 128.485 78.575 ;
        RECT 127.565 77.665 128.485 77.895 ;
        RECT 128.495 77.765 129.865 78.575 ;
        RECT 129.875 77.795 131.245 78.575 ;
        RECT 131.255 77.795 132.625 78.575 ;
        RECT 132.635 77.765 134.465 78.575 ;
        RECT 135.080 78.545 135.250 78.765 ;
        RECT 135.995 78.595 136.165 78.785 ;
        RECT 137.845 78.620 138.005 78.730 ;
        RECT 138.755 78.575 138.925 78.765 ;
        RECT 139.215 78.595 139.385 78.785 ;
        RECT 140.140 78.575 140.310 78.765 ;
        RECT 141.515 78.595 141.685 78.765 ;
        RECT 141.985 78.630 142.145 78.740 ;
        RECT 142.895 78.595 143.065 78.785 ;
        RECT 152.090 78.765 152.260 78.815 ;
        RECT 153.290 78.785 154.245 78.815 ;
        RECT 154.255 78.785 155.625 79.595 ;
        RECT 155.635 78.785 157.005 79.595 ;
        RECT 145.660 78.575 145.830 78.765 ;
        RECT 150.715 78.575 150.885 78.765 ;
        RECT 151.170 78.625 151.290 78.735 ;
        RECT 152.090 78.595 152.265 78.765 ;
        RECT 154.395 78.595 154.565 78.785 ;
        RECT 152.095 78.575 152.265 78.595 ;
        RECT 155.315 78.575 155.485 78.765 ;
        RECT 156.695 78.575 156.865 78.785 ;
        RECT 136.740 78.545 137.685 78.575 ;
        RECT 134.935 77.865 137.685 78.545 ;
        RECT 136.740 77.665 137.685 77.865 ;
        RECT 138.615 77.795 139.985 78.575 ;
        RECT 139.995 77.895 145.505 78.575 ;
        RECT 144.115 77.665 145.505 77.895 ;
        RECT 145.515 77.665 147.345 78.575 ;
        RECT 147.495 77.665 150.945 78.575 ;
        RECT 151.505 77.705 151.935 78.490 ;
        RECT 151.955 77.895 154.245 78.575 ;
        RECT 153.325 77.665 154.245 77.895 ;
        RECT 154.255 77.795 155.625 78.575 ;
        RECT 155.635 77.765 157.005 78.575 ;
      LAYER nwell ;
        RECT 22.500 74.545 157.200 77.375 ;
      LAYER pwell ;
        RECT 22.695 73.345 24.065 74.155 ;
        RECT 24.075 73.345 29.585 74.155 ;
        RECT 30.065 73.345 31.415 74.255 ;
        RECT 32.205 74.025 33.135 74.255 ;
        RECT 32.205 73.345 34.040 74.025 ;
        RECT 34.195 73.345 35.565 74.155 ;
        RECT 35.585 73.430 36.015 74.215 ;
        RECT 37.855 74.025 38.785 74.255 ;
        RECT 36.035 73.345 38.785 74.025 ;
        RECT 38.995 74.165 39.945 74.255 ;
        RECT 38.995 73.345 40.925 74.165 ;
        RECT 42.465 74.025 43.385 74.255 ;
        RECT 41.095 73.345 43.385 74.025 ;
        RECT 43.865 73.345 45.215 74.255 ;
        RECT 45.235 73.345 46.605 74.125 ;
        RECT 46.625 73.345 49.355 74.255 ;
        RECT 52.100 74.055 53.045 74.255 ;
        RECT 50.295 73.375 53.045 74.055 ;
        RECT 22.835 73.135 23.005 73.345 ;
        RECT 24.215 73.135 24.385 73.345 ;
        RECT 29.735 73.295 29.905 73.325 ;
        RECT 29.730 73.185 29.905 73.295 ;
        RECT 29.735 73.135 29.905 73.185 ;
        RECT 30.195 73.155 30.365 73.345 ;
        RECT 33.875 73.325 34.040 73.345 ;
        RECT 31.570 73.185 31.690 73.295 ;
        RECT 33.415 73.135 33.585 73.325 ;
        RECT 33.875 73.155 34.045 73.325 ;
        RECT 34.335 73.155 34.505 73.345 ;
        RECT 34.800 73.135 34.970 73.325 ;
        RECT 36.175 73.295 36.345 73.345 ;
        RECT 40.775 73.325 40.925 73.345 ;
        RECT 36.170 73.185 36.345 73.295 ;
        RECT 36.175 73.155 36.345 73.185 ;
        RECT 36.640 73.135 36.810 73.325 ;
        RECT 38.935 73.135 39.105 73.325 ;
        RECT 40.310 73.135 40.480 73.325 ;
        RECT 40.775 73.155 40.945 73.325 ;
        RECT 41.235 73.155 41.405 73.345 ;
        RECT 42.610 73.135 42.780 73.325 ;
        RECT 43.070 73.185 43.190 73.295 ;
        RECT 22.695 72.325 24.065 73.135 ;
        RECT 24.075 72.325 29.585 73.135 ;
        RECT 29.595 72.325 33.265 73.135 ;
        RECT 33.275 72.325 34.645 73.135 ;
        RECT 34.655 72.225 36.005 73.135 ;
        RECT 36.640 72.905 38.330 73.135 ;
        RECT 36.495 72.225 38.330 72.905 ;
        RECT 38.795 72.325 40.165 73.135 ;
        RECT 40.195 72.225 41.545 73.135 ;
        RECT 41.575 72.225 42.925 73.135 ;
        RECT 43.530 73.105 43.700 73.325 ;
        RECT 43.995 73.155 44.165 73.345 ;
        RECT 45.375 73.155 45.545 73.345 ;
        RECT 48.135 73.135 48.305 73.325 ;
        RECT 49.055 73.135 49.225 73.345 ;
        RECT 49.525 73.190 49.685 73.300 ;
        RECT 44.730 73.105 45.685 73.135 ;
        RECT 43.405 72.425 45.685 73.105 ;
        RECT 44.730 72.225 45.685 72.425 ;
        RECT 45.705 72.225 48.435 73.135 ;
        RECT 48.465 72.265 48.895 73.050 ;
        RECT 48.915 72.325 50.285 73.135 ;
        RECT 50.440 73.105 50.610 73.375 ;
        RECT 52.100 73.345 53.045 73.375 ;
        RECT 53.515 73.345 54.885 74.125 ;
        RECT 59.015 74.025 60.405 74.255 ;
        RECT 54.895 73.345 60.405 74.025 ;
        RECT 61.345 73.430 61.775 74.215 ;
        RECT 64.050 74.055 65.005 74.255 ;
        RECT 62.725 73.375 65.005 74.055 ;
        RECT 52.100 73.105 53.045 73.135 ;
        RECT 53.190 73.105 53.360 73.325 ;
        RECT 53.655 73.155 53.825 73.345 ;
        RECT 55.040 73.155 55.210 73.345 ;
        RECT 55.495 73.135 55.665 73.325 ;
        RECT 56.870 73.185 56.990 73.295 ;
        RECT 58.255 73.155 58.425 73.325 ;
        RECT 58.715 73.135 58.885 73.325 ;
        RECT 60.565 73.190 60.725 73.300 ;
        RECT 61.945 73.190 62.105 73.300 ;
        RECT 62.405 73.180 62.565 73.290 ;
        RECT 62.850 73.155 63.020 73.375 ;
        RECT 64.050 73.345 65.005 73.375 ;
        RECT 65.515 74.025 66.865 74.255 ;
        RECT 68.400 74.025 69.310 74.245 ;
        RECT 65.515 73.345 72.825 74.025 ;
        RECT 72.845 73.345 74.195 74.255 ;
        RECT 74.215 73.345 77.885 74.155 ;
        RECT 78.375 73.345 79.725 74.255 ;
        RECT 79.735 73.345 83.405 74.155 ;
        RECT 85.705 74.025 86.625 74.255 ;
        RECT 84.335 73.345 86.625 74.025 ;
        RECT 87.105 73.430 87.535 74.215 ;
        RECT 87.565 73.345 88.915 74.255 ;
        RECT 89.395 73.345 90.765 74.125 ;
        RECT 90.775 73.345 96.285 74.155 ;
        RECT 96.295 73.345 97.665 74.125 ;
        RECT 97.675 73.345 99.045 74.125 ;
        RECT 104.555 74.025 105.945 74.255 ;
        RECT 100.435 73.345 105.945 74.025 ;
        RECT 106.435 73.345 107.785 74.255 ;
        RECT 108.935 74.165 109.885 74.255 ;
        RECT 107.955 73.345 109.885 74.165 ;
        RECT 111.430 74.055 112.385 74.255 ;
        RECT 110.105 73.375 112.385 74.055 ;
        RECT 112.865 73.430 113.295 74.215 ;
        RECT 114.685 74.025 115.605 74.255 ;
        RECT 63.315 73.155 63.485 73.325 ;
        RECT 65.150 73.185 65.270 73.295 ;
        RECT 63.320 73.135 63.485 73.155 ;
        RECT 66.540 73.135 66.710 73.325 ;
        RECT 66.995 73.135 67.165 73.325 ;
        RECT 72.515 73.295 72.685 73.345 ;
        RECT 72.510 73.185 72.685 73.295 ;
        RECT 72.515 73.155 72.685 73.185 ;
        RECT 72.975 73.155 73.145 73.345 ;
        RECT 73.890 73.135 74.060 73.325 ;
        RECT 74.355 73.155 74.525 73.345 ;
        RECT 74.815 73.135 74.985 73.325 ;
        RECT 78.030 73.135 78.200 73.325 ;
        RECT 78.495 73.135 78.665 73.325 ;
        RECT 79.410 73.155 79.580 73.345 ;
        RECT 79.875 73.155 80.045 73.345 ;
        RECT 84.475 73.325 84.645 73.345 ;
        RECT 83.095 73.155 83.265 73.325 ;
        RECT 83.565 73.180 83.725 73.300 ;
        RECT 84.475 73.155 84.650 73.325 ;
        RECT 83.095 73.135 83.245 73.155 ;
        RECT 84.480 73.135 84.650 73.155 ;
        RECT 85.850 73.135 86.020 73.325 ;
        RECT 86.770 73.185 86.890 73.295 ;
        RECT 87.230 73.185 87.350 73.295 ;
        RECT 87.695 73.155 87.865 73.345 ;
        RECT 89.070 73.185 89.190 73.295 ;
        RECT 89.535 73.155 89.705 73.345 ;
        RECT 89.995 73.135 90.165 73.325 ;
        RECT 90.455 73.135 90.625 73.325 ;
        RECT 90.915 73.155 91.085 73.345 ;
        RECT 94.595 73.135 94.765 73.325 ;
        RECT 54.390 73.105 55.345 73.135 ;
        RECT 50.295 72.425 53.045 73.105 ;
        RECT 53.065 72.425 55.345 73.105 ;
        RECT 52.100 72.225 53.045 72.425 ;
        RECT 54.390 72.225 55.345 72.425 ;
        RECT 55.355 72.355 56.725 73.135 ;
        RECT 58.575 72.325 62.245 73.135 ;
        RECT 63.320 72.455 65.155 73.135 ;
        RECT 64.225 72.225 65.155 72.455 ;
        RECT 65.475 72.225 66.825 73.135 ;
        RECT 66.855 72.325 72.365 73.135 ;
        RECT 72.855 72.225 74.205 73.135 ;
        RECT 74.225 72.265 74.655 73.050 ;
        RECT 74.675 72.325 76.045 73.135 ;
        RECT 76.510 72.905 78.200 73.135 ;
        RECT 76.510 72.225 78.345 72.905 ;
        RECT 78.355 72.455 81.105 73.135 ;
        RECT 80.175 72.225 81.105 72.455 ;
        RECT 81.315 72.315 83.245 73.135 ;
        RECT 81.315 72.225 82.265 72.315 ;
        RECT 84.335 72.225 85.685 73.135 ;
        RECT 85.735 72.225 87.085 73.135 ;
        RECT 87.565 72.225 90.295 73.135 ;
        RECT 90.315 72.325 92.145 73.135 ;
        RECT 92.165 72.225 94.895 73.135 ;
        RECT 95.060 73.105 95.230 73.325 ;
        RECT 96.435 73.155 96.605 73.345 ;
        RECT 97.815 73.155 97.985 73.345 ;
        RECT 100.580 73.325 100.750 73.345 ;
        RECT 99.195 73.155 99.365 73.325 ;
        RECT 100.570 73.155 100.750 73.325 ;
        RECT 97.820 73.135 97.985 73.155 ;
        RECT 96.720 73.105 97.665 73.135 ;
        RECT 94.915 72.425 97.665 73.105 ;
        RECT 97.820 72.455 99.655 73.135 ;
        RECT 100.570 73.105 100.740 73.155 ;
        RECT 102.875 73.135 103.045 73.325 ;
        RECT 106.090 73.185 106.210 73.295 ;
        RECT 107.470 73.155 107.640 73.345 ;
        RECT 107.955 73.325 108.105 73.345 ;
        RECT 107.935 73.155 108.105 73.325 ;
        RECT 108.390 73.185 108.510 73.295 ;
        RECT 108.860 73.135 109.030 73.325 ;
        RECT 110.230 73.155 110.400 73.375 ;
        RECT 111.430 73.345 112.385 73.375 ;
        RECT 113.315 73.345 115.605 74.025 ;
        RECT 115.615 73.345 116.985 74.125 ;
        RECT 116.995 73.345 118.365 74.155 ;
        RECT 118.395 73.345 119.745 74.255 ;
        RECT 122.035 74.025 122.965 74.255 ;
        RECT 120.215 73.345 122.965 74.025 ;
        RECT 123.175 74.165 124.125 74.255 ;
        RECT 123.175 73.345 125.105 74.165 ;
        RECT 125.730 73.575 127.565 74.255 ;
        RECT 125.730 73.345 127.420 73.575 ;
        RECT 127.575 73.345 128.925 74.255 ;
        RECT 128.965 73.345 131.695 74.255 ;
        RECT 132.185 73.345 134.915 74.255 ;
        RECT 136.740 74.055 137.685 74.255 ;
        RECT 134.935 73.375 137.685 74.055 ;
        RECT 138.625 73.430 139.055 74.215 ;
        RECT 143.655 74.025 145.045 74.255 ;
        RECT 146.195 74.165 147.145 74.255 ;
        RECT 110.695 73.135 110.865 73.325 ;
        RECT 112.530 73.185 112.650 73.295 ;
        RECT 113.455 73.155 113.625 73.345 ;
        RECT 115.755 73.155 115.925 73.345 ;
        RECT 116.215 73.135 116.385 73.325 ;
        RECT 117.135 73.155 117.305 73.345 ;
        RECT 117.590 73.135 117.760 73.325 ;
        RECT 118.975 73.135 119.145 73.325 ;
        RECT 119.430 73.155 119.600 73.345 ;
        RECT 119.890 73.185 120.010 73.295 ;
        RECT 120.355 73.155 120.525 73.345 ;
        RECT 124.955 73.325 125.105 73.345 ;
        RECT 124.495 73.135 124.665 73.325 ;
        RECT 124.955 73.155 125.125 73.325 ;
        RECT 126.330 73.185 126.450 73.295 ;
        RECT 127.250 73.155 127.420 73.345 ;
        RECT 127.720 73.135 127.890 73.345 ;
        RECT 128.170 73.135 128.340 73.325 ;
        RECT 129.565 73.180 129.725 73.290 ;
        RECT 101.770 73.105 102.725 73.135 ;
        RECT 96.720 72.225 97.665 72.425 ;
        RECT 98.725 72.225 99.655 72.455 ;
        RECT 99.985 72.265 100.415 73.050 ;
        RECT 100.445 72.425 102.725 73.105 ;
        RECT 101.770 72.225 102.725 72.425 ;
        RECT 102.735 72.325 108.245 73.135 ;
        RECT 108.715 72.225 110.545 73.135 ;
        RECT 110.555 72.325 116.065 73.135 ;
        RECT 116.075 72.325 117.445 73.135 ;
        RECT 117.475 72.225 118.825 73.135 ;
        RECT 118.835 72.325 124.345 73.135 ;
        RECT 124.355 72.325 125.725 73.135 ;
        RECT 125.745 72.265 126.175 73.050 ;
        RECT 126.655 72.225 128.005 73.135 ;
        RECT 128.055 72.225 129.405 73.135 ;
        RECT 130.470 73.105 130.640 73.325 ;
        RECT 131.395 73.155 131.565 73.345 ;
        RECT 131.850 73.185 131.970 73.295 ;
        RECT 132.770 73.185 132.890 73.295 ;
        RECT 133.235 73.155 133.405 73.325 ;
        RECT 134.615 73.155 134.785 73.345 ;
        RECT 135.080 73.155 135.250 73.375 ;
        RECT 136.740 73.345 137.685 73.375 ;
        RECT 139.535 73.345 145.045 74.025 ;
        RECT 145.215 73.345 147.145 74.165 ;
        RECT 148.315 74.025 149.665 74.255 ;
        RECT 151.200 74.025 152.110 74.245 ;
        RECT 148.315 73.345 155.625 74.025 ;
        RECT 155.635 73.345 157.005 74.155 ;
        RECT 139.680 73.325 139.850 73.345 ;
        RECT 145.215 73.325 145.365 73.345 ;
        RECT 133.240 73.135 133.405 73.155 ;
        RECT 131.670 73.105 132.625 73.135 ;
        RECT 130.345 72.425 132.625 73.105 ;
        RECT 133.240 72.455 135.075 73.135 ;
        RECT 135.530 73.105 135.700 73.325 ;
        RECT 137.845 73.295 138.005 73.300 ;
        RECT 137.830 73.190 138.005 73.295 ;
        RECT 137.830 73.185 137.950 73.190 ;
        RECT 138.295 73.135 138.465 73.325 ;
        RECT 139.210 73.185 139.330 73.295 ;
        RECT 139.675 73.155 139.850 73.325 ;
        RECT 141.975 73.155 142.145 73.325 ;
        RECT 139.675 73.135 139.845 73.155 ;
        RECT 142.435 73.135 142.605 73.325 ;
        RECT 145.195 73.155 145.365 73.325 ;
        RECT 146.125 73.180 146.285 73.290 ;
        RECT 147.505 73.190 147.665 73.300 ;
        RECT 147.950 73.135 148.120 73.325 ;
        RECT 148.415 73.135 148.585 73.325 ;
        RECT 151.170 73.185 151.290 73.295 ;
        RECT 152.095 73.135 152.265 73.325 ;
        RECT 155.315 73.155 155.485 73.345 ;
        RECT 156.695 73.135 156.865 73.345 ;
        RECT 136.730 73.105 137.685 73.135 ;
        RECT 131.670 72.225 132.625 72.425 ;
        RECT 134.145 72.225 135.075 72.455 ;
        RECT 135.405 72.425 137.685 73.105 ;
        RECT 136.730 72.225 137.685 72.425 ;
        RECT 138.155 72.355 139.525 73.135 ;
        RECT 139.535 72.355 140.905 73.135 ;
        RECT 142.295 72.325 145.965 73.135 ;
        RECT 146.915 72.225 148.265 73.135 ;
        RECT 148.275 72.325 151.025 73.135 ;
        RECT 151.505 72.265 151.935 73.050 ;
        RECT 151.955 72.325 155.625 73.135 ;
        RECT 155.635 72.325 157.005 73.135 ;
      LAYER nwell ;
        RECT 22.500 69.105 157.200 71.935 ;
      LAYER pwell ;
        RECT 22.695 67.905 24.065 68.715 ;
        RECT 24.075 67.905 27.745 68.715 ;
        RECT 28.215 67.905 29.565 68.815 ;
        RECT 29.615 67.905 30.965 68.815 ;
        RECT 30.995 67.905 32.345 68.815 ;
        RECT 33.295 67.905 34.645 68.815 ;
        RECT 35.585 67.990 36.015 68.775 ;
        RECT 38.005 68.585 38.935 68.815 ;
        RECT 37.100 67.905 38.935 68.585 ;
        RECT 39.255 67.905 44.765 68.715 ;
        RECT 44.775 67.905 47.525 68.715 ;
        RECT 49.045 68.585 49.975 68.815 ;
        RECT 48.140 67.905 49.975 68.585 ;
        RECT 50.755 67.905 52.105 68.815 ;
        RECT 52.155 67.905 53.505 68.815 ;
        RECT 53.515 67.905 54.865 68.815 ;
        RECT 59.935 68.585 61.325 68.815 ;
        RECT 55.815 67.905 61.325 68.585 ;
        RECT 61.345 67.990 61.775 68.775 ;
        RECT 62.755 68.585 64.105 68.815 ;
        RECT 65.640 68.585 66.550 68.805 ;
        RECT 62.755 67.905 70.065 68.585 ;
        RECT 70.995 67.905 72.345 68.815 ;
        RECT 72.395 67.905 73.745 68.815 ;
        RECT 73.775 67.905 75.125 68.815 ;
        RECT 75.135 67.905 76.485 68.815 ;
        RECT 78.485 68.585 79.415 68.815 ;
        RECT 77.580 67.905 79.415 68.585 ;
        RECT 79.735 67.905 82.485 68.715 ;
        RECT 82.515 67.905 83.865 68.815 ;
        RECT 83.895 67.905 85.245 68.815 ;
        RECT 85.255 67.905 87.085 68.715 ;
        RECT 87.105 67.990 87.535 68.775 ;
        RECT 87.555 67.905 88.925 68.715 ;
        RECT 90.270 68.615 91.225 68.815 ;
        RECT 88.945 67.935 91.225 68.615 ;
        RECT 22.835 67.695 23.005 67.905 ;
        RECT 24.215 67.695 24.385 67.905 ;
        RECT 27.890 67.745 28.010 67.855 ;
        RECT 28.360 67.715 28.530 67.905 ;
        RECT 29.735 67.695 29.905 67.885 ;
        RECT 30.650 67.715 30.820 67.905 ;
        RECT 32.030 67.715 32.200 67.905 ;
        RECT 32.505 67.750 32.665 67.860 ;
        RECT 33.410 67.695 33.580 67.905 ;
        RECT 37.100 67.885 37.265 67.905 ;
        RECT 33.875 67.695 34.045 67.885 ;
        RECT 34.805 67.750 34.965 67.860 ;
        RECT 36.185 67.750 36.345 67.860 ;
        RECT 36.630 67.745 36.750 67.855 ;
        RECT 37.095 67.715 37.265 67.885 ;
        RECT 38.010 67.695 38.180 67.885 ;
        RECT 38.475 67.695 38.645 67.885 ;
        RECT 39.395 67.715 39.565 67.905 ;
        RECT 44.915 67.885 45.085 67.905 ;
        RECT 48.140 67.885 48.305 67.905 ;
        RECT 41.235 67.715 41.405 67.885 ;
        RECT 42.610 67.695 42.780 67.885 ;
        RECT 43.990 67.695 44.160 67.885 ;
        RECT 44.450 67.745 44.570 67.855 ;
        RECT 44.915 67.715 45.090 67.885 ;
        RECT 46.290 67.745 46.410 67.855 ;
        RECT 44.920 67.695 45.090 67.715 ;
        RECT 47.670 67.695 47.840 67.885 ;
        RECT 48.135 67.855 48.305 67.885 ;
        RECT 48.130 67.745 48.305 67.855 ;
        RECT 48.135 67.715 48.305 67.745 ;
        RECT 49.055 67.715 49.225 67.885 ;
        RECT 50.430 67.745 50.550 67.855 ;
        RECT 50.900 67.715 51.070 67.905 ;
        RECT 49.060 67.695 49.225 67.715 ;
        RECT 52.270 67.695 52.440 67.885 ;
        RECT 52.745 67.740 52.905 67.850 ;
        RECT 53.190 67.715 53.360 67.905 ;
        RECT 54.580 67.695 54.750 67.905 ;
        RECT 55.960 67.885 56.130 67.905 ;
        RECT 55.045 67.750 55.205 67.860 ;
        RECT 55.955 67.715 56.130 67.885 ;
        RECT 56.415 67.695 56.585 67.885 ;
        RECT 61.935 67.695 62.105 67.885 ;
        RECT 63.315 67.695 63.485 67.885 ;
        RECT 65.615 67.695 65.785 67.885 ;
        RECT 66.995 67.695 67.165 67.885 ;
        RECT 69.755 67.715 69.925 67.905 ;
        RECT 70.225 67.750 70.385 67.860 ;
        RECT 70.675 67.715 70.845 67.885 ;
        RECT 71.140 67.715 71.310 67.905 ;
        RECT 72.055 67.695 72.225 67.885 ;
        RECT 73.430 67.715 73.600 67.905 ;
        RECT 74.810 67.885 74.980 67.905 ;
        RECT 73.890 67.745 74.010 67.855 ;
        RECT 74.810 67.715 74.985 67.885 ;
        RECT 76.200 67.715 76.370 67.905 ;
        RECT 77.580 67.885 77.745 67.905 ;
        RECT 76.665 67.750 76.825 67.860 ;
        RECT 77.575 67.715 77.745 67.885 ;
        RECT 74.815 67.695 74.985 67.715 ;
        RECT 79.410 67.695 79.580 67.885 ;
        RECT 79.875 67.715 80.045 67.905 ;
        RECT 80.795 67.695 80.965 67.885 ;
        RECT 81.255 67.695 81.425 67.885 ;
        RECT 82.630 67.715 82.800 67.905 ;
        RECT 84.010 67.885 84.180 67.905 ;
        RECT 83.550 67.695 83.720 67.885 ;
        RECT 84.010 67.715 84.190 67.885 ;
        RECT 84.020 67.695 84.190 67.715 ;
        RECT 85.395 67.695 85.565 67.905 ;
        RECT 87.695 67.715 87.865 67.905 ;
        RECT 89.070 67.695 89.240 67.935 ;
        RECT 90.270 67.905 91.225 67.935 ;
        RECT 91.235 67.905 92.585 68.815 ;
        RECT 92.635 67.905 93.985 68.815 ;
        RECT 93.995 67.905 95.825 68.715 ;
        RECT 97.640 68.615 98.585 68.815 ;
        RECT 95.835 67.935 98.585 68.615 ;
        RECT 89.535 67.695 89.705 67.885 ;
        RECT 91.380 67.695 91.550 67.905 ;
        RECT 93.670 67.695 93.840 67.905 ;
        RECT 94.135 67.855 94.305 67.905 ;
        RECT 94.130 67.745 94.305 67.855 ;
        RECT 94.135 67.715 94.305 67.745 ;
        RECT 94.595 67.715 94.765 67.885 ;
        RECT 95.980 67.715 96.150 67.935 ;
        RECT 97.640 67.905 98.585 67.935 ;
        RECT 99.515 67.905 100.885 68.685 ;
        RECT 105.015 68.585 106.405 68.815 ;
        RECT 100.895 67.905 106.405 68.585 ;
        RECT 106.415 67.905 108.245 68.715 ;
        RECT 108.255 68.585 109.175 68.815 ;
        RECT 108.255 67.905 110.545 68.585 ;
        RECT 110.555 67.905 111.905 68.815 ;
        RECT 112.865 67.990 113.295 68.775 ;
        RECT 113.315 67.905 115.145 68.715 ;
        RECT 115.155 67.905 116.505 68.815 ;
        RECT 116.555 67.905 117.905 68.815 ;
        RECT 117.935 67.905 119.285 68.815 ;
        RECT 119.295 67.905 120.645 68.815 ;
        RECT 121.615 67.905 122.965 68.815 ;
        RECT 123.745 68.585 124.675 68.815 ;
        RECT 123.745 67.905 125.580 68.585 ;
        RECT 125.735 67.905 129.405 68.715 ;
        RECT 129.875 67.905 131.225 68.815 ;
        RECT 131.255 67.905 132.605 68.815 ;
        RECT 132.655 67.905 134.005 68.815 ;
        RECT 134.015 67.905 136.765 68.715 ;
        RECT 138.625 67.990 139.055 68.775 ;
        RECT 143.655 68.585 145.045 68.815 ;
        RECT 139.535 67.905 145.045 68.585 ;
        RECT 145.055 67.905 146.425 68.685 ;
        RECT 146.435 68.585 147.355 68.815 ;
        RECT 149.045 68.585 149.975 68.815 ;
        RECT 146.435 67.905 148.725 68.585 ;
        RECT 149.045 67.905 150.880 68.585 ;
        RECT 151.055 67.905 152.405 68.815 ;
        RECT 152.415 67.905 155.165 68.715 ;
        RECT 155.635 67.905 157.005 68.715 ;
        RECT 94.600 67.695 94.765 67.715 ;
        RECT 96.895 67.695 97.065 67.885 ;
        RECT 98.745 67.750 98.905 67.860 ;
        RECT 99.655 67.855 99.825 67.905 ;
        RECT 99.650 67.745 99.825 67.855 ;
        RECT 100.570 67.745 100.690 67.855 ;
        RECT 99.655 67.715 99.825 67.745 ;
        RECT 101.040 67.715 101.210 67.905 ;
        RECT 101.955 67.715 102.125 67.885 ;
        RECT 102.415 67.695 102.585 67.885 ;
        RECT 104.255 67.695 104.425 67.885 ;
        RECT 106.555 67.715 106.725 67.905 ;
        RECT 110.235 67.715 110.405 67.905 ;
        RECT 111.620 67.885 111.790 67.905 ;
        RECT 111.615 67.715 111.790 67.885 ;
        RECT 112.085 67.750 112.245 67.860 ;
        RECT 113.455 67.715 113.625 67.905 ;
        RECT 111.620 67.695 111.785 67.715 ;
        RECT 113.915 67.695 114.085 67.885 ;
        RECT 115.300 67.715 115.470 67.905 ;
        RECT 117.590 67.715 117.760 67.905 ;
        RECT 118.970 67.715 119.140 67.905 ;
        RECT 119.440 67.885 119.610 67.905 ;
        RECT 119.435 67.715 119.610 67.885 ;
        RECT 120.825 67.750 120.985 67.860 ;
        RECT 119.435 67.695 119.605 67.715 ;
        RECT 121.275 67.695 121.445 67.885 ;
        RECT 121.730 67.715 121.900 67.905 ;
        RECT 125.415 67.885 125.580 67.905 ;
        RECT 122.660 67.695 122.830 67.885 ;
        RECT 123.110 67.745 123.230 67.855 ;
        RECT 124.950 67.695 125.120 67.885 ;
        RECT 125.415 67.855 125.585 67.885 ;
        RECT 125.410 67.745 125.585 67.855 ;
        RECT 125.415 67.715 125.585 67.745 ;
        RECT 125.875 67.715 126.045 67.905 ;
        RECT 126.340 67.695 126.510 67.885 ;
        RECT 127.715 67.695 127.885 67.885 ;
        RECT 129.550 67.745 129.670 67.855 ;
        RECT 130.020 67.715 130.190 67.905 ;
        RECT 130.480 67.695 130.650 67.885 ;
        RECT 131.400 67.715 131.570 67.905 ;
        RECT 132.770 67.695 132.940 67.885 ;
        RECT 133.245 67.740 133.405 67.850 ;
        RECT 133.690 67.715 133.860 67.905 ;
        RECT 134.155 67.715 134.325 67.905 ;
        RECT 134.160 67.695 134.325 67.715 ;
        RECT 136.460 67.695 136.630 67.885 ;
        RECT 137.835 67.715 138.005 67.885 ;
        RECT 138.290 67.745 138.410 67.855 ;
        RECT 139.210 67.745 139.330 67.855 ;
        RECT 139.680 67.715 139.850 67.905 ;
        RECT 142.435 67.695 142.605 67.885 ;
        RECT 146.115 67.715 146.285 67.905 ;
        RECT 148.415 67.715 148.585 67.905 ;
        RECT 150.715 67.885 150.880 67.905 ;
        RECT 149.795 67.695 149.965 67.885 ;
        RECT 150.715 67.715 150.885 67.885 ;
        RECT 151.170 67.715 151.340 67.905 ;
        RECT 152.095 67.695 152.265 67.885 ;
        RECT 152.555 67.715 152.725 67.905 ;
        RECT 155.310 67.745 155.430 67.855 ;
        RECT 156.695 67.695 156.865 67.905 ;
        RECT 22.695 66.885 24.065 67.695 ;
        RECT 24.075 66.885 29.585 67.695 ;
        RECT 29.595 66.885 32.345 67.695 ;
        RECT 32.375 66.785 33.725 67.695 ;
        RECT 33.735 66.885 36.485 67.695 ;
        RECT 36.975 66.785 38.325 67.695 ;
        RECT 38.335 66.885 40.165 67.695 ;
        RECT 41.575 66.785 42.925 67.695 ;
        RECT 42.955 66.785 44.305 67.695 ;
        RECT 44.775 66.785 46.125 67.695 ;
        RECT 46.635 66.785 47.985 67.695 ;
        RECT 48.465 66.825 48.895 67.610 ;
        RECT 49.060 67.015 50.895 67.695 ;
        RECT 49.965 66.785 50.895 67.015 ;
        RECT 51.235 66.785 52.585 67.695 ;
        RECT 53.515 66.785 54.865 67.695 ;
        RECT 56.275 66.885 61.785 67.695 ;
        RECT 61.795 66.885 63.165 67.695 ;
        RECT 63.175 67.015 65.465 67.695 ;
        RECT 64.545 66.785 65.465 67.015 ;
        RECT 65.475 66.915 66.845 67.695 ;
        RECT 66.855 66.885 70.525 67.695 ;
        RECT 71.915 66.885 73.745 67.695 ;
        RECT 74.225 66.825 74.655 67.610 ;
        RECT 74.675 66.885 78.345 67.695 ;
        RECT 78.375 66.785 79.725 67.695 ;
        RECT 79.735 66.915 81.105 67.695 ;
        RECT 81.115 66.885 82.485 67.695 ;
        RECT 82.515 66.785 83.865 67.695 ;
        RECT 83.875 66.785 85.225 67.695 ;
        RECT 85.255 66.885 88.005 67.695 ;
        RECT 88.035 66.785 89.385 67.695 ;
        RECT 89.395 66.885 91.225 67.695 ;
        RECT 91.235 66.785 92.585 67.695 ;
        RECT 92.635 66.785 93.985 67.695 ;
        RECT 94.600 67.015 96.435 67.695 ;
        RECT 95.505 66.785 96.435 67.015 ;
        RECT 96.755 66.885 99.505 67.695 ;
        RECT 99.985 66.825 100.415 67.610 ;
        RECT 102.275 66.885 104.105 67.695 ;
        RECT 104.115 67.015 111.425 67.695 ;
        RECT 111.620 67.015 113.455 67.695 ;
        RECT 107.630 66.795 108.540 67.015 ;
        RECT 110.075 66.785 111.425 67.015 ;
        RECT 112.525 66.785 113.455 67.015 ;
        RECT 113.775 66.885 119.285 67.695 ;
        RECT 119.295 66.885 121.125 67.695 ;
        RECT 121.135 66.915 122.505 67.695 ;
        RECT 122.515 66.785 123.865 67.695 ;
        RECT 123.915 66.785 125.265 67.695 ;
        RECT 125.745 66.825 126.175 67.610 ;
        RECT 126.195 66.785 127.545 67.695 ;
        RECT 127.575 66.885 130.325 67.695 ;
        RECT 130.335 66.785 131.685 67.695 ;
        RECT 131.735 66.785 133.085 67.695 ;
        RECT 134.160 67.015 135.995 67.695 ;
        RECT 136.315 67.015 142.285 67.695 ;
        RECT 142.295 67.015 149.605 67.695 ;
        RECT 135.065 66.785 135.995 67.015 ;
        RECT 140.500 66.785 142.285 67.015 ;
        RECT 145.810 66.795 146.720 67.015 ;
        RECT 148.255 66.785 149.605 67.015 ;
        RECT 149.655 66.885 151.485 67.695 ;
        RECT 151.505 66.825 151.935 67.610 ;
        RECT 151.955 66.885 155.625 67.695 ;
        RECT 155.635 66.885 157.005 67.695 ;
      LAYER nwell ;
        RECT 22.500 63.665 157.200 66.495 ;
      LAYER pwell ;
        RECT 22.695 62.465 24.065 63.275 ;
        RECT 33.320 63.145 35.105 63.375 ;
        RECT 29.135 62.465 35.105 63.145 ;
        RECT 35.585 62.550 36.015 63.335 ;
        RECT 37.415 62.465 38.785 63.245 ;
        RECT 44.360 63.145 46.145 63.375 ;
        RECT 51.720 63.145 53.505 63.375 ;
        RECT 57.700 63.145 59.485 63.375 ;
        RECT 40.175 62.465 46.145 63.145 ;
        RECT 47.535 62.465 53.505 63.145 ;
        RECT 53.515 62.465 59.485 63.145 ;
        RECT 61.345 62.550 61.775 63.335 ;
        RECT 61.795 62.465 64.545 63.275 ;
        RECT 66.395 63.145 68.180 63.375 ;
        RECT 76.560 63.145 78.345 63.375 ;
        RECT 82.540 63.145 84.325 63.375 ;
        RECT 66.395 62.465 72.365 63.145 ;
        RECT 72.375 62.465 78.345 63.145 ;
        RECT 78.355 62.465 84.325 63.145 ;
        RECT 87.105 62.550 87.535 63.335 ;
        RECT 87.555 62.465 90.305 63.275 ;
        RECT 100.020 63.145 101.805 63.375 ;
        RECT 95.835 62.465 101.805 63.145 ;
        RECT 104.575 62.465 107.325 63.275 ;
        RECT 107.335 62.465 108.705 63.245 ;
        RECT 108.715 62.465 112.385 63.275 ;
        RECT 112.865 62.550 113.295 63.335 ;
        RECT 118.880 63.145 120.665 63.375 ;
        RECT 124.860 63.145 126.645 63.375 ;
        RECT 135.900 63.145 137.685 63.375 ;
        RECT 114.695 62.465 120.665 63.145 ;
        RECT 120.675 62.465 126.645 63.145 ;
        RECT 131.715 62.465 137.685 63.145 ;
        RECT 138.625 62.550 139.055 63.335 ;
        RECT 140.455 62.465 142.285 63.275 ;
        RECT 146.940 63.145 148.725 63.375 ;
        RECT 142.755 62.465 148.725 63.145 ;
        RECT 148.735 62.465 154.245 63.275 ;
        RECT 154.255 62.465 155.625 63.275 ;
        RECT 155.635 62.465 157.005 63.275 ;
        RECT 22.835 62.255 23.005 62.465 ;
        RECT 24.210 62.305 24.330 62.415 ;
        RECT 24.680 62.255 24.850 62.445 ;
        RECT 25.595 62.275 25.765 62.445 ;
        RECT 26.050 62.305 26.170 62.415 ;
        RECT 27.435 62.275 27.605 62.445 ;
        RECT 27.895 62.275 28.065 62.445 ;
        RECT 29.280 62.275 29.450 62.465 ;
        RECT 30.660 62.255 30.830 62.445 ;
        RECT 35.250 62.305 35.370 62.415 ;
        RECT 36.640 62.255 36.810 62.445 ;
        RECT 37.095 62.275 37.265 62.445 ;
        RECT 38.475 62.275 38.645 62.465 ;
        RECT 38.935 62.275 39.105 62.445 ;
        RECT 40.320 62.275 40.490 62.465 ;
        RECT 42.620 62.255 42.790 62.445 ;
        RECT 47.215 62.275 47.385 62.445 ;
        RECT 47.680 62.275 47.850 62.465 ;
        RECT 49.975 62.275 50.145 62.445 ;
        RECT 50.445 62.300 50.605 62.410 ;
        RECT 52.275 62.275 52.445 62.445 ;
        RECT 52.735 62.275 52.905 62.445 ;
        RECT 53.660 62.275 53.830 62.465 ;
        RECT 54.120 62.255 54.290 62.445 ;
        RECT 60.100 62.255 60.270 62.445 ;
        RECT 60.555 62.275 60.725 62.445 ;
        RECT 61.010 62.305 61.130 62.415 ;
        RECT 61.935 62.275 62.105 62.465 ;
        RECT 64.690 62.305 64.810 62.415 ;
        RECT 65.155 62.275 65.325 62.445 ;
        RECT 66.070 62.305 66.190 62.415 ;
        RECT 66.535 62.275 66.705 62.445 ;
        RECT 67.920 62.255 68.090 62.445 ;
        RECT 72.050 62.275 72.220 62.465 ;
        RECT 72.520 62.275 72.690 62.465 ;
        RECT 73.890 62.305 74.010 62.415 ;
        RECT 74.810 62.305 74.930 62.415 ;
        RECT 75.280 62.255 75.450 62.445 ;
        RECT 78.500 62.275 78.670 62.465 ;
        RECT 81.260 62.255 81.430 62.445 ;
        RECT 85.395 62.275 85.565 62.445 ;
        RECT 86.775 62.275 86.945 62.445 ;
        RECT 87.240 62.255 87.410 62.445 ;
        RECT 87.695 62.275 87.865 62.465 ;
        RECT 90.450 62.305 90.570 62.415 ;
        RECT 91.835 62.275 92.005 62.445 ;
        RECT 92.305 62.310 92.465 62.420 ;
        RECT 93.220 62.255 93.390 62.445 ;
        RECT 94.135 62.275 94.305 62.445 ;
        RECT 94.595 62.275 94.765 62.445 ;
        RECT 95.980 62.275 96.150 62.465 ;
        RECT 99.205 62.300 99.365 62.410 ;
        RECT 100.580 62.255 100.750 62.445 ;
        RECT 102.875 62.275 103.045 62.445 ;
        RECT 103.335 62.275 103.505 62.445 ;
        RECT 104.715 62.275 104.885 62.465 ;
        RECT 106.560 62.255 106.730 62.445 ;
        RECT 108.395 62.275 108.565 62.465 ;
        RECT 108.855 62.275 109.025 62.465 ;
        RECT 112.530 62.305 112.650 62.415 ;
        RECT 113.455 62.275 113.625 62.445 ;
        RECT 114.840 62.275 115.010 62.465 ;
        RECT 118.050 62.255 118.220 62.445 ;
        RECT 118.520 62.255 118.690 62.445 ;
        RECT 120.820 62.275 120.990 62.465 ;
        RECT 124.495 62.275 124.665 62.445 ;
        RECT 126.340 62.255 126.510 62.445 ;
        RECT 127.715 62.275 127.885 62.445 ;
        RECT 129.095 62.275 129.265 62.445 ;
        RECT 130.475 62.275 130.645 62.445 ;
        RECT 130.945 62.310 131.105 62.420 ;
        RECT 131.860 62.275 132.030 62.465 ;
        RECT 132.320 62.255 132.490 62.445 ;
        RECT 137.845 62.310 138.005 62.420 ;
        RECT 138.300 62.255 138.470 62.445 ;
        RECT 140.135 62.275 140.305 62.445 ;
        RECT 140.595 62.275 140.765 62.465 ;
        RECT 142.430 62.305 142.550 62.415 ;
        RECT 142.900 62.275 143.070 62.465 ;
        RECT 144.280 62.255 144.450 62.445 ;
        RECT 148.875 62.275 149.045 62.465 ;
        RECT 150.255 62.255 150.425 62.445 ;
        RECT 152.095 62.255 152.265 62.445 ;
        RECT 154.395 62.275 154.565 62.465 ;
        RECT 156.695 62.255 156.865 62.465 ;
        RECT 22.695 61.445 24.065 62.255 ;
        RECT 24.535 61.575 30.505 62.255 ;
        RECT 30.515 61.575 36.485 62.255 ;
        RECT 36.495 61.575 42.465 62.255 ;
        RECT 42.475 61.575 48.445 62.255 ;
        RECT 28.720 61.345 30.505 61.575 ;
        RECT 34.700 61.345 36.485 61.575 ;
        RECT 40.680 61.345 42.465 61.575 ;
        RECT 46.660 61.345 48.445 61.575 ;
        RECT 48.465 61.385 48.895 62.170 ;
        RECT 53.975 61.575 59.945 62.255 ;
        RECT 59.955 61.575 65.925 62.255 ;
        RECT 67.775 61.575 73.745 62.255 ;
        RECT 58.160 61.345 59.945 61.575 ;
        RECT 64.140 61.345 65.925 61.575 ;
        RECT 71.960 61.345 73.745 61.575 ;
        RECT 74.225 61.385 74.655 62.170 ;
        RECT 75.135 61.575 81.105 62.255 ;
        RECT 81.115 61.575 87.085 62.255 ;
        RECT 87.095 61.575 93.065 62.255 ;
        RECT 93.075 61.575 99.045 62.255 ;
        RECT 79.320 61.345 81.105 61.575 ;
        RECT 85.300 61.345 87.085 61.575 ;
        RECT 91.280 61.345 93.065 61.575 ;
        RECT 97.260 61.345 99.045 61.575 ;
        RECT 99.985 61.385 100.415 62.170 ;
        RECT 100.435 61.575 106.405 62.255 ;
        RECT 106.415 61.575 112.385 62.255 ;
        RECT 104.620 61.345 106.405 61.575 ;
        RECT 110.600 61.345 112.385 61.575 ;
        RECT 112.395 61.575 118.365 62.255 ;
        RECT 118.375 61.575 124.345 62.255 ;
        RECT 112.395 61.345 114.180 61.575 ;
        RECT 122.560 61.345 124.345 61.575 ;
        RECT 125.745 61.385 126.175 62.170 ;
        RECT 126.195 61.575 132.165 62.255 ;
        RECT 132.175 61.575 138.145 62.255 ;
        RECT 138.155 61.575 144.125 62.255 ;
        RECT 144.135 61.575 150.105 62.255 ;
        RECT 130.380 61.345 132.165 61.575 ;
        RECT 136.360 61.345 138.145 61.575 ;
        RECT 142.340 61.345 144.125 61.575 ;
        RECT 148.320 61.345 150.105 61.575 ;
        RECT 150.115 61.445 151.485 62.255 ;
        RECT 151.505 61.385 151.935 62.170 ;
        RECT 151.955 61.445 155.625 62.255 ;
        RECT 155.635 61.445 157.005 62.255 ;
      LAYER nwell ;
        RECT 22.500 58.225 157.200 61.055 ;
      LAYER pwell ;
        RECT 22.695 57.025 24.065 57.835 ;
        RECT 28.720 57.705 30.505 57.935 ;
        RECT 24.535 57.025 30.505 57.705 ;
        RECT 32.355 57.025 34.185 57.835 ;
        RECT 35.585 57.110 36.015 57.895 ;
        RECT 40.220 57.705 42.005 57.935 ;
        RECT 46.200 57.705 47.985 57.935 ;
        RECT 36.035 57.025 42.005 57.705 ;
        RECT 42.015 57.025 47.985 57.705 ;
        RECT 48.465 57.110 48.895 57.895 ;
        RECT 53.560 57.705 55.345 57.935 ;
        RECT 59.540 57.705 61.325 57.935 ;
        RECT 49.375 57.025 55.345 57.705 ;
        RECT 55.355 57.025 61.325 57.705 ;
        RECT 61.345 57.110 61.775 57.895 ;
        RECT 63.175 57.025 65.925 57.835 ;
        RECT 70.120 57.705 71.905 57.935 ;
        RECT 65.935 57.025 71.905 57.705 ;
        RECT 74.225 57.110 74.655 57.895 ;
        RECT 74.675 57.025 76.045 57.835 ;
        RECT 79.735 57.025 81.105 57.835 ;
        RECT 85.300 57.705 87.085 57.935 ;
        RECT 81.115 57.025 87.085 57.705 ;
        RECT 87.105 57.110 87.535 57.895 ;
        RECT 88.935 57.025 90.305 57.835 ;
        RECT 94.500 57.705 96.285 57.935 ;
        RECT 90.315 57.025 96.285 57.705 ;
        RECT 96.295 57.025 97.665 57.835 ;
        RECT 99.985 57.110 100.415 57.895 ;
        RECT 105.080 57.705 106.865 57.935 ;
        RECT 100.895 57.025 106.865 57.705 ;
        RECT 106.875 57.025 108.245 57.835 ;
        RECT 112.865 57.110 113.295 57.895 ;
        RECT 117.500 57.705 119.285 57.935 ;
        RECT 113.315 57.025 119.285 57.705 ;
        RECT 119.295 57.705 121.080 57.935 ;
        RECT 119.295 57.025 125.265 57.705 ;
        RECT 125.745 57.110 126.175 57.895 ;
        RECT 130.380 57.705 132.165 57.935 ;
        RECT 126.195 57.025 132.165 57.705 ;
        RECT 136.315 57.025 138.145 57.835 ;
        RECT 138.625 57.110 139.055 57.895 ;
        RECT 143.260 57.705 145.045 57.935 ;
        RECT 139.075 57.025 145.045 57.705 ;
        RECT 147.815 57.025 151.485 57.835 ;
        RECT 151.505 57.110 151.935 57.895 ;
        RECT 151.955 57.025 155.625 57.835 ;
        RECT 155.635 57.025 157.005 57.835 ;
        RECT 22.835 56.835 23.005 57.025 ;
        RECT 24.210 56.865 24.330 56.975 ;
        RECT 24.680 56.835 24.850 57.025 ;
        RECT 30.650 56.865 30.770 56.975 ;
        RECT 32.035 56.835 32.205 57.005 ;
        RECT 32.495 56.835 32.665 57.025 ;
        RECT 34.335 56.835 34.505 57.005 ;
        RECT 36.180 56.835 36.350 57.025 ;
        RECT 42.160 56.835 42.330 57.025 ;
        RECT 48.130 56.865 48.250 56.975 ;
        RECT 49.050 56.865 49.170 56.975 ;
        RECT 49.520 56.835 49.690 57.025 ;
        RECT 55.500 56.835 55.670 57.025 ;
        RECT 62.855 56.835 63.025 57.005 ;
        RECT 63.315 56.835 63.485 57.025 ;
        RECT 66.080 56.835 66.250 57.025 ;
        RECT 72.065 56.870 72.225 56.980 ;
        RECT 73.895 56.835 74.065 57.005 ;
        RECT 74.815 56.835 74.985 57.025 ;
        RECT 77.115 56.835 77.285 57.005 ;
        RECT 77.585 56.870 77.745 56.980 ;
        RECT 79.415 56.835 79.585 57.005 ;
        RECT 79.875 56.835 80.045 57.025 ;
        RECT 81.260 56.835 81.430 57.025 ;
        RECT 88.615 56.835 88.785 57.005 ;
        RECT 89.075 56.835 89.245 57.025 ;
        RECT 90.460 56.835 90.630 57.025 ;
        RECT 96.435 56.835 96.605 57.025 ;
        RECT 97.815 56.835 97.985 57.005 ;
        RECT 99.205 56.870 99.365 56.980 ;
        RECT 100.570 56.865 100.690 56.975 ;
        RECT 101.040 56.835 101.210 57.025 ;
        RECT 107.015 56.835 107.185 57.025 ;
        RECT 108.395 56.835 108.565 57.005 ;
        RECT 109.770 56.865 109.890 56.975 ;
        RECT 110.235 56.835 110.405 57.005 ;
        RECT 111.615 56.835 111.785 57.005 ;
        RECT 113.460 56.835 113.630 57.025 ;
        RECT 124.950 56.835 125.120 57.025 ;
        RECT 125.410 56.865 125.530 56.975 ;
        RECT 126.340 56.835 126.510 57.025 ;
        RECT 133.235 56.835 133.405 57.005 ;
        RECT 134.615 56.835 134.785 57.005 ;
        RECT 135.075 56.835 135.245 57.005 ;
        RECT 136.455 56.835 136.625 57.025 ;
        RECT 138.290 56.865 138.410 56.975 ;
        RECT 139.220 56.835 139.390 57.025 ;
        RECT 146.115 56.835 146.285 57.005 ;
        RECT 147.495 56.835 147.665 57.005 ;
        RECT 147.955 56.835 148.125 57.025 ;
        RECT 152.095 56.835 152.265 57.025 ;
        RECT 156.695 56.835 156.865 57.025 ;
        RECT 32.820 33.660 35.780 47.760 ;
        RECT 39.820 37.910 42.780 38.760 ;
        RECT 43.520 37.910 46.480 38.310 ;
        RECT 39.820 36.460 46.480 37.910 ;
        RECT 39.820 33.660 42.780 36.460 ;
        RECT 43.520 34.090 46.480 36.460 ;
        RECT 32.980 29.260 33.280 29.860 ;
        RECT 34.820 22.680 37.780 33.260 ;
        RECT 46.530 32.150 50.130 35.110 ;
        RECT 50.230 28.700 53.330 35.110 ;
        RECT 74.040 34.500 77.000 48.600 ;
        RECT 81.040 38.750 84.000 39.600 ;
        RECT 84.740 38.750 87.700 39.150 ;
        RECT 81.040 37.300 87.700 38.750 ;
        RECT 81.040 34.500 84.000 37.300 ;
        RECT 84.740 34.930 87.700 37.300 ;
        RECT 74.200 30.100 74.500 30.700 ;
        RECT 49.800 25.310 53.880 28.410 ;
        RECT 50.350 24.860 53.420 25.310 ;
        RECT 36.320 14.160 39.280 22.260 ;
        RECT 49.970 21.760 54.930 24.860 ;
        RECT 76.040 23.520 79.000 34.100 ;
        RECT 87.750 32.990 91.350 35.950 ;
        RECT 91.450 29.540 94.550 35.950 ;
        RECT 113.920 35.900 116.880 50.000 ;
        RECT 120.920 40.150 123.880 41.000 ;
        RECT 124.620 40.150 127.580 40.550 ;
        RECT 120.920 38.700 127.580 40.150 ;
        RECT 120.920 35.900 123.880 38.700 ;
        RECT 124.620 36.330 127.580 38.700 ;
        RECT 114.080 31.500 114.380 32.100 ;
        RECT 91.020 26.150 95.100 29.250 ;
        RECT 91.570 25.700 94.640 26.150 ;
        RECT 50.350 21.280 53.420 21.760 ;
        RECT 49.940 18.180 56.140 21.280 ;
        RECT 50.350 17.700 53.420 18.180 ;
        RECT 49.810 14.600 57.770 17.700 ;
        RECT 77.540 15.000 80.500 23.100 ;
        RECT 91.190 22.600 96.150 25.700 ;
        RECT 115.920 24.920 118.880 35.500 ;
        RECT 127.630 34.390 131.230 37.350 ;
        RECT 131.330 30.940 134.430 37.350 ;
        RECT 130.900 27.550 134.980 30.650 ;
        RECT 131.450 27.100 134.520 27.550 ;
        RECT 91.570 22.120 94.640 22.600 ;
        RECT 91.160 19.020 97.360 22.120 ;
        RECT 91.570 18.540 94.640 19.020 ;
        RECT 91.030 15.440 98.990 18.540 ;
        RECT 117.420 16.400 120.380 24.500 ;
        RECT 131.070 24.000 136.030 27.100 ;
        RECT 131.450 23.520 134.520 24.000 ;
        RECT 131.040 20.420 137.240 23.520 ;
        RECT 131.450 19.940 134.520 20.420 ;
        RECT 130.910 16.840 138.870 19.940 ;
        RECT 131.450 16.360 134.520 16.840 ;
        RECT 91.570 14.960 94.640 15.440 ;
        RECT 50.350 14.120 53.420 14.600 ;
        RECT 38.320 7.420 41.280 13.760 ;
        RECT 49.830 11.020 60.270 14.120 ;
        RECT 50.350 10.540 53.420 11.020 ;
        RECT 49.840 7.440 63.800 10.540 ;
        RECT 79.540 8.260 82.500 14.600 ;
        RECT 91.050 11.860 101.490 14.960 ;
        RECT 91.570 11.380 94.640 11.860 ;
        RECT 91.060 8.280 105.020 11.380 ;
        RECT 119.420 9.660 122.380 16.000 ;
        RECT 130.930 13.260 141.370 16.360 ;
        RECT 131.450 12.780 134.520 13.260 ;
        RECT 130.940 9.680 144.900 12.780 ;
      LAYER li1 ;
        RECT 22.690 209.155 157.010 209.325 ;
        RECT 22.775 208.405 23.985 209.155 ;
        RECT 24.325 208.640 24.495 209.155 ;
        RECT 24.665 208.500 24.995 208.935 ;
        RECT 25.165 208.545 25.335 209.155 ;
        RECT 24.615 208.415 24.995 208.500 ;
        RECT 25.505 208.415 25.835 208.940 ;
        RECT 26.095 208.625 26.305 209.155 ;
        RECT 26.580 208.705 27.365 208.875 ;
        RECT 27.535 208.705 27.940 208.875 ;
        RECT 22.775 207.865 23.295 208.405 ;
        RECT 24.615 208.375 24.840 208.415 ;
        RECT 23.465 207.695 23.985 208.235 ;
        RECT 22.775 206.605 23.985 207.695 ;
        RECT 24.615 207.795 24.785 208.375 ;
        RECT 25.505 208.245 25.705 208.415 ;
        RECT 26.580 208.245 26.750 208.705 ;
        RECT 24.955 207.915 25.705 208.245 ;
        RECT 25.875 207.915 26.750 208.245 ;
        RECT 24.615 207.745 24.830 207.795 ;
        RECT 24.615 207.665 25.005 207.745 ;
        RECT 24.335 206.605 24.505 207.520 ;
        RECT 24.675 206.820 25.005 207.665 ;
        RECT 25.515 207.710 25.705 207.915 ;
        RECT 25.175 206.605 25.345 207.615 ;
        RECT 25.515 207.335 26.410 207.710 ;
        RECT 25.515 206.775 25.855 207.335 ;
        RECT 26.085 206.605 26.400 207.105 ;
        RECT 26.580 207.075 26.750 207.915 ;
        RECT 26.920 208.205 27.385 208.535 ;
        RECT 27.770 208.475 27.940 208.705 ;
        RECT 28.120 208.655 28.490 209.155 ;
        RECT 28.810 208.705 29.485 208.875 ;
        RECT 29.680 208.705 30.015 208.875 ;
        RECT 26.920 207.245 27.240 208.205 ;
        RECT 27.770 208.175 28.600 208.475 ;
        RECT 27.410 207.275 27.600 207.995 ;
        RECT 27.770 207.105 27.940 208.175 ;
        RECT 28.400 208.145 28.600 208.175 ;
        RECT 28.110 207.925 28.280 207.995 ;
        RECT 28.810 207.925 28.980 208.705 ;
        RECT 29.845 208.565 30.015 208.705 ;
        RECT 30.185 208.695 30.435 209.155 ;
        RECT 28.110 207.755 28.980 207.925 ;
        RECT 29.150 208.285 29.675 208.505 ;
        RECT 29.845 208.435 30.070 208.565 ;
        RECT 28.110 207.665 28.620 207.755 ;
        RECT 26.580 206.905 27.465 207.075 ;
        RECT 27.690 206.775 27.940 207.105 ;
        RECT 28.110 206.605 28.280 207.405 ;
        RECT 28.450 207.050 28.620 207.665 ;
        RECT 29.150 207.585 29.320 208.285 ;
        RECT 28.790 207.220 29.320 207.585 ;
        RECT 29.490 207.520 29.730 208.115 ;
        RECT 29.900 207.330 30.070 208.435 ;
        RECT 30.240 207.575 30.520 208.525 ;
        RECT 29.765 207.200 30.070 207.330 ;
        RECT 28.450 206.880 29.555 207.050 ;
        RECT 29.765 206.775 30.015 207.200 ;
        RECT 30.185 206.605 30.450 207.065 ;
        RECT 30.690 206.775 30.875 208.895 ;
        RECT 31.045 208.775 31.375 209.155 ;
        RECT 31.545 208.605 31.715 208.895 ;
        RECT 31.050 208.435 31.715 208.605 ;
        RECT 31.050 207.445 31.280 208.435 ;
        RECT 31.975 208.385 35.485 209.155 ;
        RECT 35.655 208.430 35.945 209.155 ;
        RECT 36.115 208.385 37.785 209.155 ;
        RECT 38.415 208.480 38.675 208.985 ;
        RECT 38.855 208.775 39.185 209.155 ;
        RECT 39.365 208.605 39.535 208.985 ;
        RECT 39.795 208.610 45.140 209.155 ;
        RECT 31.450 207.615 31.800 208.265 ;
        RECT 31.975 207.865 33.625 208.385 ;
        RECT 33.795 207.695 35.485 208.215 ;
        RECT 36.115 207.865 36.865 208.385 ;
        RECT 31.050 207.275 31.715 207.445 ;
        RECT 31.045 206.605 31.375 207.105 ;
        RECT 31.545 206.775 31.715 207.275 ;
        RECT 31.975 206.605 35.485 207.695 ;
        RECT 35.655 206.605 35.945 207.770 ;
        RECT 37.035 207.695 37.785 208.215 ;
        RECT 36.115 206.605 37.785 207.695 ;
        RECT 38.415 207.680 38.585 208.480 ;
        RECT 38.870 208.435 39.535 208.605 ;
        RECT 38.870 208.180 39.040 208.435 ;
        RECT 38.755 207.850 39.040 208.180 ;
        RECT 39.275 207.885 39.605 208.255 ;
        RECT 38.870 207.705 39.040 207.850 ;
        RECT 41.380 207.780 41.720 208.610 ;
        RECT 45.315 208.385 47.905 209.155 ;
        RECT 48.535 208.430 48.825 209.155 ;
        RECT 49.455 208.480 49.715 208.985 ;
        RECT 49.895 208.775 50.225 209.155 ;
        RECT 50.405 208.605 50.575 208.985 ;
        RECT 50.835 208.610 56.180 209.155 ;
        RECT 38.415 206.775 38.685 207.680 ;
        RECT 38.870 207.535 39.535 207.705 ;
        RECT 38.855 206.605 39.185 207.365 ;
        RECT 39.365 206.775 39.535 207.535 ;
        RECT 43.200 207.040 43.550 208.290 ;
        RECT 45.315 207.865 46.525 208.385 ;
        RECT 46.695 207.695 47.905 208.215 ;
        RECT 39.795 206.605 45.140 207.040 ;
        RECT 45.315 206.605 47.905 207.695 ;
        RECT 48.535 206.605 48.825 207.770 ;
        RECT 49.455 207.680 49.625 208.480 ;
        RECT 49.910 208.435 50.575 208.605 ;
        RECT 49.910 208.180 50.080 208.435 ;
        RECT 49.795 207.850 50.080 208.180 ;
        RECT 50.315 207.885 50.645 208.255 ;
        RECT 49.910 207.705 50.080 207.850 ;
        RECT 52.420 207.780 52.760 208.610 ;
        RECT 56.815 208.480 57.075 208.985 ;
        RECT 57.255 208.775 57.585 209.155 ;
        RECT 57.765 208.605 57.935 208.985 ;
        RECT 49.455 206.775 49.725 207.680 ;
        RECT 49.910 207.535 50.575 207.705 ;
        RECT 49.895 206.605 50.225 207.365 ;
        RECT 50.405 206.775 50.575 207.535 ;
        RECT 54.240 207.040 54.590 208.290 ;
        RECT 56.815 207.680 56.985 208.480 ;
        RECT 57.270 208.435 57.935 208.605 ;
        RECT 57.270 208.180 57.440 208.435 ;
        RECT 58.195 208.385 60.785 209.155 ;
        RECT 61.415 208.430 61.705 209.155 ;
        RECT 57.155 207.850 57.440 208.180 ;
        RECT 57.675 207.885 58.005 208.255 ;
        RECT 58.195 207.865 59.405 208.385 ;
        RECT 61.935 208.335 62.145 209.155 ;
        RECT 62.315 208.355 62.645 208.985 ;
        RECT 57.270 207.705 57.440 207.850 ;
        RECT 50.835 206.605 56.180 207.040 ;
        RECT 56.815 206.775 57.085 207.680 ;
        RECT 57.270 207.535 57.935 207.705 ;
        RECT 59.575 207.695 60.785 208.215 ;
        RECT 57.255 206.605 57.585 207.365 ;
        RECT 57.765 206.775 57.935 207.535 ;
        RECT 58.195 206.605 60.785 207.695 ;
        RECT 61.415 206.605 61.705 207.770 ;
        RECT 62.315 207.755 62.565 208.355 ;
        RECT 62.815 208.335 63.045 209.155 ;
        RECT 64.265 208.605 64.435 208.985 ;
        RECT 64.615 208.775 64.945 209.155 ;
        RECT 64.265 208.435 64.930 208.605 ;
        RECT 65.125 208.480 65.385 208.985 ;
        RECT 62.735 207.915 63.065 208.165 ;
        RECT 64.195 207.885 64.535 208.255 ;
        RECT 64.760 208.180 64.930 208.435 ;
        RECT 64.760 207.850 65.035 208.180 ;
        RECT 61.935 206.605 62.145 207.745 ;
        RECT 62.315 206.775 62.645 207.755 ;
        RECT 62.815 206.605 63.045 207.745 ;
        RECT 64.760 207.705 64.930 207.850 ;
        RECT 64.255 207.535 64.930 207.705 ;
        RECT 65.205 207.680 65.385 208.480 ;
        RECT 65.555 208.385 67.225 209.155 ;
        RECT 67.400 208.390 67.855 209.155 ;
        RECT 68.130 208.775 69.430 208.985 ;
        RECT 69.685 208.795 70.015 209.155 ;
        RECT 69.260 208.625 69.430 208.775 ;
        RECT 70.185 208.655 70.445 208.985 ;
        RECT 65.555 207.865 66.305 208.385 ;
        RECT 66.475 207.695 67.225 208.215 ;
        RECT 68.330 208.165 68.550 208.565 ;
        RECT 67.395 207.965 67.885 208.165 ;
        RECT 68.075 207.955 68.550 208.165 ;
        RECT 68.795 208.165 69.005 208.565 ;
        RECT 69.260 208.500 70.015 208.625 ;
        RECT 69.260 208.455 70.105 208.500 ;
        RECT 69.835 208.335 70.105 208.455 ;
        RECT 68.795 207.955 69.125 208.165 ;
        RECT 69.295 207.895 69.705 208.200 ;
        RECT 64.255 206.775 64.435 207.535 ;
        RECT 64.615 206.605 64.945 207.365 ;
        RECT 65.115 206.775 65.385 207.680 ;
        RECT 65.555 206.605 67.225 207.695 ;
        RECT 67.400 207.725 68.575 207.785 ;
        RECT 69.935 207.760 70.105 208.335 ;
        RECT 69.905 207.725 70.105 207.760 ;
        RECT 67.400 207.615 70.105 207.725 ;
        RECT 67.400 206.995 67.655 207.615 ;
        RECT 68.245 207.555 70.045 207.615 ;
        RECT 68.245 207.525 68.575 207.555 ;
        RECT 70.275 207.455 70.445 208.655 ;
        RECT 67.905 207.355 68.090 207.445 ;
        RECT 68.680 207.355 69.515 207.365 ;
        RECT 67.905 207.155 69.515 207.355 ;
        RECT 67.905 207.115 68.135 207.155 ;
        RECT 67.400 206.775 67.735 206.995 ;
        RECT 68.740 206.605 69.095 206.985 ;
        RECT 69.265 206.775 69.515 207.155 ;
        RECT 69.765 206.605 70.015 207.385 ;
        RECT 70.185 206.775 70.445 207.455 ;
        RECT 70.615 208.415 71.000 208.985 ;
        RECT 71.170 208.695 71.495 209.155 ;
        RECT 72.015 208.525 72.295 208.985 ;
        RECT 70.615 207.745 70.895 208.415 ;
        RECT 71.170 208.355 72.295 208.525 ;
        RECT 71.170 208.245 71.620 208.355 ;
        RECT 71.065 207.915 71.620 208.245 ;
        RECT 72.485 208.185 72.885 208.985 ;
        RECT 73.285 208.695 73.555 209.155 ;
        RECT 73.725 208.525 74.010 208.985 ;
        RECT 70.615 206.775 71.000 207.745 ;
        RECT 71.170 207.455 71.620 207.915 ;
        RECT 71.790 207.625 72.885 208.185 ;
        RECT 71.170 207.235 72.295 207.455 ;
        RECT 71.170 206.605 71.495 207.065 ;
        RECT 72.015 206.775 72.295 207.235 ;
        RECT 72.485 206.775 72.885 207.625 ;
        RECT 73.055 208.355 74.010 208.525 ;
        RECT 74.295 208.430 74.585 209.155 ;
        RECT 74.845 208.605 75.015 208.985 ;
        RECT 75.195 208.775 75.525 209.155 ;
        RECT 74.845 208.435 75.510 208.605 ;
        RECT 75.705 208.480 75.965 208.985 ;
        RECT 73.055 207.455 73.265 208.355 ;
        RECT 73.435 207.625 74.125 208.185 ;
        RECT 74.775 207.885 75.105 208.255 ;
        RECT 75.340 208.180 75.510 208.435 ;
        RECT 75.340 207.850 75.625 208.180 ;
        RECT 73.055 207.235 74.010 207.455 ;
        RECT 73.285 206.605 73.555 207.065 ;
        RECT 73.725 206.775 74.010 207.235 ;
        RECT 74.295 206.605 74.585 207.770 ;
        RECT 75.340 207.705 75.510 207.850 ;
        RECT 74.845 207.535 75.510 207.705 ;
        RECT 75.795 207.680 75.965 208.480 ;
        RECT 74.845 206.775 75.015 207.535 ;
        RECT 75.195 206.605 75.525 207.365 ;
        RECT 75.695 206.775 75.965 207.680 ;
        RECT 76.135 208.415 76.520 208.985 ;
        RECT 76.690 208.695 77.015 209.155 ;
        RECT 77.535 208.525 77.815 208.985 ;
        RECT 76.135 207.745 76.415 208.415 ;
        RECT 76.690 208.355 77.815 208.525 ;
        RECT 76.690 208.245 77.140 208.355 ;
        RECT 76.585 207.915 77.140 208.245 ;
        RECT 78.005 208.185 78.405 208.985 ;
        RECT 78.805 208.695 79.075 209.155 ;
        RECT 79.245 208.525 79.530 208.985 ;
        RECT 76.135 206.775 76.520 207.745 ;
        RECT 76.690 207.455 77.140 207.915 ;
        RECT 77.310 207.625 78.405 208.185 ;
        RECT 76.690 207.235 77.815 207.455 ;
        RECT 76.690 206.605 77.015 207.065 ;
        RECT 77.535 206.775 77.815 207.235 ;
        RECT 78.005 206.775 78.405 207.625 ;
        RECT 78.575 208.355 79.530 208.525 ;
        RECT 79.905 208.605 80.075 208.985 ;
        RECT 80.290 208.775 80.620 209.155 ;
        RECT 79.905 208.435 80.620 208.605 ;
        RECT 78.575 207.455 78.785 208.355 ;
        RECT 78.955 207.625 79.645 208.185 ;
        RECT 79.815 207.885 80.170 208.255 ;
        RECT 80.450 208.245 80.620 208.435 ;
        RECT 80.790 208.410 81.045 208.985 ;
        RECT 80.450 207.915 80.705 208.245 ;
        RECT 80.450 207.705 80.620 207.915 ;
        RECT 79.905 207.535 80.620 207.705 ;
        RECT 80.875 207.680 81.045 208.410 ;
        RECT 81.220 208.315 81.480 209.155 ;
        RECT 81.655 208.355 82.350 208.985 ;
        RECT 82.555 208.355 82.865 209.155 ;
        RECT 83.035 208.385 86.545 209.155 ;
        RECT 87.175 208.430 87.465 209.155 ;
        RECT 87.635 208.415 88.020 208.985 ;
        RECT 88.190 208.695 88.515 209.155 ;
        RECT 89.035 208.525 89.315 208.985 ;
        RECT 81.675 207.915 82.010 208.165 ;
        RECT 82.180 207.755 82.350 208.355 ;
        RECT 82.520 207.915 82.855 208.185 ;
        RECT 83.035 207.865 84.685 208.385 ;
        RECT 78.575 207.235 79.530 207.455 ;
        RECT 78.805 206.605 79.075 207.065 ;
        RECT 79.245 206.775 79.530 207.235 ;
        RECT 79.905 206.775 80.075 207.535 ;
        RECT 80.290 206.605 80.620 207.365 ;
        RECT 80.790 206.775 81.045 207.680 ;
        RECT 81.220 206.605 81.480 207.755 ;
        RECT 81.655 206.605 81.915 207.745 ;
        RECT 82.085 206.775 82.415 207.755 ;
        RECT 82.585 206.605 82.865 207.745 ;
        RECT 84.855 207.695 86.545 208.215 ;
        RECT 83.035 206.605 86.545 207.695 ;
        RECT 87.175 206.605 87.465 207.770 ;
        RECT 87.635 207.745 87.915 208.415 ;
        RECT 88.190 208.355 89.315 208.525 ;
        RECT 88.190 208.245 88.640 208.355 ;
        RECT 88.085 207.915 88.640 208.245 ;
        RECT 89.505 208.185 89.905 208.985 ;
        RECT 90.305 208.695 90.575 209.155 ;
        RECT 90.745 208.525 91.030 208.985 ;
        RECT 87.635 206.775 88.020 207.745 ;
        RECT 88.190 207.455 88.640 207.915 ;
        RECT 88.810 207.625 89.905 208.185 ;
        RECT 88.190 207.235 89.315 207.455 ;
        RECT 88.190 206.605 88.515 207.065 ;
        RECT 89.035 206.775 89.315 207.235 ;
        RECT 89.505 206.775 89.905 207.625 ;
        RECT 90.075 208.355 91.030 208.525 ;
        RECT 91.405 208.605 91.575 208.985 ;
        RECT 91.790 208.775 92.120 209.155 ;
        RECT 91.405 208.435 92.120 208.605 ;
        RECT 90.075 207.455 90.285 208.355 ;
        RECT 90.455 207.625 91.145 208.185 ;
        RECT 91.315 207.885 91.670 208.255 ;
        RECT 91.950 208.245 92.120 208.435 ;
        RECT 92.290 208.410 92.545 208.985 ;
        RECT 91.950 207.915 92.205 208.245 ;
        RECT 91.950 207.705 92.120 207.915 ;
        RECT 91.405 207.535 92.120 207.705 ;
        RECT 92.375 207.680 92.545 208.410 ;
        RECT 92.720 208.315 92.980 209.155 ;
        RECT 93.705 208.605 93.875 208.985 ;
        RECT 94.090 208.775 94.420 209.155 ;
        RECT 93.705 208.435 94.420 208.605 ;
        RECT 93.615 207.885 93.970 208.255 ;
        RECT 94.250 208.245 94.420 208.435 ;
        RECT 94.590 208.410 94.845 208.985 ;
        RECT 94.250 207.915 94.505 208.245 ;
        RECT 90.075 207.235 91.030 207.455 ;
        RECT 90.305 206.605 90.575 207.065 ;
        RECT 90.745 206.775 91.030 207.235 ;
        RECT 91.405 206.775 91.575 207.535 ;
        RECT 91.790 206.605 92.120 207.365 ;
        RECT 92.290 206.775 92.545 207.680 ;
        RECT 92.720 206.605 92.980 207.755 ;
        RECT 94.250 207.705 94.420 207.915 ;
        RECT 93.705 207.535 94.420 207.705 ;
        RECT 94.675 207.680 94.845 208.410 ;
        RECT 95.020 208.315 95.280 209.155 ;
        RECT 95.455 208.480 95.715 208.985 ;
        RECT 95.895 208.775 96.225 209.155 ;
        RECT 96.405 208.605 96.575 208.985 ;
        RECT 93.705 206.775 93.875 207.535 ;
        RECT 94.090 206.605 94.420 207.365 ;
        RECT 94.590 206.775 94.845 207.680 ;
        RECT 95.020 206.605 95.280 207.755 ;
        RECT 95.455 207.680 95.625 208.480 ;
        RECT 95.910 208.435 96.575 208.605 ;
        RECT 95.910 208.180 96.080 208.435 ;
        RECT 96.835 208.385 99.425 209.155 ;
        RECT 100.055 208.430 100.345 209.155 ;
        RECT 101.065 208.605 101.235 208.985 ;
        RECT 101.415 208.775 101.745 209.155 ;
        RECT 101.065 208.435 101.730 208.605 ;
        RECT 101.925 208.480 102.185 208.985 ;
        RECT 95.795 207.850 96.080 208.180 ;
        RECT 96.315 207.885 96.645 208.255 ;
        RECT 96.835 207.865 98.045 208.385 ;
        RECT 95.910 207.705 96.080 207.850 ;
        RECT 95.455 206.775 95.725 207.680 ;
        RECT 95.910 207.535 96.575 207.705 ;
        RECT 98.215 207.695 99.425 208.215 ;
        RECT 100.995 207.885 101.325 208.255 ;
        RECT 101.560 208.180 101.730 208.435 ;
        RECT 101.560 207.850 101.845 208.180 ;
        RECT 95.895 206.605 96.225 207.365 ;
        RECT 96.405 206.775 96.575 207.535 ;
        RECT 96.835 206.605 99.425 207.695 ;
        RECT 100.055 206.605 100.345 207.770 ;
        RECT 101.560 207.705 101.730 207.850 ;
        RECT 101.065 207.535 101.730 207.705 ;
        RECT 102.015 207.680 102.185 208.480 ;
        RECT 102.355 208.385 104.025 209.155 ;
        RECT 104.745 208.605 104.915 208.985 ;
        RECT 105.095 208.775 105.425 209.155 ;
        RECT 104.745 208.435 105.410 208.605 ;
        RECT 105.605 208.480 105.865 208.985 ;
        RECT 102.355 207.865 103.105 208.385 ;
        RECT 103.275 207.695 104.025 208.215 ;
        RECT 104.675 207.885 105.005 208.255 ;
        RECT 105.240 208.180 105.410 208.435 ;
        RECT 105.240 207.850 105.525 208.180 ;
        RECT 105.240 207.705 105.410 207.850 ;
        RECT 101.065 206.775 101.235 207.535 ;
        RECT 101.415 206.605 101.745 207.365 ;
        RECT 101.915 206.775 102.185 207.680 ;
        RECT 102.355 206.605 104.025 207.695 ;
        RECT 104.745 207.535 105.410 207.705 ;
        RECT 105.695 207.680 105.865 208.480 ;
        RECT 106.035 208.385 107.705 209.155 ;
        RECT 108.340 208.755 108.675 209.155 ;
        RECT 108.845 208.585 109.050 208.985 ;
        RECT 109.260 208.675 109.535 209.155 ;
        RECT 109.745 208.655 110.005 208.985 ;
        RECT 108.365 208.415 109.050 208.585 ;
        RECT 106.035 207.865 106.785 208.385 ;
        RECT 106.955 207.695 107.705 208.215 ;
        RECT 104.745 206.775 104.915 207.535 ;
        RECT 105.095 206.605 105.425 207.365 ;
        RECT 105.595 206.775 105.865 207.680 ;
        RECT 106.035 206.605 107.705 207.695 ;
        RECT 108.365 207.385 108.705 208.415 ;
        RECT 108.875 207.745 109.125 208.245 ;
        RECT 109.305 207.915 109.665 208.495 ;
        RECT 109.835 207.745 110.005 208.655 ;
        RECT 110.265 208.605 110.435 208.985 ;
        RECT 110.615 208.775 110.945 209.155 ;
        RECT 110.265 208.435 110.930 208.605 ;
        RECT 111.125 208.480 111.385 208.985 ;
        RECT 110.195 207.885 110.525 208.255 ;
        RECT 110.760 208.180 110.930 208.435 ;
        RECT 108.875 207.575 110.005 207.745 ;
        RECT 110.760 207.850 111.045 208.180 ;
        RECT 110.760 207.705 110.930 207.850 ;
        RECT 108.365 207.210 109.030 207.385 ;
        RECT 108.340 206.605 108.675 207.030 ;
        RECT 108.845 206.805 109.030 207.210 ;
        RECT 109.235 206.605 109.565 207.385 ;
        RECT 109.735 206.805 110.005 207.575 ;
        RECT 110.265 207.535 110.930 207.705 ;
        RECT 111.215 207.680 111.385 208.480 ;
        RECT 111.555 208.405 112.765 209.155 ;
        RECT 112.935 208.430 113.225 209.155 ;
        RECT 111.555 207.865 112.075 208.405 ;
        RECT 113.395 208.385 115.985 209.155 ;
        RECT 116.155 208.655 116.415 208.985 ;
        RECT 116.585 208.795 116.915 209.155 ;
        RECT 117.170 208.775 118.470 208.985 ;
        RECT 112.245 207.695 112.765 208.235 ;
        RECT 113.395 207.865 114.605 208.385 ;
        RECT 110.265 206.775 110.435 207.535 ;
        RECT 110.615 206.605 110.945 207.365 ;
        RECT 111.115 206.775 111.385 207.680 ;
        RECT 111.555 206.605 112.765 207.695 ;
        RECT 112.935 206.605 113.225 207.770 ;
        RECT 114.775 207.695 115.985 208.215 ;
        RECT 113.395 206.605 115.985 207.695 ;
        RECT 116.155 207.455 116.325 208.655 ;
        RECT 117.170 208.625 117.340 208.775 ;
        RECT 116.585 208.500 117.340 208.625 ;
        RECT 116.495 208.455 117.340 208.500 ;
        RECT 116.495 208.335 116.765 208.455 ;
        RECT 116.495 207.760 116.665 208.335 ;
        RECT 116.895 207.895 117.305 208.200 ;
        RECT 117.595 208.165 117.805 208.565 ;
        RECT 117.475 207.955 117.805 208.165 ;
        RECT 118.050 208.165 118.270 208.565 ;
        RECT 118.745 208.390 119.200 209.155 ;
        RECT 119.375 208.655 119.635 208.985 ;
        RECT 119.845 208.675 120.120 209.155 ;
        RECT 118.050 207.955 118.525 208.165 ;
        RECT 118.715 207.965 119.205 208.165 ;
        RECT 116.495 207.725 116.695 207.760 ;
        RECT 118.025 207.725 119.200 207.785 ;
        RECT 116.495 207.615 119.200 207.725 ;
        RECT 116.555 207.555 118.355 207.615 ;
        RECT 118.025 207.525 118.355 207.555 ;
        RECT 116.155 206.775 116.415 207.455 ;
        RECT 116.585 206.605 116.835 207.385 ;
        RECT 117.085 207.355 117.920 207.365 ;
        RECT 118.510 207.355 118.695 207.445 ;
        RECT 117.085 207.155 118.695 207.355 ;
        RECT 117.085 206.775 117.335 207.155 ;
        RECT 118.465 207.115 118.695 207.155 ;
        RECT 118.945 206.995 119.200 207.615 ;
        RECT 117.505 206.605 117.860 206.985 ;
        RECT 118.865 206.775 119.200 206.995 ;
        RECT 119.375 207.745 119.545 208.655 ;
        RECT 120.330 208.585 120.535 208.985 ;
        RECT 120.705 208.755 121.040 209.155 ;
        RECT 119.715 207.915 120.075 208.495 ;
        RECT 120.330 208.415 121.015 208.585 ;
        RECT 120.255 207.745 120.505 208.245 ;
        RECT 119.375 207.575 120.505 207.745 ;
        RECT 119.375 206.805 119.645 207.575 ;
        RECT 120.675 207.385 121.015 208.415 ;
        RECT 119.815 206.605 120.145 207.385 ;
        RECT 120.350 207.210 121.015 207.385 ;
        RECT 121.215 208.415 121.600 208.985 ;
        RECT 121.770 208.695 122.095 209.155 ;
        RECT 122.615 208.525 122.895 208.985 ;
        RECT 121.215 207.745 121.495 208.415 ;
        RECT 121.770 208.355 122.895 208.525 ;
        RECT 121.770 208.245 122.220 208.355 ;
        RECT 121.665 207.915 122.220 208.245 ;
        RECT 123.085 208.185 123.485 208.985 ;
        RECT 123.885 208.695 124.155 209.155 ;
        RECT 124.325 208.525 124.610 208.985 ;
        RECT 120.350 206.805 120.535 207.210 ;
        RECT 120.705 206.605 121.040 207.030 ;
        RECT 121.215 206.775 121.600 207.745 ;
        RECT 121.770 207.455 122.220 207.915 ;
        RECT 122.390 207.625 123.485 208.185 ;
        RECT 121.770 207.235 122.895 207.455 ;
        RECT 121.770 206.605 122.095 207.065 ;
        RECT 122.615 206.775 122.895 207.235 ;
        RECT 123.085 206.775 123.485 207.625 ;
        RECT 123.655 208.355 124.610 208.525 ;
        RECT 125.815 208.430 126.105 209.155 ;
        RECT 123.655 207.455 123.865 208.355 ;
        RECT 126.280 208.315 126.540 209.155 ;
        RECT 126.715 208.410 126.970 208.985 ;
        RECT 127.140 208.775 127.470 209.155 ;
        RECT 127.685 208.605 127.855 208.985 ;
        RECT 127.140 208.435 127.855 208.605 ;
        RECT 128.230 208.525 128.515 208.985 ;
        RECT 128.685 208.695 128.955 209.155 ;
        RECT 124.035 207.625 124.725 208.185 ;
        RECT 123.655 207.235 124.610 207.455 ;
        RECT 123.885 206.605 124.155 207.065 ;
        RECT 124.325 206.775 124.610 207.235 ;
        RECT 125.815 206.605 126.105 207.770 ;
        RECT 126.280 206.605 126.540 207.755 ;
        RECT 126.715 207.680 126.885 208.410 ;
        RECT 127.140 208.245 127.310 208.435 ;
        RECT 128.230 208.355 129.185 208.525 ;
        RECT 127.055 207.915 127.310 208.245 ;
        RECT 127.140 207.705 127.310 207.915 ;
        RECT 127.590 207.885 127.945 208.255 ;
        RECT 126.715 206.775 126.970 207.680 ;
        RECT 127.140 207.535 127.855 207.705 ;
        RECT 128.115 207.625 128.805 208.185 ;
        RECT 127.140 206.605 127.470 207.365 ;
        RECT 127.685 206.775 127.855 207.535 ;
        RECT 128.975 207.455 129.185 208.355 ;
        RECT 128.230 207.235 129.185 207.455 ;
        RECT 129.355 208.185 129.755 208.985 ;
        RECT 129.945 208.525 130.225 208.985 ;
        RECT 130.745 208.695 131.070 209.155 ;
        RECT 129.945 208.355 131.070 208.525 ;
        RECT 131.240 208.415 131.625 208.985 ;
        RECT 130.620 208.245 131.070 208.355 ;
        RECT 129.355 207.625 130.450 208.185 ;
        RECT 130.620 207.915 131.175 208.245 ;
        RECT 128.230 206.775 128.515 207.235 ;
        RECT 128.685 206.605 128.955 207.065 ;
        RECT 129.355 206.775 129.755 207.625 ;
        RECT 130.620 207.455 131.070 207.915 ;
        RECT 131.345 207.745 131.625 208.415 ;
        RECT 131.910 208.525 132.195 208.985 ;
        RECT 132.365 208.695 132.635 209.155 ;
        RECT 131.910 208.355 132.865 208.525 ;
        RECT 129.945 207.235 131.070 207.455 ;
        RECT 129.945 206.775 130.225 207.235 ;
        RECT 130.745 206.605 131.070 207.065 ;
        RECT 131.240 206.775 131.625 207.745 ;
        RECT 131.795 207.625 132.485 208.185 ;
        RECT 132.655 207.455 132.865 208.355 ;
        RECT 131.910 207.235 132.865 207.455 ;
        RECT 133.035 208.185 133.435 208.985 ;
        RECT 133.625 208.525 133.905 208.985 ;
        RECT 134.425 208.695 134.750 209.155 ;
        RECT 133.625 208.355 134.750 208.525 ;
        RECT 134.920 208.415 135.305 208.985 ;
        RECT 134.300 208.245 134.750 208.355 ;
        RECT 133.035 207.625 134.130 208.185 ;
        RECT 134.300 207.915 134.855 208.245 ;
        RECT 131.910 206.775 132.195 207.235 ;
        RECT 132.365 206.605 132.635 207.065 ;
        RECT 133.035 206.775 133.435 207.625 ;
        RECT 134.300 207.455 134.750 207.915 ;
        RECT 135.025 207.745 135.305 208.415 ;
        RECT 133.625 207.235 134.750 207.455 ;
        RECT 133.625 206.775 133.905 207.235 ;
        RECT 134.425 206.605 134.750 207.065 ;
        RECT 134.920 206.775 135.305 207.745 ;
        RECT 135.475 208.655 135.735 208.985 ;
        RECT 135.905 208.795 136.235 209.155 ;
        RECT 136.490 208.775 137.790 208.985 ;
        RECT 135.475 207.455 135.645 208.655 ;
        RECT 136.490 208.625 136.660 208.775 ;
        RECT 135.905 208.500 136.660 208.625 ;
        RECT 135.815 208.455 136.660 208.500 ;
        RECT 135.815 208.335 136.085 208.455 ;
        RECT 135.815 207.760 135.985 208.335 ;
        RECT 136.215 207.895 136.625 208.200 ;
        RECT 136.915 208.165 137.125 208.565 ;
        RECT 136.795 207.955 137.125 208.165 ;
        RECT 137.370 208.165 137.590 208.565 ;
        RECT 138.065 208.390 138.520 209.155 ;
        RECT 138.695 208.430 138.985 209.155 ;
        RECT 139.245 208.605 139.415 208.985 ;
        RECT 139.630 208.775 139.960 209.155 ;
        RECT 139.245 208.435 139.960 208.605 ;
        RECT 137.370 207.955 137.845 208.165 ;
        RECT 138.035 207.965 138.525 208.165 ;
        RECT 139.155 207.885 139.510 208.255 ;
        RECT 139.790 208.245 139.960 208.435 ;
        RECT 140.130 208.410 140.385 208.985 ;
        RECT 139.790 207.915 140.045 208.245 ;
        RECT 135.815 207.725 136.015 207.760 ;
        RECT 137.345 207.725 138.520 207.785 ;
        RECT 135.815 207.615 138.520 207.725 ;
        RECT 135.875 207.555 137.675 207.615 ;
        RECT 137.345 207.525 137.675 207.555 ;
        RECT 135.475 206.775 135.735 207.455 ;
        RECT 135.905 206.605 136.155 207.385 ;
        RECT 136.405 207.355 137.240 207.365 ;
        RECT 137.830 207.355 138.015 207.445 ;
        RECT 136.405 207.155 138.015 207.355 ;
        RECT 136.405 206.775 136.655 207.155 ;
        RECT 137.785 207.115 138.015 207.155 ;
        RECT 138.265 206.995 138.520 207.615 ;
        RECT 136.825 206.605 137.180 206.985 ;
        RECT 138.185 206.775 138.520 206.995 ;
        RECT 138.695 206.605 138.985 207.770 ;
        RECT 139.790 207.705 139.960 207.915 ;
        RECT 139.245 207.535 139.960 207.705 ;
        RECT 140.215 207.680 140.385 208.410 ;
        RECT 140.560 208.315 140.820 209.155 ;
        RECT 140.995 208.610 146.340 209.155 ;
        RECT 142.580 207.780 142.920 208.610 ;
        RECT 146.515 208.385 150.025 209.155 ;
        RECT 150.195 208.405 151.405 209.155 ;
        RECT 151.575 208.430 151.865 209.155 ;
        RECT 152.495 208.480 152.755 208.985 ;
        RECT 152.935 208.775 153.265 209.155 ;
        RECT 153.445 208.605 153.615 208.985 ;
        RECT 139.245 206.775 139.415 207.535 ;
        RECT 139.630 206.605 139.960 207.365 ;
        RECT 140.130 206.775 140.385 207.680 ;
        RECT 140.560 206.605 140.820 207.755 ;
        RECT 144.400 207.040 144.750 208.290 ;
        RECT 146.515 207.865 148.165 208.385 ;
        RECT 148.335 207.695 150.025 208.215 ;
        RECT 150.195 207.865 150.715 208.405 ;
        RECT 150.885 207.695 151.405 208.235 ;
        RECT 140.995 206.605 146.340 207.040 ;
        RECT 146.515 206.605 150.025 207.695 ;
        RECT 150.195 206.605 151.405 207.695 ;
        RECT 151.575 206.605 151.865 207.770 ;
        RECT 152.495 207.680 152.675 208.480 ;
        RECT 152.950 208.435 153.615 208.605 ;
        RECT 152.950 208.180 153.120 208.435 ;
        RECT 153.875 208.385 155.545 209.155 ;
        RECT 155.715 208.405 156.925 209.155 ;
        RECT 152.845 207.850 153.120 208.180 ;
        RECT 153.345 207.885 153.685 208.255 ;
        RECT 153.875 207.865 154.625 208.385 ;
        RECT 152.950 207.705 153.120 207.850 ;
        RECT 152.495 206.775 152.765 207.680 ;
        RECT 152.950 207.535 153.625 207.705 ;
        RECT 154.795 207.695 155.545 208.215 ;
        RECT 152.935 206.605 153.265 207.365 ;
        RECT 153.445 206.775 153.625 207.535 ;
        RECT 153.875 206.605 155.545 207.695 ;
        RECT 155.715 207.695 156.235 208.235 ;
        RECT 156.405 207.865 156.925 208.405 ;
        RECT 155.715 206.605 156.925 207.695 ;
        RECT 22.690 206.435 157.010 206.605 ;
        RECT 22.775 205.345 23.985 206.435 ;
        RECT 24.155 205.345 27.665 206.435 ;
        RECT 27.925 205.765 28.095 206.265 ;
        RECT 28.265 205.935 28.595 206.435 ;
        RECT 27.925 205.595 28.590 205.765 ;
        RECT 22.775 204.635 23.295 205.175 ;
        RECT 23.465 204.805 23.985 205.345 ;
        RECT 24.155 204.655 25.805 205.175 ;
        RECT 25.975 204.825 27.665 205.345 ;
        RECT 27.840 204.775 28.190 205.425 ;
        RECT 22.775 203.885 23.985 204.635 ;
        RECT 24.155 203.885 27.665 204.655 ;
        RECT 28.360 204.605 28.590 205.595 ;
        RECT 27.925 204.435 28.590 204.605 ;
        RECT 27.925 204.145 28.095 204.435 ;
        RECT 28.265 203.885 28.595 204.265 ;
        RECT 28.765 204.145 28.950 206.265 ;
        RECT 29.190 205.975 29.455 206.435 ;
        RECT 29.625 205.840 29.875 206.265 ;
        RECT 30.085 205.990 31.190 206.160 ;
        RECT 29.570 205.710 29.875 205.840 ;
        RECT 29.120 204.515 29.400 205.465 ;
        RECT 29.570 204.605 29.740 205.710 ;
        RECT 29.910 204.925 30.150 205.520 ;
        RECT 30.320 205.455 30.850 205.820 ;
        RECT 30.320 204.755 30.490 205.455 ;
        RECT 31.020 205.375 31.190 205.990 ;
        RECT 31.360 205.635 31.530 206.435 ;
        RECT 31.700 205.935 31.950 206.265 ;
        RECT 32.175 205.965 33.060 206.135 ;
        RECT 31.020 205.285 31.530 205.375 ;
        RECT 29.570 204.475 29.795 204.605 ;
        RECT 29.965 204.535 30.490 204.755 ;
        RECT 30.660 205.115 31.530 205.285 ;
        RECT 29.205 203.885 29.455 204.345 ;
        RECT 29.625 204.335 29.795 204.475 ;
        RECT 30.660 204.335 30.830 205.115 ;
        RECT 31.360 205.045 31.530 205.115 ;
        RECT 31.040 204.865 31.240 204.895 ;
        RECT 31.700 204.865 31.870 205.935 ;
        RECT 32.040 205.045 32.230 205.765 ;
        RECT 31.040 204.565 31.870 204.865 ;
        RECT 32.400 204.835 32.720 205.795 ;
        RECT 29.625 204.165 29.960 204.335 ;
        RECT 30.155 204.165 30.830 204.335 ;
        RECT 31.150 203.885 31.520 204.385 ;
        RECT 31.700 204.335 31.870 204.565 ;
        RECT 32.255 204.505 32.720 204.835 ;
        RECT 32.890 205.125 33.060 205.965 ;
        RECT 33.240 205.935 33.555 206.435 ;
        RECT 33.785 205.705 34.125 206.265 ;
        RECT 33.230 205.330 34.125 205.705 ;
        RECT 34.295 205.425 34.465 206.435 ;
        RECT 33.935 205.125 34.125 205.330 ;
        RECT 34.635 205.375 34.965 206.220 ;
        RECT 35.135 205.520 35.305 206.435 ;
        RECT 34.635 205.295 35.025 205.375 ;
        RECT 34.810 205.245 35.025 205.295 ;
        RECT 35.655 205.270 35.945 206.435 ;
        RECT 36.665 205.765 36.835 206.265 ;
        RECT 37.005 205.935 37.335 206.435 ;
        RECT 36.665 205.595 37.330 205.765 ;
        RECT 32.890 204.795 33.765 205.125 ;
        RECT 33.935 204.795 34.685 205.125 ;
        RECT 32.890 204.335 33.060 204.795 ;
        RECT 33.935 204.625 34.135 204.795 ;
        RECT 34.855 204.665 35.025 205.245 ;
        RECT 36.580 204.775 36.930 205.425 ;
        RECT 34.800 204.625 35.025 204.665 ;
        RECT 31.700 204.165 32.105 204.335 ;
        RECT 32.275 204.165 33.060 204.335 ;
        RECT 33.335 203.885 33.545 204.415 ;
        RECT 33.805 204.100 34.135 204.625 ;
        RECT 34.645 204.540 35.025 204.625 ;
        RECT 34.305 203.885 34.475 204.495 ;
        RECT 34.645 204.105 34.975 204.540 ;
        RECT 35.145 203.885 35.315 204.400 ;
        RECT 35.655 203.885 35.945 204.610 ;
        RECT 37.100 204.605 37.330 205.595 ;
        RECT 36.665 204.435 37.330 204.605 ;
        RECT 36.665 204.145 36.835 204.435 ;
        RECT 37.005 203.885 37.335 204.265 ;
        RECT 37.505 204.145 37.690 206.265 ;
        RECT 37.930 205.975 38.195 206.435 ;
        RECT 38.365 205.840 38.615 206.265 ;
        RECT 38.825 205.990 39.930 206.160 ;
        RECT 38.310 205.710 38.615 205.840 ;
        RECT 37.860 204.515 38.140 205.465 ;
        RECT 38.310 204.605 38.480 205.710 ;
        RECT 38.650 204.925 38.890 205.520 ;
        RECT 39.060 205.455 39.590 205.820 ;
        RECT 39.060 204.755 39.230 205.455 ;
        RECT 39.760 205.375 39.930 205.990 ;
        RECT 40.100 205.635 40.270 206.435 ;
        RECT 40.440 205.935 40.690 206.265 ;
        RECT 40.915 205.965 41.800 206.135 ;
        RECT 39.760 205.285 40.270 205.375 ;
        RECT 38.310 204.475 38.535 204.605 ;
        RECT 38.705 204.535 39.230 204.755 ;
        RECT 39.400 205.115 40.270 205.285 ;
        RECT 37.945 203.885 38.195 204.345 ;
        RECT 38.365 204.335 38.535 204.475 ;
        RECT 39.400 204.335 39.570 205.115 ;
        RECT 40.100 205.045 40.270 205.115 ;
        RECT 39.780 204.865 39.980 204.895 ;
        RECT 40.440 204.865 40.610 205.935 ;
        RECT 40.780 205.045 40.970 205.765 ;
        RECT 39.780 204.565 40.610 204.865 ;
        RECT 41.140 204.835 41.460 205.795 ;
        RECT 38.365 204.165 38.700 204.335 ;
        RECT 38.895 204.165 39.570 204.335 ;
        RECT 39.890 203.885 40.260 204.385 ;
        RECT 40.440 204.335 40.610 204.565 ;
        RECT 40.995 204.505 41.460 204.835 ;
        RECT 41.630 205.125 41.800 205.965 ;
        RECT 41.980 205.935 42.295 206.435 ;
        RECT 42.525 205.705 42.865 206.265 ;
        RECT 41.970 205.330 42.865 205.705 ;
        RECT 43.035 205.425 43.205 206.435 ;
        RECT 42.675 205.125 42.865 205.330 ;
        RECT 43.375 205.375 43.705 206.220 ;
        RECT 44.025 205.815 44.195 206.245 ;
        RECT 44.365 205.985 44.695 206.435 ;
        RECT 44.025 205.585 44.700 205.815 ;
        RECT 43.375 205.295 43.765 205.375 ;
        RECT 43.550 205.245 43.765 205.295 ;
        RECT 41.630 204.795 42.505 205.125 ;
        RECT 42.675 204.795 43.425 205.125 ;
        RECT 41.630 204.335 41.800 204.795 ;
        RECT 42.675 204.625 42.875 204.795 ;
        RECT 43.595 204.665 43.765 205.245 ;
        RECT 43.540 204.625 43.765 204.665 ;
        RECT 40.440 204.165 40.845 204.335 ;
        RECT 41.015 204.165 41.800 204.335 ;
        RECT 42.075 203.885 42.285 204.415 ;
        RECT 42.545 204.100 42.875 204.625 ;
        RECT 43.385 204.540 43.765 204.625 ;
        RECT 43.995 204.565 44.295 205.415 ;
        RECT 44.465 204.935 44.700 205.585 ;
        RECT 44.870 205.275 45.155 206.220 ;
        RECT 45.335 205.965 46.020 206.435 ;
        RECT 45.330 205.445 46.025 205.755 ;
        RECT 46.200 205.380 46.505 206.165 ;
        RECT 44.870 205.125 45.730 205.275 ;
        RECT 44.870 205.105 46.155 205.125 ;
        RECT 44.465 204.605 45.000 204.935 ;
        RECT 45.170 204.745 46.155 205.105 ;
        RECT 43.045 203.885 43.215 204.495 ;
        RECT 43.385 204.105 43.715 204.540 ;
        RECT 44.465 204.455 44.685 204.605 ;
        RECT 43.940 203.885 44.275 204.390 ;
        RECT 44.445 204.080 44.685 204.455 ;
        RECT 45.170 204.410 45.340 204.745 ;
        RECT 46.330 204.575 46.505 205.380 ;
        RECT 44.965 204.215 45.340 204.410 ;
        RECT 44.965 204.070 45.135 204.215 ;
        RECT 45.700 203.885 46.095 204.380 ;
        RECT 46.265 204.055 46.505 204.575 ;
        RECT 46.695 205.295 46.965 206.265 ;
        RECT 47.175 205.635 47.455 206.435 ;
        RECT 47.635 205.885 48.830 206.215 ;
        RECT 47.960 205.465 48.380 205.715 ;
        RECT 47.135 205.295 48.380 205.465 ;
        RECT 46.695 204.560 46.865 205.295 ;
        RECT 47.135 205.125 47.305 205.295 ;
        RECT 48.605 205.125 48.775 205.685 ;
        RECT 49.025 205.295 49.280 206.435 ;
        RECT 49.545 205.505 49.715 206.265 ;
        RECT 49.895 205.675 50.225 206.435 ;
        RECT 49.545 205.335 50.210 205.505 ;
        RECT 50.395 205.360 50.665 206.265 ;
        RECT 50.925 205.765 51.095 206.265 ;
        RECT 51.265 205.935 51.595 206.435 ;
        RECT 50.925 205.595 51.590 205.765 ;
        RECT 50.040 205.190 50.210 205.335 ;
        RECT 47.075 204.795 47.305 205.125 ;
        RECT 48.035 204.795 48.775 205.125 ;
        RECT 48.945 204.875 49.280 205.125 ;
        RECT 47.135 204.625 47.305 204.795 ;
        RECT 48.525 204.705 48.775 204.795 ;
        RECT 49.475 204.785 49.805 205.155 ;
        RECT 50.040 204.860 50.325 205.190 ;
        RECT 46.695 204.215 46.965 204.560 ;
        RECT 47.135 204.455 47.875 204.625 ;
        RECT 48.525 204.535 49.260 204.705 ;
        RECT 50.040 204.605 50.210 204.860 ;
        RECT 47.155 203.885 47.535 204.285 ;
        RECT 47.705 204.105 47.875 204.455 ;
        RECT 48.045 203.885 48.780 204.365 ;
        RECT 48.950 204.065 49.260 204.535 ;
        RECT 49.545 204.435 50.210 204.605 ;
        RECT 50.495 204.560 50.665 205.360 ;
        RECT 50.840 204.775 51.190 205.425 ;
        RECT 51.360 204.605 51.590 205.595 ;
        RECT 49.545 204.055 49.715 204.435 ;
        RECT 49.895 203.885 50.225 204.265 ;
        RECT 50.405 204.055 50.665 204.560 ;
        RECT 50.925 204.435 51.590 204.605 ;
        RECT 50.925 204.145 51.095 204.435 ;
        RECT 51.265 203.885 51.595 204.265 ;
        RECT 51.765 204.145 51.950 206.265 ;
        RECT 52.190 205.975 52.455 206.435 ;
        RECT 52.625 205.840 52.875 206.265 ;
        RECT 53.085 205.990 54.190 206.160 ;
        RECT 52.570 205.710 52.875 205.840 ;
        RECT 52.120 204.515 52.400 205.465 ;
        RECT 52.570 204.605 52.740 205.710 ;
        RECT 52.910 204.925 53.150 205.520 ;
        RECT 53.320 205.455 53.850 205.820 ;
        RECT 53.320 204.755 53.490 205.455 ;
        RECT 54.020 205.375 54.190 205.990 ;
        RECT 54.360 205.635 54.530 206.435 ;
        RECT 54.700 205.935 54.950 206.265 ;
        RECT 55.175 205.965 56.060 206.135 ;
        RECT 54.020 205.285 54.530 205.375 ;
        RECT 52.570 204.475 52.795 204.605 ;
        RECT 52.965 204.535 53.490 204.755 ;
        RECT 53.660 205.115 54.530 205.285 ;
        RECT 52.205 203.885 52.455 204.345 ;
        RECT 52.625 204.335 52.795 204.475 ;
        RECT 53.660 204.335 53.830 205.115 ;
        RECT 54.360 205.045 54.530 205.115 ;
        RECT 54.040 204.865 54.240 204.895 ;
        RECT 54.700 204.865 54.870 205.935 ;
        RECT 55.040 205.045 55.230 205.765 ;
        RECT 54.040 204.565 54.870 204.865 ;
        RECT 55.400 204.835 55.720 205.795 ;
        RECT 52.625 204.165 52.960 204.335 ;
        RECT 53.155 204.165 53.830 204.335 ;
        RECT 54.150 203.885 54.520 204.385 ;
        RECT 54.700 204.335 54.870 204.565 ;
        RECT 55.255 204.505 55.720 204.835 ;
        RECT 55.890 205.125 56.060 205.965 ;
        RECT 56.240 205.935 56.555 206.435 ;
        RECT 56.785 205.705 57.125 206.265 ;
        RECT 56.230 205.330 57.125 205.705 ;
        RECT 57.295 205.425 57.465 206.435 ;
        RECT 56.935 205.125 57.125 205.330 ;
        RECT 57.635 205.375 57.965 206.220 ;
        RECT 58.215 205.380 58.520 206.165 ;
        RECT 58.700 205.965 59.385 206.435 ;
        RECT 58.695 205.445 59.390 205.755 ;
        RECT 57.635 205.295 58.025 205.375 ;
        RECT 57.810 205.245 58.025 205.295 ;
        RECT 55.890 204.795 56.765 205.125 ;
        RECT 56.935 204.795 57.685 205.125 ;
        RECT 55.890 204.335 56.060 204.795 ;
        RECT 56.935 204.625 57.135 204.795 ;
        RECT 57.855 204.665 58.025 205.245 ;
        RECT 57.800 204.625 58.025 204.665 ;
        RECT 54.700 204.165 55.105 204.335 ;
        RECT 55.275 204.165 56.060 204.335 ;
        RECT 56.335 203.885 56.545 204.415 ;
        RECT 56.805 204.100 57.135 204.625 ;
        RECT 57.645 204.540 58.025 204.625 ;
        RECT 58.215 204.575 58.390 205.380 ;
        RECT 59.565 205.275 59.850 206.220 ;
        RECT 60.025 205.985 60.355 206.435 ;
        RECT 60.525 205.815 60.695 206.245 ;
        RECT 58.990 205.125 59.850 205.275 ;
        RECT 58.565 205.105 59.850 205.125 ;
        RECT 60.020 205.585 60.695 205.815 ;
        RECT 58.565 204.745 59.550 205.105 ;
        RECT 60.020 204.935 60.255 205.585 ;
        RECT 57.305 203.885 57.475 204.495 ;
        RECT 57.645 204.105 57.975 204.540 ;
        RECT 58.215 204.055 58.455 204.575 ;
        RECT 59.380 204.410 59.550 204.745 ;
        RECT 59.720 204.605 60.255 204.935 ;
        RECT 60.035 204.455 60.255 204.605 ;
        RECT 60.425 204.565 60.725 205.415 ;
        RECT 61.415 205.270 61.705 206.435 ;
        RECT 62.855 205.375 63.185 206.220 ;
        RECT 63.355 205.425 63.525 206.435 ;
        RECT 63.695 205.705 64.035 206.265 ;
        RECT 64.265 205.935 64.580 206.435 ;
        RECT 64.760 205.965 65.645 206.135 ;
        RECT 62.795 205.295 63.185 205.375 ;
        RECT 63.695 205.330 64.590 205.705 ;
        RECT 62.795 205.245 63.010 205.295 ;
        RECT 62.795 204.665 62.965 205.245 ;
        RECT 63.695 205.125 63.885 205.330 ;
        RECT 64.760 205.125 64.930 205.965 ;
        RECT 65.870 205.935 66.120 206.265 ;
        RECT 63.135 204.795 63.885 205.125 ;
        RECT 64.055 204.795 64.930 205.125 ;
        RECT 62.795 204.625 63.020 204.665 ;
        RECT 63.685 204.625 63.885 204.795 ;
        RECT 58.625 203.885 59.020 204.380 ;
        RECT 59.380 204.215 59.755 204.410 ;
        RECT 59.585 204.070 59.755 204.215 ;
        RECT 60.035 204.080 60.275 204.455 ;
        RECT 60.445 203.885 60.780 204.390 ;
        RECT 61.415 203.885 61.705 204.610 ;
        RECT 62.795 204.540 63.175 204.625 ;
        RECT 62.845 204.105 63.175 204.540 ;
        RECT 63.345 203.885 63.515 204.495 ;
        RECT 63.685 204.100 64.015 204.625 ;
        RECT 64.275 203.885 64.485 204.415 ;
        RECT 64.760 204.335 64.930 204.795 ;
        RECT 65.100 204.835 65.420 205.795 ;
        RECT 65.590 205.045 65.780 205.765 ;
        RECT 65.950 204.865 66.120 205.935 ;
        RECT 66.290 205.635 66.460 206.435 ;
        RECT 66.630 205.990 67.735 206.160 ;
        RECT 66.630 205.375 66.800 205.990 ;
        RECT 67.945 205.840 68.195 206.265 ;
        RECT 68.365 205.975 68.630 206.435 ;
        RECT 66.970 205.455 67.500 205.820 ;
        RECT 67.945 205.710 68.250 205.840 ;
        RECT 66.290 205.285 66.800 205.375 ;
        RECT 66.290 205.115 67.160 205.285 ;
        RECT 66.290 205.045 66.460 205.115 ;
        RECT 66.580 204.865 66.780 204.895 ;
        RECT 65.100 204.505 65.565 204.835 ;
        RECT 65.950 204.565 66.780 204.865 ;
        RECT 65.950 204.335 66.120 204.565 ;
        RECT 64.760 204.165 65.545 204.335 ;
        RECT 65.715 204.165 66.120 204.335 ;
        RECT 66.300 203.885 66.670 204.385 ;
        RECT 66.990 204.335 67.160 205.115 ;
        RECT 67.330 204.755 67.500 205.455 ;
        RECT 67.670 204.925 67.910 205.520 ;
        RECT 67.330 204.535 67.855 204.755 ;
        RECT 68.080 204.605 68.250 205.710 ;
        RECT 68.025 204.475 68.250 204.605 ;
        RECT 68.420 204.515 68.700 205.465 ;
        RECT 68.025 204.335 68.195 204.475 ;
        RECT 66.990 204.165 67.665 204.335 ;
        RECT 67.860 204.165 68.195 204.335 ;
        RECT 68.365 203.885 68.615 204.345 ;
        RECT 68.870 204.145 69.055 206.265 ;
        RECT 69.225 205.935 69.555 206.435 ;
        RECT 69.725 205.765 69.895 206.265 ;
        RECT 69.230 205.595 69.895 205.765 ;
        RECT 69.230 204.605 69.460 205.595 ;
        RECT 69.630 204.775 69.980 205.425 ;
        RECT 70.675 205.375 71.005 206.220 ;
        RECT 71.175 205.425 71.345 206.435 ;
        RECT 71.515 205.705 71.855 206.265 ;
        RECT 72.085 205.935 72.400 206.435 ;
        RECT 72.580 205.965 73.465 206.135 ;
        RECT 70.615 205.295 71.005 205.375 ;
        RECT 71.515 205.330 72.410 205.705 ;
        RECT 70.615 205.245 70.830 205.295 ;
        RECT 70.615 204.665 70.785 205.245 ;
        RECT 71.515 205.125 71.705 205.330 ;
        RECT 72.580 205.125 72.750 205.965 ;
        RECT 73.690 205.935 73.940 206.265 ;
        RECT 70.955 204.795 71.705 205.125 ;
        RECT 71.875 204.795 72.750 205.125 ;
        RECT 70.615 204.625 70.840 204.665 ;
        RECT 71.505 204.625 71.705 204.795 ;
        RECT 69.230 204.435 69.895 204.605 ;
        RECT 70.615 204.540 70.995 204.625 ;
        RECT 69.225 203.885 69.555 204.265 ;
        RECT 69.725 204.145 69.895 204.435 ;
        RECT 70.665 204.105 70.995 204.540 ;
        RECT 71.165 203.885 71.335 204.495 ;
        RECT 71.505 204.100 71.835 204.625 ;
        RECT 72.095 203.885 72.305 204.415 ;
        RECT 72.580 204.335 72.750 204.795 ;
        RECT 72.920 204.835 73.240 205.795 ;
        RECT 73.410 205.045 73.600 205.765 ;
        RECT 73.770 204.865 73.940 205.935 ;
        RECT 74.110 205.635 74.280 206.435 ;
        RECT 74.450 205.990 75.555 206.160 ;
        RECT 74.450 205.375 74.620 205.990 ;
        RECT 75.765 205.840 76.015 206.265 ;
        RECT 76.185 205.975 76.450 206.435 ;
        RECT 74.790 205.455 75.320 205.820 ;
        RECT 75.765 205.710 76.070 205.840 ;
        RECT 74.110 205.285 74.620 205.375 ;
        RECT 74.110 205.115 74.980 205.285 ;
        RECT 74.110 205.045 74.280 205.115 ;
        RECT 74.400 204.865 74.600 204.895 ;
        RECT 72.920 204.505 73.385 204.835 ;
        RECT 73.770 204.565 74.600 204.865 ;
        RECT 73.770 204.335 73.940 204.565 ;
        RECT 72.580 204.165 73.365 204.335 ;
        RECT 73.535 204.165 73.940 204.335 ;
        RECT 74.120 203.885 74.490 204.385 ;
        RECT 74.810 204.335 74.980 205.115 ;
        RECT 75.150 204.755 75.320 205.455 ;
        RECT 75.490 204.925 75.730 205.520 ;
        RECT 75.150 204.535 75.675 204.755 ;
        RECT 75.900 204.605 76.070 205.710 ;
        RECT 75.845 204.475 76.070 204.605 ;
        RECT 76.240 204.515 76.520 205.465 ;
        RECT 75.845 204.335 76.015 204.475 ;
        RECT 74.810 204.165 75.485 204.335 ;
        RECT 75.680 204.165 76.015 204.335 ;
        RECT 76.185 203.885 76.435 204.345 ;
        RECT 76.690 204.145 76.875 206.265 ;
        RECT 77.045 205.935 77.375 206.435 ;
        RECT 77.545 205.765 77.715 206.265 ;
        RECT 77.050 205.595 77.715 205.765 ;
        RECT 78.065 205.765 78.235 206.265 ;
        RECT 78.405 205.935 78.735 206.435 ;
        RECT 78.065 205.595 78.730 205.765 ;
        RECT 77.050 204.605 77.280 205.595 ;
        RECT 77.450 204.775 77.800 205.425 ;
        RECT 77.980 204.775 78.330 205.425 ;
        RECT 78.500 204.605 78.730 205.595 ;
        RECT 77.050 204.435 77.715 204.605 ;
        RECT 77.045 203.885 77.375 204.265 ;
        RECT 77.545 204.145 77.715 204.435 ;
        RECT 78.065 204.435 78.730 204.605 ;
        RECT 78.065 204.145 78.235 204.435 ;
        RECT 78.405 203.885 78.735 204.265 ;
        RECT 78.905 204.145 79.090 206.265 ;
        RECT 79.330 205.975 79.595 206.435 ;
        RECT 79.765 205.840 80.015 206.265 ;
        RECT 80.225 205.990 81.330 206.160 ;
        RECT 79.710 205.710 80.015 205.840 ;
        RECT 79.260 204.515 79.540 205.465 ;
        RECT 79.710 204.605 79.880 205.710 ;
        RECT 80.050 204.925 80.290 205.520 ;
        RECT 80.460 205.455 80.990 205.820 ;
        RECT 80.460 204.755 80.630 205.455 ;
        RECT 81.160 205.375 81.330 205.990 ;
        RECT 81.500 205.635 81.670 206.435 ;
        RECT 81.840 205.935 82.090 206.265 ;
        RECT 82.315 205.965 83.200 206.135 ;
        RECT 81.160 205.285 81.670 205.375 ;
        RECT 79.710 204.475 79.935 204.605 ;
        RECT 80.105 204.535 80.630 204.755 ;
        RECT 80.800 205.115 81.670 205.285 ;
        RECT 79.345 203.885 79.595 204.345 ;
        RECT 79.765 204.335 79.935 204.475 ;
        RECT 80.800 204.335 80.970 205.115 ;
        RECT 81.500 205.045 81.670 205.115 ;
        RECT 81.180 204.865 81.380 204.895 ;
        RECT 81.840 204.865 82.010 205.935 ;
        RECT 82.180 205.045 82.370 205.765 ;
        RECT 81.180 204.565 82.010 204.865 ;
        RECT 82.540 204.835 82.860 205.795 ;
        RECT 79.765 204.165 80.100 204.335 ;
        RECT 80.295 204.165 80.970 204.335 ;
        RECT 81.290 203.885 81.660 204.385 ;
        RECT 81.840 204.335 82.010 204.565 ;
        RECT 82.395 204.505 82.860 204.835 ;
        RECT 83.030 205.125 83.200 205.965 ;
        RECT 83.380 205.935 83.695 206.435 ;
        RECT 83.925 205.705 84.265 206.265 ;
        RECT 83.370 205.330 84.265 205.705 ;
        RECT 84.435 205.425 84.605 206.435 ;
        RECT 84.075 205.125 84.265 205.330 ;
        RECT 84.775 205.375 85.105 206.220 ;
        RECT 84.775 205.295 85.165 205.375 ;
        RECT 85.335 205.295 85.615 206.435 ;
        RECT 84.950 205.245 85.165 205.295 ;
        RECT 85.785 205.285 86.115 206.265 ;
        RECT 86.285 205.295 86.545 206.435 ;
        RECT 83.030 204.795 83.905 205.125 ;
        RECT 84.075 204.795 84.825 205.125 ;
        RECT 83.030 204.335 83.200 204.795 ;
        RECT 84.075 204.625 84.275 204.795 ;
        RECT 84.995 204.665 85.165 205.245 ;
        RECT 85.345 204.855 85.680 205.125 ;
        RECT 85.850 204.685 86.020 205.285 ;
        RECT 87.175 205.270 87.465 206.435 ;
        RECT 87.635 205.345 88.845 206.435 ;
        RECT 89.105 205.765 89.275 206.265 ;
        RECT 89.445 205.935 89.775 206.435 ;
        RECT 89.105 205.595 89.770 205.765 ;
        RECT 86.190 204.875 86.525 205.125 ;
        RECT 84.940 204.625 85.165 204.665 ;
        RECT 81.840 204.165 82.245 204.335 ;
        RECT 82.415 204.165 83.200 204.335 ;
        RECT 83.475 203.885 83.685 204.415 ;
        RECT 83.945 204.100 84.275 204.625 ;
        RECT 84.785 204.540 85.165 204.625 ;
        RECT 84.445 203.885 84.615 204.495 ;
        RECT 84.785 204.105 85.115 204.540 ;
        RECT 85.335 203.885 85.645 204.685 ;
        RECT 85.850 204.055 86.545 204.685 ;
        RECT 87.635 204.635 88.155 205.175 ;
        RECT 88.325 204.805 88.845 205.345 ;
        RECT 89.020 204.775 89.370 205.425 ;
        RECT 87.175 203.885 87.465 204.610 ;
        RECT 87.635 203.885 88.845 204.635 ;
        RECT 89.540 204.605 89.770 205.595 ;
        RECT 89.105 204.435 89.770 204.605 ;
        RECT 89.105 204.145 89.275 204.435 ;
        RECT 89.445 203.885 89.775 204.265 ;
        RECT 89.945 204.145 90.130 206.265 ;
        RECT 90.370 205.975 90.635 206.435 ;
        RECT 90.805 205.840 91.055 206.265 ;
        RECT 91.265 205.990 92.370 206.160 ;
        RECT 90.750 205.710 91.055 205.840 ;
        RECT 90.300 204.515 90.580 205.465 ;
        RECT 90.750 204.605 90.920 205.710 ;
        RECT 91.090 204.925 91.330 205.520 ;
        RECT 91.500 205.455 92.030 205.820 ;
        RECT 91.500 204.755 91.670 205.455 ;
        RECT 92.200 205.375 92.370 205.990 ;
        RECT 92.540 205.635 92.710 206.435 ;
        RECT 92.880 205.935 93.130 206.265 ;
        RECT 93.355 205.965 94.240 206.135 ;
        RECT 92.200 205.285 92.710 205.375 ;
        RECT 90.750 204.475 90.975 204.605 ;
        RECT 91.145 204.535 91.670 204.755 ;
        RECT 91.840 205.115 92.710 205.285 ;
        RECT 90.385 203.885 90.635 204.345 ;
        RECT 90.805 204.335 90.975 204.475 ;
        RECT 91.840 204.335 92.010 205.115 ;
        RECT 92.540 205.045 92.710 205.115 ;
        RECT 92.220 204.865 92.420 204.895 ;
        RECT 92.880 204.865 93.050 205.935 ;
        RECT 93.220 205.045 93.410 205.765 ;
        RECT 92.220 204.565 93.050 204.865 ;
        RECT 93.580 204.835 93.900 205.795 ;
        RECT 90.805 204.165 91.140 204.335 ;
        RECT 91.335 204.165 92.010 204.335 ;
        RECT 92.330 203.885 92.700 204.385 ;
        RECT 92.880 204.335 93.050 204.565 ;
        RECT 93.435 204.505 93.900 204.835 ;
        RECT 94.070 205.125 94.240 205.965 ;
        RECT 94.420 205.935 94.735 206.435 ;
        RECT 94.965 205.705 95.305 206.265 ;
        RECT 94.410 205.330 95.305 205.705 ;
        RECT 95.475 205.425 95.645 206.435 ;
        RECT 95.115 205.125 95.305 205.330 ;
        RECT 95.815 205.375 96.145 206.220 ;
        RECT 95.815 205.295 96.205 205.375 ;
        RECT 96.435 205.295 96.645 206.435 ;
        RECT 95.990 205.245 96.205 205.295 ;
        RECT 94.070 204.795 94.945 205.125 ;
        RECT 95.115 204.795 95.865 205.125 ;
        RECT 94.070 204.335 94.240 204.795 ;
        RECT 95.115 204.625 95.315 204.795 ;
        RECT 96.035 204.665 96.205 205.245 ;
        RECT 96.815 205.285 97.145 206.265 ;
        RECT 97.315 205.295 97.545 206.435 ;
        RECT 98.675 205.295 98.950 206.265 ;
        RECT 99.160 205.635 99.440 206.435 ;
        RECT 99.610 205.925 101.225 206.255 ;
        RECT 99.610 205.585 100.785 205.755 ;
        RECT 99.610 205.465 99.780 205.585 ;
        RECT 99.120 205.295 99.780 205.465 ;
        RECT 95.980 204.625 96.205 204.665 ;
        RECT 92.880 204.165 93.285 204.335 ;
        RECT 93.455 204.165 94.240 204.335 ;
        RECT 94.515 203.885 94.725 204.415 ;
        RECT 94.985 204.100 95.315 204.625 ;
        RECT 95.825 204.540 96.205 204.625 ;
        RECT 95.485 203.885 95.655 204.495 ;
        RECT 95.825 204.105 96.155 204.540 ;
        RECT 96.435 203.885 96.645 204.705 ;
        RECT 96.815 204.685 97.065 205.285 ;
        RECT 97.235 204.875 97.565 205.125 ;
        RECT 96.815 204.055 97.145 204.685 ;
        RECT 97.315 203.885 97.545 204.705 ;
        RECT 98.675 204.560 98.845 205.295 ;
        RECT 99.120 205.125 99.290 205.295 ;
        RECT 100.040 205.125 100.285 205.415 ;
        RECT 100.455 205.295 100.785 205.585 ;
        RECT 101.045 205.125 101.215 205.685 ;
        RECT 101.465 205.295 101.725 206.435 ;
        RECT 101.905 205.455 102.235 206.265 ;
        RECT 102.405 205.635 102.645 206.435 ;
        RECT 101.905 205.285 102.620 205.455 ;
        RECT 99.015 204.795 99.290 205.125 ;
        RECT 99.460 204.795 100.285 205.125 ;
        RECT 100.500 204.795 101.215 205.125 ;
        RECT 101.385 204.875 101.720 205.125 ;
        RECT 101.900 204.875 102.280 205.115 ;
        RECT 102.450 205.045 102.620 205.285 ;
        RECT 102.825 205.415 102.995 206.265 ;
        RECT 103.165 205.635 103.495 206.435 ;
        RECT 103.665 205.415 103.835 206.265 ;
        RECT 102.825 205.245 103.835 205.415 ;
        RECT 104.005 205.285 104.335 206.435 ;
        RECT 105.175 205.375 105.505 206.220 ;
        RECT 105.675 205.425 105.845 206.435 ;
        RECT 106.015 205.705 106.355 206.265 ;
        RECT 106.585 205.935 106.900 206.435 ;
        RECT 107.080 205.965 107.965 206.135 ;
        RECT 105.115 205.295 105.505 205.375 ;
        RECT 106.015 205.330 106.910 205.705 ;
        RECT 102.450 204.875 102.950 205.045 ;
        RECT 99.120 204.625 99.290 204.795 ;
        RECT 100.965 204.705 101.215 204.795 ;
        RECT 102.450 204.705 102.620 204.875 ;
        RECT 103.340 204.735 103.835 205.245 ;
        RECT 103.335 204.705 103.835 204.735 ;
        RECT 98.675 204.215 98.950 204.560 ;
        RECT 99.120 204.455 100.785 204.625 ;
        RECT 99.140 203.885 99.515 204.285 ;
        RECT 99.685 204.105 99.855 204.455 ;
        RECT 100.025 203.885 100.355 204.285 ;
        RECT 100.525 204.055 100.785 204.455 ;
        RECT 100.965 204.285 101.295 204.705 ;
        RECT 101.465 203.885 101.725 204.705 ;
        RECT 101.985 204.535 102.620 204.705 ;
        RECT 102.825 204.535 103.835 204.705 ;
        RECT 105.115 205.245 105.330 205.295 ;
        RECT 101.985 204.055 102.155 204.535 ;
        RECT 102.335 203.885 102.575 204.365 ;
        RECT 102.825 204.055 102.995 204.535 ;
        RECT 103.165 203.885 103.495 204.365 ;
        RECT 103.665 204.055 103.835 204.535 ;
        RECT 104.005 203.885 104.335 204.685 ;
        RECT 105.115 204.665 105.285 205.245 ;
        RECT 106.015 205.125 106.205 205.330 ;
        RECT 107.080 205.125 107.250 205.965 ;
        RECT 108.190 205.935 108.440 206.265 ;
        RECT 105.455 204.795 106.205 205.125 ;
        RECT 106.375 204.795 107.250 205.125 ;
        RECT 105.115 204.625 105.340 204.665 ;
        RECT 106.005 204.625 106.205 204.795 ;
        RECT 105.115 204.540 105.495 204.625 ;
        RECT 105.165 204.105 105.495 204.540 ;
        RECT 105.665 203.885 105.835 204.495 ;
        RECT 106.005 204.100 106.335 204.625 ;
        RECT 106.595 203.885 106.805 204.415 ;
        RECT 107.080 204.335 107.250 204.795 ;
        RECT 107.420 204.835 107.740 205.795 ;
        RECT 107.910 205.045 108.100 205.765 ;
        RECT 108.270 204.865 108.440 205.935 ;
        RECT 108.610 205.635 108.780 206.435 ;
        RECT 108.950 205.990 110.055 206.160 ;
        RECT 108.950 205.375 109.120 205.990 ;
        RECT 110.265 205.840 110.515 206.265 ;
        RECT 110.685 205.975 110.950 206.435 ;
        RECT 109.290 205.455 109.820 205.820 ;
        RECT 110.265 205.710 110.570 205.840 ;
        RECT 108.610 205.285 109.120 205.375 ;
        RECT 108.610 205.115 109.480 205.285 ;
        RECT 108.610 205.045 108.780 205.115 ;
        RECT 108.900 204.865 109.100 204.895 ;
        RECT 107.420 204.505 107.885 204.835 ;
        RECT 108.270 204.565 109.100 204.865 ;
        RECT 108.270 204.335 108.440 204.565 ;
        RECT 107.080 204.165 107.865 204.335 ;
        RECT 108.035 204.165 108.440 204.335 ;
        RECT 108.620 203.885 108.990 204.385 ;
        RECT 109.310 204.335 109.480 205.115 ;
        RECT 109.650 204.755 109.820 205.455 ;
        RECT 109.990 204.925 110.230 205.520 ;
        RECT 109.650 204.535 110.175 204.755 ;
        RECT 110.400 204.605 110.570 205.710 ;
        RECT 110.345 204.475 110.570 204.605 ;
        RECT 110.740 204.515 111.020 205.465 ;
        RECT 110.345 204.335 110.515 204.475 ;
        RECT 109.310 204.165 109.985 204.335 ;
        RECT 110.180 204.165 110.515 204.335 ;
        RECT 110.685 203.885 110.935 204.345 ;
        RECT 111.190 204.145 111.375 206.265 ;
        RECT 111.545 205.935 111.875 206.435 ;
        RECT 112.045 205.765 112.215 206.265 ;
        RECT 111.550 205.595 112.215 205.765 ;
        RECT 111.550 204.605 111.780 205.595 ;
        RECT 111.950 204.775 112.300 205.425 ;
        RECT 112.935 205.270 113.225 206.435 ;
        RECT 113.395 205.345 115.985 206.435 ;
        RECT 116.705 205.765 116.875 206.265 ;
        RECT 117.045 205.935 117.375 206.435 ;
        RECT 116.705 205.595 117.370 205.765 ;
        RECT 113.395 204.655 114.605 205.175 ;
        RECT 114.775 204.825 115.985 205.345 ;
        RECT 116.620 204.775 116.970 205.425 ;
        RECT 111.550 204.435 112.215 204.605 ;
        RECT 111.545 203.885 111.875 204.265 ;
        RECT 112.045 204.145 112.215 204.435 ;
        RECT 112.935 203.885 113.225 204.610 ;
        RECT 113.395 203.885 115.985 204.655 ;
        RECT 117.140 204.605 117.370 205.595 ;
        RECT 116.705 204.435 117.370 204.605 ;
        RECT 116.705 204.145 116.875 204.435 ;
        RECT 117.045 203.885 117.375 204.265 ;
        RECT 117.545 204.145 117.730 206.265 ;
        RECT 117.970 205.975 118.235 206.435 ;
        RECT 118.405 205.840 118.655 206.265 ;
        RECT 118.865 205.990 119.970 206.160 ;
        RECT 118.350 205.710 118.655 205.840 ;
        RECT 117.900 204.515 118.180 205.465 ;
        RECT 118.350 204.605 118.520 205.710 ;
        RECT 118.690 204.925 118.930 205.520 ;
        RECT 119.100 205.455 119.630 205.820 ;
        RECT 119.100 204.755 119.270 205.455 ;
        RECT 119.800 205.375 119.970 205.990 ;
        RECT 120.140 205.635 120.310 206.435 ;
        RECT 120.480 205.935 120.730 206.265 ;
        RECT 120.955 205.965 121.840 206.135 ;
        RECT 119.800 205.285 120.310 205.375 ;
        RECT 118.350 204.475 118.575 204.605 ;
        RECT 118.745 204.535 119.270 204.755 ;
        RECT 119.440 205.115 120.310 205.285 ;
        RECT 117.985 203.885 118.235 204.345 ;
        RECT 118.405 204.335 118.575 204.475 ;
        RECT 119.440 204.335 119.610 205.115 ;
        RECT 120.140 205.045 120.310 205.115 ;
        RECT 119.820 204.865 120.020 204.895 ;
        RECT 120.480 204.865 120.650 205.935 ;
        RECT 120.820 205.045 121.010 205.765 ;
        RECT 119.820 204.565 120.650 204.865 ;
        RECT 121.180 204.835 121.500 205.795 ;
        RECT 118.405 204.165 118.740 204.335 ;
        RECT 118.935 204.165 119.610 204.335 ;
        RECT 119.930 203.885 120.300 204.385 ;
        RECT 120.480 204.335 120.650 204.565 ;
        RECT 121.035 204.505 121.500 204.835 ;
        RECT 121.670 205.125 121.840 205.965 ;
        RECT 122.020 205.935 122.335 206.435 ;
        RECT 122.565 205.705 122.905 206.265 ;
        RECT 122.010 205.330 122.905 205.705 ;
        RECT 123.075 205.425 123.245 206.435 ;
        RECT 122.715 205.125 122.905 205.330 ;
        RECT 123.415 205.375 123.745 206.220 ;
        RECT 124.065 205.505 124.235 206.265 ;
        RECT 124.450 205.675 124.780 206.435 ;
        RECT 123.415 205.295 123.805 205.375 ;
        RECT 124.065 205.335 124.780 205.505 ;
        RECT 124.950 205.360 125.205 206.265 ;
        RECT 123.590 205.245 123.805 205.295 ;
        RECT 121.670 204.795 122.545 205.125 ;
        RECT 122.715 204.795 123.465 205.125 ;
        RECT 121.670 204.335 121.840 204.795 ;
        RECT 122.715 204.625 122.915 204.795 ;
        RECT 123.635 204.665 123.805 205.245 ;
        RECT 123.975 204.785 124.330 205.155 ;
        RECT 124.610 205.125 124.780 205.335 ;
        RECT 124.610 204.795 124.865 205.125 ;
        RECT 123.580 204.625 123.805 204.665 ;
        RECT 120.480 204.165 120.885 204.335 ;
        RECT 121.055 204.165 121.840 204.335 ;
        RECT 122.115 203.885 122.325 204.415 ;
        RECT 122.585 204.100 122.915 204.625 ;
        RECT 123.425 204.540 123.805 204.625 ;
        RECT 124.610 204.605 124.780 204.795 ;
        RECT 125.035 204.630 125.205 205.360 ;
        RECT 125.380 205.285 125.640 206.435 ;
        RECT 126.365 205.765 126.535 206.265 ;
        RECT 126.705 205.935 127.035 206.435 ;
        RECT 126.365 205.595 127.030 205.765 ;
        RECT 126.280 204.775 126.630 205.425 ;
        RECT 123.085 203.885 123.255 204.495 ;
        RECT 123.425 204.105 123.755 204.540 ;
        RECT 124.065 204.435 124.780 204.605 ;
        RECT 124.065 204.055 124.235 204.435 ;
        RECT 124.450 203.885 124.780 204.265 ;
        RECT 124.950 204.055 125.205 204.630 ;
        RECT 125.380 203.885 125.640 204.725 ;
        RECT 126.800 204.605 127.030 205.595 ;
        RECT 126.365 204.435 127.030 204.605 ;
        RECT 126.365 204.145 126.535 204.435 ;
        RECT 126.705 203.885 127.035 204.265 ;
        RECT 127.205 204.145 127.390 206.265 ;
        RECT 127.630 205.975 127.895 206.435 ;
        RECT 128.065 205.840 128.315 206.265 ;
        RECT 128.525 205.990 129.630 206.160 ;
        RECT 128.010 205.710 128.315 205.840 ;
        RECT 127.560 204.515 127.840 205.465 ;
        RECT 128.010 204.605 128.180 205.710 ;
        RECT 128.350 204.925 128.590 205.520 ;
        RECT 128.760 205.455 129.290 205.820 ;
        RECT 128.760 204.755 128.930 205.455 ;
        RECT 129.460 205.375 129.630 205.990 ;
        RECT 129.800 205.635 129.970 206.435 ;
        RECT 130.140 205.935 130.390 206.265 ;
        RECT 130.615 205.965 131.500 206.135 ;
        RECT 129.460 205.285 129.970 205.375 ;
        RECT 128.010 204.475 128.235 204.605 ;
        RECT 128.405 204.535 128.930 204.755 ;
        RECT 129.100 205.115 129.970 205.285 ;
        RECT 127.645 203.885 127.895 204.345 ;
        RECT 128.065 204.335 128.235 204.475 ;
        RECT 129.100 204.335 129.270 205.115 ;
        RECT 129.800 205.045 129.970 205.115 ;
        RECT 129.480 204.865 129.680 204.895 ;
        RECT 130.140 204.865 130.310 205.935 ;
        RECT 130.480 205.045 130.670 205.765 ;
        RECT 129.480 204.565 130.310 204.865 ;
        RECT 130.840 204.835 131.160 205.795 ;
        RECT 128.065 204.165 128.400 204.335 ;
        RECT 128.595 204.165 129.270 204.335 ;
        RECT 129.590 203.885 129.960 204.385 ;
        RECT 130.140 204.335 130.310 204.565 ;
        RECT 130.695 204.505 131.160 204.835 ;
        RECT 131.330 205.125 131.500 205.965 ;
        RECT 131.680 205.935 131.995 206.435 ;
        RECT 132.225 205.705 132.565 206.265 ;
        RECT 131.670 205.330 132.565 205.705 ;
        RECT 132.735 205.425 132.905 206.435 ;
        RECT 132.375 205.125 132.565 205.330 ;
        RECT 133.075 205.375 133.405 206.220 ;
        RECT 133.635 205.585 133.895 206.265 ;
        RECT 134.065 205.655 134.315 206.435 ;
        RECT 134.565 205.885 134.815 206.265 ;
        RECT 134.985 206.055 135.340 206.435 ;
        RECT 136.345 206.045 136.680 206.265 ;
        RECT 135.945 205.885 136.175 205.925 ;
        RECT 134.565 205.685 136.175 205.885 ;
        RECT 134.565 205.675 135.400 205.685 ;
        RECT 135.990 205.595 136.175 205.685 ;
        RECT 133.075 205.295 133.465 205.375 ;
        RECT 133.250 205.245 133.465 205.295 ;
        RECT 131.330 204.795 132.205 205.125 ;
        RECT 132.375 204.795 133.125 205.125 ;
        RECT 131.330 204.335 131.500 204.795 ;
        RECT 132.375 204.625 132.575 204.795 ;
        RECT 133.295 204.665 133.465 205.245 ;
        RECT 133.240 204.625 133.465 204.665 ;
        RECT 130.140 204.165 130.545 204.335 ;
        RECT 130.715 204.165 131.500 204.335 ;
        RECT 131.775 203.885 131.985 204.415 ;
        RECT 132.245 204.100 132.575 204.625 ;
        RECT 133.085 204.540 133.465 204.625 ;
        RECT 132.745 203.885 132.915 204.495 ;
        RECT 133.085 204.105 133.415 204.540 ;
        RECT 133.635 204.395 133.805 205.585 ;
        RECT 135.505 205.485 135.835 205.515 ;
        RECT 134.035 205.425 135.835 205.485 ;
        RECT 136.425 205.425 136.680 206.045 ;
        RECT 133.975 205.315 136.680 205.425 ;
        RECT 133.975 205.280 134.175 205.315 ;
        RECT 133.975 204.705 134.145 205.280 ;
        RECT 135.505 205.255 136.680 205.315 ;
        RECT 136.895 205.295 137.125 206.435 ;
        RECT 137.295 205.285 137.625 206.265 ;
        RECT 137.795 205.295 138.005 206.435 ;
        RECT 134.375 204.840 134.785 205.145 ;
        RECT 134.955 204.875 135.285 205.085 ;
        RECT 133.975 204.585 134.245 204.705 ;
        RECT 133.975 204.540 134.820 204.585 ;
        RECT 134.065 204.415 134.820 204.540 ;
        RECT 135.075 204.475 135.285 204.875 ;
        RECT 135.530 204.875 136.005 205.085 ;
        RECT 136.195 204.875 136.685 205.075 ;
        RECT 136.875 204.875 137.205 205.125 ;
        RECT 135.530 204.475 135.750 204.875 ;
        RECT 133.635 204.385 133.865 204.395 ;
        RECT 133.635 204.055 133.895 204.385 ;
        RECT 134.650 204.265 134.820 204.415 ;
        RECT 134.065 203.885 134.395 204.245 ;
        RECT 134.650 204.055 135.950 204.265 ;
        RECT 136.225 203.885 136.680 204.650 ;
        RECT 136.895 203.885 137.125 204.705 ;
        RECT 137.375 204.685 137.625 205.285 ;
        RECT 138.695 205.270 138.985 206.435 ;
        RECT 139.155 206.005 139.495 206.265 ;
        RECT 137.295 204.055 137.625 204.685 ;
        RECT 137.795 203.885 138.005 204.705 ;
        RECT 138.695 203.885 138.985 204.610 ;
        RECT 139.155 204.605 139.415 206.005 ;
        RECT 139.665 205.635 139.995 206.435 ;
        RECT 140.460 205.465 140.710 206.265 ;
        RECT 140.895 205.715 141.225 206.435 ;
        RECT 141.445 205.465 141.695 206.265 ;
        RECT 141.865 206.055 142.200 206.435 ;
        RECT 139.605 205.295 141.795 205.465 ;
        RECT 139.605 205.125 139.920 205.295 ;
        RECT 139.590 204.875 139.920 205.125 ;
        RECT 139.155 204.095 139.495 204.605 ;
        RECT 139.665 203.885 139.935 204.685 ;
        RECT 140.115 204.155 140.395 205.125 ;
        RECT 140.575 204.155 140.875 205.125 ;
        RECT 141.055 204.160 141.405 205.125 ;
        RECT 141.625 204.385 141.795 205.295 ;
        RECT 141.965 204.565 142.205 205.875 ;
        RECT 142.375 205.295 142.655 206.435 ;
        RECT 142.825 205.285 143.155 206.265 ;
        RECT 143.325 205.295 143.585 206.435 ;
        RECT 143.815 205.295 144.025 206.435 ;
        RECT 144.195 205.285 144.525 206.265 ;
        RECT 144.695 205.295 144.925 206.435 ;
        RECT 145.135 206.000 150.480 206.435 ;
        RECT 142.890 205.245 143.065 205.285 ;
        RECT 142.385 204.855 142.720 205.125 ;
        RECT 142.890 204.685 143.060 205.245 ;
        RECT 143.230 204.875 143.565 205.125 ;
        RECT 141.625 204.055 142.120 204.385 ;
        RECT 142.375 203.885 142.685 204.685 ;
        RECT 142.890 204.055 143.585 204.685 ;
        RECT 143.815 203.885 144.025 204.705 ;
        RECT 144.195 204.685 144.445 205.285 ;
        RECT 144.615 204.875 144.945 205.125 ;
        RECT 144.195 204.055 144.525 204.685 ;
        RECT 144.695 203.885 144.925 204.705 ;
        RECT 146.720 204.430 147.060 205.260 ;
        RECT 148.540 204.750 148.890 206.000 ;
        RECT 150.655 205.345 154.165 206.435 ;
        RECT 154.335 205.345 155.545 206.435 ;
        RECT 150.655 204.655 152.305 205.175 ;
        RECT 152.475 204.825 154.165 205.345 ;
        RECT 145.135 203.885 150.480 204.430 ;
        RECT 150.655 203.885 154.165 204.655 ;
        RECT 154.335 204.635 154.855 205.175 ;
        RECT 155.025 204.805 155.545 205.345 ;
        RECT 155.715 205.345 156.925 206.435 ;
        RECT 155.715 204.805 156.235 205.345 ;
        RECT 156.405 204.635 156.925 205.175 ;
        RECT 154.335 203.885 155.545 204.635 ;
        RECT 155.715 203.885 156.925 204.635 ;
        RECT 22.690 203.715 157.010 203.885 ;
        RECT 22.775 202.965 23.985 203.715 ;
        RECT 24.155 203.170 29.500 203.715 ;
        RECT 22.775 202.425 23.295 202.965 ;
        RECT 23.465 202.255 23.985 202.795 ;
        RECT 25.740 202.340 26.080 203.170 ;
        RECT 29.765 203.165 29.935 203.455 ;
        RECT 30.105 203.335 30.435 203.715 ;
        RECT 29.765 202.995 30.430 203.165 ;
        RECT 22.775 201.165 23.985 202.255 ;
        RECT 27.560 201.600 27.910 202.850 ;
        RECT 29.680 202.175 30.030 202.825 ;
        RECT 30.200 202.005 30.430 202.995 ;
        RECT 29.765 201.835 30.430 202.005 ;
        RECT 24.155 201.165 29.500 201.600 ;
        RECT 29.765 201.335 29.935 201.835 ;
        RECT 30.105 201.165 30.435 201.665 ;
        RECT 30.605 201.335 30.790 203.455 ;
        RECT 31.045 203.255 31.295 203.715 ;
        RECT 31.465 203.265 31.800 203.435 ;
        RECT 31.995 203.265 32.670 203.435 ;
        RECT 31.465 203.125 31.635 203.265 ;
        RECT 30.960 202.135 31.240 203.085 ;
        RECT 31.410 202.995 31.635 203.125 ;
        RECT 31.410 201.890 31.580 202.995 ;
        RECT 31.805 202.845 32.330 203.065 ;
        RECT 31.750 202.080 31.990 202.675 ;
        RECT 32.160 202.145 32.330 202.845 ;
        RECT 32.500 202.485 32.670 203.265 ;
        RECT 32.990 203.215 33.360 203.715 ;
        RECT 33.540 203.265 33.945 203.435 ;
        RECT 34.115 203.265 34.900 203.435 ;
        RECT 33.540 203.035 33.710 203.265 ;
        RECT 32.880 202.735 33.710 203.035 ;
        RECT 34.095 202.765 34.560 203.095 ;
        RECT 32.880 202.705 33.080 202.735 ;
        RECT 33.200 202.485 33.370 202.555 ;
        RECT 32.500 202.315 33.370 202.485 ;
        RECT 32.860 202.225 33.370 202.315 ;
        RECT 31.410 201.760 31.715 201.890 ;
        RECT 32.160 201.780 32.690 202.145 ;
        RECT 31.030 201.165 31.295 201.625 ;
        RECT 31.465 201.335 31.715 201.760 ;
        RECT 32.860 201.610 33.030 202.225 ;
        RECT 31.925 201.440 33.030 201.610 ;
        RECT 33.200 201.165 33.370 201.965 ;
        RECT 33.540 201.665 33.710 202.735 ;
        RECT 33.880 201.835 34.070 202.555 ;
        RECT 34.240 201.805 34.560 202.765 ;
        RECT 34.730 202.805 34.900 203.265 ;
        RECT 35.175 203.185 35.385 203.715 ;
        RECT 35.645 202.975 35.975 203.500 ;
        RECT 36.145 203.105 36.315 203.715 ;
        RECT 36.485 203.060 36.815 203.495 ;
        RECT 36.985 203.200 37.155 203.715 ;
        RECT 36.485 202.975 36.865 203.060 ;
        RECT 35.775 202.805 35.975 202.975 ;
        RECT 36.640 202.935 36.865 202.975 ;
        RECT 34.730 202.475 35.605 202.805 ;
        RECT 35.775 202.475 36.525 202.805 ;
        RECT 33.540 201.335 33.790 201.665 ;
        RECT 34.730 201.635 34.900 202.475 ;
        RECT 35.775 202.270 35.965 202.475 ;
        RECT 36.695 202.355 36.865 202.935 ;
        RECT 37.495 202.895 37.755 203.715 ;
        RECT 37.925 202.895 38.255 203.315 ;
        RECT 38.435 203.230 39.225 203.495 ;
        RECT 38.005 202.805 38.255 202.895 ;
        RECT 36.650 202.305 36.865 202.355 ;
        RECT 35.070 201.895 35.965 202.270 ;
        RECT 36.475 202.225 36.865 202.305 ;
        RECT 34.015 201.465 34.900 201.635 ;
        RECT 35.080 201.165 35.395 201.665 ;
        RECT 35.625 201.335 35.965 201.895 ;
        RECT 36.135 201.165 36.305 202.175 ;
        RECT 36.475 201.380 36.805 202.225 ;
        RECT 36.975 201.165 37.145 202.080 ;
        RECT 37.495 201.845 37.835 202.725 ;
        RECT 38.005 202.555 38.800 202.805 ;
        RECT 37.495 201.165 37.755 201.675 ;
        RECT 38.005 201.335 38.175 202.555 ;
        RECT 38.970 202.375 39.225 203.230 ;
        RECT 39.395 203.075 39.595 203.495 ;
        RECT 39.785 203.255 40.115 203.715 ;
        RECT 39.395 202.555 39.805 203.075 ;
        RECT 40.285 203.065 40.545 203.545 ;
        RECT 39.975 202.375 40.205 202.805 ;
        RECT 38.415 202.205 40.205 202.375 ;
        RECT 38.415 201.840 38.665 202.205 ;
        RECT 38.835 201.845 39.165 202.035 ;
        RECT 39.385 201.910 40.100 202.205 ;
        RECT 40.375 202.035 40.545 203.065 ;
        RECT 41.175 202.915 41.485 203.715 ;
        RECT 41.690 202.915 42.385 203.545 ;
        RECT 42.720 203.205 42.960 203.715 ;
        RECT 43.140 203.205 43.420 203.535 ;
        RECT 43.650 203.205 43.865 203.715 ;
        RECT 41.185 202.475 41.520 202.745 ;
        RECT 41.690 202.355 41.860 202.915 ;
        RECT 42.030 202.475 42.365 202.725 ;
        RECT 42.615 202.475 42.970 203.035 ;
        RECT 41.690 202.315 41.865 202.355 ;
        RECT 38.835 201.670 39.030 201.845 ;
        RECT 38.415 201.165 39.030 201.670 ;
        RECT 39.200 201.335 39.675 201.675 ;
        RECT 39.845 201.165 40.060 201.710 ;
        RECT 40.270 201.335 40.545 202.035 ;
        RECT 41.175 201.165 41.455 202.305 ;
        RECT 41.625 201.335 41.955 202.315 ;
        RECT 43.140 202.305 43.310 203.205 ;
        RECT 43.480 202.475 43.745 203.035 ;
        RECT 44.035 202.975 44.650 203.545 ;
        RECT 43.995 202.305 44.165 202.805 ;
        RECT 42.125 201.165 42.385 202.305 ;
        RECT 42.740 202.135 44.165 202.305 ;
        RECT 42.740 201.960 43.130 202.135 ;
        RECT 43.615 201.165 43.945 201.965 ;
        RECT 44.335 201.955 44.650 202.975 ;
        RECT 44.115 201.335 44.650 201.955 ;
        RECT 44.855 202.975 45.320 203.520 ;
        RECT 44.855 202.015 45.025 202.975 ;
        RECT 45.825 202.895 45.995 203.715 ;
        RECT 46.165 203.065 46.495 203.545 ;
        RECT 46.665 203.325 47.015 203.715 ;
        RECT 47.185 203.145 47.415 203.545 ;
        RECT 46.905 203.065 47.415 203.145 ;
        RECT 46.165 202.975 47.415 203.065 ;
        RECT 47.585 202.975 47.905 203.455 ;
        RECT 48.535 202.990 48.825 203.715 ;
        RECT 49.195 203.085 49.525 203.445 ;
        RECT 50.145 203.255 50.395 203.715 ;
        RECT 50.565 203.255 51.125 203.545 ;
        RECT 46.165 202.895 47.075 202.975 ;
        RECT 45.195 202.355 45.440 202.805 ;
        RECT 45.700 202.525 46.395 202.725 ;
        RECT 46.565 202.555 47.165 202.725 ;
        RECT 46.565 202.355 46.735 202.555 ;
        RECT 47.395 202.385 47.565 202.805 ;
        RECT 45.195 202.185 46.735 202.355 ;
        RECT 46.905 202.215 47.565 202.385 ;
        RECT 46.905 202.015 47.075 202.215 ;
        RECT 47.735 202.045 47.905 202.975 ;
        RECT 49.195 202.895 50.585 203.085 ;
        RECT 50.415 202.805 50.585 202.895 ;
        RECT 49.010 202.475 49.685 202.725 ;
        RECT 49.905 202.475 50.245 202.725 ;
        RECT 50.415 202.475 50.705 202.805 ;
        RECT 44.855 201.845 47.075 202.015 ;
        RECT 47.245 201.845 47.905 202.045 ;
        RECT 44.855 201.165 45.155 201.675 ;
        RECT 45.325 201.335 45.655 201.845 ;
        RECT 47.245 201.675 47.415 201.845 ;
        RECT 45.825 201.165 46.455 201.675 ;
        RECT 47.035 201.505 47.415 201.675 ;
        RECT 47.585 201.165 47.885 201.675 ;
        RECT 48.535 201.165 48.825 202.330 ;
        RECT 49.010 202.115 49.275 202.475 ;
        RECT 50.415 202.225 50.585 202.475 ;
        RECT 49.645 202.055 50.585 202.225 ;
        RECT 49.195 201.165 49.475 201.835 ;
        RECT 49.645 201.505 49.945 202.055 ;
        RECT 50.875 201.885 51.125 203.255 ;
        RECT 51.295 202.945 53.885 203.715 ;
        RECT 54.060 202.975 54.395 203.715 ;
        RECT 51.295 202.425 52.505 202.945 ;
        RECT 54.565 202.805 54.780 203.500 ;
        RECT 54.970 202.975 55.320 203.500 ;
        RECT 55.490 202.975 56.185 203.545 ;
        RECT 55.115 202.805 55.320 202.975 ;
        RECT 52.675 202.255 53.885 202.775 ;
        RECT 54.080 202.475 54.365 202.805 ;
        RECT 54.565 202.475 54.945 202.805 ;
        RECT 55.115 202.475 55.425 202.805 ;
        RECT 55.595 202.305 55.765 202.975 ;
        RECT 56.375 202.905 56.625 203.715 ;
        RECT 56.795 203.075 57.125 203.495 ;
        RECT 57.295 203.245 57.985 203.715 ;
        RECT 58.155 203.325 59.325 203.545 ;
        RECT 59.540 203.245 59.710 203.715 ;
        RECT 59.915 203.325 61.085 203.545 ;
        RECT 58.555 203.075 58.905 203.155 ;
        RECT 60.335 203.075 60.665 203.155 ;
        RECT 56.795 202.935 60.665 203.075 ;
        RECT 56.875 202.895 60.665 202.935 ;
        RECT 60.835 202.895 61.085 203.325 ;
        RECT 61.255 202.895 61.425 203.715 ;
        RECT 62.395 202.895 62.605 203.715 ;
        RECT 62.775 202.915 63.105 203.545 ;
        RECT 50.145 201.165 50.475 201.885 ;
        RECT 50.665 201.335 51.125 201.885 ;
        RECT 51.295 201.165 53.885 202.255 ;
        RECT 54.055 201.165 54.315 202.305 ;
        RECT 54.485 202.135 55.765 202.305 ;
        RECT 55.945 202.135 56.185 202.805 ;
        RECT 56.360 202.185 56.690 202.725 ;
        RECT 54.485 201.335 54.815 202.135 ;
        RECT 54.985 201.165 55.155 201.965 ;
        RECT 55.355 201.335 55.685 202.135 ;
        RECT 55.885 201.165 56.165 201.965 ;
        RECT 56.360 201.505 56.705 202.005 ;
        RECT 56.875 201.675 57.125 202.895 ;
        RECT 57.775 202.355 58.310 202.725 ;
        RECT 58.480 202.525 59.035 202.725 ;
        RECT 59.205 202.355 59.535 202.725 ;
        RECT 57.295 202.015 57.545 202.305 ;
        RECT 57.775 202.185 59.535 202.355 ;
        RECT 59.705 202.355 60.035 202.725 ;
        RECT 60.255 202.525 60.750 202.725 ;
        RECT 60.920 202.525 61.705 202.725 ;
        RECT 60.920 202.355 61.090 202.525 ;
        RECT 59.705 202.185 61.090 202.355 ;
        RECT 61.260 202.015 61.465 202.345 ;
        RECT 62.775 202.315 63.025 202.915 ;
        RECT 63.275 202.895 63.505 203.715 ;
        RECT 63.830 203.085 64.115 203.545 ;
        RECT 64.285 203.255 64.555 203.715 ;
        RECT 63.830 202.915 64.785 203.085 ;
        RECT 63.195 202.475 63.525 202.725 ;
        RECT 57.295 201.845 59.285 202.015 ;
        RECT 57.295 201.505 57.545 201.845 ;
        RECT 58.195 201.675 58.445 201.845 ;
        RECT 59.035 201.675 59.285 201.845 ;
        RECT 59.495 201.845 61.465 202.015 ;
        RECT 56.360 201.335 57.545 201.505 ;
        RECT 57.775 201.505 58.025 201.675 ;
        RECT 58.615 201.505 58.865 201.675 ;
        RECT 59.495 201.505 59.745 201.845 ;
        RECT 57.775 201.335 59.745 201.505 ;
        RECT 59.955 201.165 60.205 201.675 ;
        RECT 60.375 201.335 60.625 201.845 ;
        RECT 60.795 201.165 61.045 201.675 ;
        RECT 61.260 201.335 61.465 201.845 ;
        RECT 62.395 201.165 62.605 202.305 ;
        RECT 62.775 201.335 63.105 202.315 ;
        RECT 63.275 201.165 63.505 202.305 ;
        RECT 63.715 202.185 64.405 202.745 ;
        RECT 64.575 202.015 64.785 202.915 ;
        RECT 63.830 201.795 64.785 202.015 ;
        RECT 64.955 202.745 65.355 203.545 ;
        RECT 65.545 203.085 65.825 203.545 ;
        RECT 66.345 203.255 66.670 203.715 ;
        RECT 65.545 202.915 66.670 203.085 ;
        RECT 66.840 202.975 67.225 203.545 ;
        RECT 66.220 202.805 66.670 202.915 ;
        RECT 64.955 202.185 66.050 202.745 ;
        RECT 66.220 202.475 66.775 202.805 ;
        RECT 63.830 201.335 64.115 201.795 ;
        RECT 64.285 201.165 64.555 201.625 ;
        RECT 64.955 201.335 65.355 202.185 ;
        RECT 66.220 202.015 66.670 202.475 ;
        RECT 66.945 202.305 67.225 202.975 ;
        RECT 67.455 202.895 67.665 203.715 ;
        RECT 67.835 202.915 68.165 203.545 ;
        RECT 67.835 202.315 68.085 202.915 ;
        RECT 68.335 202.895 68.565 203.715 ;
        RECT 68.775 202.965 69.985 203.715 ;
        RECT 68.255 202.475 68.585 202.725 ;
        RECT 68.775 202.425 69.295 202.965 ;
        RECT 70.160 202.950 70.615 203.715 ;
        RECT 70.890 203.335 72.190 203.545 ;
        RECT 72.445 203.355 72.775 203.715 ;
        RECT 72.020 203.185 72.190 203.335 ;
        RECT 72.945 203.215 73.205 203.545 ;
        RECT 65.545 201.795 66.670 202.015 ;
        RECT 65.545 201.335 65.825 201.795 ;
        RECT 66.345 201.165 66.670 201.625 ;
        RECT 66.840 201.335 67.225 202.305 ;
        RECT 67.455 201.165 67.665 202.305 ;
        RECT 67.835 201.335 68.165 202.315 ;
        RECT 68.335 201.165 68.565 202.305 ;
        RECT 69.465 202.255 69.985 202.795 ;
        RECT 71.090 202.725 71.310 203.125 ;
        RECT 70.155 202.525 70.645 202.725 ;
        RECT 70.835 202.515 71.310 202.725 ;
        RECT 71.555 202.725 71.765 203.125 ;
        RECT 72.020 203.060 72.775 203.185 ;
        RECT 72.020 203.015 72.865 203.060 ;
        RECT 72.595 202.895 72.865 203.015 ;
        RECT 71.555 202.515 71.885 202.725 ;
        RECT 72.055 202.455 72.465 202.760 ;
        RECT 68.775 201.165 69.985 202.255 ;
        RECT 70.160 202.285 71.335 202.345 ;
        RECT 72.695 202.320 72.865 202.895 ;
        RECT 72.665 202.285 72.865 202.320 ;
        RECT 70.160 202.175 72.865 202.285 ;
        RECT 70.160 201.555 70.415 202.175 ;
        RECT 71.005 202.115 72.805 202.175 ;
        RECT 71.005 202.085 71.335 202.115 ;
        RECT 73.035 202.015 73.205 203.215 ;
        RECT 74.295 202.990 74.585 203.715 ;
        RECT 74.845 203.165 75.015 203.455 ;
        RECT 75.185 203.335 75.515 203.715 ;
        RECT 74.845 202.995 75.510 203.165 ;
        RECT 70.665 201.915 70.850 202.005 ;
        RECT 71.440 201.915 72.275 201.925 ;
        RECT 70.665 201.715 72.275 201.915 ;
        RECT 70.665 201.675 70.895 201.715 ;
        RECT 70.160 201.335 70.495 201.555 ;
        RECT 71.500 201.165 71.855 201.545 ;
        RECT 72.025 201.335 72.275 201.715 ;
        RECT 72.525 201.165 72.775 201.945 ;
        RECT 72.945 201.335 73.205 202.015 ;
        RECT 74.295 201.165 74.585 202.330 ;
        RECT 74.760 202.175 75.110 202.825 ;
        RECT 75.280 202.005 75.510 202.995 ;
        RECT 74.845 201.835 75.510 202.005 ;
        RECT 74.845 201.335 75.015 201.835 ;
        RECT 75.185 201.165 75.515 201.665 ;
        RECT 75.685 201.335 75.870 203.455 ;
        RECT 76.125 203.255 76.375 203.715 ;
        RECT 76.545 203.265 76.880 203.435 ;
        RECT 77.075 203.265 77.750 203.435 ;
        RECT 76.545 203.125 76.715 203.265 ;
        RECT 76.040 202.135 76.320 203.085 ;
        RECT 76.490 202.995 76.715 203.125 ;
        RECT 76.490 201.890 76.660 202.995 ;
        RECT 76.885 202.845 77.410 203.065 ;
        RECT 76.830 202.080 77.070 202.675 ;
        RECT 77.240 202.145 77.410 202.845 ;
        RECT 77.580 202.485 77.750 203.265 ;
        RECT 78.070 203.215 78.440 203.715 ;
        RECT 78.620 203.265 79.025 203.435 ;
        RECT 79.195 203.265 79.980 203.435 ;
        RECT 78.620 203.035 78.790 203.265 ;
        RECT 77.960 202.735 78.790 203.035 ;
        RECT 79.175 202.765 79.640 203.095 ;
        RECT 77.960 202.705 78.160 202.735 ;
        RECT 78.280 202.485 78.450 202.555 ;
        RECT 77.580 202.315 78.450 202.485 ;
        RECT 77.940 202.225 78.450 202.315 ;
        RECT 76.490 201.760 76.795 201.890 ;
        RECT 77.240 201.780 77.770 202.145 ;
        RECT 76.110 201.165 76.375 201.625 ;
        RECT 76.545 201.335 76.795 201.760 ;
        RECT 77.940 201.610 78.110 202.225 ;
        RECT 77.005 201.440 78.110 201.610 ;
        RECT 78.280 201.165 78.450 201.965 ;
        RECT 78.620 201.665 78.790 202.735 ;
        RECT 78.960 201.835 79.150 202.555 ;
        RECT 79.320 201.805 79.640 202.765 ;
        RECT 79.810 202.805 79.980 203.265 ;
        RECT 80.255 203.185 80.465 203.715 ;
        RECT 80.725 202.975 81.055 203.500 ;
        RECT 81.225 203.105 81.395 203.715 ;
        RECT 81.565 203.060 81.895 203.495 ;
        RECT 82.125 203.335 82.455 203.715 ;
        RECT 82.625 203.215 82.835 203.545 ;
        RECT 83.125 203.215 83.345 203.545 ;
        RECT 81.565 202.975 81.945 203.060 ;
        RECT 80.855 202.805 81.055 202.975 ;
        RECT 81.720 202.935 81.945 202.975 ;
        RECT 79.810 202.475 80.685 202.805 ;
        RECT 80.855 202.475 81.605 202.805 ;
        RECT 78.620 201.335 78.870 201.665 ;
        RECT 79.810 201.635 79.980 202.475 ;
        RECT 80.855 202.270 81.045 202.475 ;
        RECT 81.775 202.355 81.945 202.935 ;
        RECT 81.730 202.305 81.945 202.355 ;
        RECT 80.150 201.895 81.045 202.270 ;
        RECT 81.555 202.225 81.945 202.305 ;
        RECT 79.095 201.465 79.980 201.635 ;
        RECT 80.160 201.165 80.475 201.665 ;
        RECT 80.705 201.335 81.045 201.895 ;
        RECT 81.215 201.165 81.385 202.175 ;
        RECT 81.555 201.380 81.885 202.225 ;
        RECT 82.165 202.170 82.365 203.060 ;
        RECT 82.665 202.805 82.835 203.215 ;
        RECT 82.665 202.475 83.005 202.805 ;
        RECT 82.665 201.970 82.835 202.475 ;
        RECT 83.175 202.140 83.345 203.215 ;
        RECT 82.205 201.800 82.835 201.970 ;
        RECT 83.045 201.885 83.345 202.140 ;
        RECT 83.555 202.055 83.775 203.380 ;
        RECT 83.990 202.105 84.305 203.380 ;
        RECT 84.790 203.335 85.120 203.715 ;
        RECT 85.290 203.160 85.575 203.545 ;
        RECT 85.745 203.335 86.080 203.715 ;
        RECT 86.360 203.245 86.530 203.715 ;
        RECT 84.475 202.185 84.805 203.155 ;
        RECT 85.290 202.975 86.085 203.160 ;
        RECT 86.700 203.075 87.030 203.545 ;
        RECT 87.200 203.245 87.370 203.715 ;
        RECT 87.540 203.075 87.790 203.545 ;
        RECT 87.970 203.315 88.350 203.715 ;
        RECT 88.570 203.145 88.740 203.495 ;
        RECT 88.910 203.315 89.240 203.715 ;
        RECT 89.440 203.145 89.610 203.495 ;
        RECT 89.940 203.215 90.190 203.715 ;
        RECT 85.025 202.475 85.285 202.805 ;
        RECT 85.025 202.005 85.195 202.475 ;
        RECT 85.455 202.265 86.085 202.975 ;
        RECT 84.470 201.885 85.195 202.005 ;
        RECT 83.045 201.835 85.195 201.885 ;
        RECT 85.370 202.055 86.085 202.265 ;
        RECT 86.255 202.895 87.790 203.075 ;
        RECT 87.960 202.975 89.770 203.145 ;
        RECT 86.255 202.345 86.500 202.895 ;
        RECT 87.960 202.725 88.130 202.975 ;
        RECT 86.670 202.555 88.130 202.725 ;
        RECT 88.300 202.355 88.470 202.805 ;
        RECT 86.255 202.175 87.830 202.345 ;
        RECT 88.035 202.185 88.470 202.355 ;
        RECT 88.700 202.350 89.030 202.805 ;
        RECT 82.205 201.335 82.375 201.800 ;
        RECT 83.045 201.715 84.640 201.835 ;
        RECT 82.545 201.165 82.875 201.605 ;
        RECT 83.045 201.335 83.215 201.715 ;
        RECT 83.585 201.165 84.255 201.545 ;
        RECT 84.470 201.335 84.640 201.715 ;
        RECT 84.870 201.165 85.200 201.605 ;
        RECT 85.370 201.335 85.575 202.055 ;
        RECT 85.745 201.165 86.080 201.885 ;
        RECT 86.320 201.165 86.570 202.005 ;
        RECT 86.740 201.335 86.990 202.175 ;
        RECT 87.160 201.165 87.410 202.005 ;
        RECT 87.580 201.335 87.830 202.175 ;
        RECT 88.700 202.015 88.910 202.350 ;
        RECT 89.260 202.180 89.430 202.805 ;
        RECT 88.055 201.165 88.305 202.005 ;
        RECT 88.590 201.425 88.910 202.015 ;
        RECT 89.080 201.425 89.430 202.180 ;
        RECT 89.600 202.305 89.770 202.975 ;
        RECT 89.940 202.475 90.225 203.045 ;
        RECT 90.855 202.915 91.165 203.715 ;
        RECT 91.370 202.915 92.065 203.545 ;
        RECT 92.400 203.205 92.640 203.715 ;
        RECT 92.820 203.205 93.100 203.535 ;
        RECT 93.330 203.205 93.545 203.715 ;
        RECT 90.865 202.475 91.200 202.745 ;
        RECT 91.370 202.315 91.540 202.915 ;
        RECT 91.710 202.475 92.045 202.725 ;
        RECT 92.295 202.475 92.650 203.035 ;
        RECT 89.600 202.135 90.195 202.305 ;
        RECT 89.860 201.350 90.195 202.135 ;
        RECT 90.855 201.165 91.135 202.305 ;
        RECT 91.305 201.335 91.635 202.315 ;
        RECT 92.820 202.305 92.990 203.205 ;
        RECT 93.160 202.475 93.425 203.035 ;
        RECT 93.715 202.975 94.330 203.545 ;
        RECT 94.535 203.335 95.425 203.505 ;
        RECT 93.675 202.305 93.845 202.805 ;
        RECT 91.805 201.165 92.065 202.305 ;
        RECT 92.420 202.135 93.845 202.305 ;
        RECT 92.420 201.960 92.810 202.135 ;
        RECT 93.295 201.165 93.625 201.965 ;
        RECT 94.015 201.955 94.330 202.975 ;
        RECT 94.535 202.780 95.085 203.165 ;
        RECT 95.255 202.610 95.425 203.335 ;
        RECT 94.535 202.540 95.425 202.610 ;
        RECT 95.595 203.010 95.815 203.495 ;
        RECT 95.985 203.175 96.235 203.715 ;
        RECT 96.405 203.065 96.665 203.545 ;
        RECT 97.755 203.335 98.645 203.505 ;
        RECT 95.595 202.585 95.925 203.010 ;
        RECT 94.535 202.515 95.430 202.540 ;
        RECT 94.535 202.500 95.440 202.515 ;
        RECT 94.535 202.485 95.445 202.500 ;
        RECT 94.535 202.480 95.455 202.485 ;
        RECT 94.535 202.470 95.460 202.480 ;
        RECT 94.535 202.460 95.465 202.470 ;
        RECT 94.535 202.455 95.475 202.460 ;
        RECT 94.535 202.445 95.485 202.455 ;
        RECT 94.535 202.440 95.495 202.445 ;
        RECT 94.535 201.990 94.795 202.440 ;
        RECT 95.160 202.435 95.495 202.440 ;
        RECT 95.160 202.430 95.510 202.435 ;
        RECT 95.160 202.420 95.525 202.430 ;
        RECT 95.160 202.415 95.550 202.420 ;
        RECT 96.095 202.415 96.325 202.810 ;
        RECT 95.160 202.410 96.325 202.415 ;
        RECT 95.190 202.375 96.325 202.410 ;
        RECT 95.225 202.350 96.325 202.375 ;
        RECT 95.255 202.320 96.325 202.350 ;
        RECT 95.275 202.290 96.325 202.320 ;
        RECT 95.295 202.260 96.325 202.290 ;
        RECT 95.365 202.250 96.325 202.260 ;
        RECT 95.390 202.240 96.325 202.250 ;
        RECT 95.410 202.225 96.325 202.240 ;
        RECT 95.430 202.210 96.325 202.225 ;
        RECT 95.435 202.200 96.220 202.210 ;
        RECT 95.450 202.165 96.220 202.200 ;
        RECT 93.795 201.335 94.330 201.955 ;
        RECT 94.965 201.845 95.295 202.090 ;
        RECT 95.465 201.915 96.220 202.165 ;
        RECT 96.495 202.035 96.665 203.065 ;
        RECT 97.755 202.780 98.305 203.165 ;
        RECT 98.475 202.610 98.645 203.335 ;
        RECT 94.965 201.820 95.150 201.845 ;
        RECT 94.535 201.720 95.150 201.820 ;
        RECT 94.535 201.165 95.140 201.720 ;
        RECT 95.315 201.335 95.795 201.675 ;
        RECT 95.965 201.165 96.220 201.710 ;
        RECT 96.390 201.335 96.665 202.035 ;
        RECT 97.755 202.540 98.645 202.610 ;
        RECT 98.815 203.035 99.035 203.495 ;
        RECT 99.205 203.175 99.455 203.715 ;
        RECT 99.625 203.065 99.885 203.545 ;
        RECT 98.815 203.010 99.065 203.035 ;
        RECT 98.815 202.585 99.145 203.010 ;
        RECT 97.755 202.515 98.650 202.540 ;
        RECT 97.755 202.500 98.660 202.515 ;
        RECT 97.755 202.485 98.665 202.500 ;
        RECT 97.755 202.480 98.675 202.485 ;
        RECT 97.755 202.470 98.680 202.480 ;
        RECT 97.755 202.460 98.685 202.470 ;
        RECT 97.755 202.455 98.695 202.460 ;
        RECT 97.755 202.445 98.705 202.455 ;
        RECT 97.755 202.440 98.715 202.445 ;
        RECT 97.755 201.990 98.015 202.440 ;
        RECT 98.380 202.435 98.715 202.440 ;
        RECT 98.380 202.430 98.730 202.435 ;
        RECT 98.380 202.420 98.745 202.430 ;
        RECT 98.380 202.415 98.770 202.420 ;
        RECT 99.315 202.415 99.545 202.810 ;
        RECT 98.380 202.410 99.545 202.415 ;
        RECT 98.410 202.375 99.545 202.410 ;
        RECT 98.445 202.350 99.545 202.375 ;
        RECT 98.475 202.320 99.545 202.350 ;
        RECT 98.495 202.290 99.545 202.320 ;
        RECT 98.515 202.260 99.545 202.290 ;
        RECT 98.585 202.250 99.545 202.260 ;
        RECT 98.610 202.240 99.545 202.250 ;
        RECT 98.630 202.225 99.545 202.240 ;
        RECT 98.650 202.210 99.545 202.225 ;
        RECT 98.655 202.200 99.440 202.210 ;
        RECT 98.670 202.165 99.440 202.200 ;
        RECT 98.185 201.845 98.515 202.090 ;
        RECT 98.685 201.915 99.440 202.165 ;
        RECT 99.715 202.035 99.885 203.065 ;
        RECT 100.055 202.990 100.345 203.715 ;
        RECT 100.600 203.215 101.095 203.545 ;
        RECT 98.185 201.820 98.370 201.845 ;
        RECT 97.755 201.720 98.370 201.820 ;
        RECT 97.755 201.165 98.360 201.720 ;
        RECT 98.535 201.335 99.015 201.675 ;
        RECT 99.185 201.165 99.440 201.710 ;
        RECT 99.610 201.335 99.885 202.035 ;
        RECT 100.055 201.165 100.345 202.330 ;
        RECT 100.515 201.725 100.755 203.035 ;
        RECT 100.925 202.305 101.095 203.215 ;
        RECT 101.315 202.475 101.665 203.440 ;
        RECT 101.845 202.475 102.145 203.445 ;
        RECT 102.325 202.475 102.605 203.445 ;
        RECT 102.785 202.915 103.055 203.715 ;
        RECT 103.225 202.995 103.565 203.505 ;
        RECT 102.800 202.475 103.130 202.725 ;
        RECT 102.800 202.305 103.115 202.475 ;
        RECT 100.925 202.135 103.115 202.305 ;
        RECT 100.520 201.165 100.855 201.545 ;
        RECT 101.025 201.335 101.275 202.135 ;
        RECT 101.495 201.165 101.825 201.885 ;
        RECT 102.010 201.335 102.260 202.135 ;
        RECT 102.725 201.165 103.055 201.965 ;
        RECT 103.305 201.595 103.565 202.995 ;
        RECT 103.225 201.335 103.565 201.595 ;
        RECT 103.735 203.065 103.995 203.545 ;
        RECT 104.165 203.255 104.495 203.715 ;
        RECT 104.685 203.075 104.885 203.495 ;
        RECT 103.735 202.035 103.905 203.065 ;
        RECT 104.075 202.375 104.305 202.805 ;
        RECT 104.475 202.555 104.885 203.075 ;
        RECT 105.055 203.230 105.845 203.495 ;
        RECT 105.055 202.375 105.310 203.230 ;
        RECT 106.025 202.895 106.355 203.315 ;
        RECT 106.525 202.895 106.785 203.715 ;
        RECT 107.465 203.060 107.795 203.495 ;
        RECT 107.965 203.105 108.135 203.715 ;
        RECT 107.415 202.975 107.795 203.060 ;
        RECT 108.305 202.975 108.635 203.500 ;
        RECT 108.895 203.185 109.105 203.715 ;
        RECT 109.380 203.265 110.165 203.435 ;
        RECT 110.335 203.265 110.740 203.435 ;
        RECT 107.415 202.935 107.640 202.975 ;
        RECT 106.025 202.805 106.275 202.895 ;
        RECT 105.480 202.555 106.275 202.805 ;
        RECT 104.075 202.205 105.865 202.375 ;
        RECT 103.735 201.335 104.010 202.035 ;
        RECT 104.180 201.910 104.895 202.205 ;
        RECT 105.115 201.845 105.445 202.035 ;
        RECT 104.220 201.165 104.435 201.710 ;
        RECT 104.605 201.335 105.080 201.675 ;
        RECT 105.250 201.670 105.445 201.845 ;
        RECT 105.615 201.840 105.865 202.205 ;
        RECT 105.250 201.165 105.865 201.670 ;
        RECT 106.105 201.335 106.275 202.555 ;
        RECT 106.445 201.845 106.785 202.725 ;
        RECT 107.415 202.355 107.585 202.935 ;
        RECT 108.305 202.805 108.505 202.975 ;
        RECT 109.380 202.805 109.550 203.265 ;
        RECT 107.755 202.475 108.505 202.805 ;
        RECT 108.675 202.475 109.550 202.805 ;
        RECT 107.415 202.305 107.630 202.355 ;
        RECT 107.415 202.225 107.805 202.305 ;
        RECT 106.525 201.165 106.785 201.675 ;
        RECT 107.475 201.380 107.805 202.225 ;
        RECT 108.315 202.270 108.505 202.475 ;
        RECT 107.975 201.165 108.145 202.175 ;
        RECT 108.315 201.895 109.210 202.270 ;
        RECT 108.315 201.335 108.655 201.895 ;
        RECT 108.885 201.165 109.200 201.665 ;
        RECT 109.380 201.635 109.550 202.475 ;
        RECT 109.720 202.765 110.185 203.095 ;
        RECT 110.570 203.035 110.740 203.265 ;
        RECT 110.920 203.215 111.290 203.715 ;
        RECT 111.610 203.265 112.285 203.435 ;
        RECT 112.480 203.265 112.815 203.435 ;
        RECT 109.720 201.805 110.040 202.765 ;
        RECT 110.570 202.735 111.400 203.035 ;
        RECT 110.210 201.835 110.400 202.555 ;
        RECT 110.570 201.665 110.740 202.735 ;
        RECT 111.200 202.705 111.400 202.735 ;
        RECT 110.910 202.485 111.080 202.555 ;
        RECT 111.610 202.485 111.780 203.265 ;
        RECT 112.645 203.125 112.815 203.265 ;
        RECT 112.985 203.255 113.235 203.715 ;
        RECT 110.910 202.315 111.780 202.485 ;
        RECT 111.950 202.845 112.475 203.065 ;
        RECT 112.645 202.995 112.870 203.125 ;
        RECT 110.910 202.225 111.420 202.315 ;
        RECT 109.380 201.465 110.265 201.635 ;
        RECT 110.490 201.335 110.740 201.665 ;
        RECT 110.910 201.165 111.080 201.965 ;
        RECT 111.250 201.610 111.420 202.225 ;
        RECT 111.950 202.145 112.120 202.845 ;
        RECT 111.590 201.780 112.120 202.145 ;
        RECT 112.290 202.080 112.530 202.675 ;
        RECT 112.700 201.890 112.870 202.995 ;
        RECT 113.040 202.135 113.320 203.085 ;
        RECT 112.565 201.760 112.870 201.890 ;
        RECT 111.250 201.440 112.355 201.610 ;
        RECT 112.565 201.335 112.815 201.760 ;
        RECT 112.985 201.165 113.250 201.625 ;
        RECT 113.490 201.335 113.675 203.455 ;
        RECT 113.845 203.335 114.175 203.715 ;
        RECT 114.345 203.165 114.515 203.455 ;
        RECT 113.850 202.995 114.515 203.165 ;
        RECT 113.850 202.005 114.080 202.995 ;
        RECT 114.775 202.945 116.445 203.715 ;
        RECT 117.165 203.165 117.335 203.455 ;
        RECT 117.505 203.335 117.835 203.715 ;
        RECT 117.165 202.995 117.830 203.165 ;
        RECT 114.250 202.175 114.600 202.825 ;
        RECT 114.775 202.425 115.525 202.945 ;
        RECT 115.695 202.255 116.445 202.775 ;
        RECT 113.850 201.835 114.515 202.005 ;
        RECT 113.845 201.165 114.175 201.665 ;
        RECT 114.345 201.335 114.515 201.835 ;
        RECT 114.775 201.165 116.445 202.255 ;
        RECT 117.080 202.175 117.430 202.825 ;
        RECT 117.600 202.005 117.830 202.995 ;
        RECT 117.165 201.835 117.830 202.005 ;
        RECT 117.165 201.335 117.335 201.835 ;
        RECT 117.505 201.165 117.835 201.665 ;
        RECT 118.005 201.335 118.190 203.455 ;
        RECT 118.445 203.255 118.695 203.715 ;
        RECT 118.865 203.265 119.200 203.435 ;
        RECT 119.395 203.265 120.070 203.435 ;
        RECT 118.865 203.125 119.035 203.265 ;
        RECT 118.360 202.135 118.640 203.085 ;
        RECT 118.810 202.995 119.035 203.125 ;
        RECT 118.810 201.890 118.980 202.995 ;
        RECT 119.205 202.845 119.730 203.065 ;
        RECT 119.150 202.080 119.390 202.675 ;
        RECT 119.560 202.145 119.730 202.845 ;
        RECT 119.900 202.485 120.070 203.265 ;
        RECT 120.390 203.215 120.760 203.715 ;
        RECT 120.940 203.265 121.345 203.435 ;
        RECT 121.515 203.265 122.300 203.435 ;
        RECT 120.940 203.035 121.110 203.265 ;
        RECT 120.280 202.735 121.110 203.035 ;
        RECT 121.495 202.765 121.960 203.095 ;
        RECT 120.280 202.705 120.480 202.735 ;
        RECT 120.600 202.485 120.770 202.555 ;
        RECT 119.900 202.315 120.770 202.485 ;
        RECT 120.260 202.225 120.770 202.315 ;
        RECT 118.810 201.760 119.115 201.890 ;
        RECT 119.560 201.780 120.090 202.145 ;
        RECT 118.430 201.165 118.695 201.625 ;
        RECT 118.865 201.335 119.115 201.760 ;
        RECT 120.260 201.610 120.430 202.225 ;
        RECT 119.325 201.440 120.430 201.610 ;
        RECT 120.600 201.165 120.770 201.965 ;
        RECT 120.940 201.665 121.110 202.735 ;
        RECT 121.280 201.835 121.470 202.555 ;
        RECT 121.640 201.805 121.960 202.765 ;
        RECT 122.130 202.805 122.300 203.265 ;
        RECT 122.575 203.185 122.785 203.715 ;
        RECT 123.045 202.975 123.375 203.500 ;
        RECT 123.545 203.105 123.715 203.715 ;
        RECT 123.885 203.060 124.215 203.495 ;
        RECT 123.885 202.975 124.265 203.060 ;
        RECT 123.175 202.805 123.375 202.975 ;
        RECT 124.040 202.935 124.265 202.975 ;
        RECT 122.130 202.475 123.005 202.805 ;
        RECT 123.175 202.475 123.925 202.805 ;
        RECT 120.940 201.335 121.190 201.665 ;
        RECT 122.130 201.635 122.300 202.475 ;
        RECT 123.175 202.270 123.365 202.475 ;
        RECT 124.095 202.355 124.265 202.935 ;
        RECT 124.435 202.965 125.645 203.715 ;
        RECT 125.815 202.990 126.105 203.715 ;
        RECT 126.325 203.060 126.655 203.495 ;
        RECT 126.825 203.105 126.995 203.715 ;
        RECT 126.275 202.975 126.655 203.060 ;
        RECT 127.165 202.975 127.495 203.500 ;
        RECT 127.755 203.185 127.965 203.715 ;
        RECT 128.240 203.265 129.025 203.435 ;
        RECT 129.195 203.265 129.600 203.435 ;
        RECT 124.435 202.425 124.955 202.965 ;
        RECT 126.275 202.935 126.500 202.975 ;
        RECT 124.050 202.305 124.265 202.355 ;
        RECT 122.470 201.895 123.365 202.270 ;
        RECT 123.875 202.225 124.265 202.305 ;
        RECT 125.125 202.255 125.645 202.795 ;
        RECT 126.275 202.355 126.445 202.935 ;
        RECT 127.165 202.805 127.365 202.975 ;
        RECT 128.240 202.805 128.410 203.265 ;
        RECT 126.615 202.475 127.365 202.805 ;
        RECT 127.535 202.475 128.410 202.805 ;
        RECT 121.415 201.465 122.300 201.635 ;
        RECT 122.480 201.165 122.795 201.665 ;
        RECT 123.025 201.335 123.365 201.895 ;
        RECT 123.535 201.165 123.705 202.175 ;
        RECT 123.875 201.380 124.205 202.225 ;
        RECT 124.435 201.165 125.645 202.255 ;
        RECT 125.815 201.165 126.105 202.330 ;
        RECT 126.275 202.305 126.490 202.355 ;
        RECT 126.275 202.225 126.665 202.305 ;
        RECT 126.335 201.380 126.665 202.225 ;
        RECT 127.175 202.270 127.365 202.475 ;
        RECT 126.835 201.165 127.005 202.175 ;
        RECT 127.175 201.895 128.070 202.270 ;
        RECT 127.175 201.335 127.515 201.895 ;
        RECT 127.745 201.165 128.060 201.665 ;
        RECT 128.240 201.635 128.410 202.475 ;
        RECT 128.580 202.765 129.045 203.095 ;
        RECT 129.430 203.035 129.600 203.265 ;
        RECT 129.780 203.215 130.150 203.715 ;
        RECT 130.470 203.265 131.145 203.435 ;
        RECT 131.340 203.265 131.675 203.435 ;
        RECT 128.580 201.805 128.900 202.765 ;
        RECT 129.430 202.735 130.260 203.035 ;
        RECT 129.070 201.835 129.260 202.555 ;
        RECT 129.430 201.665 129.600 202.735 ;
        RECT 130.060 202.705 130.260 202.735 ;
        RECT 129.770 202.485 129.940 202.555 ;
        RECT 130.470 202.485 130.640 203.265 ;
        RECT 131.505 203.125 131.675 203.265 ;
        RECT 131.845 203.255 132.095 203.715 ;
        RECT 129.770 202.315 130.640 202.485 ;
        RECT 130.810 202.845 131.335 203.065 ;
        RECT 131.505 202.995 131.730 203.125 ;
        RECT 129.770 202.225 130.280 202.315 ;
        RECT 128.240 201.465 129.125 201.635 ;
        RECT 129.350 201.335 129.600 201.665 ;
        RECT 129.770 201.165 129.940 201.965 ;
        RECT 130.110 201.610 130.280 202.225 ;
        RECT 130.810 202.145 130.980 202.845 ;
        RECT 130.450 201.780 130.980 202.145 ;
        RECT 131.150 202.080 131.390 202.675 ;
        RECT 131.560 201.890 131.730 202.995 ;
        RECT 131.900 202.135 132.180 203.085 ;
        RECT 131.425 201.760 131.730 201.890 ;
        RECT 130.110 201.440 131.215 201.610 ;
        RECT 131.425 201.335 131.675 201.760 ;
        RECT 131.845 201.165 132.110 201.625 ;
        RECT 132.350 201.335 132.535 203.455 ;
        RECT 132.705 203.335 133.035 203.715 ;
        RECT 133.205 203.165 133.375 203.455 ;
        RECT 132.710 202.995 133.375 203.165 ;
        RECT 132.710 202.005 132.940 202.995 ;
        RECT 133.635 202.975 133.975 203.545 ;
        RECT 134.170 203.050 134.340 203.715 ;
        RECT 134.620 203.375 134.840 203.420 ;
        RECT 134.615 203.205 134.840 203.375 ;
        RECT 135.010 203.235 135.455 203.405 ;
        RECT 134.620 203.065 134.840 203.205 ;
        RECT 133.110 202.175 133.460 202.825 ;
        RECT 133.635 202.015 133.810 202.975 ;
        RECT 134.620 202.895 135.115 203.065 ;
        RECT 133.980 202.355 134.150 202.805 ;
        RECT 134.320 202.525 134.770 202.725 ;
        RECT 134.940 202.700 135.115 202.895 ;
        RECT 135.285 202.445 135.455 203.235 ;
        RECT 135.625 203.110 135.875 203.480 ;
        RECT 135.705 202.725 135.875 203.110 ;
        RECT 136.045 203.075 136.295 203.480 ;
        RECT 136.465 203.245 136.635 203.715 ;
        RECT 136.805 203.075 137.145 203.480 ;
        RECT 136.045 202.895 137.145 203.075 ;
        RECT 137.475 203.155 137.805 203.545 ;
        RECT 137.975 203.325 139.160 203.495 ;
        RECT 139.420 203.245 139.590 203.715 ;
        RECT 137.475 202.975 137.985 203.155 ;
        RECT 135.705 202.555 135.900 202.725 ;
        RECT 133.980 202.185 134.375 202.355 ;
        RECT 135.285 202.305 135.560 202.445 ;
        RECT 133.635 202.005 133.865 202.015 ;
        RECT 132.710 201.835 133.375 202.005 ;
        RECT 132.705 201.165 133.035 201.665 ;
        RECT 133.205 201.335 133.375 201.835 ;
        RECT 133.635 201.335 133.895 202.005 ;
        RECT 134.205 201.915 134.375 202.185 ;
        RECT 134.545 202.085 135.560 202.305 ;
        RECT 135.730 202.305 135.900 202.555 ;
        RECT 136.070 202.475 136.630 202.725 ;
        RECT 135.730 201.915 136.285 202.305 ;
        RECT 134.205 201.745 136.285 201.915 ;
        RECT 134.065 201.165 134.395 201.565 ;
        RECT 135.265 201.165 135.665 201.565 ;
        RECT 135.955 201.510 136.285 201.745 ;
        RECT 136.455 201.375 136.630 202.475 ;
        RECT 136.800 202.155 137.145 202.725 ;
        RECT 137.315 202.515 137.645 202.805 ;
        RECT 137.815 202.345 137.985 202.975 ;
        RECT 138.390 203.065 138.775 203.155 ;
        RECT 139.760 203.065 140.090 203.530 ;
        RECT 138.390 202.895 140.090 203.065 ;
        RECT 140.260 202.895 140.430 203.715 ;
        RECT 140.600 202.895 141.285 203.535 ;
        RECT 138.155 202.515 138.485 202.725 ;
        RECT 138.665 202.475 139.045 202.725 ;
        RECT 139.235 202.695 139.720 202.725 ;
        RECT 139.215 202.525 139.720 202.695 ;
        RECT 137.470 202.175 138.555 202.345 ;
        RECT 136.800 201.165 137.145 201.985 ;
        RECT 137.470 201.335 137.770 202.175 ;
        RECT 137.965 201.165 138.215 202.005 ;
        RECT 138.385 201.925 138.555 202.175 ;
        RECT 138.725 202.095 139.045 202.475 ;
        RECT 139.235 202.515 139.720 202.525 ;
        RECT 139.910 202.515 140.360 202.725 ;
        RECT 140.530 202.515 140.865 202.725 ;
        RECT 139.235 202.095 139.610 202.515 ;
        RECT 140.530 202.345 140.700 202.515 ;
        RECT 139.780 202.175 140.700 202.345 ;
        RECT 139.780 201.925 139.950 202.175 ;
        RECT 138.385 201.755 139.950 201.925 ;
        RECT 138.805 201.335 139.610 201.755 ;
        RECT 140.120 201.165 140.450 202.005 ;
        RECT 141.035 201.925 141.285 202.895 ;
        RECT 140.620 201.335 141.285 201.925 ;
        RECT 141.455 202.975 141.795 203.545 ;
        RECT 141.990 203.050 142.160 203.715 ;
        RECT 142.440 203.375 142.660 203.420 ;
        RECT 142.435 203.205 142.660 203.375 ;
        RECT 142.830 203.235 143.275 203.405 ;
        RECT 142.440 203.065 142.660 203.205 ;
        RECT 141.455 202.005 141.630 202.975 ;
        RECT 142.440 202.895 142.935 203.065 ;
        RECT 141.800 202.355 141.970 202.805 ;
        RECT 142.140 202.525 142.590 202.725 ;
        RECT 142.760 202.700 142.935 202.895 ;
        RECT 143.105 202.445 143.275 203.235 ;
        RECT 143.445 203.110 143.695 203.480 ;
        RECT 143.525 202.725 143.695 203.110 ;
        RECT 143.865 203.075 144.115 203.480 ;
        RECT 144.285 203.245 144.455 203.715 ;
        RECT 144.625 203.075 144.965 203.480 ;
        RECT 143.865 202.895 144.965 203.075 ;
        RECT 145.135 203.040 145.405 203.385 ;
        RECT 145.595 203.315 145.975 203.715 ;
        RECT 146.145 203.145 146.315 203.495 ;
        RECT 146.485 203.235 147.220 203.715 ;
        RECT 143.525 202.555 143.720 202.725 ;
        RECT 141.800 202.185 142.195 202.355 ;
        RECT 143.105 202.305 143.380 202.445 ;
        RECT 141.455 201.335 141.715 202.005 ;
        RECT 142.025 201.915 142.195 202.185 ;
        RECT 142.365 202.085 143.380 202.305 ;
        RECT 143.550 202.305 143.720 202.555 ;
        RECT 143.890 202.475 144.450 202.725 ;
        RECT 143.550 201.915 144.105 202.305 ;
        RECT 142.025 201.745 144.105 201.915 ;
        RECT 141.885 201.165 142.215 201.565 ;
        RECT 143.085 201.165 143.485 201.565 ;
        RECT 143.775 201.510 144.105 201.745 ;
        RECT 144.275 201.375 144.450 202.475 ;
        RECT 144.620 202.155 144.965 202.725 ;
        RECT 145.135 202.305 145.305 203.040 ;
        RECT 145.575 202.975 146.315 203.145 ;
        RECT 147.390 203.065 147.700 203.535 ;
        RECT 145.575 202.805 145.745 202.975 ;
        RECT 146.965 202.895 147.700 203.065 ;
        RECT 147.895 202.945 151.405 203.715 ;
        RECT 151.575 202.990 151.865 203.715 ;
        RECT 152.035 202.945 155.545 203.715 ;
        RECT 155.715 202.965 156.925 203.715 ;
        RECT 146.965 202.805 147.215 202.895 ;
        RECT 145.515 202.475 145.745 202.805 ;
        RECT 146.475 202.475 147.215 202.805 ;
        RECT 147.385 202.475 147.720 202.725 ;
        RECT 145.575 202.305 145.745 202.475 ;
        RECT 144.620 201.165 144.965 201.985 ;
        RECT 145.135 201.335 145.405 202.305 ;
        RECT 145.575 202.135 146.820 202.305 ;
        RECT 145.615 201.165 145.895 201.965 ;
        RECT 146.400 201.885 146.820 202.135 ;
        RECT 147.045 201.915 147.215 202.475 ;
        RECT 147.895 202.425 149.545 202.945 ;
        RECT 146.075 201.385 147.270 201.715 ;
        RECT 147.465 201.165 147.720 202.305 ;
        RECT 149.715 202.255 151.405 202.775 ;
        RECT 152.035 202.425 153.685 202.945 ;
        RECT 147.895 201.165 151.405 202.255 ;
        RECT 151.575 201.165 151.865 202.330 ;
        RECT 153.855 202.255 155.545 202.775 ;
        RECT 152.035 201.165 155.545 202.255 ;
        RECT 155.715 202.255 156.235 202.795 ;
        RECT 156.405 202.425 156.925 202.965 ;
        RECT 155.715 201.165 156.925 202.255 ;
        RECT 22.690 200.995 157.010 201.165 ;
        RECT 22.775 199.905 23.985 200.995 ;
        RECT 24.155 200.560 29.500 200.995 ;
        RECT 29.675 200.560 35.020 200.995 ;
        RECT 22.775 199.195 23.295 199.735 ;
        RECT 23.465 199.365 23.985 199.905 ;
        RECT 22.775 198.445 23.985 199.195 ;
        RECT 25.740 198.990 26.080 199.820 ;
        RECT 27.560 199.310 27.910 200.560 ;
        RECT 31.260 198.990 31.600 199.820 ;
        RECT 33.080 199.310 33.430 200.560 ;
        RECT 35.655 199.830 35.945 200.995 ;
        RECT 36.115 199.905 37.785 200.995 ;
        RECT 36.115 199.215 36.865 199.735 ;
        RECT 37.035 199.385 37.785 199.905 ;
        RECT 38.425 200.025 38.755 200.810 ;
        RECT 38.425 199.855 39.105 200.025 ;
        RECT 39.285 199.855 39.615 200.995 ;
        RECT 40.775 199.855 40.985 200.995 ;
        RECT 38.415 199.435 38.765 199.685 ;
        RECT 38.935 199.255 39.105 199.855 ;
        RECT 41.155 199.845 41.485 200.825 ;
        RECT 41.655 199.855 41.885 200.995 ;
        RECT 42.095 199.855 42.355 200.995 ;
        RECT 42.525 199.845 42.855 200.825 ;
        RECT 43.025 199.855 43.305 200.995 ;
        RECT 43.935 200.440 44.540 200.995 ;
        RECT 44.715 200.485 45.195 200.825 ;
        RECT 45.365 200.450 45.620 200.995 ;
        RECT 43.935 200.340 44.550 200.440 ;
        RECT 44.365 200.315 44.550 200.340 ;
        RECT 39.275 199.435 39.625 199.685 ;
        RECT 24.155 198.445 29.500 198.990 ;
        RECT 29.675 198.445 35.020 198.990 ;
        RECT 35.655 198.445 35.945 199.170 ;
        RECT 36.115 198.445 37.785 199.215 ;
        RECT 38.435 198.445 38.675 199.255 ;
        RECT 38.845 198.615 39.175 199.255 ;
        RECT 39.345 198.445 39.615 199.255 ;
        RECT 40.775 198.445 40.985 199.265 ;
        RECT 41.155 199.245 41.405 199.845 ;
        RECT 41.575 199.435 41.905 199.685 ;
        RECT 42.115 199.435 42.450 199.685 ;
        RECT 41.155 198.615 41.485 199.245 ;
        RECT 41.655 198.445 41.885 199.265 ;
        RECT 42.620 199.245 42.790 199.845 ;
        RECT 43.935 199.720 44.195 200.170 ;
        RECT 44.365 200.070 44.695 200.315 ;
        RECT 44.865 199.995 45.620 200.245 ;
        RECT 45.790 200.125 46.065 200.825 ;
        RECT 44.850 199.960 45.620 199.995 ;
        RECT 44.835 199.950 45.620 199.960 ;
        RECT 44.830 199.935 45.725 199.950 ;
        RECT 44.810 199.920 45.725 199.935 ;
        RECT 44.790 199.910 45.725 199.920 ;
        RECT 44.765 199.900 45.725 199.910 ;
        RECT 44.695 199.870 45.725 199.900 ;
        RECT 44.675 199.840 45.725 199.870 ;
        RECT 44.655 199.810 45.725 199.840 ;
        RECT 44.625 199.785 45.725 199.810 ;
        RECT 44.590 199.750 45.725 199.785 ;
        RECT 44.560 199.745 45.725 199.750 ;
        RECT 44.560 199.740 44.950 199.745 ;
        RECT 44.560 199.730 44.925 199.740 ;
        RECT 44.560 199.725 44.910 199.730 ;
        RECT 44.560 199.720 44.895 199.725 ;
        RECT 43.935 199.715 44.895 199.720 ;
        RECT 43.935 199.705 44.885 199.715 ;
        RECT 43.935 199.700 44.875 199.705 ;
        RECT 43.935 199.690 44.865 199.700 ;
        RECT 42.960 199.415 43.295 199.685 ;
        RECT 43.935 199.680 44.860 199.690 ;
        RECT 43.935 199.675 44.855 199.680 ;
        RECT 43.935 199.660 44.845 199.675 ;
        RECT 43.935 199.645 44.840 199.660 ;
        RECT 43.935 199.620 44.830 199.645 ;
        RECT 43.935 199.550 44.825 199.620 ;
        RECT 42.095 198.615 42.790 199.245 ;
        RECT 42.995 198.445 43.305 199.245 ;
        RECT 43.935 198.995 44.485 199.380 ;
        RECT 44.655 198.825 44.825 199.550 ;
        RECT 43.935 198.655 44.825 198.825 ;
        RECT 44.995 199.150 45.325 199.575 ;
        RECT 45.495 199.350 45.725 199.745 ;
        RECT 44.995 198.665 45.215 199.150 ;
        RECT 45.895 199.095 46.065 200.125 ;
        RECT 46.325 200.065 46.495 200.825 ;
        RECT 46.675 200.235 47.005 200.995 ;
        RECT 46.325 199.895 46.990 200.065 ;
        RECT 47.175 199.920 47.445 200.825 ;
        RECT 46.820 199.750 46.990 199.895 ;
        RECT 46.255 199.345 46.585 199.715 ;
        RECT 46.820 199.420 47.105 199.750 ;
        RECT 46.820 199.165 46.990 199.420 ;
        RECT 45.385 198.445 45.635 198.985 ;
        RECT 45.805 198.615 46.065 199.095 ;
        RECT 46.325 198.995 46.990 199.165 ;
        RECT 47.275 199.120 47.445 199.920 ;
        RECT 47.615 199.905 51.125 200.995 ;
        RECT 46.325 198.615 46.495 198.995 ;
        RECT 46.675 198.445 47.005 198.825 ;
        RECT 47.185 198.615 47.445 199.120 ;
        RECT 47.615 199.215 49.265 199.735 ;
        RECT 49.435 199.385 51.125 199.905 ;
        RECT 51.755 199.815 52.075 200.995 ;
        RECT 52.245 199.975 52.445 200.765 ;
        RECT 52.770 200.165 53.155 200.825 ;
        RECT 53.550 200.235 54.335 200.995 ;
        RECT 52.745 200.065 53.155 200.165 ;
        RECT 52.245 199.805 52.575 199.975 ;
        RECT 52.745 199.855 54.355 200.065 ;
        RECT 52.395 199.685 52.575 199.805 ;
        RECT 51.755 199.435 52.220 199.635 ;
        RECT 52.395 199.435 52.725 199.685 ;
        RECT 52.895 199.635 53.360 199.685 ;
        RECT 52.895 199.465 53.365 199.635 ;
        RECT 52.895 199.435 53.360 199.465 ;
        RECT 53.555 199.435 53.910 199.685 ;
        RECT 54.080 199.255 54.355 199.855 ;
        RECT 47.615 198.445 51.125 199.215 ;
        RECT 51.755 199.055 52.935 199.225 ;
        RECT 51.755 198.640 52.095 199.055 ;
        RECT 52.265 198.445 52.435 198.885 ;
        RECT 52.605 198.835 52.935 199.055 ;
        RECT 53.105 199.075 54.355 199.255 ;
        RECT 53.105 199.005 53.470 199.075 ;
        RECT 52.605 198.655 53.855 198.835 ;
        RECT 54.125 198.445 54.295 198.905 ;
        RECT 54.525 198.725 54.805 200.825 ;
        RECT 54.975 198.725 55.255 200.825 ;
        RECT 55.445 200.235 56.230 200.995 ;
        RECT 56.625 200.165 57.010 200.825 ;
        RECT 56.625 200.065 57.035 200.165 ;
        RECT 55.425 199.855 57.035 200.065 ;
        RECT 57.335 199.975 57.535 200.765 ;
        RECT 55.425 199.255 55.700 199.855 ;
        RECT 57.205 199.805 57.535 199.975 ;
        RECT 57.705 199.815 58.025 200.995 ;
        RECT 57.205 199.685 57.385 199.805 ;
        RECT 55.870 199.435 56.225 199.685 ;
        RECT 56.420 199.635 56.885 199.685 ;
        RECT 56.415 199.465 56.885 199.635 ;
        RECT 56.420 199.435 56.885 199.465 ;
        RECT 57.055 199.435 57.385 199.685 ;
        RECT 57.560 199.435 58.025 199.635 ;
        RECT 55.425 199.075 56.675 199.255 ;
        RECT 56.310 199.005 56.675 199.075 ;
        RECT 56.845 199.055 58.025 199.225 ;
        RECT 55.485 198.445 55.655 198.905 ;
        RECT 56.845 198.835 57.175 199.055 ;
        RECT 55.925 198.655 57.175 198.835 ;
        RECT 57.345 198.445 57.515 198.885 ;
        RECT 57.685 198.640 58.025 199.055 ;
        RECT 58.195 198.725 58.475 200.825 ;
        RECT 58.665 200.235 59.450 200.995 ;
        RECT 59.845 200.165 60.230 200.825 ;
        RECT 59.845 200.065 60.255 200.165 ;
        RECT 58.645 199.855 60.255 200.065 ;
        RECT 60.555 199.975 60.755 200.765 ;
        RECT 58.645 199.255 58.920 199.855 ;
        RECT 60.425 199.805 60.755 199.975 ;
        RECT 60.925 199.815 61.245 200.995 ;
        RECT 61.415 199.830 61.705 200.995 ;
        RECT 61.875 199.905 63.085 200.995 ;
        RECT 60.425 199.685 60.605 199.805 ;
        RECT 59.090 199.435 59.445 199.685 ;
        RECT 59.640 199.635 60.105 199.685 ;
        RECT 59.635 199.465 60.105 199.635 ;
        RECT 59.640 199.435 60.105 199.465 ;
        RECT 60.275 199.435 60.605 199.685 ;
        RECT 60.780 199.435 61.245 199.635 ;
        RECT 58.645 199.075 59.895 199.255 ;
        RECT 59.530 199.005 59.895 199.075 ;
        RECT 60.065 199.055 61.245 199.225 ;
        RECT 61.875 199.195 62.395 199.735 ;
        RECT 62.565 199.365 63.085 199.905 ;
        RECT 63.255 200.145 63.515 200.825 ;
        RECT 63.685 200.215 63.935 200.995 ;
        RECT 64.185 200.445 64.435 200.825 ;
        RECT 64.605 200.615 64.960 200.995 ;
        RECT 65.965 200.605 66.300 200.825 ;
        RECT 65.565 200.445 65.795 200.485 ;
        RECT 64.185 200.245 65.795 200.445 ;
        RECT 64.185 200.235 65.020 200.245 ;
        RECT 65.610 200.155 65.795 200.245 ;
        RECT 58.705 198.445 58.875 198.905 ;
        RECT 60.065 198.835 60.395 199.055 ;
        RECT 59.145 198.655 60.395 198.835 ;
        RECT 60.565 198.445 60.735 198.885 ;
        RECT 60.905 198.640 61.245 199.055 ;
        RECT 61.415 198.445 61.705 199.170 ;
        RECT 61.875 198.445 63.085 199.195 ;
        RECT 63.255 198.945 63.425 200.145 ;
        RECT 65.125 200.045 65.455 200.075 ;
        RECT 63.655 199.985 65.455 200.045 ;
        RECT 66.045 199.985 66.300 200.605 ;
        RECT 66.565 200.250 66.835 200.995 ;
        RECT 67.465 200.990 73.740 200.995 ;
        RECT 67.005 200.080 67.295 200.820 ;
        RECT 67.465 200.265 67.720 200.990 ;
        RECT 67.905 200.095 68.165 200.820 ;
        RECT 68.335 200.265 68.580 200.990 ;
        RECT 68.765 200.095 69.025 200.820 ;
        RECT 69.195 200.265 69.440 200.990 ;
        RECT 69.625 200.095 69.885 200.820 ;
        RECT 70.055 200.265 70.300 200.990 ;
        RECT 70.470 200.095 70.730 200.820 ;
        RECT 70.900 200.265 71.160 200.990 ;
        RECT 71.330 200.095 71.590 200.820 ;
        RECT 71.760 200.265 72.020 200.990 ;
        RECT 72.190 200.095 72.450 200.820 ;
        RECT 72.620 200.265 72.880 200.990 ;
        RECT 73.050 200.095 73.310 200.820 ;
        RECT 73.480 200.195 73.740 200.990 ;
        RECT 67.905 200.080 73.310 200.095 ;
        RECT 63.595 199.875 66.300 199.985 ;
        RECT 63.595 199.840 63.795 199.875 ;
        RECT 63.595 199.265 63.765 199.840 ;
        RECT 65.125 199.815 66.300 199.875 ;
        RECT 66.565 199.855 73.310 200.080 ;
        RECT 63.995 199.400 64.405 199.705 ;
        RECT 64.575 199.435 64.905 199.645 ;
        RECT 63.595 199.145 63.865 199.265 ;
        RECT 63.595 199.100 64.440 199.145 ;
        RECT 63.685 198.975 64.440 199.100 ;
        RECT 64.695 199.035 64.905 199.435 ;
        RECT 65.150 199.435 65.625 199.645 ;
        RECT 65.815 199.435 66.305 199.635 ;
        RECT 65.150 199.035 65.370 199.435 ;
        RECT 66.565 199.265 67.730 199.855 ;
        RECT 73.910 199.685 74.160 200.820 ;
        RECT 74.340 200.185 74.600 200.995 ;
        RECT 74.775 199.685 75.020 200.825 ;
        RECT 75.200 200.185 75.495 200.995 ;
        RECT 75.675 199.905 78.265 200.995 ;
        RECT 67.900 199.435 75.020 199.685 ;
        RECT 63.255 198.615 63.515 198.945 ;
        RECT 64.270 198.825 64.440 198.975 ;
        RECT 63.685 198.445 64.015 198.805 ;
        RECT 64.270 198.615 65.570 198.825 ;
        RECT 65.845 198.445 66.300 199.210 ;
        RECT 66.565 199.095 73.310 199.265 ;
        RECT 66.565 198.445 66.865 198.925 ;
        RECT 67.035 198.640 67.295 199.095 ;
        RECT 67.465 198.445 67.725 198.925 ;
        RECT 67.905 198.640 68.165 199.095 ;
        RECT 68.335 198.445 68.585 198.925 ;
        RECT 68.765 198.640 69.025 199.095 ;
        RECT 69.195 198.445 69.445 198.925 ;
        RECT 69.625 198.640 69.885 199.095 ;
        RECT 70.055 198.445 70.300 198.925 ;
        RECT 70.470 198.640 70.745 199.095 ;
        RECT 70.915 198.445 71.160 198.925 ;
        RECT 71.330 198.640 71.590 199.095 ;
        RECT 71.760 198.445 72.020 198.925 ;
        RECT 72.190 198.640 72.450 199.095 ;
        RECT 72.620 198.445 72.880 198.925 ;
        RECT 73.050 198.640 73.310 199.095 ;
        RECT 73.480 198.445 73.740 199.005 ;
        RECT 73.910 198.625 74.160 199.435 ;
        RECT 74.340 198.445 74.600 198.970 ;
        RECT 74.770 198.625 75.020 199.435 ;
        RECT 75.190 199.125 75.505 199.685 ;
        RECT 75.675 199.215 76.885 199.735 ;
        RECT 77.055 199.385 78.265 199.905 ;
        RECT 78.435 200.145 78.695 200.825 ;
        RECT 78.865 200.215 79.115 200.995 ;
        RECT 79.365 200.445 79.615 200.825 ;
        RECT 79.785 200.615 80.140 200.995 ;
        RECT 81.145 200.605 81.480 200.825 ;
        RECT 80.745 200.445 80.975 200.485 ;
        RECT 79.365 200.245 80.975 200.445 ;
        RECT 79.365 200.235 80.200 200.245 ;
        RECT 80.790 200.155 80.975 200.245 ;
        RECT 75.200 198.445 75.505 198.955 ;
        RECT 75.675 198.445 78.265 199.215 ;
        RECT 78.435 198.955 78.605 200.145 ;
        RECT 80.305 200.045 80.635 200.075 ;
        RECT 78.835 199.985 80.635 200.045 ;
        RECT 81.225 199.985 81.480 200.605 ;
        RECT 78.775 199.875 81.480 199.985 ;
        RECT 78.775 199.840 78.975 199.875 ;
        RECT 78.775 199.265 78.945 199.840 ;
        RECT 80.305 199.815 81.480 199.875 ;
        RECT 81.655 199.855 82.040 200.825 ;
        RECT 82.210 200.535 82.535 200.995 ;
        RECT 83.055 200.365 83.335 200.825 ;
        RECT 82.210 200.145 83.335 200.365 ;
        RECT 79.175 199.400 79.585 199.705 ;
        RECT 79.755 199.435 80.085 199.645 ;
        RECT 78.775 199.145 79.045 199.265 ;
        RECT 78.775 199.100 79.620 199.145 ;
        RECT 78.865 198.975 79.620 199.100 ;
        RECT 79.875 199.035 80.085 199.435 ;
        RECT 80.330 199.435 80.805 199.645 ;
        RECT 80.995 199.435 81.485 199.635 ;
        RECT 80.330 199.035 80.550 199.435 ;
        RECT 78.435 198.945 78.665 198.955 ;
        RECT 78.435 198.615 78.695 198.945 ;
        RECT 79.450 198.825 79.620 198.975 ;
        RECT 78.865 198.445 79.195 198.805 ;
        RECT 79.450 198.615 80.750 198.825 ;
        RECT 81.025 198.445 81.480 199.210 ;
        RECT 81.655 199.185 81.935 199.855 ;
        RECT 82.210 199.685 82.660 200.145 ;
        RECT 83.525 199.975 83.925 200.825 ;
        RECT 84.325 200.535 84.595 200.995 ;
        RECT 84.765 200.365 85.050 200.825 ;
        RECT 82.105 199.355 82.660 199.685 ;
        RECT 82.830 199.415 83.925 199.975 ;
        RECT 82.210 199.245 82.660 199.355 ;
        RECT 81.655 198.615 82.040 199.185 ;
        RECT 82.210 199.075 83.335 199.245 ;
        RECT 82.210 198.445 82.535 198.905 ;
        RECT 83.055 198.615 83.335 199.075 ;
        RECT 83.525 198.615 83.925 199.415 ;
        RECT 84.095 200.145 85.050 200.365 ;
        RECT 84.095 199.245 84.305 200.145 ;
        RECT 84.475 199.415 85.165 199.975 ;
        RECT 85.335 199.905 87.005 200.995 ;
        RECT 84.095 199.075 85.050 199.245 ;
        RECT 84.325 198.445 84.595 198.905 ;
        RECT 84.765 198.615 85.050 199.075 ;
        RECT 85.335 199.215 86.085 199.735 ;
        RECT 86.255 199.385 87.005 199.905 ;
        RECT 87.175 199.830 87.465 200.995 ;
        RECT 87.725 200.085 87.895 200.815 ;
        RECT 88.075 200.265 88.405 200.995 ;
        RECT 88.575 200.085 88.765 200.815 ;
        RECT 87.725 199.885 88.765 200.085 ;
        RECT 88.935 199.705 89.265 200.815 ;
        RECT 89.455 200.585 89.785 200.995 ;
        RECT 89.955 200.405 90.215 200.795 ;
        RECT 87.670 199.355 87.960 199.705 ;
        RECT 88.155 199.355 88.550 199.705 ;
        RECT 88.730 199.405 89.265 199.705 ;
        RECT 89.455 200.205 90.215 200.405 ;
        RECT 89.455 199.525 89.795 200.205 ;
        RECT 85.335 198.445 87.005 199.215 ;
        RECT 87.175 198.445 87.465 199.170 ;
        RECT 87.655 198.445 87.985 199.175 ;
        RECT 88.155 198.735 88.365 199.355 ;
        RECT 88.730 199.155 88.975 199.405 ;
        RECT 88.545 198.625 88.975 199.155 ;
        RECT 89.155 198.445 89.385 199.225 ;
        RECT 89.565 199.075 89.795 199.525 ;
        RECT 89.975 199.335 90.205 200.025 ;
        RECT 90.395 199.905 93.905 200.995 ;
        RECT 90.395 199.215 92.045 199.735 ;
        RECT 92.215 199.385 93.905 199.905 ;
        RECT 94.535 199.855 94.815 200.995 ;
        RECT 94.985 199.845 95.315 200.825 ;
        RECT 95.485 199.855 95.745 200.995 ;
        RECT 95.915 199.905 97.125 200.995 ;
        RECT 94.545 199.415 94.880 199.685 ;
        RECT 95.050 199.295 95.220 199.845 ;
        RECT 95.390 199.435 95.725 199.685 ;
        RECT 95.050 199.245 95.225 199.295 ;
        RECT 89.565 198.625 89.945 199.075 ;
        RECT 90.395 198.445 93.905 199.215 ;
        RECT 94.535 198.445 94.845 199.245 ;
        RECT 95.050 198.615 95.745 199.245 ;
        RECT 95.915 199.195 96.435 199.735 ;
        RECT 96.605 199.365 97.125 199.905 ;
        RECT 97.355 199.855 97.565 200.995 ;
        RECT 97.735 199.845 98.065 200.825 ;
        RECT 98.235 199.855 98.465 200.995 ;
        RECT 98.715 199.855 98.945 200.995 ;
        RECT 99.115 199.845 99.445 200.825 ;
        RECT 99.615 199.855 99.825 200.995 ;
        RECT 100.055 199.905 103.565 200.995 ;
        RECT 103.735 200.485 103.995 200.995 ;
        RECT 95.915 198.445 97.125 199.195 ;
        RECT 97.355 198.445 97.565 199.265 ;
        RECT 97.735 199.245 97.985 199.845 ;
        RECT 98.155 199.435 98.485 199.685 ;
        RECT 98.695 199.435 99.025 199.685 ;
        RECT 97.735 198.615 98.065 199.245 ;
        RECT 98.235 198.445 98.465 199.265 ;
        RECT 98.715 198.445 98.945 199.265 ;
        RECT 99.195 199.245 99.445 199.845 ;
        RECT 99.115 198.615 99.445 199.245 ;
        RECT 99.615 198.445 99.825 199.265 ;
        RECT 100.055 199.215 101.705 199.735 ;
        RECT 101.875 199.385 103.565 199.905 ;
        RECT 103.735 199.435 104.075 200.315 ;
        RECT 104.245 199.605 104.415 200.825 ;
        RECT 104.655 200.490 105.270 200.995 ;
        RECT 104.655 199.955 104.905 200.320 ;
        RECT 105.075 200.315 105.270 200.490 ;
        RECT 105.440 200.485 105.915 200.825 ;
        RECT 106.085 200.450 106.300 200.995 ;
        RECT 105.075 200.125 105.405 200.315 ;
        RECT 105.625 199.955 106.340 200.250 ;
        RECT 106.510 200.125 106.785 200.825 ;
        RECT 104.655 199.785 106.445 199.955 ;
        RECT 104.245 199.355 105.040 199.605 ;
        RECT 104.245 199.265 104.495 199.355 ;
        RECT 100.055 198.445 103.565 199.215 ;
        RECT 103.735 198.445 103.995 199.265 ;
        RECT 104.165 198.845 104.495 199.265 ;
        RECT 105.210 198.930 105.465 199.785 ;
        RECT 104.675 198.665 105.465 198.930 ;
        RECT 105.635 199.085 106.045 199.605 ;
        RECT 106.215 199.355 106.445 199.785 ;
        RECT 106.615 199.095 106.785 200.125 ;
        RECT 107.140 200.025 107.530 200.200 ;
        RECT 108.015 200.195 108.345 200.995 ;
        RECT 108.515 200.205 109.050 200.825 ;
        RECT 107.140 199.855 108.565 200.025 ;
        RECT 107.015 199.125 107.370 199.685 ;
        RECT 105.635 198.665 105.835 199.085 ;
        RECT 106.025 198.445 106.355 198.905 ;
        RECT 106.525 198.615 106.785 199.095 ;
        RECT 107.540 198.955 107.710 199.855 ;
        RECT 107.880 199.125 108.145 199.685 ;
        RECT 108.395 199.355 108.565 199.855 ;
        RECT 108.735 199.185 109.050 200.205 ;
        RECT 109.720 200.605 110.055 200.825 ;
        RECT 111.060 200.615 111.415 200.995 ;
        RECT 109.720 199.985 109.975 200.605 ;
        RECT 110.225 200.445 110.455 200.485 ;
        RECT 111.585 200.445 111.835 200.825 ;
        RECT 110.225 200.245 111.835 200.445 ;
        RECT 110.225 200.155 110.410 200.245 ;
        RECT 111.000 200.235 111.835 200.245 ;
        RECT 112.085 200.215 112.335 200.995 ;
        RECT 112.505 200.145 112.765 200.825 ;
        RECT 110.565 200.045 110.895 200.075 ;
        RECT 110.565 199.985 112.365 200.045 ;
        RECT 109.720 199.875 112.425 199.985 ;
        RECT 109.720 199.815 110.895 199.875 ;
        RECT 112.225 199.840 112.425 199.875 ;
        RECT 109.715 199.435 110.205 199.635 ;
        RECT 110.395 199.435 110.870 199.645 ;
        RECT 107.120 198.445 107.360 198.955 ;
        RECT 107.540 198.625 107.820 198.955 ;
        RECT 108.050 198.445 108.265 198.955 ;
        RECT 108.435 198.615 109.050 199.185 ;
        RECT 109.720 198.445 110.175 199.210 ;
        RECT 110.650 199.035 110.870 199.435 ;
        RECT 111.115 199.435 111.445 199.645 ;
        RECT 111.115 199.035 111.325 199.435 ;
        RECT 111.615 199.400 112.025 199.705 ;
        RECT 112.255 199.265 112.425 199.840 ;
        RECT 112.155 199.145 112.425 199.265 ;
        RECT 111.580 199.100 112.425 199.145 ;
        RECT 111.580 198.975 112.335 199.100 ;
        RECT 111.580 198.825 111.750 198.975 ;
        RECT 112.595 198.945 112.765 200.145 ;
        RECT 112.935 199.830 113.225 200.995 ;
        RECT 113.485 200.065 113.655 200.825 ;
        RECT 113.835 200.235 114.165 200.995 ;
        RECT 113.485 199.895 114.150 200.065 ;
        RECT 114.335 199.920 114.605 200.825 ;
        RECT 113.980 199.750 114.150 199.895 ;
        RECT 113.415 199.345 113.745 199.715 ;
        RECT 113.980 199.420 114.265 199.750 ;
        RECT 110.450 198.615 111.750 198.825 ;
        RECT 112.005 198.445 112.335 198.805 ;
        RECT 112.505 198.615 112.765 198.945 ;
        RECT 112.935 198.445 113.225 199.170 ;
        RECT 113.980 199.165 114.150 199.420 ;
        RECT 113.485 198.995 114.150 199.165 ;
        RECT 114.435 199.120 114.605 199.920 ;
        RECT 114.780 200.605 115.115 200.825 ;
        RECT 116.120 200.615 116.475 200.995 ;
        RECT 114.780 199.985 115.035 200.605 ;
        RECT 115.285 200.445 115.515 200.485 ;
        RECT 116.645 200.445 116.895 200.825 ;
        RECT 115.285 200.245 116.895 200.445 ;
        RECT 115.285 200.155 115.470 200.245 ;
        RECT 116.060 200.235 116.895 200.245 ;
        RECT 117.145 200.215 117.395 200.995 ;
        RECT 117.565 200.145 117.825 200.825 ;
        RECT 115.625 200.045 115.955 200.075 ;
        RECT 115.625 199.985 117.425 200.045 ;
        RECT 114.780 199.875 117.485 199.985 ;
        RECT 114.780 199.815 115.955 199.875 ;
        RECT 117.285 199.840 117.485 199.875 ;
        RECT 114.775 199.435 115.265 199.635 ;
        RECT 115.455 199.435 115.930 199.645 ;
        RECT 113.485 198.615 113.655 198.995 ;
        RECT 113.835 198.445 114.165 198.825 ;
        RECT 114.345 198.615 114.605 199.120 ;
        RECT 114.780 198.445 115.235 199.210 ;
        RECT 115.710 199.035 115.930 199.435 ;
        RECT 116.175 199.435 116.505 199.645 ;
        RECT 116.175 199.035 116.385 199.435 ;
        RECT 116.675 199.400 117.085 199.705 ;
        RECT 117.315 199.265 117.485 199.840 ;
        RECT 117.215 199.145 117.485 199.265 ;
        RECT 116.640 199.100 117.485 199.145 ;
        RECT 116.640 198.975 117.395 199.100 ;
        RECT 116.640 198.825 116.810 198.975 ;
        RECT 117.655 198.945 117.825 200.145 ;
        RECT 117.995 199.905 119.665 200.995 ;
        RECT 115.510 198.615 116.810 198.825 ;
        RECT 117.065 198.445 117.395 198.805 ;
        RECT 117.565 198.615 117.825 198.945 ;
        RECT 117.995 199.215 118.745 199.735 ;
        RECT 118.915 199.385 119.665 199.905 ;
        RECT 119.835 199.855 120.220 200.825 ;
        RECT 120.390 200.535 120.715 200.995 ;
        RECT 121.235 200.365 121.515 200.825 ;
        RECT 120.390 200.145 121.515 200.365 ;
        RECT 117.995 198.445 119.665 199.215 ;
        RECT 119.835 199.185 120.115 199.855 ;
        RECT 120.390 199.685 120.840 200.145 ;
        RECT 121.705 199.975 122.105 200.825 ;
        RECT 122.505 200.535 122.775 200.995 ;
        RECT 122.945 200.365 123.230 200.825 ;
        RECT 120.285 199.355 120.840 199.685 ;
        RECT 121.010 199.415 122.105 199.975 ;
        RECT 120.390 199.245 120.840 199.355 ;
        RECT 119.835 198.615 120.220 199.185 ;
        RECT 120.390 199.075 121.515 199.245 ;
        RECT 120.390 198.445 120.715 198.905 ;
        RECT 121.235 198.615 121.515 199.075 ;
        RECT 121.705 198.615 122.105 199.415 ;
        RECT 122.275 200.145 123.230 200.365 ;
        RECT 122.275 199.245 122.485 200.145 ;
        RECT 122.655 199.415 123.345 199.975 ;
        RECT 123.515 199.855 123.900 200.825 ;
        RECT 124.070 200.535 124.395 200.995 ;
        RECT 124.915 200.365 125.195 200.825 ;
        RECT 124.070 200.145 125.195 200.365 ;
        RECT 122.275 199.075 123.230 199.245 ;
        RECT 122.505 198.445 122.775 198.905 ;
        RECT 122.945 198.615 123.230 199.075 ;
        RECT 123.515 199.185 123.795 199.855 ;
        RECT 124.070 199.685 124.520 200.145 ;
        RECT 125.385 199.975 125.785 200.825 ;
        RECT 126.185 200.535 126.455 200.995 ;
        RECT 126.625 200.365 126.910 200.825 ;
        RECT 123.965 199.355 124.520 199.685 ;
        RECT 124.690 199.415 125.785 199.975 ;
        RECT 124.070 199.245 124.520 199.355 ;
        RECT 123.515 198.615 123.900 199.185 ;
        RECT 124.070 199.075 125.195 199.245 ;
        RECT 124.070 198.445 124.395 198.905 ;
        RECT 124.915 198.615 125.195 199.075 ;
        RECT 125.385 198.615 125.785 199.415 ;
        RECT 125.955 200.145 126.910 200.365 ;
        RECT 125.955 199.245 126.165 200.145 ;
        RECT 126.335 199.415 127.025 199.975 ;
        RECT 127.195 199.920 127.465 200.825 ;
        RECT 127.635 200.235 127.965 200.995 ;
        RECT 128.145 200.065 128.315 200.825 ;
        RECT 128.575 200.560 133.920 200.995 ;
        RECT 125.955 199.075 126.910 199.245 ;
        RECT 126.185 198.445 126.455 198.905 ;
        RECT 126.625 198.615 126.910 199.075 ;
        RECT 127.195 199.120 127.365 199.920 ;
        RECT 127.650 199.895 128.315 200.065 ;
        RECT 127.650 199.750 127.820 199.895 ;
        RECT 127.535 199.420 127.820 199.750 ;
        RECT 127.650 199.165 127.820 199.420 ;
        RECT 128.055 199.345 128.385 199.715 ;
        RECT 127.195 198.615 127.455 199.120 ;
        RECT 127.650 198.995 128.315 199.165 ;
        RECT 127.635 198.445 127.965 198.825 ;
        RECT 128.145 198.615 128.315 198.995 ;
        RECT 130.160 198.990 130.500 199.820 ;
        RECT 131.980 199.310 132.330 200.560 ;
        RECT 134.095 199.905 137.605 200.995 ;
        RECT 134.095 199.215 135.745 199.735 ;
        RECT 135.915 199.385 137.605 199.905 ;
        RECT 138.695 199.830 138.985 200.995 ;
        RECT 139.155 200.485 139.415 200.995 ;
        RECT 139.155 199.435 139.495 200.315 ;
        RECT 139.665 199.605 139.835 200.825 ;
        RECT 140.075 200.490 140.690 200.995 ;
        RECT 140.075 199.955 140.325 200.320 ;
        RECT 140.495 200.315 140.690 200.490 ;
        RECT 140.860 200.485 141.335 200.825 ;
        RECT 141.505 200.450 141.720 200.995 ;
        RECT 140.495 200.125 140.825 200.315 ;
        RECT 141.045 199.955 141.760 200.250 ;
        RECT 141.930 200.125 142.205 200.825 ;
        RECT 140.075 199.785 141.865 199.955 ;
        RECT 139.665 199.355 140.460 199.605 ;
        RECT 139.665 199.265 139.915 199.355 ;
        RECT 128.575 198.445 133.920 198.990 ;
        RECT 134.095 198.445 137.605 199.215 ;
        RECT 138.695 198.445 138.985 199.170 ;
        RECT 139.155 198.445 139.415 199.265 ;
        RECT 139.585 198.845 139.915 199.265 ;
        RECT 140.630 198.930 140.885 199.785 ;
        RECT 140.095 198.665 140.885 198.930 ;
        RECT 141.055 199.085 141.465 199.605 ;
        RECT 141.635 199.355 141.865 199.785 ;
        RECT 142.035 199.095 142.205 200.125 ;
        RECT 141.055 198.665 141.255 199.085 ;
        RECT 141.445 198.445 141.775 198.905 ;
        RECT 141.945 198.615 142.205 199.095 ;
        RECT 142.395 199.940 142.700 200.725 ;
        RECT 142.880 200.525 143.565 200.995 ;
        RECT 142.875 200.005 143.570 200.315 ;
        RECT 142.395 199.135 142.570 199.940 ;
        RECT 143.745 199.835 144.030 200.780 ;
        RECT 144.205 200.545 144.535 200.995 ;
        RECT 144.705 200.375 144.875 200.805 ;
        RECT 143.170 199.685 144.030 199.835 ;
        RECT 142.745 199.665 144.030 199.685 ;
        RECT 144.200 200.145 144.875 200.375 ;
        RECT 142.745 199.305 143.730 199.665 ;
        RECT 144.200 199.495 144.435 200.145 ;
        RECT 142.395 198.615 142.635 199.135 ;
        RECT 143.560 198.970 143.730 199.305 ;
        RECT 143.900 199.165 144.435 199.495 ;
        RECT 144.215 199.015 144.435 199.165 ;
        RECT 144.605 199.125 144.905 199.975 ;
        RECT 145.135 199.905 146.345 200.995 ;
        RECT 146.575 199.935 146.905 200.780 ;
        RECT 147.075 199.985 147.245 200.995 ;
        RECT 147.415 200.265 147.755 200.825 ;
        RECT 147.985 200.495 148.300 200.995 ;
        RECT 148.480 200.525 149.365 200.695 ;
        RECT 145.135 199.195 145.655 199.735 ;
        RECT 145.825 199.365 146.345 199.905 ;
        RECT 146.515 199.855 146.905 199.935 ;
        RECT 147.415 199.890 148.310 200.265 ;
        RECT 146.515 199.805 146.730 199.855 ;
        RECT 146.515 199.225 146.685 199.805 ;
        RECT 147.415 199.685 147.605 199.890 ;
        RECT 148.480 199.685 148.650 200.525 ;
        RECT 149.590 200.495 149.840 200.825 ;
        RECT 146.855 199.355 147.605 199.685 ;
        RECT 147.775 199.355 148.650 199.685 ;
        RECT 142.805 198.445 143.200 198.940 ;
        RECT 143.560 198.775 143.935 198.970 ;
        RECT 143.765 198.630 143.935 198.775 ;
        RECT 144.215 198.640 144.455 199.015 ;
        RECT 144.625 198.445 144.960 198.950 ;
        RECT 145.135 198.445 146.345 199.195 ;
        RECT 146.515 199.185 146.740 199.225 ;
        RECT 147.405 199.185 147.605 199.355 ;
        RECT 146.515 199.100 146.895 199.185 ;
        RECT 146.565 198.665 146.895 199.100 ;
        RECT 147.065 198.445 147.235 199.055 ;
        RECT 147.405 198.660 147.735 199.185 ;
        RECT 147.995 198.445 148.205 198.975 ;
        RECT 148.480 198.895 148.650 199.355 ;
        RECT 148.820 199.395 149.140 200.355 ;
        RECT 149.310 199.605 149.500 200.325 ;
        RECT 149.670 199.425 149.840 200.495 ;
        RECT 150.010 200.195 150.180 200.995 ;
        RECT 150.350 200.550 151.455 200.720 ;
        RECT 150.350 199.935 150.520 200.550 ;
        RECT 151.665 200.400 151.915 200.825 ;
        RECT 152.085 200.535 152.350 200.995 ;
        RECT 150.690 200.015 151.220 200.380 ;
        RECT 151.665 200.270 151.970 200.400 ;
        RECT 150.010 199.845 150.520 199.935 ;
        RECT 150.010 199.675 150.880 199.845 ;
        RECT 150.010 199.605 150.180 199.675 ;
        RECT 150.300 199.425 150.500 199.455 ;
        RECT 148.820 199.065 149.285 199.395 ;
        RECT 149.670 199.125 150.500 199.425 ;
        RECT 149.670 198.895 149.840 199.125 ;
        RECT 148.480 198.725 149.265 198.895 ;
        RECT 149.435 198.725 149.840 198.895 ;
        RECT 150.020 198.445 150.390 198.945 ;
        RECT 150.710 198.895 150.880 199.675 ;
        RECT 151.050 199.315 151.220 200.015 ;
        RECT 151.390 199.485 151.630 200.080 ;
        RECT 151.050 199.095 151.575 199.315 ;
        RECT 151.800 199.165 151.970 200.270 ;
        RECT 151.745 199.035 151.970 199.165 ;
        RECT 152.140 199.075 152.420 200.025 ;
        RECT 151.745 198.895 151.915 199.035 ;
        RECT 150.710 198.725 151.385 198.895 ;
        RECT 151.580 198.725 151.915 198.895 ;
        RECT 152.085 198.445 152.335 198.905 ;
        RECT 152.590 198.705 152.775 200.825 ;
        RECT 152.945 200.495 153.275 200.995 ;
        RECT 153.445 200.325 153.615 200.825 ;
        RECT 152.950 200.155 153.615 200.325 ;
        RECT 152.950 199.165 153.180 200.155 ;
        RECT 153.350 199.335 153.700 199.985 ;
        RECT 153.875 199.905 155.545 200.995 ;
        RECT 153.875 199.215 154.625 199.735 ;
        RECT 154.795 199.385 155.545 199.905 ;
        RECT 155.715 199.905 156.925 200.995 ;
        RECT 155.715 199.365 156.235 199.905 ;
        RECT 152.950 198.995 153.615 199.165 ;
        RECT 152.945 198.445 153.275 198.825 ;
        RECT 153.445 198.705 153.615 198.995 ;
        RECT 153.875 198.445 155.545 199.215 ;
        RECT 156.405 199.195 156.925 199.735 ;
        RECT 155.715 198.445 156.925 199.195 ;
        RECT 22.690 198.275 157.010 198.445 ;
        RECT 22.775 197.525 23.985 198.275 ;
        RECT 22.775 196.985 23.295 197.525 ;
        RECT 24.155 197.505 27.665 198.275 ;
        RECT 27.835 197.525 29.045 198.275 ;
        RECT 29.305 197.725 29.475 198.015 ;
        RECT 29.645 197.895 29.975 198.275 ;
        RECT 29.305 197.555 29.970 197.725 ;
        RECT 23.465 196.815 23.985 197.355 ;
        RECT 24.155 196.985 25.805 197.505 ;
        RECT 25.975 196.815 27.665 197.335 ;
        RECT 27.835 196.985 28.355 197.525 ;
        RECT 28.525 196.815 29.045 197.355 ;
        RECT 22.775 195.725 23.985 196.815 ;
        RECT 24.155 195.725 27.665 196.815 ;
        RECT 27.835 195.725 29.045 196.815 ;
        RECT 29.220 196.735 29.570 197.385 ;
        RECT 29.740 196.565 29.970 197.555 ;
        RECT 29.305 196.395 29.970 196.565 ;
        RECT 29.305 195.895 29.475 196.395 ;
        RECT 29.645 195.725 29.975 196.225 ;
        RECT 30.145 195.895 30.330 198.015 ;
        RECT 30.585 197.815 30.835 198.275 ;
        RECT 31.005 197.825 31.340 197.995 ;
        RECT 31.535 197.825 32.210 197.995 ;
        RECT 31.005 197.685 31.175 197.825 ;
        RECT 30.500 196.695 30.780 197.645 ;
        RECT 30.950 197.555 31.175 197.685 ;
        RECT 30.950 196.450 31.120 197.555 ;
        RECT 31.345 197.405 31.870 197.625 ;
        RECT 31.290 196.640 31.530 197.235 ;
        RECT 31.700 196.705 31.870 197.405 ;
        RECT 32.040 197.045 32.210 197.825 ;
        RECT 32.530 197.775 32.900 198.275 ;
        RECT 33.080 197.825 33.485 197.995 ;
        RECT 33.655 197.825 34.440 197.995 ;
        RECT 33.080 197.595 33.250 197.825 ;
        RECT 32.420 197.295 33.250 197.595 ;
        RECT 33.635 197.325 34.100 197.655 ;
        RECT 32.420 197.265 32.620 197.295 ;
        RECT 32.740 197.045 32.910 197.115 ;
        RECT 32.040 196.875 32.910 197.045 ;
        RECT 32.400 196.785 32.910 196.875 ;
        RECT 30.950 196.320 31.255 196.450 ;
        RECT 31.700 196.340 32.230 196.705 ;
        RECT 30.570 195.725 30.835 196.185 ;
        RECT 31.005 195.895 31.255 196.320 ;
        RECT 32.400 196.170 32.570 196.785 ;
        RECT 31.465 196.000 32.570 196.170 ;
        RECT 32.740 195.725 32.910 196.525 ;
        RECT 33.080 196.225 33.250 197.295 ;
        RECT 33.420 196.395 33.610 197.115 ;
        RECT 33.780 196.365 34.100 197.325 ;
        RECT 34.270 197.365 34.440 197.825 ;
        RECT 34.715 197.745 34.925 198.275 ;
        RECT 35.185 197.535 35.515 198.060 ;
        RECT 35.685 197.665 35.855 198.275 ;
        RECT 36.025 197.620 36.355 198.055 ;
        RECT 36.025 197.535 36.405 197.620 ;
        RECT 37.515 197.545 37.805 198.275 ;
        RECT 35.315 197.365 35.515 197.535 ;
        RECT 36.180 197.495 36.405 197.535 ;
        RECT 34.270 197.035 35.145 197.365 ;
        RECT 35.315 197.035 36.065 197.365 ;
        RECT 33.080 195.895 33.330 196.225 ;
        RECT 34.270 196.195 34.440 197.035 ;
        RECT 35.315 196.830 35.505 197.035 ;
        RECT 36.235 196.915 36.405 197.495 ;
        RECT 37.505 197.035 37.805 197.365 ;
        RECT 37.985 197.345 38.215 197.985 ;
        RECT 38.395 197.725 38.705 198.095 ;
        RECT 38.885 197.905 39.555 198.275 ;
        RECT 38.395 197.525 39.625 197.725 ;
        RECT 37.985 197.035 38.510 197.345 ;
        RECT 38.690 197.035 39.155 197.345 ;
        RECT 36.190 196.865 36.405 196.915 ;
        RECT 34.610 196.455 35.505 196.830 ;
        RECT 36.015 196.785 36.405 196.865 ;
        RECT 39.335 196.855 39.625 197.525 ;
        RECT 33.555 196.025 34.440 196.195 ;
        RECT 34.620 195.725 34.935 196.225 ;
        RECT 35.165 195.895 35.505 196.455 ;
        RECT 35.675 195.725 35.845 196.735 ;
        RECT 36.015 195.940 36.345 196.785 ;
        RECT 37.515 196.615 38.675 196.855 ;
        RECT 37.515 195.905 37.775 196.615 ;
        RECT 37.945 195.725 38.275 196.435 ;
        RECT 38.445 195.905 38.675 196.615 ;
        RECT 38.855 196.635 39.625 196.855 ;
        RECT 38.855 195.905 39.125 196.635 ;
        RECT 39.305 195.725 39.645 196.455 ;
        RECT 39.815 195.905 40.075 198.095 ;
        RECT 40.255 197.625 40.515 198.105 ;
        RECT 40.685 197.735 40.935 198.275 ;
        RECT 40.255 196.595 40.425 197.625 ;
        RECT 41.105 197.595 41.325 198.055 ;
        RECT 41.075 197.570 41.325 197.595 ;
        RECT 40.595 196.975 40.825 197.370 ;
        RECT 40.995 197.145 41.325 197.570 ;
        RECT 41.495 197.895 42.385 198.065 ;
        RECT 41.495 197.170 41.665 197.895 ;
        RECT 42.555 197.730 47.900 198.275 ;
        RECT 41.835 197.340 42.385 197.725 ;
        RECT 41.495 197.100 42.385 197.170 ;
        RECT 41.490 197.075 42.385 197.100 ;
        RECT 41.480 197.060 42.385 197.075 ;
        RECT 41.475 197.045 42.385 197.060 ;
        RECT 41.465 197.040 42.385 197.045 ;
        RECT 41.460 197.030 42.385 197.040 ;
        RECT 41.455 197.020 42.385 197.030 ;
        RECT 41.445 197.015 42.385 197.020 ;
        RECT 41.435 197.005 42.385 197.015 ;
        RECT 41.425 197.000 42.385 197.005 ;
        RECT 41.425 196.995 41.760 197.000 ;
        RECT 41.410 196.990 41.760 196.995 ;
        RECT 41.395 196.980 41.760 196.990 ;
        RECT 41.370 196.975 41.760 196.980 ;
        RECT 40.595 196.970 41.760 196.975 ;
        RECT 40.595 196.935 41.730 196.970 ;
        RECT 40.595 196.910 41.695 196.935 ;
        RECT 40.595 196.880 41.665 196.910 ;
        RECT 40.595 196.850 41.645 196.880 ;
        RECT 40.595 196.820 41.625 196.850 ;
        RECT 40.595 196.810 41.555 196.820 ;
        RECT 40.595 196.800 41.530 196.810 ;
        RECT 40.595 196.785 41.510 196.800 ;
        RECT 40.595 196.770 41.490 196.785 ;
        RECT 40.700 196.760 41.485 196.770 ;
        RECT 40.700 196.725 41.470 196.760 ;
        RECT 40.255 195.895 40.530 196.595 ;
        RECT 40.700 196.475 41.455 196.725 ;
        RECT 41.625 196.405 41.955 196.650 ;
        RECT 42.125 196.550 42.385 197.000 ;
        RECT 44.140 196.900 44.480 197.730 ;
        RECT 48.535 197.550 48.825 198.275 ;
        RECT 49.085 197.725 49.255 198.015 ;
        RECT 49.425 197.895 49.755 198.275 ;
        RECT 49.085 197.555 49.750 197.725 ;
        RECT 41.770 196.380 41.955 196.405 ;
        RECT 41.770 196.280 42.385 196.380 ;
        RECT 40.700 195.725 40.955 196.270 ;
        RECT 41.125 195.895 41.605 196.235 ;
        RECT 41.780 195.725 42.385 196.280 ;
        RECT 45.960 196.160 46.310 197.410 ;
        RECT 42.555 195.725 47.900 196.160 ;
        RECT 48.535 195.725 48.825 196.890 ;
        RECT 49.000 196.735 49.350 197.385 ;
        RECT 49.520 196.565 49.750 197.555 ;
        RECT 49.085 196.395 49.750 196.565 ;
        RECT 49.085 195.895 49.255 196.395 ;
        RECT 49.425 195.725 49.755 196.225 ;
        RECT 49.925 195.895 50.110 198.015 ;
        RECT 50.365 197.815 50.615 198.275 ;
        RECT 50.785 197.825 51.120 197.995 ;
        RECT 51.315 197.825 51.990 197.995 ;
        RECT 50.785 197.685 50.955 197.825 ;
        RECT 50.280 196.695 50.560 197.645 ;
        RECT 50.730 197.555 50.955 197.685 ;
        RECT 50.730 196.450 50.900 197.555 ;
        RECT 51.125 197.405 51.650 197.625 ;
        RECT 51.070 196.640 51.310 197.235 ;
        RECT 51.480 196.705 51.650 197.405 ;
        RECT 51.820 197.045 51.990 197.825 ;
        RECT 52.310 197.775 52.680 198.275 ;
        RECT 52.860 197.825 53.265 197.995 ;
        RECT 53.435 197.825 54.220 197.995 ;
        RECT 52.860 197.595 53.030 197.825 ;
        RECT 52.200 197.295 53.030 197.595 ;
        RECT 53.415 197.325 53.880 197.655 ;
        RECT 52.200 197.265 52.400 197.295 ;
        RECT 52.520 197.045 52.690 197.115 ;
        RECT 51.820 196.875 52.690 197.045 ;
        RECT 52.180 196.785 52.690 196.875 ;
        RECT 50.730 196.320 51.035 196.450 ;
        RECT 51.480 196.340 52.010 196.705 ;
        RECT 50.350 195.725 50.615 196.185 ;
        RECT 50.785 195.895 51.035 196.320 ;
        RECT 52.180 196.170 52.350 196.785 ;
        RECT 51.245 196.000 52.350 196.170 ;
        RECT 52.520 195.725 52.690 196.525 ;
        RECT 52.860 196.225 53.030 197.295 ;
        RECT 53.200 196.395 53.390 197.115 ;
        RECT 53.560 196.365 53.880 197.325 ;
        RECT 54.050 197.365 54.220 197.825 ;
        RECT 54.495 197.745 54.705 198.275 ;
        RECT 54.965 197.535 55.295 198.060 ;
        RECT 55.465 197.665 55.635 198.275 ;
        RECT 55.805 197.620 56.135 198.055 ;
        RECT 55.805 197.535 56.185 197.620 ;
        RECT 55.095 197.365 55.295 197.535 ;
        RECT 55.960 197.495 56.185 197.535 ;
        RECT 54.050 197.035 54.925 197.365 ;
        RECT 55.095 197.035 55.845 197.365 ;
        RECT 52.860 195.895 53.110 196.225 ;
        RECT 54.050 196.195 54.220 197.035 ;
        RECT 55.095 196.830 55.285 197.035 ;
        RECT 56.015 196.915 56.185 197.495 ;
        RECT 56.355 197.475 57.050 198.105 ;
        RECT 57.255 197.475 57.565 198.275 ;
        RECT 57.735 197.475 58.430 198.105 ;
        RECT 58.635 197.475 58.945 198.275 ;
        RECT 59.115 197.505 61.705 198.275 ;
        RECT 56.375 197.035 56.710 197.285 ;
        RECT 55.970 196.865 56.185 196.915 ;
        RECT 56.880 196.875 57.050 197.475 ;
        RECT 57.220 197.035 57.555 197.305 ;
        RECT 57.755 197.035 58.090 197.285 ;
        RECT 58.260 196.875 58.430 197.475 ;
        RECT 58.600 197.035 58.935 197.305 ;
        RECT 59.115 196.985 60.325 197.505 ;
        RECT 61.935 197.455 62.145 198.275 ;
        RECT 62.315 197.475 62.645 198.105 ;
        RECT 54.390 196.455 55.285 196.830 ;
        RECT 55.795 196.785 56.185 196.865 ;
        RECT 53.335 196.025 54.220 196.195 ;
        RECT 54.400 195.725 54.715 196.225 ;
        RECT 54.945 195.895 55.285 196.455 ;
        RECT 55.455 195.725 55.625 196.735 ;
        RECT 55.795 195.940 56.125 196.785 ;
        RECT 56.355 195.725 56.615 196.865 ;
        RECT 56.785 195.895 57.115 196.875 ;
        RECT 57.285 195.725 57.565 196.865 ;
        RECT 57.735 195.725 57.995 196.865 ;
        RECT 58.165 195.895 58.495 196.875 ;
        RECT 58.665 195.725 58.945 196.865 ;
        RECT 60.495 196.815 61.705 197.335 ;
        RECT 62.315 196.875 62.565 197.475 ;
        RECT 62.815 197.455 63.045 198.275 ;
        RECT 63.345 197.725 63.515 198.015 ;
        RECT 63.685 197.895 64.015 198.275 ;
        RECT 63.345 197.555 64.010 197.725 ;
        RECT 62.735 197.035 63.065 197.285 ;
        RECT 59.115 195.725 61.705 196.815 ;
        RECT 61.935 195.725 62.145 196.865 ;
        RECT 62.315 195.895 62.645 196.875 ;
        RECT 62.815 195.725 63.045 196.865 ;
        RECT 63.260 196.735 63.610 197.385 ;
        RECT 63.780 196.565 64.010 197.555 ;
        RECT 63.345 196.395 64.010 196.565 ;
        RECT 63.345 195.895 63.515 196.395 ;
        RECT 63.685 195.725 64.015 196.225 ;
        RECT 64.185 195.895 64.370 198.015 ;
        RECT 64.625 197.815 64.875 198.275 ;
        RECT 65.045 197.825 65.380 197.995 ;
        RECT 65.575 197.825 66.250 197.995 ;
        RECT 65.045 197.685 65.215 197.825 ;
        RECT 64.540 196.695 64.820 197.645 ;
        RECT 64.990 197.555 65.215 197.685 ;
        RECT 64.990 196.450 65.160 197.555 ;
        RECT 65.385 197.405 65.910 197.625 ;
        RECT 65.330 196.640 65.570 197.235 ;
        RECT 65.740 196.705 65.910 197.405 ;
        RECT 66.080 197.045 66.250 197.825 ;
        RECT 66.570 197.775 66.940 198.275 ;
        RECT 67.120 197.825 67.525 197.995 ;
        RECT 67.695 197.825 68.480 197.995 ;
        RECT 67.120 197.595 67.290 197.825 ;
        RECT 66.460 197.295 67.290 197.595 ;
        RECT 67.675 197.325 68.140 197.655 ;
        RECT 66.460 197.265 66.660 197.295 ;
        RECT 66.780 197.045 66.950 197.115 ;
        RECT 66.080 196.875 66.950 197.045 ;
        RECT 66.440 196.785 66.950 196.875 ;
        RECT 64.990 196.320 65.295 196.450 ;
        RECT 65.740 196.340 66.270 196.705 ;
        RECT 64.610 195.725 64.875 196.185 ;
        RECT 65.045 195.895 65.295 196.320 ;
        RECT 66.440 196.170 66.610 196.785 ;
        RECT 65.505 196.000 66.610 196.170 ;
        RECT 66.780 195.725 66.950 196.525 ;
        RECT 67.120 196.225 67.290 197.295 ;
        RECT 67.460 196.395 67.650 197.115 ;
        RECT 67.820 196.365 68.140 197.325 ;
        RECT 68.310 197.365 68.480 197.825 ;
        RECT 68.755 197.745 68.965 198.275 ;
        RECT 69.225 197.535 69.555 198.060 ;
        RECT 69.725 197.665 69.895 198.275 ;
        RECT 70.065 197.620 70.395 198.055 ;
        RECT 70.065 197.535 70.445 197.620 ;
        RECT 69.355 197.365 69.555 197.535 ;
        RECT 70.220 197.495 70.445 197.535 ;
        RECT 68.310 197.035 69.185 197.365 ;
        RECT 69.355 197.035 70.105 197.365 ;
        RECT 67.120 195.895 67.370 196.225 ;
        RECT 68.310 196.195 68.480 197.035 ;
        RECT 69.355 196.830 69.545 197.035 ;
        RECT 70.275 196.915 70.445 197.495 ;
        RECT 70.230 196.865 70.445 196.915 ;
        RECT 68.650 196.455 69.545 196.830 ;
        RECT 70.055 196.785 70.445 196.865 ;
        RECT 70.615 197.535 71.000 198.105 ;
        RECT 71.170 197.815 71.495 198.275 ;
        RECT 72.015 197.645 72.295 198.105 ;
        RECT 70.615 196.865 70.895 197.535 ;
        RECT 71.170 197.475 72.295 197.645 ;
        RECT 71.170 197.365 71.620 197.475 ;
        RECT 71.065 197.035 71.620 197.365 ;
        RECT 72.485 197.305 72.885 198.105 ;
        RECT 73.285 197.815 73.555 198.275 ;
        RECT 73.725 197.645 74.010 198.105 ;
        RECT 67.595 196.025 68.480 196.195 ;
        RECT 68.660 195.725 68.975 196.225 ;
        RECT 69.205 195.895 69.545 196.455 ;
        RECT 69.715 195.725 69.885 196.735 ;
        RECT 70.055 195.940 70.385 196.785 ;
        RECT 70.615 195.895 71.000 196.865 ;
        RECT 71.170 196.575 71.620 197.035 ;
        RECT 71.790 196.745 72.885 197.305 ;
        RECT 71.170 196.355 72.295 196.575 ;
        RECT 71.170 195.725 71.495 196.185 ;
        RECT 72.015 195.895 72.295 196.355 ;
        RECT 72.485 195.895 72.885 196.745 ;
        RECT 73.055 197.475 74.010 197.645 ;
        RECT 74.295 197.550 74.585 198.275 ;
        RECT 74.845 197.725 75.015 198.015 ;
        RECT 75.185 197.895 75.515 198.275 ;
        RECT 74.845 197.555 75.510 197.725 ;
        RECT 73.055 196.575 73.265 197.475 ;
        RECT 73.435 196.745 74.125 197.305 ;
        RECT 73.055 196.355 74.010 196.575 ;
        RECT 73.285 195.725 73.555 196.185 ;
        RECT 73.725 195.895 74.010 196.355 ;
        RECT 74.295 195.725 74.585 196.890 ;
        RECT 74.760 196.735 75.110 197.385 ;
        RECT 75.280 196.565 75.510 197.555 ;
        RECT 74.845 196.395 75.510 196.565 ;
        RECT 74.845 195.895 75.015 196.395 ;
        RECT 75.185 195.725 75.515 196.225 ;
        RECT 75.685 195.895 75.870 198.015 ;
        RECT 76.125 197.815 76.375 198.275 ;
        RECT 76.545 197.825 76.880 197.995 ;
        RECT 77.075 197.825 77.750 197.995 ;
        RECT 76.545 197.685 76.715 197.825 ;
        RECT 76.040 196.695 76.320 197.645 ;
        RECT 76.490 197.555 76.715 197.685 ;
        RECT 76.490 196.450 76.660 197.555 ;
        RECT 76.885 197.405 77.410 197.625 ;
        RECT 76.830 196.640 77.070 197.235 ;
        RECT 77.240 196.705 77.410 197.405 ;
        RECT 77.580 197.045 77.750 197.825 ;
        RECT 78.070 197.775 78.440 198.275 ;
        RECT 78.620 197.825 79.025 197.995 ;
        RECT 79.195 197.825 79.980 197.995 ;
        RECT 78.620 197.595 78.790 197.825 ;
        RECT 77.960 197.295 78.790 197.595 ;
        RECT 79.175 197.325 79.640 197.655 ;
        RECT 77.960 197.265 78.160 197.295 ;
        RECT 78.280 197.045 78.450 197.115 ;
        RECT 77.580 196.875 78.450 197.045 ;
        RECT 77.940 196.785 78.450 196.875 ;
        RECT 76.490 196.320 76.795 196.450 ;
        RECT 77.240 196.340 77.770 196.705 ;
        RECT 76.110 195.725 76.375 196.185 ;
        RECT 76.545 195.895 76.795 196.320 ;
        RECT 77.940 196.170 78.110 196.785 ;
        RECT 77.005 196.000 78.110 196.170 ;
        RECT 78.280 195.725 78.450 196.525 ;
        RECT 78.620 196.225 78.790 197.295 ;
        RECT 78.960 196.395 79.150 197.115 ;
        RECT 79.320 196.365 79.640 197.325 ;
        RECT 79.810 197.365 79.980 197.825 ;
        RECT 80.255 197.745 80.465 198.275 ;
        RECT 80.725 197.535 81.055 198.060 ;
        RECT 81.225 197.665 81.395 198.275 ;
        RECT 81.565 197.620 81.895 198.055 ;
        RECT 81.565 197.535 81.945 197.620 ;
        RECT 80.855 197.365 81.055 197.535 ;
        RECT 81.720 197.495 81.945 197.535 ;
        RECT 79.810 197.035 80.685 197.365 ;
        RECT 80.855 197.035 81.605 197.365 ;
        RECT 78.620 195.895 78.870 196.225 ;
        RECT 79.810 196.195 79.980 197.035 ;
        RECT 80.855 196.830 81.045 197.035 ;
        RECT 81.775 196.915 81.945 197.495 ;
        RECT 82.115 197.505 83.785 198.275 ;
        RECT 84.045 197.725 84.215 198.015 ;
        RECT 84.385 197.895 84.715 198.275 ;
        RECT 84.045 197.555 84.710 197.725 ;
        RECT 82.115 196.985 82.865 197.505 ;
        RECT 81.730 196.865 81.945 196.915 ;
        RECT 80.150 196.455 81.045 196.830 ;
        RECT 81.555 196.785 81.945 196.865 ;
        RECT 83.035 196.815 83.785 197.335 ;
        RECT 79.095 196.025 79.980 196.195 ;
        RECT 80.160 195.725 80.475 196.225 ;
        RECT 80.705 195.895 81.045 196.455 ;
        RECT 81.215 195.725 81.385 196.735 ;
        RECT 81.555 195.940 81.885 196.785 ;
        RECT 82.115 195.725 83.785 196.815 ;
        RECT 83.960 196.735 84.310 197.385 ;
        RECT 84.480 196.565 84.710 197.555 ;
        RECT 84.045 196.395 84.710 196.565 ;
        RECT 84.045 195.895 84.215 196.395 ;
        RECT 84.385 195.725 84.715 196.225 ;
        RECT 84.885 195.895 85.070 198.015 ;
        RECT 85.325 197.815 85.575 198.275 ;
        RECT 85.745 197.825 86.080 197.995 ;
        RECT 86.275 197.825 86.950 197.995 ;
        RECT 85.745 197.685 85.915 197.825 ;
        RECT 85.240 196.695 85.520 197.645 ;
        RECT 85.690 197.555 85.915 197.685 ;
        RECT 85.690 196.450 85.860 197.555 ;
        RECT 86.085 197.405 86.610 197.625 ;
        RECT 86.030 196.640 86.270 197.235 ;
        RECT 86.440 196.705 86.610 197.405 ;
        RECT 86.780 197.045 86.950 197.825 ;
        RECT 87.270 197.775 87.640 198.275 ;
        RECT 87.820 197.825 88.225 197.995 ;
        RECT 88.395 197.825 89.180 197.995 ;
        RECT 87.820 197.595 87.990 197.825 ;
        RECT 87.160 197.295 87.990 197.595 ;
        RECT 88.375 197.325 88.840 197.655 ;
        RECT 87.160 197.265 87.360 197.295 ;
        RECT 87.480 197.045 87.650 197.115 ;
        RECT 86.780 196.875 87.650 197.045 ;
        RECT 87.140 196.785 87.650 196.875 ;
        RECT 85.690 196.320 85.995 196.450 ;
        RECT 86.440 196.340 86.970 196.705 ;
        RECT 85.310 195.725 85.575 196.185 ;
        RECT 85.745 195.895 85.995 196.320 ;
        RECT 87.140 196.170 87.310 196.785 ;
        RECT 86.205 196.000 87.310 196.170 ;
        RECT 87.480 195.725 87.650 196.525 ;
        RECT 87.820 196.225 87.990 197.295 ;
        RECT 88.160 196.395 88.350 197.115 ;
        RECT 88.520 196.365 88.840 197.325 ;
        RECT 89.010 197.365 89.180 197.825 ;
        RECT 89.455 197.745 89.665 198.275 ;
        RECT 89.925 197.535 90.255 198.060 ;
        RECT 90.425 197.665 90.595 198.275 ;
        RECT 90.765 197.620 91.095 198.055 ;
        RECT 90.765 197.535 91.145 197.620 ;
        RECT 90.055 197.365 90.255 197.535 ;
        RECT 90.920 197.495 91.145 197.535 ;
        RECT 89.010 197.035 89.885 197.365 ;
        RECT 90.055 197.035 90.805 197.365 ;
        RECT 87.820 195.895 88.070 196.225 ;
        RECT 89.010 196.195 89.180 197.035 ;
        RECT 90.055 196.830 90.245 197.035 ;
        RECT 90.975 196.915 91.145 197.495 ;
        RECT 90.930 196.865 91.145 196.915 ;
        RECT 89.350 196.455 90.245 196.830 ;
        RECT 90.755 196.785 91.145 196.865 ;
        RECT 91.315 197.535 91.700 198.105 ;
        RECT 91.870 197.815 92.195 198.275 ;
        RECT 92.715 197.645 92.995 198.105 ;
        RECT 91.315 196.865 91.595 197.535 ;
        RECT 91.870 197.475 92.995 197.645 ;
        RECT 91.870 197.365 92.320 197.475 ;
        RECT 91.765 197.035 92.320 197.365 ;
        RECT 93.185 197.305 93.585 198.105 ;
        RECT 93.985 197.815 94.255 198.275 ;
        RECT 94.425 197.645 94.710 198.105 ;
        RECT 88.295 196.025 89.180 196.195 ;
        RECT 89.360 195.725 89.675 196.225 ;
        RECT 89.905 195.895 90.245 196.455 ;
        RECT 90.415 195.725 90.585 196.735 ;
        RECT 90.755 195.940 91.085 196.785 ;
        RECT 91.315 195.895 91.700 196.865 ;
        RECT 91.870 196.575 92.320 197.035 ;
        RECT 92.490 196.745 93.585 197.305 ;
        RECT 91.870 196.355 92.995 196.575 ;
        RECT 91.870 195.725 92.195 196.185 ;
        RECT 92.715 195.895 92.995 196.355 ;
        RECT 93.185 195.895 93.585 196.745 ;
        RECT 93.755 197.475 94.710 197.645 ;
        RECT 94.995 197.600 95.265 197.945 ;
        RECT 95.455 197.875 95.835 198.275 ;
        RECT 96.005 197.705 96.175 198.055 ;
        RECT 96.345 197.795 97.080 198.275 ;
        RECT 93.755 196.575 93.965 197.475 ;
        RECT 94.135 196.745 94.825 197.305 ;
        RECT 94.995 196.865 95.165 197.600 ;
        RECT 95.435 197.535 96.175 197.705 ;
        RECT 97.250 197.625 97.560 198.095 ;
        RECT 95.435 197.365 95.605 197.535 ;
        RECT 96.825 197.455 97.560 197.625 ;
        RECT 97.755 197.475 98.065 198.275 ;
        RECT 98.270 197.475 98.965 198.105 ;
        RECT 100.055 197.550 100.345 198.275 ;
        RECT 101.435 197.895 102.325 198.065 ;
        RECT 96.825 197.365 97.075 197.455 ;
        RECT 95.375 197.035 95.605 197.365 ;
        RECT 96.335 197.035 97.075 197.365 ;
        RECT 97.245 197.035 97.580 197.285 ;
        RECT 97.765 197.035 98.100 197.305 ;
        RECT 95.435 196.865 95.605 197.035 ;
        RECT 93.755 196.355 94.710 196.575 ;
        RECT 93.985 195.725 94.255 196.185 ;
        RECT 94.425 195.895 94.710 196.355 ;
        RECT 94.995 195.895 95.265 196.865 ;
        RECT 95.435 196.695 96.680 196.865 ;
        RECT 95.475 195.725 95.755 196.525 ;
        RECT 96.260 196.445 96.680 196.695 ;
        RECT 96.905 196.475 97.075 197.035 ;
        RECT 98.270 196.875 98.440 197.475 ;
        RECT 101.435 197.340 101.985 197.725 ;
        RECT 98.610 197.035 98.945 197.285 ;
        RECT 102.155 197.170 102.325 197.895 ;
        RECT 101.435 197.100 102.325 197.170 ;
        RECT 102.495 197.570 102.715 198.055 ;
        RECT 102.885 197.735 103.135 198.275 ;
        RECT 103.305 197.625 103.565 198.105 ;
        RECT 102.495 197.145 102.825 197.570 ;
        RECT 101.435 197.075 102.330 197.100 ;
        RECT 101.435 197.060 102.340 197.075 ;
        RECT 101.435 197.045 102.345 197.060 ;
        RECT 101.435 197.040 102.355 197.045 ;
        RECT 101.435 197.030 102.360 197.040 ;
        RECT 101.435 197.020 102.365 197.030 ;
        RECT 101.435 197.015 102.375 197.020 ;
        RECT 101.435 197.005 102.385 197.015 ;
        RECT 101.435 197.000 102.395 197.005 ;
        RECT 95.935 195.945 97.130 196.275 ;
        RECT 97.325 195.725 97.580 196.865 ;
        RECT 97.755 195.725 98.035 196.865 ;
        RECT 98.205 195.895 98.535 196.875 ;
        RECT 98.705 195.725 98.965 196.865 ;
        RECT 100.055 195.725 100.345 196.890 ;
        RECT 101.435 196.550 101.695 197.000 ;
        RECT 102.060 196.995 102.395 197.000 ;
        RECT 102.060 196.990 102.410 196.995 ;
        RECT 102.060 196.980 102.425 196.990 ;
        RECT 102.060 196.975 102.450 196.980 ;
        RECT 102.995 196.975 103.225 197.370 ;
        RECT 102.060 196.970 103.225 196.975 ;
        RECT 102.090 196.935 103.225 196.970 ;
        RECT 102.125 196.910 103.225 196.935 ;
        RECT 102.155 196.880 103.225 196.910 ;
        RECT 102.175 196.850 103.225 196.880 ;
        RECT 102.195 196.820 103.225 196.850 ;
        RECT 102.265 196.810 103.225 196.820 ;
        RECT 102.290 196.800 103.225 196.810 ;
        RECT 102.310 196.785 103.225 196.800 ;
        RECT 102.330 196.770 103.225 196.785 ;
        RECT 102.335 196.760 103.120 196.770 ;
        RECT 102.350 196.725 103.120 196.760 ;
        RECT 101.865 196.405 102.195 196.650 ;
        RECT 102.365 196.475 103.120 196.725 ;
        RECT 103.395 196.595 103.565 197.625 ;
        RECT 104.195 197.455 104.455 198.275 ;
        RECT 104.625 197.455 104.955 197.875 ;
        RECT 105.135 197.790 105.925 198.055 ;
        RECT 104.705 197.365 104.955 197.455 ;
        RECT 101.865 196.380 102.050 196.405 ;
        RECT 101.435 196.280 102.050 196.380 ;
        RECT 101.435 195.725 102.040 196.280 ;
        RECT 102.215 195.895 102.695 196.235 ;
        RECT 102.865 195.725 103.120 196.270 ;
        RECT 103.290 195.895 103.565 196.595 ;
        RECT 104.195 196.405 104.535 197.285 ;
        RECT 104.705 197.115 105.500 197.365 ;
        RECT 104.195 195.725 104.455 196.235 ;
        RECT 104.705 195.895 104.875 197.115 ;
        RECT 105.670 196.935 105.925 197.790 ;
        RECT 106.095 197.635 106.295 198.055 ;
        RECT 106.485 197.815 106.815 198.275 ;
        RECT 106.095 197.115 106.505 197.635 ;
        RECT 106.985 197.625 107.245 198.105 ;
        RECT 107.580 197.765 107.820 198.275 ;
        RECT 108.000 197.765 108.280 198.095 ;
        RECT 108.510 197.765 108.725 198.275 ;
        RECT 106.675 196.935 106.905 197.365 ;
        RECT 105.115 196.765 106.905 196.935 ;
        RECT 105.115 196.400 105.365 196.765 ;
        RECT 105.535 196.405 105.865 196.595 ;
        RECT 106.085 196.470 106.800 196.765 ;
        RECT 107.075 196.595 107.245 197.625 ;
        RECT 107.475 197.035 107.830 197.595 ;
        RECT 108.000 196.865 108.170 197.765 ;
        RECT 108.340 197.035 108.605 197.595 ;
        RECT 108.895 197.535 109.510 198.105 ;
        RECT 109.765 197.620 110.095 198.055 ;
        RECT 110.265 197.665 110.435 198.275 ;
        RECT 108.855 196.865 109.025 197.365 ;
        RECT 105.535 196.230 105.730 196.405 ;
        RECT 105.115 195.725 105.730 196.230 ;
        RECT 105.900 195.895 106.375 196.235 ;
        RECT 106.545 195.725 106.760 196.270 ;
        RECT 106.970 195.895 107.245 196.595 ;
        RECT 107.600 196.695 109.025 196.865 ;
        RECT 107.600 196.520 107.990 196.695 ;
        RECT 108.475 195.725 108.805 196.525 ;
        RECT 109.195 196.515 109.510 197.535 ;
        RECT 109.715 197.535 110.095 197.620 ;
        RECT 110.605 197.535 110.935 198.060 ;
        RECT 111.195 197.745 111.405 198.275 ;
        RECT 111.680 197.825 112.465 197.995 ;
        RECT 112.635 197.825 113.040 197.995 ;
        RECT 109.715 197.495 109.940 197.535 ;
        RECT 109.715 196.915 109.885 197.495 ;
        RECT 110.605 197.365 110.805 197.535 ;
        RECT 111.680 197.365 111.850 197.825 ;
        RECT 110.055 197.035 110.805 197.365 ;
        RECT 110.975 197.035 111.850 197.365 ;
        RECT 109.715 196.865 109.930 196.915 ;
        RECT 109.715 196.785 110.105 196.865 ;
        RECT 108.975 195.895 109.510 196.515 ;
        RECT 109.775 195.940 110.105 196.785 ;
        RECT 110.615 196.830 110.805 197.035 ;
        RECT 110.275 195.725 110.445 196.735 ;
        RECT 110.615 196.455 111.510 196.830 ;
        RECT 110.615 195.895 110.955 196.455 ;
        RECT 111.185 195.725 111.500 196.225 ;
        RECT 111.680 196.195 111.850 197.035 ;
        RECT 112.020 197.325 112.485 197.655 ;
        RECT 112.870 197.595 113.040 197.825 ;
        RECT 113.220 197.775 113.590 198.275 ;
        RECT 113.910 197.825 114.585 197.995 ;
        RECT 114.780 197.825 115.115 197.995 ;
        RECT 112.020 196.365 112.340 197.325 ;
        RECT 112.870 197.295 113.700 197.595 ;
        RECT 112.510 196.395 112.700 197.115 ;
        RECT 112.870 196.225 113.040 197.295 ;
        RECT 113.500 197.265 113.700 197.295 ;
        RECT 113.210 197.045 113.380 197.115 ;
        RECT 113.910 197.045 114.080 197.825 ;
        RECT 114.945 197.685 115.115 197.825 ;
        RECT 115.285 197.815 115.535 198.275 ;
        RECT 113.210 196.875 114.080 197.045 ;
        RECT 114.250 197.405 114.775 197.625 ;
        RECT 114.945 197.555 115.170 197.685 ;
        RECT 113.210 196.785 113.720 196.875 ;
        RECT 111.680 196.025 112.565 196.195 ;
        RECT 112.790 195.895 113.040 196.225 ;
        RECT 113.210 195.725 113.380 196.525 ;
        RECT 113.550 196.170 113.720 196.785 ;
        RECT 114.250 196.705 114.420 197.405 ;
        RECT 113.890 196.340 114.420 196.705 ;
        RECT 114.590 196.640 114.830 197.235 ;
        RECT 115.000 196.450 115.170 197.555 ;
        RECT 115.340 196.695 115.620 197.645 ;
        RECT 114.865 196.320 115.170 196.450 ;
        RECT 113.550 196.000 114.655 196.170 ;
        RECT 114.865 195.895 115.115 196.320 ;
        RECT 115.285 195.725 115.550 196.185 ;
        RECT 115.790 195.895 115.975 198.015 ;
        RECT 116.145 197.895 116.475 198.275 ;
        RECT 116.645 197.725 116.815 198.015 ;
        RECT 116.150 197.555 116.815 197.725 ;
        RECT 117.625 197.725 117.795 198.015 ;
        RECT 117.965 197.895 118.295 198.275 ;
        RECT 117.625 197.555 118.290 197.725 ;
        RECT 116.150 196.565 116.380 197.555 ;
        RECT 116.550 196.735 116.900 197.385 ;
        RECT 117.540 196.735 117.890 197.385 ;
        RECT 118.060 196.565 118.290 197.555 ;
        RECT 116.150 196.395 116.815 196.565 ;
        RECT 116.145 195.725 116.475 196.225 ;
        RECT 116.645 195.895 116.815 196.395 ;
        RECT 117.625 196.395 118.290 196.565 ;
        RECT 117.625 195.895 117.795 196.395 ;
        RECT 117.965 195.725 118.295 196.225 ;
        RECT 118.465 195.895 118.650 198.015 ;
        RECT 118.905 197.815 119.155 198.275 ;
        RECT 119.325 197.825 119.660 197.995 ;
        RECT 119.855 197.825 120.530 197.995 ;
        RECT 119.325 197.685 119.495 197.825 ;
        RECT 118.820 196.695 119.100 197.645 ;
        RECT 119.270 197.555 119.495 197.685 ;
        RECT 119.270 196.450 119.440 197.555 ;
        RECT 119.665 197.405 120.190 197.625 ;
        RECT 119.610 196.640 119.850 197.235 ;
        RECT 120.020 196.705 120.190 197.405 ;
        RECT 120.360 197.045 120.530 197.825 ;
        RECT 120.850 197.775 121.220 198.275 ;
        RECT 121.400 197.825 121.805 197.995 ;
        RECT 121.975 197.825 122.760 197.995 ;
        RECT 121.400 197.595 121.570 197.825 ;
        RECT 120.740 197.295 121.570 197.595 ;
        RECT 121.955 197.325 122.420 197.655 ;
        RECT 120.740 197.265 120.940 197.295 ;
        RECT 121.060 197.045 121.230 197.115 ;
        RECT 120.360 196.875 121.230 197.045 ;
        RECT 120.720 196.785 121.230 196.875 ;
        RECT 119.270 196.320 119.575 196.450 ;
        RECT 120.020 196.340 120.550 196.705 ;
        RECT 118.890 195.725 119.155 196.185 ;
        RECT 119.325 195.895 119.575 196.320 ;
        RECT 120.720 196.170 120.890 196.785 ;
        RECT 119.785 196.000 120.890 196.170 ;
        RECT 121.060 195.725 121.230 196.525 ;
        RECT 121.400 196.225 121.570 197.295 ;
        RECT 121.740 196.395 121.930 197.115 ;
        RECT 122.100 196.365 122.420 197.325 ;
        RECT 122.590 197.365 122.760 197.825 ;
        RECT 123.035 197.745 123.245 198.275 ;
        RECT 123.505 197.535 123.835 198.060 ;
        RECT 124.005 197.665 124.175 198.275 ;
        RECT 124.345 197.620 124.675 198.055 ;
        RECT 124.345 197.535 124.725 197.620 ;
        RECT 125.815 197.550 126.105 198.275 ;
        RECT 126.365 197.725 126.535 198.015 ;
        RECT 126.705 197.895 127.035 198.275 ;
        RECT 126.365 197.555 127.030 197.725 ;
        RECT 123.635 197.365 123.835 197.535 ;
        RECT 124.500 197.495 124.725 197.535 ;
        RECT 122.590 197.035 123.465 197.365 ;
        RECT 123.635 197.035 124.385 197.365 ;
        RECT 121.400 195.895 121.650 196.225 ;
        RECT 122.590 196.195 122.760 197.035 ;
        RECT 123.635 196.830 123.825 197.035 ;
        RECT 124.555 196.915 124.725 197.495 ;
        RECT 124.510 196.865 124.725 196.915 ;
        RECT 122.930 196.455 123.825 196.830 ;
        RECT 124.335 196.785 124.725 196.865 ;
        RECT 121.875 196.025 122.760 196.195 ;
        RECT 122.940 195.725 123.255 196.225 ;
        RECT 123.485 195.895 123.825 196.455 ;
        RECT 123.995 195.725 124.165 196.735 ;
        RECT 124.335 195.940 124.665 196.785 ;
        RECT 125.815 195.725 126.105 196.890 ;
        RECT 126.280 196.735 126.630 197.385 ;
        RECT 126.800 196.565 127.030 197.555 ;
        RECT 126.365 196.395 127.030 196.565 ;
        RECT 126.365 195.895 126.535 196.395 ;
        RECT 126.705 195.725 127.035 196.225 ;
        RECT 127.205 195.895 127.390 198.015 ;
        RECT 127.645 197.815 127.895 198.275 ;
        RECT 128.065 197.825 128.400 197.995 ;
        RECT 128.595 197.825 129.270 197.995 ;
        RECT 128.065 197.685 128.235 197.825 ;
        RECT 127.560 196.695 127.840 197.645 ;
        RECT 128.010 197.555 128.235 197.685 ;
        RECT 128.010 196.450 128.180 197.555 ;
        RECT 128.405 197.405 128.930 197.625 ;
        RECT 128.350 196.640 128.590 197.235 ;
        RECT 128.760 196.705 128.930 197.405 ;
        RECT 129.100 197.045 129.270 197.825 ;
        RECT 129.590 197.775 129.960 198.275 ;
        RECT 130.140 197.825 130.545 197.995 ;
        RECT 130.715 197.825 131.500 197.995 ;
        RECT 130.140 197.595 130.310 197.825 ;
        RECT 129.480 197.295 130.310 197.595 ;
        RECT 130.695 197.325 131.160 197.655 ;
        RECT 129.480 197.265 129.680 197.295 ;
        RECT 129.800 197.045 129.970 197.115 ;
        RECT 129.100 196.875 129.970 197.045 ;
        RECT 129.460 196.785 129.970 196.875 ;
        RECT 128.010 196.320 128.315 196.450 ;
        RECT 128.760 196.340 129.290 196.705 ;
        RECT 127.630 195.725 127.895 196.185 ;
        RECT 128.065 195.895 128.315 196.320 ;
        RECT 129.460 196.170 129.630 196.785 ;
        RECT 128.525 196.000 129.630 196.170 ;
        RECT 129.800 195.725 129.970 196.525 ;
        RECT 130.140 196.225 130.310 197.295 ;
        RECT 130.480 196.395 130.670 197.115 ;
        RECT 130.840 196.365 131.160 197.325 ;
        RECT 131.330 197.365 131.500 197.825 ;
        RECT 131.775 197.745 131.985 198.275 ;
        RECT 132.245 197.535 132.575 198.060 ;
        RECT 132.745 197.665 132.915 198.275 ;
        RECT 133.085 197.620 133.415 198.055 ;
        RECT 133.085 197.535 133.465 197.620 ;
        RECT 132.375 197.365 132.575 197.535 ;
        RECT 133.240 197.495 133.465 197.535 ;
        RECT 131.330 197.035 132.205 197.365 ;
        RECT 132.375 197.035 133.125 197.365 ;
        RECT 130.140 195.895 130.390 196.225 ;
        RECT 131.330 196.195 131.500 197.035 ;
        RECT 132.375 196.830 132.565 197.035 ;
        RECT 133.295 196.915 133.465 197.495 ;
        RECT 133.250 196.865 133.465 196.915 ;
        RECT 131.670 196.455 132.565 196.830 ;
        RECT 133.075 196.785 133.465 196.865 ;
        RECT 134.555 197.600 134.815 198.105 ;
        RECT 134.995 197.895 135.325 198.275 ;
        RECT 135.505 197.725 135.675 198.105 ;
        RECT 135.935 197.730 141.280 198.275 ;
        RECT 134.555 196.800 134.725 197.600 ;
        RECT 135.010 197.555 135.675 197.725 ;
        RECT 135.010 197.300 135.180 197.555 ;
        RECT 134.895 196.970 135.180 197.300 ;
        RECT 135.415 197.005 135.745 197.375 ;
        RECT 135.010 196.825 135.180 196.970 ;
        RECT 137.520 196.900 137.860 197.730 ;
        RECT 141.455 197.525 142.665 198.275 ;
        RECT 142.925 197.725 143.095 198.105 ;
        RECT 143.275 197.895 143.605 198.275 ;
        RECT 142.925 197.555 143.590 197.725 ;
        RECT 143.785 197.600 144.045 198.105 ;
        RECT 130.615 196.025 131.500 196.195 ;
        RECT 131.680 195.725 131.995 196.225 ;
        RECT 132.225 195.895 132.565 196.455 ;
        RECT 132.735 195.725 132.905 196.735 ;
        RECT 133.075 195.940 133.405 196.785 ;
        RECT 134.555 195.895 134.825 196.800 ;
        RECT 135.010 196.655 135.675 196.825 ;
        RECT 134.995 195.725 135.325 196.485 ;
        RECT 135.505 195.895 135.675 196.655 ;
        RECT 139.340 196.160 139.690 197.410 ;
        RECT 141.455 196.985 141.975 197.525 ;
        RECT 142.145 196.815 142.665 197.355 ;
        RECT 142.855 197.005 143.185 197.375 ;
        RECT 143.420 197.300 143.590 197.555 ;
        RECT 143.420 196.970 143.705 197.300 ;
        RECT 143.420 196.825 143.590 196.970 ;
        RECT 135.935 195.725 141.280 196.160 ;
        RECT 141.455 195.725 142.665 196.815 ;
        RECT 142.925 196.655 143.590 196.825 ;
        RECT 143.875 196.800 144.045 197.600 ;
        RECT 142.925 195.895 143.095 196.655 ;
        RECT 143.275 195.725 143.605 196.485 ;
        RECT 143.775 195.895 144.045 196.800 ;
        RECT 144.215 197.625 144.475 198.105 ;
        RECT 144.645 197.735 144.895 198.275 ;
        RECT 144.215 196.595 144.385 197.625 ;
        RECT 145.065 197.570 145.285 198.055 ;
        RECT 144.555 196.975 144.785 197.370 ;
        RECT 144.955 197.145 145.285 197.570 ;
        RECT 145.455 197.895 146.345 198.065 ;
        RECT 145.455 197.170 145.625 197.895 ;
        RECT 145.795 197.340 146.345 197.725 ;
        RECT 146.515 197.475 146.825 198.275 ;
        RECT 147.030 197.475 147.725 198.105 ;
        RECT 145.455 197.100 146.345 197.170 ;
        RECT 145.450 197.075 146.345 197.100 ;
        RECT 145.440 197.060 146.345 197.075 ;
        RECT 145.435 197.045 146.345 197.060 ;
        RECT 145.425 197.040 146.345 197.045 ;
        RECT 145.420 197.030 146.345 197.040 ;
        RECT 146.525 197.035 146.860 197.305 ;
        RECT 145.415 197.020 146.345 197.030 ;
        RECT 145.405 197.015 146.345 197.020 ;
        RECT 145.395 197.005 146.345 197.015 ;
        RECT 145.385 197.000 146.345 197.005 ;
        RECT 145.385 196.995 145.720 197.000 ;
        RECT 145.370 196.990 145.720 196.995 ;
        RECT 145.355 196.980 145.720 196.990 ;
        RECT 145.330 196.975 145.720 196.980 ;
        RECT 144.555 196.970 145.720 196.975 ;
        RECT 144.555 196.935 145.690 196.970 ;
        RECT 144.555 196.910 145.655 196.935 ;
        RECT 144.555 196.880 145.625 196.910 ;
        RECT 144.555 196.850 145.605 196.880 ;
        RECT 144.555 196.820 145.585 196.850 ;
        RECT 144.555 196.810 145.515 196.820 ;
        RECT 144.555 196.800 145.490 196.810 ;
        RECT 144.555 196.785 145.470 196.800 ;
        RECT 144.555 196.770 145.450 196.785 ;
        RECT 144.660 196.760 145.445 196.770 ;
        RECT 144.660 196.725 145.430 196.760 ;
        RECT 144.215 195.895 144.490 196.595 ;
        RECT 144.660 196.475 145.415 196.725 ;
        RECT 145.585 196.405 145.915 196.650 ;
        RECT 146.085 196.550 146.345 197.000 ;
        RECT 147.030 196.875 147.200 197.475 ;
        RECT 147.935 197.455 148.165 198.275 ;
        RECT 148.335 197.475 148.665 198.105 ;
        RECT 147.370 197.035 147.705 197.285 ;
        RECT 147.915 197.035 148.245 197.285 ;
        RECT 148.415 196.875 148.665 197.475 ;
        RECT 148.835 197.455 149.045 198.275 ;
        RECT 149.365 197.725 149.535 198.105 ;
        RECT 149.715 197.895 150.045 198.275 ;
        RECT 149.365 197.555 150.030 197.725 ;
        RECT 150.225 197.600 150.485 198.105 ;
        RECT 149.295 197.005 149.625 197.375 ;
        RECT 149.860 197.300 150.030 197.555 ;
        RECT 145.730 196.380 145.915 196.405 ;
        RECT 145.730 196.280 146.345 196.380 ;
        RECT 144.660 195.725 144.915 196.270 ;
        RECT 145.085 195.895 145.565 196.235 ;
        RECT 145.740 195.725 146.345 196.280 ;
        RECT 146.515 195.725 146.795 196.865 ;
        RECT 146.965 195.895 147.295 196.875 ;
        RECT 147.465 195.725 147.725 196.865 ;
        RECT 147.935 195.725 148.165 196.865 ;
        RECT 148.335 195.895 148.665 196.875 ;
        RECT 149.860 196.970 150.145 197.300 ;
        RECT 148.835 195.725 149.045 196.865 ;
        RECT 149.860 196.825 150.030 196.970 ;
        RECT 149.365 196.655 150.030 196.825 ;
        RECT 150.315 196.800 150.485 197.600 ;
        RECT 151.575 197.550 151.865 198.275 ;
        RECT 152.035 197.505 155.545 198.275 ;
        RECT 155.715 197.525 156.925 198.275 ;
        RECT 152.035 196.985 153.685 197.505 ;
        RECT 149.365 195.895 149.535 196.655 ;
        RECT 149.715 195.725 150.045 196.485 ;
        RECT 150.215 195.895 150.485 196.800 ;
        RECT 151.575 195.725 151.865 196.890 ;
        RECT 153.855 196.815 155.545 197.335 ;
        RECT 152.035 195.725 155.545 196.815 ;
        RECT 155.715 196.815 156.235 197.355 ;
        RECT 156.405 196.985 156.925 197.525 ;
        RECT 155.715 195.725 156.925 196.815 ;
        RECT 22.690 195.555 157.010 195.725 ;
        RECT 22.775 194.465 23.985 195.555 ;
        RECT 24.155 195.120 29.500 195.555 ;
        RECT 22.775 193.755 23.295 194.295 ;
        RECT 23.465 193.925 23.985 194.465 ;
        RECT 22.775 193.005 23.985 193.755 ;
        RECT 25.740 193.550 26.080 194.380 ;
        RECT 27.560 193.870 27.910 195.120 ;
        RECT 29.675 194.465 30.885 195.555 ;
        RECT 29.675 193.755 30.195 194.295 ;
        RECT 30.365 193.925 30.885 194.465 ;
        RECT 31.055 194.480 31.325 195.385 ;
        RECT 31.495 194.795 31.825 195.555 ;
        RECT 32.005 194.625 32.175 195.385 ;
        RECT 24.155 193.005 29.500 193.550 ;
        RECT 29.675 193.005 30.885 193.755 ;
        RECT 31.055 193.680 31.225 194.480 ;
        RECT 31.510 194.455 32.175 194.625 ;
        RECT 32.435 194.480 32.705 195.385 ;
        RECT 32.875 194.795 33.205 195.555 ;
        RECT 33.385 194.625 33.555 195.385 ;
        RECT 31.510 194.310 31.680 194.455 ;
        RECT 31.395 193.980 31.680 194.310 ;
        RECT 31.510 193.725 31.680 193.980 ;
        RECT 31.915 193.905 32.245 194.275 ;
        RECT 31.055 193.175 31.315 193.680 ;
        RECT 31.510 193.555 32.175 193.725 ;
        RECT 31.495 193.005 31.825 193.385 ;
        RECT 32.005 193.175 32.175 193.555 ;
        RECT 32.435 193.680 32.605 194.480 ;
        RECT 32.890 194.455 33.555 194.625 ;
        RECT 32.890 194.310 33.060 194.455 ;
        RECT 33.820 194.415 34.075 195.555 ;
        RECT 34.245 194.585 34.575 195.385 ;
        RECT 34.745 194.755 34.975 195.555 ;
        RECT 35.145 194.585 35.475 195.385 ;
        RECT 34.245 194.415 35.475 194.585 ;
        RECT 32.775 193.980 33.060 194.310 ;
        RECT 32.890 193.725 33.060 193.980 ;
        RECT 33.295 193.905 33.625 194.275 ;
        RECT 32.435 193.175 32.695 193.680 ;
        RECT 32.890 193.555 33.555 193.725 ;
        RECT 33.840 193.665 34.060 194.245 ;
        RECT 32.875 193.005 33.205 193.385 ;
        RECT 33.385 193.175 33.555 193.555 ;
        RECT 34.245 193.515 34.425 194.415 ;
        RECT 35.655 194.390 35.945 195.555 ;
        RECT 36.125 194.745 36.420 195.555 ;
        RECT 36.600 194.245 36.845 195.385 ;
        RECT 37.020 194.745 37.280 195.555 ;
        RECT 37.880 195.550 44.155 195.555 ;
        RECT 37.460 194.245 37.710 195.380 ;
        RECT 37.880 194.755 38.140 195.550 ;
        RECT 38.310 194.655 38.570 195.380 ;
        RECT 38.740 194.825 39.000 195.550 ;
        RECT 39.170 194.655 39.430 195.380 ;
        RECT 39.600 194.825 39.860 195.550 ;
        RECT 40.030 194.655 40.290 195.380 ;
        RECT 40.460 194.825 40.720 195.550 ;
        RECT 40.890 194.655 41.150 195.380 ;
        RECT 41.320 194.825 41.565 195.550 ;
        RECT 41.735 194.655 41.995 195.380 ;
        RECT 42.180 194.825 42.425 195.550 ;
        RECT 42.595 194.655 42.855 195.380 ;
        RECT 43.040 194.825 43.285 195.550 ;
        RECT 43.455 194.655 43.715 195.380 ;
        RECT 43.900 194.825 44.155 195.550 ;
        RECT 38.310 194.640 43.715 194.655 ;
        RECT 44.325 194.640 44.615 195.380 ;
        RECT 44.785 194.810 45.055 195.555 ;
        RECT 45.315 195.120 50.660 195.555 ;
        RECT 38.310 194.415 45.055 194.640 ;
        RECT 34.595 193.685 34.970 194.245 ;
        RECT 35.175 193.915 35.485 194.245 ;
        RECT 35.145 193.515 35.475 193.745 ;
        RECT 33.820 193.005 34.075 193.495 ;
        RECT 34.245 193.175 35.475 193.515 ;
        RECT 35.655 193.005 35.945 193.730 ;
        RECT 36.115 193.685 36.430 194.245 ;
        RECT 36.600 193.995 43.720 194.245 ;
        RECT 36.115 193.005 36.420 193.515 ;
        RECT 36.600 193.185 36.850 193.995 ;
        RECT 37.020 193.005 37.280 193.530 ;
        RECT 37.460 193.185 37.710 193.995 ;
        RECT 43.890 193.825 45.055 194.415 ;
        RECT 38.310 193.655 45.055 193.825 ;
        RECT 37.880 193.005 38.140 193.565 ;
        RECT 38.310 193.200 38.570 193.655 ;
        RECT 38.740 193.005 39.000 193.485 ;
        RECT 39.170 193.200 39.430 193.655 ;
        RECT 39.600 193.005 39.860 193.485 ;
        RECT 40.030 193.200 40.290 193.655 ;
        RECT 40.460 193.005 40.705 193.485 ;
        RECT 40.875 193.200 41.150 193.655 ;
        RECT 41.320 193.005 41.565 193.485 ;
        RECT 41.735 193.200 41.995 193.655 ;
        RECT 42.175 193.005 42.425 193.485 ;
        RECT 42.595 193.200 42.855 193.655 ;
        RECT 43.035 193.005 43.285 193.485 ;
        RECT 43.455 193.200 43.715 193.655 ;
        RECT 43.895 193.005 44.155 193.485 ;
        RECT 44.325 193.200 44.585 193.655 ;
        RECT 46.900 193.550 47.240 194.380 ;
        RECT 48.720 193.870 49.070 195.120 ;
        RECT 50.835 194.465 52.505 195.555 ;
        RECT 50.835 193.775 51.585 194.295 ;
        RECT 51.755 193.945 52.505 194.465 ;
        RECT 53.140 194.415 53.460 195.555 ;
        RECT 53.640 194.245 53.835 195.295 ;
        RECT 54.015 194.705 54.345 195.385 ;
        RECT 54.545 194.755 54.800 195.555 ;
        RECT 54.015 194.425 54.365 194.705 ;
        RECT 53.200 194.195 53.460 194.245 ;
        RECT 53.195 194.025 53.460 194.195 ;
        RECT 53.200 193.915 53.460 194.025 ;
        RECT 53.640 193.915 54.025 194.245 ;
        RECT 54.195 194.045 54.365 194.425 ;
        RECT 54.555 194.215 54.800 194.575 ;
        RECT 54.975 194.465 58.485 195.555 ;
        RECT 54.195 193.875 54.715 194.045 ;
        RECT 44.755 193.005 45.055 193.485 ;
        RECT 45.315 193.005 50.660 193.550 ;
        RECT 50.835 193.005 52.505 193.775 ;
        RECT 53.140 193.535 54.355 193.705 ;
        RECT 53.140 193.185 53.430 193.535 ;
        RECT 53.625 193.005 53.955 193.365 ;
        RECT 54.125 193.230 54.355 193.535 ;
        RECT 54.545 193.310 54.715 193.875 ;
        RECT 54.975 193.775 56.625 194.295 ;
        RECT 56.795 193.945 58.485 194.465 ;
        RECT 58.655 194.835 59.115 195.385 ;
        RECT 59.305 194.835 59.635 195.555 ;
        RECT 54.975 193.005 58.485 193.775 ;
        RECT 58.655 193.465 58.905 194.835 ;
        RECT 59.835 194.665 60.135 195.215 ;
        RECT 60.305 194.885 60.585 195.555 ;
        RECT 59.195 194.495 60.135 194.665 ;
        RECT 59.195 194.245 59.365 194.495 ;
        RECT 60.505 194.245 60.770 194.605 ;
        RECT 61.415 194.390 61.705 195.555 ;
        RECT 62.395 194.415 62.605 195.555 ;
        RECT 62.775 194.405 63.105 195.385 ;
        RECT 63.275 194.415 63.505 195.555 ;
        RECT 64.175 194.705 64.435 195.385 ;
        RECT 64.605 194.775 64.855 195.555 ;
        RECT 65.105 195.005 65.355 195.385 ;
        RECT 65.525 195.175 65.880 195.555 ;
        RECT 66.885 195.165 67.220 195.385 ;
        RECT 66.485 195.005 66.715 195.045 ;
        RECT 65.105 194.805 66.715 195.005 ;
        RECT 65.105 194.795 65.940 194.805 ;
        RECT 66.530 194.715 66.715 194.805 ;
        RECT 59.075 193.915 59.365 194.245 ;
        RECT 59.535 193.995 59.875 194.245 ;
        RECT 60.095 193.995 60.770 194.245 ;
        RECT 59.195 193.825 59.365 193.915 ;
        RECT 59.195 193.635 60.585 193.825 ;
        RECT 58.655 193.175 59.215 193.465 ;
        RECT 59.385 193.005 59.635 193.465 ;
        RECT 60.255 193.275 60.585 193.635 ;
        RECT 61.415 193.005 61.705 193.730 ;
        RECT 62.395 193.005 62.605 193.825 ;
        RECT 62.775 193.805 63.025 194.405 ;
        RECT 63.195 193.995 63.525 194.245 ;
        RECT 62.775 193.175 63.105 193.805 ;
        RECT 63.275 193.005 63.505 193.825 ;
        RECT 64.175 193.515 64.345 194.705 ;
        RECT 66.045 194.605 66.375 194.635 ;
        RECT 64.575 194.545 66.375 194.605 ;
        RECT 66.965 194.545 67.220 195.165 ;
        RECT 67.485 194.885 67.655 195.385 ;
        RECT 67.825 195.055 68.155 195.555 ;
        RECT 67.485 194.715 68.150 194.885 ;
        RECT 64.515 194.435 67.220 194.545 ;
        RECT 64.515 194.400 64.715 194.435 ;
        RECT 64.515 193.825 64.685 194.400 ;
        RECT 66.045 194.375 67.220 194.435 ;
        RECT 64.915 193.960 65.325 194.265 ;
        RECT 65.495 193.995 65.825 194.205 ;
        RECT 64.515 193.705 64.785 193.825 ;
        RECT 64.515 193.660 65.360 193.705 ;
        RECT 64.605 193.535 65.360 193.660 ;
        RECT 65.615 193.595 65.825 193.995 ;
        RECT 66.070 193.995 66.545 194.205 ;
        RECT 66.735 193.995 67.225 194.195 ;
        RECT 66.070 193.595 66.290 193.995 ;
        RECT 67.400 193.895 67.750 194.545 ;
        RECT 64.175 193.505 64.405 193.515 ;
        RECT 64.175 193.175 64.435 193.505 ;
        RECT 65.190 193.385 65.360 193.535 ;
        RECT 64.605 193.005 64.935 193.365 ;
        RECT 65.190 193.175 66.490 193.385 ;
        RECT 66.765 193.005 67.220 193.770 ;
        RECT 67.920 193.725 68.150 194.715 ;
        RECT 67.485 193.555 68.150 193.725 ;
        RECT 67.485 193.265 67.655 193.555 ;
        RECT 67.825 193.005 68.155 193.385 ;
        RECT 68.325 193.265 68.510 195.385 ;
        RECT 68.750 195.095 69.015 195.555 ;
        RECT 69.185 194.960 69.435 195.385 ;
        RECT 69.645 195.110 70.750 195.280 ;
        RECT 69.130 194.830 69.435 194.960 ;
        RECT 68.680 193.635 68.960 194.585 ;
        RECT 69.130 193.725 69.300 194.830 ;
        RECT 69.470 194.045 69.710 194.640 ;
        RECT 69.880 194.575 70.410 194.940 ;
        RECT 69.880 193.875 70.050 194.575 ;
        RECT 70.580 194.495 70.750 195.110 ;
        RECT 70.920 194.755 71.090 195.555 ;
        RECT 71.260 195.055 71.510 195.385 ;
        RECT 71.735 195.085 72.620 195.255 ;
        RECT 70.580 194.405 71.090 194.495 ;
        RECT 69.130 193.595 69.355 193.725 ;
        RECT 69.525 193.655 70.050 193.875 ;
        RECT 70.220 194.235 71.090 194.405 ;
        RECT 68.765 193.005 69.015 193.465 ;
        RECT 69.185 193.455 69.355 193.595 ;
        RECT 70.220 193.455 70.390 194.235 ;
        RECT 70.920 194.165 71.090 194.235 ;
        RECT 70.600 193.985 70.800 194.015 ;
        RECT 71.260 193.985 71.430 195.055 ;
        RECT 71.600 194.165 71.790 194.885 ;
        RECT 70.600 193.685 71.430 193.985 ;
        RECT 71.960 193.955 72.280 194.915 ;
        RECT 69.185 193.285 69.520 193.455 ;
        RECT 69.715 193.285 70.390 193.455 ;
        RECT 70.710 193.005 71.080 193.505 ;
        RECT 71.260 193.455 71.430 193.685 ;
        RECT 71.815 193.625 72.280 193.955 ;
        RECT 72.450 194.245 72.620 195.085 ;
        RECT 72.800 195.055 73.115 195.555 ;
        RECT 73.345 194.825 73.685 195.385 ;
        RECT 72.790 194.450 73.685 194.825 ;
        RECT 73.855 194.545 74.025 195.555 ;
        RECT 73.495 194.245 73.685 194.450 ;
        RECT 74.195 194.495 74.525 195.340 ;
        RECT 74.195 194.415 74.585 194.495 ;
        RECT 74.370 194.365 74.585 194.415 ;
        RECT 72.450 193.915 73.325 194.245 ;
        RECT 73.495 193.915 74.245 194.245 ;
        RECT 72.450 193.455 72.620 193.915 ;
        RECT 73.495 193.745 73.695 193.915 ;
        RECT 74.415 193.785 74.585 194.365 ;
        RECT 74.360 193.745 74.585 193.785 ;
        RECT 71.260 193.285 71.665 193.455 ;
        RECT 71.835 193.285 72.620 193.455 ;
        RECT 72.895 193.005 73.105 193.535 ;
        RECT 73.365 193.220 73.695 193.745 ;
        RECT 74.205 193.660 74.585 193.745 ;
        RECT 74.755 194.415 75.140 195.385 ;
        RECT 75.310 195.095 75.635 195.555 ;
        RECT 76.155 194.925 76.435 195.385 ;
        RECT 75.310 194.705 76.435 194.925 ;
        RECT 74.755 193.745 75.035 194.415 ;
        RECT 75.310 194.245 75.760 194.705 ;
        RECT 76.625 194.535 77.025 195.385 ;
        RECT 77.425 195.095 77.695 195.555 ;
        RECT 77.865 194.925 78.150 195.385 ;
        RECT 75.205 193.915 75.760 194.245 ;
        RECT 75.930 193.975 77.025 194.535 ;
        RECT 75.310 193.805 75.760 193.915 ;
        RECT 73.865 193.005 74.035 193.615 ;
        RECT 74.205 193.225 74.535 193.660 ;
        RECT 74.755 193.175 75.140 193.745 ;
        RECT 75.310 193.635 76.435 193.805 ;
        RECT 75.310 193.005 75.635 193.465 ;
        RECT 76.155 193.175 76.435 193.635 ;
        RECT 76.625 193.175 77.025 193.975 ;
        RECT 77.195 194.705 78.150 194.925 ;
        RECT 77.195 193.805 77.405 194.705 ;
        RECT 77.575 193.975 78.265 194.535 ;
        RECT 78.435 194.465 79.645 195.555 ;
        RECT 77.195 193.635 78.150 193.805 ;
        RECT 77.425 193.005 77.695 193.465 ;
        RECT 77.865 193.175 78.150 193.635 ;
        RECT 78.435 193.755 78.955 194.295 ;
        RECT 79.125 193.925 79.645 194.465 ;
        RECT 79.815 194.415 80.200 195.385 ;
        RECT 80.370 195.095 80.695 195.555 ;
        RECT 81.215 194.925 81.495 195.385 ;
        RECT 80.370 194.705 81.495 194.925 ;
        RECT 78.435 193.005 79.645 193.755 ;
        RECT 79.815 193.745 80.095 194.415 ;
        RECT 80.370 194.245 80.820 194.705 ;
        RECT 81.685 194.535 82.085 195.385 ;
        RECT 82.485 195.095 82.755 195.555 ;
        RECT 82.925 194.925 83.210 195.385 ;
        RECT 80.265 193.915 80.820 194.245 ;
        RECT 80.990 193.975 82.085 194.535 ;
        RECT 80.370 193.805 80.820 193.915 ;
        RECT 79.815 193.175 80.200 193.745 ;
        RECT 80.370 193.635 81.495 193.805 ;
        RECT 80.370 193.005 80.695 193.465 ;
        RECT 81.215 193.175 81.495 193.635 ;
        RECT 81.685 193.175 82.085 193.975 ;
        RECT 82.255 194.705 83.210 194.925 ;
        RECT 83.495 194.705 83.755 195.385 ;
        RECT 83.925 194.775 84.175 195.555 ;
        RECT 84.425 195.005 84.675 195.385 ;
        RECT 84.845 195.175 85.200 195.555 ;
        RECT 86.205 195.165 86.540 195.385 ;
        RECT 85.805 195.005 86.035 195.045 ;
        RECT 84.425 194.805 86.035 195.005 ;
        RECT 84.425 194.795 85.260 194.805 ;
        RECT 85.850 194.715 86.035 194.805 ;
        RECT 82.255 193.805 82.465 194.705 ;
        RECT 82.635 193.975 83.325 194.535 ;
        RECT 82.255 193.635 83.210 193.805 ;
        RECT 82.485 193.005 82.755 193.465 ;
        RECT 82.925 193.175 83.210 193.635 ;
        RECT 83.495 193.505 83.665 194.705 ;
        RECT 85.365 194.605 85.695 194.635 ;
        RECT 83.895 194.545 85.695 194.605 ;
        RECT 86.285 194.545 86.540 195.165 ;
        RECT 83.835 194.435 86.540 194.545 ;
        RECT 83.835 194.400 84.035 194.435 ;
        RECT 83.835 193.825 84.005 194.400 ;
        RECT 85.365 194.375 86.540 194.435 ;
        RECT 87.175 194.390 87.465 195.555 ;
        RECT 87.675 194.415 87.905 195.555 ;
        RECT 88.075 194.405 88.405 195.385 ;
        RECT 88.575 194.415 88.785 195.555 ;
        RECT 89.015 194.465 92.525 195.555 ;
        RECT 84.235 193.960 84.645 194.265 ;
        RECT 84.815 193.995 85.145 194.205 ;
        RECT 83.835 193.705 84.105 193.825 ;
        RECT 83.835 193.660 84.680 193.705 ;
        RECT 83.925 193.535 84.680 193.660 ;
        RECT 84.935 193.595 85.145 193.995 ;
        RECT 85.390 193.995 85.865 194.205 ;
        RECT 86.055 193.995 86.545 194.195 ;
        RECT 87.655 193.995 87.985 194.245 ;
        RECT 85.390 193.595 85.610 193.995 ;
        RECT 83.495 193.175 83.755 193.505 ;
        RECT 84.510 193.385 84.680 193.535 ;
        RECT 83.925 193.005 84.255 193.365 ;
        RECT 84.510 193.175 85.810 193.385 ;
        RECT 86.085 193.005 86.540 193.770 ;
        RECT 87.175 193.005 87.465 193.730 ;
        RECT 87.675 193.005 87.905 193.825 ;
        RECT 88.155 193.805 88.405 194.405 ;
        RECT 88.075 193.175 88.405 193.805 ;
        RECT 88.575 193.005 88.785 193.825 ;
        RECT 89.015 193.775 90.665 194.295 ;
        RECT 90.835 193.945 92.525 194.465 ;
        RECT 93.310 194.545 93.610 195.385 ;
        RECT 93.805 194.715 94.055 195.555 ;
        RECT 94.645 194.965 95.450 195.385 ;
        RECT 94.225 194.795 95.790 194.965 ;
        RECT 94.225 194.545 94.395 194.795 ;
        RECT 93.310 194.375 94.395 194.545 ;
        RECT 93.155 193.915 93.485 194.205 ;
        RECT 89.015 193.005 92.525 193.775 ;
        RECT 93.655 193.745 93.825 194.375 ;
        RECT 94.565 194.245 94.885 194.625 ;
        RECT 93.995 193.995 94.325 194.205 ;
        RECT 94.505 193.995 94.885 194.245 ;
        RECT 95.075 194.205 95.450 194.625 ;
        RECT 95.620 194.545 95.790 194.795 ;
        RECT 95.960 194.715 96.290 195.555 ;
        RECT 96.460 194.795 97.125 195.385 ;
        RECT 95.620 194.375 96.540 194.545 ;
        RECT 96.370 194.205 96.540 194.375 ;
        RECT 95.075 194.195 95.560 194.205 ;
        RECT 95.055 194.025 95.560 194.195 ;
        RECT 95.075 193.995 95.560 194.025 ;
        RECT 95.750 193.995 96.200 194.205 ;
        RECT 96.370 193.995 96.705 194.205 ;
        RECT 96.875 193.825 97.125 194.795 ;
        RECT 93.315 193.565 93.825 193.745 ;
        RECT 94.230 193.655 95.930 193.825 ;
        RECT 94.230 193.565 94.615 193.655 ;
        RECT 93.315 193.175 93.645 193.565 ;
        RECT 93.815 193.225 95.000 193.395 ;
        RECT 95.260 193.005 95.430 193.475 ;
        RECT 95.600 193.190 95.930 193.655 ;
        RECT 96.100 193.005 96.270 193.825 ;
        RECT 96.440 193.185 97.125 193.825 ;
        RECT 97.295 194.715 97.555 195.385 ;
        RECT 97.725 195.155 98.055 195.555 ;
        RECT 98.925 195.155 99.325 195.555 ;
        RECT 99.615 194.975 99.945 195.210 ;
        RECT 97.865 194.805 99.945 194.975 ;
        RECT 97.295 193.745 97.470 194.715 ;
        RECT 97.865 194.535 98.035 194.805 ;
        RECT 97.640 194.365 98.035 194.535 ;
        RECT 98.205 194.415 99.220 194.635 ;
        RECT 97.640 193.915 97.810 194.365 ;
        RECT 98.945 194.275 99.220 194.415 ;
        RECT 99.390 194.415 99.945 194.805 ;
        RECT 97.980 193.995 98.430 194.195 ;
        RECT 98.600 193.825 98.775 194.020 ;
        RECT 97.295 193.175 97.635 193.745 ;
        RECT 97.830 193.005 98.000 193.670 ;
        RECT 98.280 193.655 98.775 193.825 ;
        RECT 98.280 193.515 98.500 193.655 ;
        RECT 98.275 193.345 98.500 193.515 ;
        RECT 98.945 193.485 99.115 194.275 ;
        RECT 99.390 194.165 99.560 194.415 ;
        RECT 100.115 194.245 100.290 195.345 ;
        RECT 100.460 194.735 100.805 195.555 ;
        RECT 102.100 194.585 102.430 195.385 ;
        RECT 102.600 194.755 102.930 195.555 ;
        RECT 103.230 194.585 103.560 195.385 ;
        RECT 104.205 194.755 104.455 195.555 ;
        RECT 99.365 193.995 99.560 194.165 ;
        RECT 99.730 193.995 100.290 194.245 ;
        RECT 100.460 193.995 100.805 194.565 ;
        RECT 102.100 194.415 104.535 194.585 ;
        RECT 104.725 194.415 104.895 195.555 ;
        RECT 105.065 194.415 105.405 195.385 ;
        RECT 105.665 194.885 105.835 195.385 ;
        RECT 106.005 195.055 106.335 195.555 ;
        RECT 105.665 194.715 106.330 194.885 ;
        RECT 101.895 193.995 102.245 194.245 ;
        RECT 99.365 193.610 99.535 193.995 ;
        RECT 98.280 193.300 98.500 193.345 ;
        RECT 98.670 193.315 99.115 193.485 ;
        RECT 99.285 193.240 99.535 193.610 ;
        RECT 99.705 193.645 100.805 193.825 ;
        RECT 102.430 193.785 102.600 194.415 ;
        RECT 102.770 193.995 103.100 194.195 ;
        RECT 103.270 193.995 103.600 194.195 ;
        RECT 103.770 193.995 104.190 194.195 ;
        RECT 104.365 194.165 104.535 194.415 ;
        RECT 104.365 193.995 105.060 194.165 ;
        RECT 105.230 193.855 105.405 194.415 ;
        RECT 105.580 193.895 105.930 194.545 ;
        RECT 99.705 193.240 99.955 193.645 ;
        RECT 100.125 193.005 100.295 193.475 ;
        RECT 100.465 193.240 100.805 193.645 ;
        RECT 102.100 193.175 102.600 193.785 ;
        RECT 103.230 193.655 104.455 193.825 ;
        RECT 105.175 193.805 105.405 193.855 ;
        RECT 103.230 193.175 103.560 193.655 ;
        RECT 103.730 193.005 103.955 193.465 ;
        RECT 104.125 193.175 104.455 193.655 ;
        RECT 104.645 193.005 104.895 193.805 ;
        RECT 105.065 193.175 105.405 193.805 ;
        RECT 106.100 193.725 106.330 194.715 ;
        RECT 105.665 193.555 106.330 193.725 ;
        RECT 105.665 193.265 105.835 193.555 ;
        RECT 106.005 193.005 106.335 193.385 ;
        RECT 106.505 193.265 106.690 195.385 ;
        RECT 106.930 195.095 107.195 195.555 ;
        RECT 107.365 194.960 107.615 195.385 ;
        RECT 107.825 195.110 108.930 195.280 ;
        RECT 107.310 194.830 107.615 194.960 ;
        RECT 106.860 193.635 107.140 194.585 ;
        RECT 107.310 193.725 107.480 194.830 ;
        RECT 107.650 194.045 107.890 194.640 ;
        RECT 108.060 194.575 108.590 194.940 ;
        RECT 108.060 193.875 108.230 194.575 ;
        RECT 108.760 194.495 108.930 195.110 ;
        RECT 109.100 194.755 109.270 195.555 ;
        RECT 109.440 195.055 109.690 195.385 ;
        RECT 109.915 195.085 110.800 195.255 ;
        RECT 108.760 194.405 109.270 194.495 ;
        RECT 107.310 193.595 107.535 193.725 ;
        RECT 107.705 193.655 108.230 193.875 ;
        RECT 108.400 194.235 109.270 194.405 ;
        RECT 106.945 193.005 107.195 193.465 ;
        RECT 107.365 193.455 107.535 193.595 ;
        RECT 108.400 193.455 108.570 194.235 ;
        RECT 109.100 194.165 109.270 194.235 ;
        RECT 108.780 193.985 108.980 194.015 ;
        RECT 109.440 193.985 109.610 195.055 ;
        RECT 109.780 194.165 109.970 194.885 ;
        RECT 108.780 193.685 109.610 193.985 ;
        RECT 110.140 193.955 110.460 194.915 ;
        RECT 107.365 193.285 107.700 193.455 ;
        RECT 107.895 193.285 108.570 193.455 ;
        RECT 108.890 193.005 109.260 193.505 ;
        RECT 109.440 193.455 109.610 193.685 ;
        RECT 109.995 193.625 110.460 193.955 ;
        RECT 110.630 194.245 110.800 195.085 ;
        RECT 110.980 195.055 111.295 195.555 ;
        RECT 111.525 194.825 111.865 195.385 ;
        RECT 110.970 194.450 111.865 194.825 ;
        RECT 112.035 194.545 112.205 195.555 ;
        RECT 111.675 194.245 111.865 194.450 ;
        RECT 112.375 194.495 112.705 195.340 ;
        RECT 112.375 194.415 112.765 194.495 ;
        RECT 112.550 194.365 112.765 194.415 ;
        RECT 112.935 194.390 113.225 195.555 ;
        RECT 113.395 195.120 118.740 195.555 ;
        RECT 110.630 193.915 111.505 194.245 ;
        RECT 111.675 193.915 112.425 194.245 ;
        RECT 110.630 193.455 110.800 193.915 ;
        RECT 111.675 193.745 111.875 193.915 ;
        RECT 112.595 193.785 112.765 194.365 ;
        RECT 112.540 193.745 112.765 193.785 ;
        RECT 109.440 193.285 109.845 193.455 ;
        RECT 110.015 193.285 110.800 193.455 ;
        RECT 111.075 193.005 111.285 193.535 ;
        RECT 111.545 193.220 111.875 193.745 ;
        RECT 112.385 193.660 112.765 193.745 ;
        RECT 112.045 193.005 112.215 193.615 ;
        RECT 112.385 193.225 112.715 193.660 ;
        RECT 112.935 193.005 113.225 193.730 ;
        RECT 114.980 193.550 115.320 194.380 ;
        RECT 116.800 193.870 117.150 195.120 ;
        RECT 119.005 194.810 119.275 195.555 ;
        RECT 119.905 195.550 126.180 195.555 ;
        RECT 119.445 194.640 119.735 195.380 ;
        RECT 119.905 194.825 120.160 195.550 ;
        RECT 120.345 194.655 120.605 195.380 ;
        RECT 120.775 194.825 121.020 195.550 ;
        RECT 121.205 194.655 121.465 195.380 ;
        RECT 121.635 194.825 121.880 195.550 ;
        RECT 122.065 194.655 122.325 195.380 ;
        RECT 122.495 194.825 122.740 195.550 ;
        RECT 122.910 194.655 123.170 195.380 ;
        RECT 123.340 194.825 123.600 195.550 ;
        RECT 123.770 194.655 124.030 195.380 ;
        RECT 124.200 194.825 124.460 195.550 ;
        RECT 124.630 194.655 124.890 195.380 ;
        RECT 125.060 194.825 125.320 195.550 ;
        RECT 125.490 194.655 125.750 195.380 ;
        RECT 125.920 194.755 126.180 195.550 ;
        RECT 120.345 194.640 125.750 194.655 ;
        RECT 119.005 194.415 125.750 194.640 ;
        RECT 119.005 193.855 120.170 194.415 ;
        RECT 126.350 194.245 126.600 195.380 ;
        RECT 126.780 194.745 127.040 195.555 ;
        RECT 127.215 194.245 127.460 195.385 ;
        RECT 127.640 194.745 127.935 195.555 ;
        RECT 128.115 194.685 128.390 195.385 ;
        RECT 128.600 195.010 128.815 195.555 ;
        RECT 128.985 195.045 129.460 195.385 ;
        RECT 129.630 195.050 130.245 195.555 ;
        RECT 129.630 194.875 129.825 195.050 ;
        RECT 120.340 193.995 127.460 194.245 ;
        RECT 118.975 193.825 120.170 193.855 ;
        RECT 118.975 193.685 125.750 193.825 ;
        RECT 119.005 193.655 125.750 193.685 ;
        RECT 113.395 193.005 118.740 193.550 ;
        RECT 119.005 193.005 119.305 193.485 ;
        RECT 119.475 193.200 119.735 193.655 ;
        RECT 119.905 193.005 120.165 193.485 ;
        RECT 120.345 193.200 120.605 193.655 ;
        RECT 120.775 193.005 121.025 193.485 ;
        RECT 121.205 193.200 121.465 193.655 ;
        RECT 121.635 193.005 121.885 193.485 ;
        RECT 122.065 193.200 122.325 193.655 ;
        RECT 122.495 193.005 122.740 193.485 ;
        RECT 122.910 193.200 123.185 193.655 ;
        RECT 123.355 193.005 123.600 193.485 ;
        RECT 123.770 193.200 124.030 193.655 ;
        RECT 124.200 193.005 124.460 193.485 ;
        RECT 124.630 193.200 124.890 193.655 ;
        RECT 125.060 193.005 125.320 193.485 ;
        RECT 125.490 193.200 125.750 193.655 ;
        RECT 125.920 193.005 126.180 193.565 ;
        RECT 126.350 193.185 126.600 193.995 ;
        RECT 126.780 193.005 127.040 193.530 ;
        RECT 127.210 193.185 127.460 193.995 ;
        RECT 127.630 193.685 127.945 194.245 ;
        RECT 128.115 193.655 128.285 194.685 ;
        RECT 128.560 194.515 129.275 194.810 ;
        RECT 129.495 194.685 129.825 194.875 ;
        RECT 129.995 194.515 130.245 194.880 ;
        RECT 128.455 194.345 130.245 194.515 ;
        RECT 128.455 193.915 128.685 194.345 ;
        RECT 127.640 193.005 127.945 193.515 ;
        RECT 128.115 193.175 128.375 193.655 ;
        RECT 128.855 193.645 129.265 194.165 ;
        RECT 128.545 193.005 128.875 193.465 ;
        RECT 129.065 193.225 129.265 193.645 ;
        RECT 129.435 193.490 129.690 194.345 ;
        RECT 130.485 194.165 130.655 195.385 ;
        RECT 130.905 195.045 131.165 195.555 ;
        RECT 131.425 194.885 131.595 195.385 ;
        RECT 131.765 195.055 132.095 195.555 ;
        RECT 129.860 193.915 130.655 194.165 ;
        RECT 130.825 193.995 131.165 194.875 ;
        RECT 131.425 194.715 132.090 194.885 ;
        RECT 130.405 193.825 130.655 193.915 ;
        RECT 131.340 193.895 131.690 194.545 ;
        RECT 129.435 193.225 130.225 193.490 ;
        RECT 130.405 193.405 130.735 193.825 ;
        RECT 130.905 193.005 131.165 193.825 ;
        RECT 131.860 193.725 132.090 194.715 ;
        RECT 131.425 193.555 132.090 193.725 ;
        RECT 131.425 193.265 131.595 193.555 ;
        RECT 131.765 193.005 132.095 193.385 ;
        RECT 132.265 193.265 132.450 195.385 ;
        RECT 132.690 195.095 132.955 195.555 ;
        RECT 133.125 194.960 133.375 195.385 ;
        RECT 133.585 195.110 134.690 195.280 ;
        RECT 133.070 194.830 133.375 194.960 ;
        RECT 132.620 193.635 132.900 194.585 ;
        RECT 133.070 193.725 133.240 194.830 ;
        RECT 133.410 194.045 133.650 194.640 ;
        RECT 133.820 194.575 134.350 194.940 ;
        RECT 133.820 193.875 133.990 194.575 ;
        RECT 134.520 194.495 134.690 195.110 ;
        RECT 134.860 194.755 135.030 195.555 ;
        RECT 135.200 195.055 135.450 195.385 ;
        RECT 135.675 195.085 136.560 195.255 ;
        RECT 134.520 194.405 135.030 194.495 ;
        RECT 133.070 193.595 133.295 193.725 ;
        RECT 133.465 193.655 133.990 193.875 ;
        RECT 134.160 194.235 135.030 194.405 ;
        RECT 132.705 193.005 132.955 193.465 ;
        RECT 133.125 193.455 133.295 193.595 ;
        RECT 134.160 193.455 134.330 194.235 ;
        RECT 134.860 194.165 135.030 194.235 ;
        RECT 134.540 193.985 134.740 194.015 ;
        RECT 135.200 193.985 135.370 195.055 ;
        RECT 135.540 194.165 135.730 194.885 ;
        RECT 134.540 193.685 135.370 193.985 ;
        RECT 135.900 193.955 136.220 194.915 ;
        RECT 133.125 193.285 133.460 193.455 ;
        RECT 133.655 193.285 134.330 193.455 ;
        RECT 134.650 193.005 135.020 193.505 ;
        RECT 135.200 193.455 135.370 193.685 ;
        RECT 135.755 193.625 136.220 193.955 ;
        RECT 136.390 194.245 136.560 195.085 ;
        RECT 136.740 195.055 137.055 195.555 ;
        RECT 137.285 194.825 137.625 195.385 ;
        RECT 136.730 194.450 137.625 194.825 ;
        RECT 137.795 194.545 137.965 195.555 ;
        RECT 137.435 194.245 137.625 194.450 ;
        RECT 138.135 194.495 138.465 195.340 ;
        RECT 138.135 194.415 138.525 194.495 ;
        RECT 138.310 194.365 138.525 194.415 ;
        RECT 138.695 194.390 138.985 195.555 ;
        RECT 139.160 194.605 139.425 195.375 ;
        RECT 139.595 194.835 139.925 195.555 ;
        RECT 140.115 195.015 140.375 195.375 ;
        RECT 140.545 195.185 140.875 195.555 ;
        RECT 141.045 195.015 141.305 195.375 ;
        RECT 140.115 194.785 141.305 195.015 ;
        RECT 141.875 194.605 142.165 195.375 ;
        RECT 136.390 193.915 137.265 194.245 ;
        RECT 137.435 193.915 138.185 194.245 ;
        RECT 136.390 193.455 136.560 193.915 ;
        RECT 137.435 193.745 137.635 193.915 ;
        RECT 138.355 193.785 138.525 194.365 ;
        RECT 138.300 193.745 138.525 193.785 ;
        RECT 135.200 193.285 135.605 193.455 ;
        RECT 135.775 193.285 136.560 193.455 ;
        RECT 136.835 193.005 137.045 193.535 ;
        RECT 137.305 193.220 137.635 193.745 ;
        RECT 138.145 193.660 138.525 193.745 ;
        RECT 137.805 193.005 137.975 193.615 ;
        RECT 138.145 193.225 138.475 193.660 ;
        RECT 138.695 193.005 138.985 193.730 ;
        RECT 139.160 193.185 139.495 194.605 ;
        RECT 139.670 194.425 142.165 194.605 ;
        RECT 143.020 194.585 143.410 194.760 ;
        RECT 143.895 194.755 144.225 195.555 ;
        RECT 144.395 194.765 144.930 195.385 ;
        RECT 145.135 195.045 145.395 195.555 ;
        RECT 139.670 193.735 139.895 194.425 ;
        RECT 143.020 194.415 144.445 194.585 ;
        RECT 140.095 193.915 140.375 194.245 ;
        RECT 140.555 193.915 141.130 194.245 ;
        RECT 141.310 193.915 141.745 194.245 ;
        RECT 141.925 193.915 142.195 194.245 ;
        RECT 139.670 193.545 142.155 193.735 ;
        RECT 142.895 193.685 143.250 194.245 ;
        RECT 139.675 193.005 140.420 193.375 ;
        RECT 140.985 193.185 141.240 193.545 ;
        RECT 141.420 193.005 141.750 193.375 ;
        RECT 141.930 193.185 142.155 193.545 ;
        RECT 143.420 193.515 143.590 194.415 ;
        RECT 143.760 193.685 144.025 194.245 ;
        RECT 144.275 193.915 144.445 194.415 ;
        RECT 144.615 193.745 144.930 194.765 ;
        RECT 145.135 193.995 145.475 194.875 ;
        RECT 145.645 194.165 145.815 195.385 ;
        RECT 146.055 195.050 146.670 195.555 ;
        RECT 146.055 194.515 146.305 194.880 ;
        RECT 146.475 194.875 146.670 195.050 ;
        RECT 146.840 195.045 147.315 195.385 ;
        RECT 147.485 195.010 147.700 195.555 ;
        RECT 146.475 194.685 146.805 194.875 ;
        RECT 147.025 194.515 147.740 194.810 ;
        RECT 147.910 194.685 148.185 195.385 ;
        RECT 146.055 194.345 147.845 194.515 ;
        RECT 145.645 193.915 146.440 194.165 ;
        RECT 145.645 193.825 145.895 193.915 ;
        RECT 143.000 193.005 143.240 193.515 ;
        RECT 143.420 193.185 143.700 193.515 ;
        RECT 143.930 193.005 144.145 193.515 ;
        RECT 144.315 193.175 144.930 193.745 ;
        RECT 145.135 193.005 145.395 193.825 ;
        RECT 145.565 193.405 145.895 193.825 ;
        RECT 146.610 193.490 146.865 194.345 ;
        RECT 146.075 193.225 146.865 193.490 ;
        RECT 147.035 193.645 147.445 194.165 ;
        RECT 147.615 193.915 147.845 194.345 ;
        RECT 148.015 193.655 148.185 194.685 ;
        RECT 148.415 194.495 148.745 195.340 ;
        RECT 148.915 194.545 149.085 195.555 ;
        RECT 149.255 194.825 149.595 195.385 ;
        RECT 149.825 195.055 150.140 195.555 ;
        RECT 150.320 195.085 151.205 195.255 ;
        RECT 148.355 194.415 148.745 194.495 ;
        RECT 149.255 194.450 150.150 194.825 ;
        RECT 148.355 194.365 148.570 194.415 ;
        RECT 148.355 193.785 148.525 194.365 ;
        RECT 149.255 194.245 149.445 194.450 ;
        RECT 150.320 194.245 150.490 195.085 ;
        RECT 151.430 195.055 151.680 195.385 ;
        RECT 148.695 193.915 149.445 194.245 ;
        RECT 149.615 193.915 150.490 194.245 ;
        RECT 148.355 193.745 148.580 193.785 ;
        RECT 149.245 193.745 149.445 193.915 ;
        RECT 148.355 193.660 148.735 193.745 ;
        RECT 147.035 193.225 147.235 193.645 ;
        RECT 147.425 193.005 147.755 193.465 ;
        RECT 147.925 193.175 148.185 193.655 ;
        RECT 148.405 193.225 148.735 193.660 ;
        RECT 148.905 193.005 149.075 193.615 ;
        RECT 149.245 193.220 149.575 193.745 ;
        RECT 149.835 193.005 150.045 193.535 ;
        RECT 150.320 193.455 150.490 193.915 ;
        RECT 150.660 193.955 150.980 194.915 ;
        RECT 151.150 194.165 151.340 194.885 ;
        RECT 151.510 193.985 151.680 195.055 ;
        RECT 151.850 194.755 152.020 195.555 ;
        RECT 152.190 195.110 153.295 195.280 ;
        RECT 152.190 194.495 152.360 195.110 ;
        RECT 153.505 194.960 153.755 195.385 ;
        RECT 153.925 195.095 154.190 195.555 ;
        RECT 152.530 194.575 153.060 194.940 ;
        RECT 153.505 194.830 153.810 194.960 ;
        RECT 151.850 194.405 152.360 194.495 ;
        RECT 151.850 194.235 152.720 194.405 ;
        RECT 151.850 194.165 152.020 194.235 ;
        RECT 152.140 193.985 152.340 194.015 ;
        RECT 150.660 193.625 151.125 193.955 ;
        RECT 151.510 193.685 152.340 193.985 ;
        RECT 151.510 193.455 151.680 193.685 ;
        RECT 150.320 193.285 151.105 193.455 ;
        RECT 151.275 193.285 151.680 193.455 ;
        RECT 151.860 193.005 152.230 193.505 ;
        RECT 152.550 193.455 152.720 194.235 ;
        RECT 152.890 193.875 153.060 194.575 ;
        RECT 153.230 194.045 153.470 194.640 ;
        RECT 152.890 193.655 153.415 193.875 ;
        RECT 153.640 193.725 153.810 194.830 ;
        RECT 153.585 193.595 153.810 193.725 ;
        RECT 153.980 193.635 154.260 194.585 ;
        RECT 153.585 193.455 153.755 193.595 ;
        RECT 152.550 193.285 153.225 193.455 ;
        RECT 153.420 193.285 153.755 193.455 ;
        RECT 153.925 193.005 154.175 193.465 ;
        RECT 154.430 193.265 154.615 195.385 ;
        RECT 154.785 195.055 155.115 195.555 ;
        RECT 155.285 194.885 155.455 195.385 ;
        RECT 154.790 194.715 155.455 194.885 ;
        RECT 154.790 193.725 155.020 194.715 ;
        RECT 155.190 193.895 155.540 194.545 ;
        RECT 155.715 194.465 156.925 195.555 ;
        RECT 155.715 193.925 156.235 194.465 ;
        RECT 156.405 193.755 156.925 194.295 ;
        RECT 154.790 193.555 155.455 193.725 ;
        RECT 154.785 193.005 155.115 193.385 ;
        RECT 155.285 193.265 155.455 193.555 ;
        RECT 155.715 193.005 156.925 193.755 ;
        RECT 22.690 192.835 157.010 193.005 ;
        RECT 22.775 192.085 23.985 192.835 ;
        RECT 24.155 192.290 29.500 192.835 ;
        RECT 22.775 191.545 23.295 192.085 ;
        RECT 23.465 191.375 23.985 191.915 ;
        RECT 25.740 191.460 26.080 192.290 ;
        RECT 29.675 192.085 30.885 192.835 ;
        RECT 31.145 192.285 31.315 192.575 ;
        RECT 31.485 192.455 31.815 192.835 ;
        RECT 31.145 192.115 31.810 192.285 ;
        RECT 22.775 190.285 23.985 191.375 ;
        RECT 27.560 190.720 27.910 191.970 ;
        RECT 29.675 191.545 30.195 192.085 ;
        RECT 30.365 191.375 30.885 191.915 ;
        RECT 24.155 190.285 29.500 190.720 ;
        RECT 29.675 190.285 30.885 191.375 ;
        RECT 31.060 191.295 31.410 191.945 ;
        RECT 31.580 191.125 31.810 192.115 ;
        RECT 31.145 190.955 31.810 191.125 ;
        RECT 31.145 190.455 31.315 190.955 ;
        RECT 31.485 190.285 31.815 190.785 ;
        RECT 31.985 190.455 32.170 192.575 ;
        RECT 32.425 192.375 32.675 192.835 ;
        RECT 32.845 192.385 33.180 192.555 ;
        RECT 33.375 192.385 34.050 192.555 ;
        RECT 32.845 192.245 33.015 192.385 ;
        RECT 32.340 191.255 32.620 192.205 ;
        RECT 32.790 192.115 33.015 192.245 ;
        RECT 32.790 191.010 32.960 192.115 ;
        RECT 33.185 191.965 33.710 192.185 ;
        RECT 33.130 191.200 33.370 191.795 ;
        RECT 33.540 191.265 33.710 191.965 ;
        RECT 33.880 191.605 34.050 192.385 ;
        RECT 34.370 192.335 34.740 192.835 ;
        RECT 34.920 192.385 35.325 192.555 ;
        RECT 35.495 192.385 36.280 192.555 ;
        RECT 34.920 192.155 35.090 192.385 ;
        RECT 34.260 191.855 35.090 192.155 ;
        RECT 35.475 191.885 35.940 192.215 ;
        RECT 34.260 191.825 34.460 191.855 ;
        RECT 34.580 191.605 34.750 191.675 ;
        RECT 33.880 191.435 34.750 191.605 ;
        RECT 34.240 191.345 34.750 191.435 ;
        RECT 32.790 190.880 33.095 191.010 ;
        RECT 33.540 190.900 34.070 191.265 ;
        RECT 32.410 190.285 32.675 190.745 ;
        RECT 32.845 190.455 33.095 190.880 ;
        RECT 34.240 190.730 34.410 191.345 ;
        RECT 33.305 190.560 34.410 190.730 ;
        RECT 34.580 190.285 34.750 191.085 ;
        RECT 34.920 190.785 35.090 191.855 ;
        RECT 35.260 190.955 35.450 191.675 ;
        RECT 35.620 190.925 35.940 191.885 ;
        RECT 36.110 191.925 36.280 192.385 ;
        RECT 36.555 192.305 36.765 192.835 ;
        RECT 37.025 192.095 37.355 192.620 ;
        RECT 37.525 192.225 37.695 192.835 ;
        RECT 37.865 192.180 38.195 192.615 ;
        RECT 38.415 192.185 38.675 192.665 ;
        RECT 38.845 192.295 39.095 192.835 ;
        RECT 37.865 192.095 38.245 192.180 ;
        RECT 37.155 191.925 37.355 192.095 ;
        RECT 38.020 192.055 38.245 192.095 ;
        RECT 36.110 191.595 36.985 191.925 ;
        RECT 37.155 191.595 37.905 191.925 ;
        RECT 34.920 190.455 35.170 190.785 ;
        RECT 36.110 190.755 36.280 191.595 ;
        RECT 37.155 191.390 37.345 191.595 ;
        RECT 38.075 191.475 38.245 192.055 ;
        RECT 38.030 191.425 38.245 191.475 ;
        RECT 36.450 191.015 37.345 191.390 ;
        RECT 37.855 191.345 38.245 191.425 ;
        RECT 35.395 190.585 36.280 190.755 ;
        RECT 36.460 190.285 36.775 190.785 ;
        RECT 37.005 190.455 37.345 191.015 ;
        RECT 37.515 190.285 37.685 191.295 ;
        RECT 37.855 190.500 38.185 191.345 ;
        RECT 38.415 191.155 38.585 192.185 ;
        RECT 39.265 192.130 39.485 192.615 ;
        RECT 38.755 191.535 38.985 191.930 ;
        RECT 39.155 191.705 39.485 192.130 ;
        RECT 39.655 192.455 40.545 192.625 ;
        RECT 39.655 191.730 39.825 192.455 ;
        RECT 39.995 191.900 40.545 192.285 ;
        RECT 40.750 192.095 41.365 192.665 ;
        RECT 41.535 192.325 41.750 192.835 ;
        RECT 41.980 192.325 42.260 192.655 ;
        RECT 42.440 192.325 42.680 192.835 ;
        RECT 39.655 191.660 40.545 191.730 ;
        RECT 39.650 191.635 40.545 191.660 ;
        RECT 39.640 191.620 40.545 191.635 ;
        RECT 39.635 191.605 40.545 191.620 ;
        RECT 39.625 191.600 40.545 191.605 ;
        RECT 39.620 191.590 40.545 191.600 ;
        RECT 39.615 191.580 40.545 191.590 ;
        RECT 39.605 191.575 40.545 191.580 ;
        RECT 39.595 191.565 40.545 191.575 ;
        RECT 39.585 191.560 40.545 191.565 ;
        RECT 39.585 191.555 39.920 191.560 ;
        RECT 39.570 191.550 39.920 191.555 ;
        RECT 39.555 191.540 39.920 191.550 ;
        RECT 39.530 191.535 39.920 191.540 ;
        RECT 38.755 191.530 39.920 191.535 ;
        RECT 38.755 191.495 39.890 191.530 ;
        RECT 38.755 191.470 39.855 191.495 ;
        RECT 38.755 191.440 39.825 191.470 ;
        RECT 38.755 191.410 39.805 191.440 ;
        RECT 38.755 191.380 39.785 191.410 ;
        RECT 38.755 191.370 39.715 191.380 ;
        RECT 38.755 191.360 39.690 191.370 ;
        RECT 38.755 191.345 39.670 191.360 ;
        RECT 38.755 191.330 39.650 191.345 ;
        RECT 38.860 191.320 39.645 191.330 ;
        RECT 38.860 191.285 39.630 191.320 ;
        RECT 38.415 190.455 38.690 191.155 ;
        RECT 38.860 191.035 39.615 191.285 ;
        RECT 39.785 190.965 40.115 191.210 ;
        RECT 40.285 191.110 40.545 191.560 ;
        RECT 39.930 190.940 40.115 190.965 ;
        RECT 40.750 191.075 41.065 192.095 ;
        RECT 41.235 191.425 41.405 191.925 ;
        RECT 41.655 191.595 41.920 192.155 ;
        RECT 42.090 191.425 42.260 192.325 ;
        RECT 42.430 191.595 42.785 192.155 ;
        RECT 43.015 192.035 43.710 192.665 ;
        RECT 43.915 192.035 44.225 192.835 ;
        RECT 44.395 192.065 46.065 192.835 ;
        RECT 46.325 192.285 46.495 192.665 ;
        RECT 46.675 192.455 47.005 192.835 ;
        RECT 46.325 192.115 46.990 192.285 ;
        RECT 47.185 192.160 47.445 192.665 ;
        RECT 43.035 191.595 43.370 191.845 ;
        RECT 43.540 191.475 43.710 192.035 ;
        RECT 43.880 191.595 44.215 191.865 ;
        RECT 44.395 191.545 45.145 192.065 ;
        RECT 43.535 191.435 43.710 191.475 ;
        RECT 41.235 191.255 42.660 191.425 ;
        RECT 39.930 190.840 40.545 190.940 ;
        RECT 38.860 190.285 39.115 190.830 ;
        RECT 39.285 190.455 39.765 190.795 ;
        RECT 39.940 190.285 40.545 190.840 ;
        RECT 40.750 190.455 41.285 191.075 ;
        RECT 41.455 190.285 41.785 191.085 ;
        RECT 42.270 191.080 42.660 191.255 ;
        RECT 43.015 190.285 43.275 191.425 ;
        RECT 43.445 190.455 43.775 191.435 ;
        RECT 43.945 190.285 44.225 191.425 ;
        RECT 45.315 191.375 46.065 191.895 ;
        RECT 46.255 191.565 46.585 191.935 ;
        RECT 46.820 191.860 46.990 192.115 ;
        RECT 46.820 191.530 47.105 191.860 ;
        RECT 46.820 191.385 46.990 191.530 ;
        RECT 44.395 190.285 46.065 191.375 ;
        RECT 46.325 191.215 46.990 191.385 ;
        RECT 47.275 191.360 47.445 192.160 ;
        RECT 48.535 192.110 48.825 192.835 ;
        RECT 49.085 192.285 49.255 192.575 ;
        RECT 49.425 192.455 49.755 192.835 ;
        RECT 49.085 192.115 49.750 192.285 ;
        RECT 46.325 190.455 46.495 191.215 ;
        RECT 46.675 190.285 47.005 191.045 ;
        RECT 47.175 190.455 47.445 191.360 ;
        RECT 48.535 190.285 48.825 191.450 ;
        RECT 49.000 191.295 49.350 191.945 ;
        RECT 49.520 191.125 49.750 192.115 ;
        RECT 49.085 190.955 49.750 191.125 ;
        RECT 49.085 190.455 49.255 190.955 ;
        RECT 49.425 190.285 49.755 190.785 ;
        RECT 49.925 190.455 50.110 192.575 ;
        RECT 50.365 192.375 50.615 192.835 ;
        RECT 50.785 192.385 51.120 192.555 ;
        RECT 51.315 192.385 51.990 192.555 ;
        RECT 50.785 192.245 50.955 192.385 ;
        RECT 50.280 191.255 50.560 192.205 ;
        RECT 50.730 192.115 50.955 192.245 ;
        RECT 50.730 191.010 50.900 192.115 ;
        RECT 51.125 191.965 51.650 192.185 ;
        RECT 51.070 191.200 51.310 191.795 ;
        RECT 51.480 191.265 51.650 191.965 ;
        RECT 51.820 191.605 51.990 192.385 ;
        RECT 52.310 192.335 52.680 192.835 ;
        RECT 52.860 192.385 53.265 192.555 ;
        RECT 53.435 192.385 54.220 192.555 ;
        RECT 52.860 192.155 53.030 192.385 ;
        RECT 52.200 191.855 53.030 192.155 ;
        RECT 53.415 191.885 53.880 192.215 ;
        RECT 52.200 191.825 52.400 191.855 ;
        RECT 52.520 191.605 52.690 191.675 ;
        RECT 51.820 191.435 52.690 191.605 ;
        RECT 52.180 191.345 52.690 191.435 ;
        RECT 50.730 190.880 51.035 191.010 ;
        RECT 51.480 190.900 52.010 191.265 ;
        RECT 50.350 190.285 50.615 190.745 ;
        RECT 50.785 190.455 51.035 190.880 ;
        RECT 52.180 190.730 52.350 191.345 ;
        RECT 51.245 190.560 52.350 190.730 ;
        RECT 52.520 190.285 52.690 191.085 ;
        RECT 52.860 190.785 53.030 191.855 ;
        RECT 53.200 190.955 53.390 191.675 ;
        RECT 53.560 190.925 53.880 191.885 ;
        RECT 54.050 191.925 54.220 192.385 ;
        RECT 54.495 192.305 54.705 192.835 ;
        RECT 54.965 192.095 55.295 192.620 ;
        RECT 55.465 192.225 55.635 192.835 ;
        RECT 55.805 192.180 56.135 192.615 ;
        RECT 55.805 192.095 56.185 192.180 ;
        RECT 55.095 191.925 55.295 192.095 ;
        RECT 55.960 192.055 56.185 192.095 ;
        RECT 54.050 191.595 54.925 191.925 ;
        RECT 55.095 191.595 55.845 191.925 ;
        RECT 52.860 190.455 53.110 190.785 ;
        RECT 54.050 190.755 54.220 191.595 ;
        RECT 55.095 191.390 55.285 191.595 ;
        RECT 56.015 191.475 56.185 192.055 ;
        RECT 55.970 191.425 56.185 191.475 ;
        RECT 54.390 191.015 55.285 191.390 ;
        RECT 55.795 191.345 56.185 191.425 ;
        RECT 53.335 190.585 54.220 190.755 ;
        RECT 54.400 190.285 54.715 190.785 ;
        RECT 54.945 190.455 55.285 191.015 ;
        RECT 55.455 190.285 55.625 191.295 ;
        RECT 55.795 190.500 56.125 191.345 ;
        RECT 57.275 190.455 57.555 192.555 ;
        RECT 57.785 192.375 57.955 192.835 ;
        RECT 58.225 192.445 59.475 192.625 ;
        RECT 58.610 192.205 58.975 192.275 ;
        RECT 57.725 192.025 58.975 192.205 ;
        RECT 59.145 192.225 59.475 192.445 ;
        RECT 59.645 192.395 59.815 192.835 ;
        RECT 59.985 192.225 60.325 192.640 ;
        RECT 59.145 192.055 60.325 192.225 ;
        RECT 61.420 192.070 61.875 192.835 ;
        RECT 62.150 192.455 63.450 192.665 ;
        RECT 63.705 192.475 64.035 192.835 ;
        RECT 63.280 192.305 63.450 192.455 ;
        RECT 64.205 192.335 64.465 192.665 ;
        RECT 64.235 192.325 64.465 192.335 ;
        RECT 57.725 191.425 58.000 192.025 ;
        RECT 62.350 191.845 62.570 192.245 ;
        RECT 58.170 191.595 58.525 191.845 ;
        RECT 58.720 191.815 59.185 191.845 ;
        RECT 58.715 191.645 59.185 191.815 ;
        RECT 58.720 191.595 59.185 191.645 ;
        RECT 59.355 191.595 59.685 191.845 ;
        RECT 59.860 191.645 60.325 191.845 ;
        RECT 61.415 191.645 61.905 191.845 ;
        RECT 62.095 191.635 62.570 191.845 ;
        RECT 62.815 191.845 63.025 192.245 ;
        RECT 63.280 192.180 64.035 192.305 ;
        RECT 63.280 192.135 64.125 192.180 ;
        RECT 63.855 192.015 64.125 192.135 ;
        RECT 62.815 191.635 63.145 191.845 ;
        RECT 59.505 191.475 59.685 191.595 ;
        RECT 63.315 191.575 63.725 191.880 ;
        RECT 57.725 191.215 59.335 191.425 ;
        RECT 59.505 191.305 59.835 191.475 ;
        RECT 58.925 191.115 59.335 191.215 ;
        RECT 57.745 190.285 58.530 191.045 ;
        RECT 58.925 190.455 59.310 191.115 ;
        RECT 59.635 190.515 59.835 191.305 ;
        RECT 60.005 190.285 60.325 191.465 ;
        RECT 61.420 191.405 62.595 191.465 ;
        RECT 63.955 191.440 64.125 192.015 ;
        RECT 63.925 191.405 64.125 191.440 ;
        RECT 61.420 191.295 64.125 191.405 ;
        RECT 61.420 190.675 61.675 191.295 ;
        RECT 62.265 191.235 64.065 191.295 ;
        RECT 62.265 191.205 62.595 191.235 ;
        RECT 64.295 191.135 64.465 192.325 ;
        RECT 64.750 192.205 65.035 192.665 ;
        RECT 65.205 192.375 65.475 192.835 ;
        RECT 64.750 192.035 65.705 192.205 ;
        RECT 64.635 191.305 65.325 191.865 ;
        RECT 65.495 191.135 65.705 192.035 ;
        RECT 61.925 191.035 62.110 191.125 ;
        RECT 62.700 191.035 63.535 191.045 ;
        RECT 61.925 190.835 63.535 191.035 ;
        RECT 61.925 190.795 62.155 190.835 ;
        RECT 61.420 190.455 61.755 190.675 ;
        RECT 62.760 190.285 63.115 190.665 ;
        RECT 63.285 190.455 63.535 190.835 ;
        RECT 63.785 190.285 64.035 191.065 ;
        RECT 64.205 190.455 64.465 191.135 ;
        RECT 64.750 190.915 65.705 191.135 ;
        RECT 65.875 191.865 66.275 192.665 ;
        RECT 66.465 192.205 66.745 192.665 ;
        RECT 67.265 192.375 67.590 192.835 ;
        RECT 66.465 192.035 67.590 192.205 ;
        RECT 67.760 192.095 68.145 192.665 ;
        RECT 67.140 191.925 67.590 192.035 ;
        RECT 65.875 191.305 66.970 191.865 ;
        RECT 67.140 191.595 67.695 191.925 ;
        RECT 64.750 190.455 65.035 190.915 ;
        RECT 65.205 190.285 65.475 190.745 ;
        RECT 65.875 190.455 66.275 191.305 ;
        RECT 67.140 191.135 67.590 191.595 ;
        RECT 67.865 191.425 68.145 192.095 ;
        RECT 66.465 190.915 67.590 191.135 ;
        RECT 66.465 190.455 66.745 190.915 ;
        RECT 67.265 190.285 67.590 190.745 ;
        RECT 67.760 190.455 68.145 191.425 ;
        RECT 68.315 192.335 68.575 192.665 ;
        RECT 68.745 192.475 69.075 192.835 ;
        RECT 69.330 192.455 70.630 192.665 ;
        RECT 68.315 192.325 68.545 192.335 ;
        RECT 68.315 191.135 68.485 192.325 ;
        RECT 69.330 192.305 69.500 192.455 ;
        RECT 68.745 192.180 69.500 192.305 ;
        RECT 68.655 192.135 69.500 192.180 ;
        RECT 68.655 192.015 68.925 192.135 ;
        RECT 68.655 191.440 68.825 192.015 ;
        RECT 69.055 191.575 69.465 191.880 ;
        RECT 69.755 191.845 69.965 192.245 ;
        RECT 69.635 191.635 69.965 191.845 ;
        RECT 70.210 191.845 70.430 192.245 ;
        RECT 70.905 192.070 71.360 192.835 ;
        RECT 71.595 192.015 71.805 192.835 ;
        RECT 71.975 192.035 72.305 192.665 ;
        RECT 70.210 191.635 70.685 191.845 ;
        RECT 70.875 191.645 71.365 191.845 ;
        RECT 68.655 191.405 68.855 191.440 ;
        RECT 70.185 191.405 71.360 191.465 ;
        RECT 71.975 191.435 72.225 192.035 ;
        RECT 72.475 192.015 72.705 192.835 ;
        RECT 72.915 192.085 74.125 192.835 ;
        RECT 74.295 192.110 74.585 192.835 ;
        RECT 74.845 192.285 75.015 192.575 ;
        RECT 75.185 192.455 75.515 192.835 ;
        RECT 74.845 192.115 75.510 192.285 ;
        RECT 72.395 191.595 72.725 191.845 ;
        RECT 72.915 191.545 73.435 192.085 ;
        RECT 68.655 191.295 71.360 191.405 ;
        RECT 68.715 191.235 70.515 191.295 ;
        RECT 70.185 191.205 70.515 191.235 ;
        RECT 68.315 190.455 68.575 191.135 ;
        RECT 68.745 190.285 68.995 191.065 ;
        RECT 69.245 191.035 70.080 191.045 ;
        RECT 70.670 191.035 70.855 191.125 ;
        RECT 69.245 190.835 70.855 191.035 ;
        RECT 69.245 190.455 69.495 190.835 ;
        RECT 70.625 190.795 70.855 190.835 ;
        RECT 71.105 190.675 71.360 191.295 ;
        RECT 69.665 190.285 70.020 190.665 ;
        RECT 71.025 190.455 71.360 190.675 ;
        RECT 71.595 190.285 71.805 191.425 ;
        RECT 71.975 190.455 72.305 191.435 ;
        RECT 72.475 190.285 72.705 191.425 ;
        RECT 73.605 191.375 74.125 191.915 ;
        RECT 72.915 190.285 74.125 191.375 ;
        RECT 74.295 190.285 74.585 191.450 ;
        RECT 74.760 191.295 75.110 191.945 ;
        RECT 75.280 191.125 75.510 192.115 ;
        RECT 74.845 190.955 75.510 191.125 ;
        RECT 74.845 190.455 75.015 190.955 ;
        RECT 75.185 190.285 75.515 190.785 ;
        RECT 75.685 190.455 75.870 192.575 ;
        RECT 76.125 192.375 76.375 192.835 ;
        RECT 76.545 192.385 76.880 192.555 ;
        RECT 77.075 192.385 77.750 192.555 ;
        RECT 76.545 192.245 76.715 192.385 ;
        RECT 76.040 191.255 76.320 192.205 ;
        RECT 76.490 192.115 76.715 192.245 ;
        RECT 76.490 191.010 76.660 192.115 ;
        RECT 76.885 191.965 77.410 192.185 ;
        RECT 76.830 191.200 77.070 191.795 ;
        RECT 77.240 191.265 77.410 191.965 ;
        RECT 77.580 191.605 77.750 192.385 ;
        RECT 78.070 192.335 78.440 192.835 ;
        RECT 78.620 192.385 79.025 192.555 ;
        RECT 79.195 192.385 79.980 192.555 ;
        RECT 78.620 192.155 78.790 192.385 ;
        RECT 77.960 191.855 78.790 192.155 ;
        RECT 79.175 191.885 79.640 192.215 ;
        RECT 77.960 191.825 78.160 191.855 ;
        RECT 78.280 191.605 78.450 191.675 ;
        RECT 77.580 191.435 78.450 191.605 ;
        RECT 77.940 191.345 78.450 191.435 ;
        RECT 76.490 190.880 76.795 191.010 ;
        RECT 77.240 190.900 77.770 191.265 ;
        RECT 76.110 190.285 76.375 190.745 ;
        RECT 76.545 190.455 76.795 190.880 ;
        RECT 77.940 190.730 78.110 191.345 ;
        RECT 77.005 190.560 78.110 190.730 ;
        RECT 78.280 190.285 78.450 191.085 ;
        RECT 78.620 190.785 78.790 191.855 ;
        RECT 78.960 190.955 79.150 191.675 ;
        RECT 79.320 190.925 79.640 191.885 ;
        RECT 79.810 191.925 79.980 192.385 ;
        RECT 80.255 192.305 80.465 192.835 ;
        RECT 80.725 192.095 81.055 192.620 ;
        RECT 81.225 192.225 81.395 192.835 ;
        RECT 81.565 192.180 81.895 192.615 ;
        RECT 81.565 192.095 81.945 192.180 ;
        RECT 80.855 191.925 81.055 192.095 ;
        RECT 81.720 192.055 81.945 192.095 ;
        RECT 79.810 191.595 80.685 191.925 ;
        RECT 80.855 191.595 81.605 191.925 ;
        RECT 78.620 190.455 78.870 190.785 ;
        RECT 79.810 190.755 79.980 191.595 ;
        RECT 80.855 191.390 81.045 191.595 ;
        RECT 81.775 191.475 81.945 192.055 ;
        RECT 82.115 192.065 83.785 192.835 ;
        RECT 84.045 192.285 84.215 192.575 ;
        RECT 84.385 192.455 84.715 192.835 ;
        RECT 84.045 192.115 84.710 192.285 ;
        RECT 82.115 191.545 82.865 192.065 ;
        RECT 81.730 191.425 81.945 191.475 ;
        RECT 80.150 191.015 81.045 191.390 ;
        RECT 81.555 191.345 81.945 191.425 ;
        RECT 83.035 191.375 83.785 191.895 ;
        RECT 79.095 190.585 79.980 190.755 ;
        RECT 80.160 190.285 80.475 190.785 ;
        RECT 80.705 190.455 81.045 191.015 ;
        RECT 81.215 190.285 81.385 191.295 ;
        RECT 81.555 190.500 81.885 191.345 ;
        RECT 82.115 190.285 83.785 191.375 ;
        RECT 83.960 191.295 84.310 191.945 ;
        RECT 84.480 191.125 84.710 192.115 ;
        RECT 84.045 190.955 84.710 191.125 ;
        RECT 84.045 190.455 84.215 190.955 ;
        RECT 84.385 190.285 84.715 190.785 ;
        RECT 84.885 190.455 85.070 192.575 ;
        RECT 85.325 192.375 85.575 192.835 ;
        RECT 85.745 192.385 86.080 192.555 ;
        RECT 86.275 192.385 86.950 192.555 ;
        RECT 85.745 192.245 85.915 192.385 ;
        RECT 85.240 191.255 85.520 192.205 ;
        RECT 85.690 192.115 85.915 192.245 ;
        RECT 85.690 191.010 85.860 192.115 ;
        RECT 86.085 191.965 86.610 192.185 ;
        RECT 86.030 191.200 86.270 191.795 ;
        RECT 86.440 191.265 86.610 191.965 ;
        RECT 86.780 191.605 86.950 192.385 ;
        RECT 87.270 192.335 87.640 192.835 ;
        RECT 87.820 192.385 88.225 192.555 ;
        RECT 88.395 192.385 89.180 192.555 ;
        RECT 87.820 192.155 87.990 192.385 ;
        RECT 87.160 191.855 87.990 192.155 ;
        RECT 88.375 191.885 88.840 192.215 ;
        RECT 87.160 191.825 87.360 191.855 ;
        RECT 87.480 191.605 87.650 191.675 ;
        RECT 86.780 191.435 87.650 191.605 ;
        RECT 87.140 191.345 87.650 191.435 ;
        RECT 85.690 190.880 85.995 191.010 ;
        RECT 86.440 190.900 86.970 191.265 ;
        RECT 85.310 190.285 85.575 190.745 ;
        RECT 85.745 190.455 85.995 190.880 ;
        RECT 87.140 190.730 87.310 191.345 ;
        RECT 86.205 190.560 87.310 190.730 ;
        RECT 87.480 190.285 87.650 191.085 ;
        RECT 87.820 190.785 87.990 191.855 ;
        RECT 88.160 190.955 88.350 191.675 ;
        RECT 88.520 190.925 88.840 191.885 ;
        RECT 89.010 191.925 89.180 192.385 ;
        RECT 89.455 192.305 89.665 192.835 ;
        RECT 89.925 192.095 90.255 192.620 ;
        RECT 90.425 192.225 90.595 192.835 ;
        RECT 90.765 192.180 91.095 192.615 ;
        RECT 92.235 192.195 92.575 192.600 ;
        RECT 92.745 192.365 92.915 192.835 ;
        RECT 93.085 192.195 93.335 192.600 ;
        RECT 90.765 192.095 91.145 192.180 ;
        RECT 90.055 191.925 90.255 192.095 ;
        RECT 90.920 192.055 91.145 192.095 ;
        RECT 89.010 191.595 89.885 191.925 ;
        RECT 90.055 191.595 90.805 191.925 ;
        RECT 87.820 190.455 88.070 190.785 ;
        RECT 89.010 190.755 89.180 191.595 ;
        RECT 90.055 191.390 90.245 191.595 ;
        RECT 90.975 191.475 91.145 192.055 ;
        RECT 92.235 192.015 93.335 192.195 ;
        RECT 93.505 192.230 93.755 192.600 ;
        RECT 93.925 192.355 94.370 192.525 ;
        RECT 94.540 192.495 94.760 192.540 ;
        RECT 93.505 191.845 93.675 192.230 ;
        RECT 90.930 191.425 91.145 191.475 ;
        RECT 89.350 191.015 90.245 191.390 ;
        RECT 90.755 191.345 91.145 191.425 ;
        RECT 88.295 190.585 89.180 190.755 ;
        RECT 89.360 190.285 89.675 190.785 ;
        RECT 89.905 190.455 90.245 191.015 ;
        RECT 90.415 190.285 90.585 191.295 ;
        RECT 90.755 190.500 91.085 191.345 ;
        RECT 92.235 191.275 92.580 191.845 ;
        RECT 92.750 191.595 93.310 191.845 ;
        RECT 93.480 191.675 93.675 191.845 ;
        RECT 92.235 190.285 92.580 191.105 ;
        RECT 92.750 190.495 92.925 191.595 ;
        RECT 93.480 191.425 93.650 191.675 ;
        RECT 93.925 191.565 94.095 192.355 ;
        RECT 94.540 192.325 94.765 192.495 ;
        RECT 94.540 192.185 94.760 192.325 ;
        RECT 94.265 192.015 94.760 192.185 ;
        RECT 95.040 192.170 95.210 192.835 ;
        RECT 95.405 192.095 95.745 192.665 ;
        RECT 94.265 191.820 94.440 192.015 ;
        RECT 94.610 191.645 95.060 191.845 ;
        RECT 93.095 191.035 93.650 191.425 ;
        RECT 93.820 191.425 94.095 191.565 ;
        RECT 95.230 191.475 95.400 191.925 ;
        RECT 93.820 191.205 94.835 191.425 ;
        RECT 95.005 191.305 95.400 191.475 ;
        RECT 95.005 191.035 95.175 191.305 ;
        RECT 95.570 191.135 95.745 192.095 ;
        RECT 95.915 192.015 96.175 192.835 ;
        RECT 96.345 192.015 96.675 192.435 ;
        RECT 96.855 192.350 97.645 192.615 ;
        RECT 96.425 191.925 96.675 192.015 ;
        RECT 95.515 191.125 95.745 191.135 ;
        RECT 93.095 190.865 95.175 191.035 ;
        RECT 93.095 190.630 93.425 190.865 ;
        RECT 93.715 190.285 94.115 190.685 ;
        RECT 94.985 190.285 95.315 190.685 ;
        RECT 95.485 190.455 95.745 191.125 ;
        RECT 95.915 190.965 96.255 191.845 ;
        RECT 96.425 191.675 97.220 191.925 ;
        RECT 95.915 190.285 96.175 190.795 ;
        RECT 96.425 190.455 96.595 191.675 ;
        RECT 97.390 191.495 97.645 192.350 ;
        RECT 97.815 192.195 98.015 192.615 ;
        RECT 98.205 192.375 98.535 192.835 ;
        RECT 97.815 191.675 98.225 192.195 ;
        RECT 98.705 192.185 98.965 192.665 ;
        RECT 98.395 191.495 98.625 191.925 ;
        RECT 96.835 191.325 98.625 191.495 ;
        RECT 96.835 190.960 97.085 191.325 ;
        RECT 97.255 190.965 97.585 191.155 ;
        RECT 97.805 191.030 98.520 191.325 ;
        RECT 98.795 191.155 98.965 192.185 ;
        RECT 100.055 192.110 100.345 192.835 ;
        RECT 100.515 192.065 102.185 192.835 ;
        RECT 102.815 192.455 103.705 192.625 ;
        RECT 100.515 191.545 101.265 192.065 ;
        RECT 102.815 191.900 103.365 192.285 ;
        RECT 97.255 190.790 97.450 190.965 ;
        RECT 96.835 190.285 97.450 190.790 ;
        RECT 97.620 190.455 98.095 190.795 ;
        RECT 98.265 190.285 98.480 190.830 ;
        RECT 98.690 190.455 98.965 191.155 ;
        RECT 100.055 190.285 100.345 191.450 ;
        RECT 101.435 191.375 102.185 191.895 ;
        RECT 103.535 191.730 103.705 192.455 ;
        RECT 100.515 190.285 102.185 191.375 ;
        RECT 102.815 191.660 103.705 191.730 ;
        RECT 103.875 192.130 104.095 192.615 ;
        RECT 104.265 192.295 104.515 192.835 ;
        RECT 104.685 192.185 104.945 192.665 ;
        RECT 103.875 191.705 104.205 192.130 ;
        RECT 102.815 191.635 103.710 191.660 ;
        RECT 102.815 191.620 103.720 191.635 ;
        RECT 102.815 191.605 103.725 191.620 ;
        RECT 102.815 191.600 103.735 191.605 ;
        RECT 102.815 191.590 103.740 191.600 ;
        RECT 102.815 191.580 103.745 191.590 ;
        RECT 102.815 191.575 103.755 191.580 ;
        RECT 102.815 191.565 103.765 191.575 ;
        RECT 102.815 191.560 103.775 191.565 ;
        RECT 102.815 191.110 103.075 191.560 ;
        RECT 103.440 191.555 103.775 191.560 ;
        RECT 103.440 191.550 103.790 191.555 ;
        RECT 103.440 191.540 103.805 191.550 ;
        RECT 103.440 191.535 103.830 191.540 ;
        RECT 104.375 191.535 104.605 191.930 ;
        RECT 103.440 191.530 104.605 191.535 ;
        RECT 103.470 191.495 104.605 191.530 ;
        RECT 103.505 191.470 104.605 191.495 ;
        RECT 103.535 191.440 104.605 191.470 ;
        RECT 103.555 191.410 104.605 191.440 ;
        RECT 103.575 191.380 104.605 191.410 ;
        RECT 103.645 191.370 104.605 191.380 ;
        RECT 103.670 191.360 104.605 191.370 ;
        RECT 103.690 191.345 104.605 191.360 ;
        RECT 103.710 191.330 104.605 191.345 ;
        RECT 103.715 191.320 104.500 191.330 ;
        RECT 103.730 191.285 104.500 191.320 ;
        RECT 103.245 190.965 103.575 191.210 ;
        RECT 103.745 191.035 104.500 191.285 ;
        RECT 104.775 191.155 104.945 192.185 ;
        RECT 103.245 190.940 103.430 190.965 ;
        RECT 102.815 190.840 103.430 190.940 ;
        RECT 102.815 190.285 103.420 190.840 ;
        RECT 103.595 190.455 104.075 190.795 ;
        RECT 104.245 190.285 104.500 190.830 ;
        RECT 104.670 190.455 104.945 191.155 ;
        RECT 105.115 192.095 105.500 192.665 ;
        RECT 105.670 192.375 105.995 192.835 ;
        RECT 106.515 192.205 106.795 192.665 ;
        RECT 105.115 191.425 105.395 192.095 ;
        RECT 105.670 192.035 106.795 192.205 ;
        RECT 105.670 191.925 106.120 192.035 ;
        RECT 105.565 191.595 106.120 191.925 ;
        RECT 106.985 191.865 107.385 192.665 ;
        RECT 107.785 192.375 108.055 192.835 ;
        RECT 108.225 192.205 108.510 192.665 ;
        RECT 105.115 190.455 105.500 191.425 ;
        RECT 105.670 191.135 106.120 191.595 ;
        RECT 106.290 191.305 107.385 191.865 ;
        RECT 105.670 190.915 106.795 191.135 ;
        RECT 105.670 190.285 105.995 190.745 ;
        RECT 106.515 190.455 106.795 190.915 ;
        RECT 106.985 190.455 107.385 191.305 ;
        RECT 107.555 192.035 108.510 192.205 ;
        RECT 107.555 191.135 107.765 192.035 ;
        RECT 108.855 192.015 109.065 192.835 ;
        RECT 109.235 192.035 109.565 192.665 ;
        RECT 107.935 191.305 108.625 191.865 ;
        RECT 109.235 191.435 109.485 192.035 ;
        RECT 109.735 192.015 109.965 192.835 ;
        RECT 111.145 192.180 111.475 192.615 ;
        RECT 111.645 192.225 111.815 192.835 ;
        RECT 111.095 192.095 111.475 192.180 ;
        RECT 111.985 192.095 112.315 192.620 ;
        RECT 112.575 192.305 112.785 192.835 ;
        RECT 113.060 192.385 113.845 192.555 ;
        RECT 114.015 192.385 114.420 192.555 ;
        RECT 111.095 192.055 111.320 192.095 ;
        RECT 109.655 191.595 109.985 191.845 ;
        RECT 111.095 191.475 111.265 192.055 ;
        RECT 111.985 191.925 112.185 192.095 ;
        RECT 113.060 191.925 113.230 192.385 ;
        RECT 111.435 191.595 112.185 191.925 ;
        RECT 112.355 191.595 113.230 191.925 ;
        RECT 107.555 190.915 108.510 191.135 ;
        RECT 107.785 190.285 108.055 190.745 ;
        RECT 108.225 190.455 108.510 190.915 ;
        RECT 108.855 190.285 109.065 191.425 ;
        RECT 109.235 190.455 109.565 191.435 ;
        RECT 111.095 191.425 111.310 191.475 ;
        RECT 109.735 190.285 109.965 191.425 ;
        RECT 111.095 191.345 111.485 191.425 ;
        RECT 111.155 190.500 111.485 191.345 ;
        RECT 111.995 191.390 112.185 191.595 ;
        RECT 111.655 190.285 111.825 191.295 ;
        RECT 111.995 191.015 112.890 191.390 ;
        RECT 111.995 190.455 112.335 191.015 ;
        RECT 112.565 190.285 112.880 190.785 ;
        RECT 113.060 190.755 113.230 191.595 ;
        RECT 113.400 191.885 113.865 192.215 ;
        RECT 114.250 192.155 114.420 192.385 ;
        RECT 114.600 192.335 114.970 192.835 ;
        RECT 115.290 192.385 115.965 192.555 ;
        RECT 116.160 192.385 116.495 192.555 ;
        RECT 113.400 190.925 113.720 191.885 ;
        RECT 114.250 191.855 115.080 192.155 ;
        RECT 113.890 190.955 114.080 191.675 ;
        RECT 114.250 190.785 114.420 191.855 ;
        RECT 114.880 191.825 115.080 191.855 ;
        RECT 114.590 191.605 114.760 191.675 ;
        RECT 115.290 191.605 115.460 192.385 ;
        RECT 116.325 192.245 116.495 192.385 ;
        RECT 116.665 192.375 116.915 192.835 ;
        RECT 114.590 191.435 115.460 191.605 ;
        RECT 115.630 191.965 116.155 192.185 ;
        RECT 116.325 192.115 116.550 192.245 ;
        RECT 114.590 191.345 115.100 191.435 ;
        RECT 113.060 190.585 113.945 190.755 ;
        RECT 114.170 190.455 114.420 190.785 ;
        RECT 114.590 190.285 114.760 191.085 ;
        RECT 114.930 190.730 115.100 191.345 ;
        RECT 115.630 191.265 115.800 191.965 ;
        RECT 115.270 190.900 115.800 191.265 ;
        RECT 115.970 191.200 116.210 191.795 ;
        RECT 116.380 191.010 116.550 192.115 ;
        RECT 116.720 191.255 117.000 192.205 ;
        RECT 116.245 190.880 116.550 191.010 ;
        RECT 114.930 190.560 116.035 190.730 ;
        RECT 116.245 190.455 116.495 190.880 ;
        RECT 116.665 190.285 116.930 190.745 ;
        RECT 117.170 190.455 117.355 192.575 ;
        RECT 117.525 192.455 117.855 192.835 ;
        RECT 118.025 192.285 118.195 192.575 ;
        RECT 117.530 192.115 118.195 192.285 ;
        RECT 118.455 192.335 118.715 192.665 ;
        RECT 118.885 192.475 119.215 192.835 ;
        RECT 119.470 192.455 120.770 192.665 ;
        RECT 117.530 191.125 117.760 192.115 ;
        RECT 117.930 191.295 118.280 191.945 ;
        RECT 118.455 191.135 118.625 192.335 ;
        RECT 119.470 192.305 119.640 192.455 ;
        RECT 118.885 192.180 119.640 192.305 ;
        RECT 118.795 192.135 119.640 192.180 ;
        RECT 118.795 192.015 119.065 192.135 ;
        RECT 118.795 191.440 118.965 192.015 ;
        RECT 119.195 191.575 119.605 191.880 ;
        RECT 119.895 191.845 120.105 192.245 ;
        RECT 119.775 191.635 120.105 191.845 ;
        RECT 120.350 191.845 120.570 192.245 ;
        RECT 121.045 192.070 121.500 192.835 ;
        RECT 121.675 192.065 125.185 192.835 ;
        RECT 125.815 192.110 126.105 192.835 ;
        RECT 126.275 192.095 126.660 192.665 ;
        RECT 126.830 192.375 127.155 192.835 ;
        RECT 127.675 192.205 127.955 192.665 ;
        RECT 120.350 191.635 120.825 191.845 ;
        RECT 121.015 191.645 121.505 191.845 ;
        RECT 121.675 191.545 123.325 192.065 ;
        RECT 118.795 191.405 118.995 191.440 ;
        RECT 120.325 191.405 121.500 191.465 ;
        RECT 118.795 191.295 121.500 191.405 ;
        RECT 123.495 191.375 125.185 191.895 ;
        RECT 118.855 191.235 120.655 191.295 ;
        RECT 120.325 191.205 120.655 191.235 ;
        RECT 117.530 190.955 118.195 191.125 ;
        RECT 117.525 190.285 117.855 190.785 ;
        RECT 118.025 190.455 118.195 190.955 ;
        RECT 118.455 190.455 118.715 191.135 ;
        RECT 118.885 190.285 119.135 191.065 ;
        RECT 119.385 191.035 120.220 191.045 ;
        RECT 120.810 191.035 120.995 191.125 ;
        RECT 119.385 190.835 120.995 191.035 ;
        RECT 119.385 190.455 119.635 190.835 ;
        RECT 120.765 190.795 120.995 190.835 ;
        RECT 121.245 190.675 121.500 191.295 ;
        RECT 119.805 190.285 120.160 190.665 ;
        RECT 121.165 190.455 121.500 190.675 ;
        RECT 121.675 190.285 125.185 191.375 ;
        RECT 125.815 190.285 126.105 191.450 ;
        RECT 126.275 191.425 126.555 192.095 ;
        RECT 126.830 192.035 127.955 192.205 ;
        RECT 126.830 191.925 127.280 192.035 ;
        RECT 126.725 191.595 127.280 191.925 ;
        RECT 128.145 191.865 128.545 192.665 ;
        RECT 128.945 192.375 129.215 192.835 ;
        RECT 129.385 192.205 129.670 192.665 ;
        RECT 126.275 190.455 126.660 191.425 ;
        RECT 126.830 191.135 127.280 191.595 ;
        RECT 127.450 191.305 128.545 191.865 ;
        RECT 126.830 190.915 127.955 191.135 ;
        RECT 126.830 190.285 127.155 190.745 ;
        RECT 127.675 190.455 127.955 190.915 ;
        RECT 128.145 190.455 128.545 191.305 ;
        RECT 128.715 192.035 129.670 192.205 ;
        RECT 129.955 192.035 130.265 192.835 ;
        RECT 130.470 192.035 131.165 192.665 ;
        RECT 128.715 191.135 128.925 192.035 ;
        RECT 130.470 191.985 130.645 192.035 ;
        RECT 131.795 192.015 132.055 192.835 ;
        RECT 132.225 192.015 132.555 192.435 ;
        RECT 132.735 192.350 133.525 192.615 ;
        RECT 129.095 191.305 129.785 191.865 ;
        RECT 129.965 191.595 130.300 191.865 ;
        RECT 130.470 191.435 130.640 191.985 ;
        RECT 132.305 191.925 132.555 192.015 ;
        RECT 130.810 191.595 131.145 191.845 ;
        RECT 128.715 190.915 129.670 191.135 ;
        RECT 128.945 190.285 129.215 190.745 ;
        RECT 129.385 190.455 129.670 190.915 ;
        RECT 129.955 190.285 130.235 191.425 ;
        RECT 130.405 190.455 130.735 191.435 ;
        RECT 130.905 190.285 131.165 191.425 ;
        RECT 131.795 190.965 132.135 191.845 ;
        RECT 132.305 191.675 133.100 191.925 ;
        RECT 131.795 190.285 132.055 190.795 ;
        RECT 132.305 190.455 132.475 191.675 ;
        RECT 133.270 191.495 133.525 192.350 ;
        RECT 133.695 192.195 133.895 192.615 ;
        RECT 134.085 192.375 134.415 192.835 ;
        RECT 133.695 191.675 134.105 192.195 ;
        RECT 134.585 192.185 134.845 192.665 ;
        RECT 134.275 191.495 134.505 191.925 ;
        RECT 132.715 191.325 134.505 191.495 ;
        RECT 132.715 190.960 132.965 191.325 ;
        RECT 133.135 190.965 133.465 191.155 ;
        RECT 133.685 191.030 134.400 191.325 ;
        RECT 134.675 191.155 134.845 192.185 ;
        RECT 135.055 192.015 135.285 192.835 ;
        RECT 135.455 192.035 135.785 192.665 ;
        RECT 135.035 191.595 135.365 191.845 ;
        RECT 135.535 191.435 135.785 192.035 ;
        RECT 135.955 192.015 136.165 192.835 ;
        RECT 136.395 192.065 139.905 192.835 ;
        RECT 140.075 192.085 141.285 192.835 ;
        RECT 136.395 191.545 138.045 192.065 ;
        RECT 133.135 190.790 133.330 190.965 ;
        RECT 132.715 190.285 133.330 190.790 ;
        RECT 133.500 190.455 133.975 190.795 ;
        RECT 134.145 190.285 134.360 190.830 ;
        RECT 134.570 190.455 134.845 191.155 ;
        RECT 135.055 190.285 135.285 191.425 ;
        RECT 135.455 190.455 135.785 191.435 ;
        RECT 135.955 190.285 136.165 191.425 ;
        RECT 138.215 191.375 139.905 191.895 ;
        RECT 140.075 191.545 140.595 192.085 ;
        RECT 141.515 192.015 141.725 192.835 ;
        RECT 141.895 192.035 142.225 192.665 ;
        RECT 140.765 191.375 141.285 191.915 ;
        RECT 141.895 191.435 142.145 192.035 ;
        RECT 142.395 192.015 142.625 192.835 ;
        RECT 142.920 192.335 143.415 192.665 ;
        RECT 142.315 191.595 142.645 191.845 ;
        RECT 136.395 190.285 139.905 191.375 ;
        RECT 140.075 190.285 141.285 191.375 ;
        RECT 141.515 190.285 141.725 191.425 ;
        RECT 141.895 190.455 142.225 191.435 ;
        RECT 142.395 190.285 142.625 191.425 ;
        RECT 142.835 190.845 143.075 192.155 ;
        RECT 143.245 191.425 143.415 192.335 ;
        RECT 143.635 191.595 143.985 192.560 ;
        RECT 144.165 191.595 144.465 192.565 ;
        RECT 144.645 191.595 144.925 192.565 ;
        RECT 145.105 192.035 145.375 192.835 ;
        RECT 145.545 192.115 145.885 192.625 ;
        RECT 145.120 191.595 145.450 191.845 ;
        RECT 145.120 191.425 145.435 191.595 ;
        RECT 143.245 191.255 145.435 191.425 ;
        RECT 142.840 190.285 143.175 190.665 ;
        RECT 143.345 190.455 143.595 191.255 ;
        RECT 143.815 190.285 144.145 191.005 ;
        RECT 144.330 190.455 144.580 191.255 ;
        RECT 145.045 190.285 145.375 191.085 ;
        RECT 145.625 190.715 145.885 192.115 ;
        RECT 145.545 190.455 145.885 190.715 ;
        RECT 146.055 192.185 146.315 192.665 ;
        RECT 146.485 192.295 146.735 192.835 ;
        RECT 146.055 191.155 146.225 192.185 ;
        RECT 146.905 192.130 147.125 192.615 ;
        RECT 146.395 191.535 146.625 191.930 ;
        RECT 146.795 191.705 147.125 192.130 ;
        RECT 147.295 192.455 148.185 192.625 ;
        RECT 147.295 191.730 147.465 192.455 ;
        RECT 147.635 191.900 148.185 192.285 ;
        RECT 148.355 192.035 149.050 192.665 ;
        RECT 149.255 192.035 149.565 192.835 ;
        RECT 149.735 192.065 151.405 192.835 ;
        RECT 151.575 192.110 151.865 192.835 ;
        RECT 152.035 192.065 155.545 192.835 ;
        RECT 155.715 192.085 156.925 192.835 ;
        RECT 147.295 191.660 148.185 191.730 ;
        RECT 147.290 191.635 148.185 191.660 ;
        RECT 147.280 191.620 148.185 191.635 ;
        RECT 147.275 191.605 148.185 191.620 ;
        RECT 147.265 191.600 148.185 191.605 ;
        RECT 147.260 191.590 148.185 191.600 ;
        RECT 148.375 191.595 148.710 191.845 ;
        RECT 147.255 191.580 148.185 191.590 ;
        RECT 147.245 191.575 148.185 191.580 ;
        RECT 147.235 191.565 148.185 191.575 ;
        RECT 147.225 191.560 148.185 191.565 ;
        RECT 147.225 191.555 147.560 191.560 ;
        RECT 147.210 191.550 147.560 191.555 ;
        RECT 147.195 191.540 147.560 191.550 ;
        RECT 147.170 191.535 147.560 191.540 ;
        RECT 146.395 191.530 147.560 191.535 ;
        RECT 146.395 191.495 147.530 191.530 ;
        RECT 146.395 191.470 147.495 191.495 ;
        RECT 146.395 191.440 147.465 191.470 ;
        RECT 146.395 191.410 147.445 191.440 ;
        RECT 146.395 191.380 147.425 191.410 ;
        RECT 146.395 191.370 147.355 191.380 ;
        RECT 146.395 191.360 147.330 191.370 ;
        RECT 146.395 191.345 147.310 191.360 ;
        RECT 146.395 191.330 147.290 191.345 ;
        RECT 146.500 191.320 147.285 191.330 ;
        RECT 146.500 191.285 147.270 191.320 ;
        RECT 146.055 190.455 146.330 191.155 ;
        RECT 146.500 191.035 147.255 191.285 ;
        RECT 147.425 190.965 147.755 191.210 ;
        RECT 147.925 191.110 148.185 191.560 ;
        RECT 148.880 191.435 149.050 192.035 ;
        RECT 149.220 191.595 149.555 191.865 ;
        RECT 149.735 191.545 150.485 192.065 ;
        RECT 147.570 190.940 147.755 190.965 ;
        RECT 147.570 190.840 148.185 190.940 ;
        RECT 146.500 190.285 146.755 190.830 ;
        RECT 146.925 190.455 147.405 190.795 ;
        RECT 147.580 190.285 148.185 190.840 ;
        RECT 148.355 190.285 148.615 191.425 ;
        RECT 148.785 190.455 149.115 191.435 ;
        RECT 149.285 190.285 149.565 191.425 ;
        RECT 150.655 191.375 151.405 191.895 ;
        RECT 152.035 191.545 153.685 192.065 ;
        RECT 149.735 190.285 151.405 191.375 ;
        RECT 151.575 190.285 151.865 191.450 ;
        RECT 153.855 191.375 155.545 191.895 ;
        RECT 152.035 190.285 155.545 191.375 ;
        RECT 155.715 191.375 156.235 191.915 ;
        RECT 156.405 191.545 156.925 192.085 ;
        RECT 155.715 190.285 156.925 191.375 ;
        RECT 22.690 190.115 157.010 190.285 ;
        RECT 22.775 189.025 23.985 190.115 ;
        RECT 24.155 189.680 29.500 190.115 ;
        RECT 22.775 188.315 23.295 188.855 ;
        RECT 23.465 188.485 23.985 189.025 ;
        RECT 22.775 187.565 23.985 188.315 ;
        RECT 25.740 188.110 26.080 188.940 ;
        RECT 27.560 188.430 27.910 189.680 ;
        RECT 29.675 189.025 30.885 190.115 ;
        RECT 29.675 188.315 30.195 188.855 ;
        RECT 30.365 188.485 30.885 189.025 ;
        RECT 31.240 189.145 31.630 189.320 ;
        RECT 32.115 189.315 32.445 190.115 ;
        RECT 32.615 189.325 33.150 189.945 ;
        RECT 31.240 188.975 32.665 189.145 ;
        RECT 24.155 187.565 29.500 188.110 ;
        RECT 29.675 187.565 30.885 188.315 ;
        RECT 31.115 188.245 31.470 188.805 ;
        RECT 31.640 188.075 31.810 188.975 ;
        RECT 31.980 188.245 32.245 188.805 ;
        RECT 32.495 188.475 32.665 188.975 ;
        RECT 32.835 188.305 33.150 189.325 ;
        RECT 33.355 189.025 35.025 190.115 ;
        RECT 31.220 187.565 31.460 188.075 ;
        RECT 31.640 187.745 31.920 188.075 ;
        RECT 32.150 187.565 32.365 188.075 ;
        RECT 32.535 187.735 33.150 188.305 ;
        RECT 33.355 188.335 34.105 188.855 ;
        RECT 34.275 188.505 35.025 189.025 ;
        RECT 35.655 188.950 35.945 190.115 ;
        RECT 36.115 189.680 41.460 190.115 ;
        RECT 33.355 187.565 35.025 188.335 ;
        RECT 35.655 187.565 35.945 188.290 ;
        RECT 37.700 188.110 38.040 188.940 ;
        RECT 39.520 188.430 39.870 189.680 ;
        RECT 41.635 189.025 43.305 190.115 ;
        RECT 43.475 189.605 43.735 190.115 ;
        RECT 41.635 188.335 42.385 188.855 ;
        RECT 42.555 188.505 43.305 189.025 ;
        RECT 43.475 188.555 43.815 189.435 ;
        RECT 43.985 188.725 44.155 189.945 ;
        RECT 44.395 189.610 45.010 190.115 ;
        RECT 44.395 189.075 44.645 189.440 ;
        RECT 44.815 189.435 45.010 189.610 ;
        RECT 45.180 189.605 45.655 189.945 ;
        RECT 45.825 189.570 46.040 190.115 ;
        RECT 44.815 189.245 45.145 189.435 ;
        RECT 45.365 189.075 46.080 189.370 ;
        RECT 46.250 189.245 46.525 189.945 ;
        RECT 44.395 188.905 46.185 189.075 ;
        RECT 43.985 188.475 44.780 188.725 ;
        RECT 43.985 188.385 44.235 188.475 ;
        RECT 36.115 187.565 41.460 188.110 ;
        RECT 41.635 187.565 43.305 188.335 ;
        RECT 43.475 187.565 43.735 188.385 ;
        RECT 43.905 187.965 44.235 188.385 ;
        RECT 44.950 188.050 45.205 188.905 ;
        RECT 44.415 187.785 45.205 188.050 ;
        RECT 45.375 188.205 45.785 188.725 ;
        RECT 45.955 188.475 46.185 188.905 ;
        RECT 46.355 188.215 46.525 189.245 ;
        RECT 45.375 187.785 45.575 188.205 ;
        RECT 45.765 187.565 46.095 188.025 ;
        RECT 46.265 187.735 46.525 188.215 ;
        RECT 46.695 189.245 46.970 189.945 ;
        RECT 47.140 189.570 47.395 190.115 ;
        RECT 47.565 189.605 48.045 189.945 ;
        RECT 48.220 189.560 48.825 190.115 ;
        RECT 48.210 189.460 48.825 189.560 ;
        RECT 48.210 189.435 48.395 189.460 ;
        RECT 46.695 188.215 46.865 189.245 ;
        RECT 47.140 189.115 47.895 189.365 ;
        RECT 48.065 189.190 48.395 189.435 ;
        RECT 47.140 189.080 47.910 189.115 ;
        RECT 47.140 189.070 47.925 189.080 ;
        RECT 47.035 189.055 47.930 189.070 ;
        RECT 47.035 189.040 47.950 189.055 ;
        RECT 47.035 189.030 47.970 189.040 ;
        RECT 47.035 189.020 47.995 189.030 ;
        RECT 47.035 188.990 48.065 189.020 ;
        RECT 47.035 188.960 48.085 188.990 ;
        RECT 47.035 188.930 48.105 188.960 ;
        RECT 47.035 188.905 48.135 188.930 ;
        RECT 47.035 188.870 48.170 188.905 ;
        RECT 47.035 188.865 48.200 188.870 ;
        RECT 47.035 188.470 47.265 188.865 ;
        RECT 47.810 188.860 48.200 188.865 ;
        RECT 47.835 188.850 48.200 188.860 ;
        RECT 47.850 188.845 48.200 188.850 ;
        RECT 47.865 188.840 48.200 188.845 ;
        RECT 48.565 188.840 48.825 189.290 ;
        RECT 49.180 189.145 49.570 189.320 ;
        RECT 50.055 189.315 50.385 190.115 ;
        RECT 50.555 189.325 51.090 189.945 ;
        RECT 49.180 188.975 50.605 189.145 ;
        RECT 47.865 188.835 48.825 188.840 ;
        RECT 47.875 188.825 48.825 188.835 ;
        RECT 47.885 188.820 48.825 188.825 ;
        RECT 47.895 188.810 48.825 188.820 ;
        RECT 47.900 188.800 48.825 188.810 ;
        RECT 47.905 188.795 48.825 188.800 ;
        RECT 47.915 188.780 48.825 188.795 ;
        RECT 47.920 188.765 48.825 188.780 ;
        RECT 47.930 188.740 48.825 188.765 ;
        RECT 47.435 188.270 47.765 188.695 ;
        RECT 47.515 188.245 47.765 188.270 ;
        RECT 46.695 187.735 46.955 188.215 ;
        RECT 47.125 187.565 47.375 188.105 ;
        RECT 47.545 187.785 47.765 188.245 ;
        RECT 47.935 188.670 48.825 188.740 ;
        RECT 47.935 187.945 48.105 188.670 ;
        RECT 48.275 188.115 48.825 188.500 ;
        RECT 49.055 188.245 49.410 188.805 ;
        RECT 49.580 188.075 49.750 188.975 ;
        RECT 49.920 188.245 50.185 188.805 ;
        RECT 50.435 188.475 50.605 188.975 ;
        RECT 50.775 188.305 51.090 189.325 ;
        RECT 51.295 189.025 52.965 190.115 ;
        RECT 47.935 187.775 48.825 187.945 ;
        RECT 49.160 187.565 49.400 188.075 ;
        RECT 49.580 187.745 49.860 188.075 ;
        RECT 50.090 187.565 50.305 188.075 ;
        RECT 50.475 187.735 51.090 188.305 ;
        RECT 51.295 188.335 52.045 188.855 ;
        RECT 52.215 188.505 52.965 189.025 ;
        RECT 53.595 188.975 53.980 189.935 ;
        RECT 54.195 189.315 54.485 190.115 ;
        RECT 54.655 189.775 56.020 189.945 ;
        RECT 54.655 189.145 54.825 189.775 ;
        RECT 54.150 188.975 54.825 189.145 ;
        RECT 51.295 187.565 52.965 188.335 ;
        RECT 53.595 188.305 53.770 188.975 ;
        RECT 54.150 188.805 54.320 188.975 ;
        RECT 54.995 188.805 55.320 189.605 ;
        RECT 55.690 189.565 56.020 189.775 ;
        RECT 55.690 189.315 56.645 189.565 ;
        RECT 53.955 188.555 54.320 188.805 ;
        RECT 54.515 188.555 54.765 188.805 ;
        RECT 53.955 188.475 54.145 188.555 ;
        RECT 54.515 188.475 54.685 188.555 ;
        RECT 54.975 188.475 55.320 188.805 ;
        RECT 55.490 188.475 55.765 189.140 ;
        RECT 55.950 188.475 56.305 189.140 ;
        RECT 56.475 188.305 56.645 189.315 ;
        RECT 56.815 188.975 57.105 190.115 ;
        RECT 57.275 188.975 57.550 189.945 ;
        RECT 57.760 189.315 58.040 190.115 ;
        RECT 58.210 189.605 59.825 189.935 ;
        RECT 58.210 189.265 59.385 189.435 ;
        RECT 58.210 189.145 58.380 189.265 ;
        RECT 57.720 188.975 58.380 189.145 ;
        RECT 56.830 188.475 57.105 188.805 ;
        RECT 53.595 187.735 54.105 188.305 ;
        RECT 54.650 188.135 56.050 188.305 ;
        RECT 54.275 187.565 54.445 188.125 ;
        RECT 54.650 187.735 54.980 188.135 ;
        RECT 55.155 187.565 55.485 187.965 ;
        RECT 55.720 187.945 56.050 188.135 ;
        RECT 56.220 188.115 56.645 188.305 ;
        RECT 57.275 188.240 57.445 188.975 ;
        RECT 57.720 188.805 57.890 188.975 ;
        RECT 58.640 188.805 58.885 189.095 ;
        RECT 59.055 188.975 59.385 189.265 ;
        RECT 59.645 188.805 59.815 189.365 ;
        RECT 60.065 188.975 60.325 190.115 ;
        RECT 61.415 188.950 61.705 190.115 ;
        RECT 61.875 189.395 62.335 189.945 ;
        RECT 62.525 189.395 62.855 190.115 ;
        RECT 57.615 188.475 57.890 188.805 ;
        RECT 58.060 188.475 58.885 188.805 ;
        RECT 59.100 188.475 59.815 188.805 ;
        RECT 59.985 188.555 60.320 188.805 ;
        RECT 57.720 188.305 57.890 188.475 ;
        RECT 59.565 188.385 59.815 188.475 ;
        RECT 56.815 187.945 57.105 188.215 ;
        RECT 55.720 187.735 57.105 187.945 ;
        RECT 57.275 187.895 57.550 188.240 ;
        RECT 57.720 188.135 59.385 188.305 ;
        RECT 57.740 187.565 58.115 187.965 ;
        RECT 58.285 187.785 58.455 188.135 ;
        RECT 58.625 187.565 58.955 187.965 ;
        RECT 59.125 187.735 59.385 188.135 ;
        RECT 59.565 187.965 59.895 188.385 ;
        RECT 60.065 187.565 60.325 188.385 ;
        RECT 61.415 187.565 61.705 188.290 ;
        RECT 61.875 188.025 62.125 189.395 ;
        RECT 63.055 189.225 63.355 189.775 ;
        RECT 63.525 189.445 63.805 190.115 ;
        RECT 62.415 189.055 63.355 189.225 ;
        RECT 62.415 188.805 62.585 189.055 ;
        RECT 63.725 188.805 63.990 189.165 ;
        RECT 64.695 189.055 65.025 189.900 ;
        RECT 65.195 189.105 65.365 190.115 ;
        RECT 65.535 189.385 65.875 189.945 ;
        RECT 66.105 189.615 66.420 190.115 ;
        RECT 66.600 189.645 67.485 189.815 ;
        RECT 62.295 188.475 62.585 188.805 ;
        RECT 62.755 188.555 63.095 188.805 ;
        RECT 63.315 188.555 63.990 188.805 ;
        RECT 64.635 188.975 65.025 189.055 ;
        RECT 65.535 189.010 66.430 189.385 ;
        RECT 64.635 188.925 64.850 188.975 ;
        RECT 62.415 188.385 62.585 188.475 ;
        RECT 62.415 188.195 63.805 188.385 ;
        RECT 64.635 188.345 64.805 188.925 ;
        RECT 65.535 188.805 65.725 189.010 ;
        RECT 66.600 188.805 66.770 189.645 ;
        RECT 67.710 189.615 67.960 189.945 ;
        RECT 64.975 188.475 65.725 188.805 ;
        RECT 65.895 188.475 66.770 188.805 ;
        RECT 64.635 188.305 64.860 188.345 ;
        RECT 65.525 188.305 65.725 188.475 ;
        RECT 64.635 188.220 65.015 188.305 ;
        RECT 61.875 187.735 62.435 188.025 ;
        RECT 62.605 187.565 62.855 188.025 ;
        RECT 63.475 187.835 63.805 188.195 ;
        RECT 64.685 187.785 65.015 188.220 ;
        RECT 65.185 187.565 65.355 188.175 ;
        RECT 65.525 187.780 65.855 188.305 ;
        RECT 66.115 187.565 66.325 188.095 ;
        RECT 66.600 188.015 66.770 188.475 ;
        RECT 66.940 188.515 67.260 189.475 ;
        RECT 67.430 188.725 67.620 189.445 ;
        RECT 67.790 188.545 67.960 189.615 ;
        RECT 68.130 189.315 68.300 190.115 ;
        RECT 68.470 189.670 69.575 189.840 ;
        RECT 68.470 189.055 68.640 189.670 ;
        RECT 69.785 189.520 70.035 189.945 ;
        RECT 70.205 189.655 70.470 190.115 ;
        RECT 68.810 189.135 69.340 189.500 ;
        RECT 69.785 189.390 70.090 189.520 ;
        RECT 68.130 188.965 68.640 189.055 ;
        RECT 68.130 188.795 69.000 188.965 ;
        RECT 68.130 188.725 68.300 188.795 ;
        RECT 68.420 188.545 68.620 188.575 ;
        RECT 66.940 188.185 67.405 188.515 ;
        RECT 67.790 188.245 68.620 188.545 ;
        RECT 67.790 188.015 67.960 188.245 ;
        RECT 66.600 187.845 67.385 188.015 ;
        RECT 67.555 187.845 67.960 188.015 ;
        RECT 68.140 187.565 68.510 188.065 ;
        RECT 68.830 188.015 69.000 188.795 ;
        RECT 69.170 188.435 69.340 189.135 ;
        RECT 69.510 188.605 69.750 189.200 ;
        RECT 69.170 188.215 69.695 188.435 ;
        RECT 69.920 188.285 70.090 189.390 ;
        RECT 69.865 188.155 70.090 188.285 ;
        RECT 70.260 188.195 70.540 189.145 ;
        RECT 69.865 188.015 70.035 188.155 ;
        RECT 68.830 187.845 69.505 188.015 ;
        RECT 69.700 187.845 70.035 188.015 ;
        RECT 70.205 187.565 70.455 188.025 ;
        RECT 70.710 187.825 70.895 189.945 ;
        RECT 71.065 189.615 71.395 190.115 ;
        RECT 71.565 189.445 71.735 189.945 ;
        RECT 71.070 189.275 71.735 189.445 ;
        RECT 71.070 188.285 71.300 189.275 ;
        RECT 71.470 188.455 71.820 189.105 ;
        RECT 71.995 189.025 74.585 190.115 ;
        RECT 71.995 188.335 73.205 188.855 ;
        RECT 73.375 188.505 74.585 189.025 ;
        RECT 74.755 189.265 75.015 189.945 ;
        RECT 75.185 189.335 75.435 190.115 ;
        RECT 75.685 189.565 75.935 189.945 ;
        RECT 76.105 189.735 76.460 190.115 ;
        RECT 77.465 189.725 77.800 189.945 ;
        RECT 77.065 189.565 77.295 189.605 ;
        RECT 75.685 189.365 77.295 189.565 ;
        RECT 75.685 189.355 76.520 189.365 ;
        RECT 77.110 189.275 77.295 189.365 ;
        RECT 71.070 188.115 71.735 188.285 ;
        RECT 71.065 187.565 71.395 187.945 ;
        RECT 71.565 187.825 71.735 188.115 ;
        RECT 71.995 187.565 74.585 188.335 ;
        RECT 74.755 188.065 74.925 189.265 ;
        RECT 76.625 189.165 76.955 189.195 ;
        RECT 75.155 189.105 76.955 189.165 ;
        RECT 77.545 189.105 77.800 189.725 ;
        RECT 77.985 189.305 78.280 190.115 ;
        RECT 75.095 188.995 77.800 189.105 ;
        RECT 75.095 188.960 75.295 188.995 ;
        RECT 75.095 188.385 75.265 188.960 ;
        RECT 76.625 188.935 77.800 188.995 ;
        RECT 75.495 188.520 75.905 188.825 ;
        RECT 78.460 188.805 78.705 189.945 ;
        RECT 78.880 189.305 79.140 190.115 ;
        RECT 79.740 190.110 86.015 190.115 ;
        RECT 79.320 188.805 79.570 189.940 ;
        RECT 79.740 189.315 80.000 190.110 ;
        RECT 80.170 189.215 80.430 189.940 ;
        RECT 80.600 189.385 80.860 190.110 ;
        RECT 81.030 189.215 81.290 189.940 ;
        RECT 81.460 189.385 81.720 190.110 ;
        RECT 81.890 189.215 82.150 189.940 ;
        RECT 82.320 189.385 82.580 190.110 ;
        RECT 82.750 189.215 83.010 189.940 ;
        RECT 83.180 189.385 83.425 190.110 ;
        RECT 83.595 189.215 83.855 189.940 ;
        RECT 84.040 189.385 84.285 190.110 ;
        RECT 84.455 189.215 84.715 189.940 ;
        RECT 84.900 189.385 85.145 190.110 ;
        RECT 85.315 189.215 85.575 189.940 ;
        RECT 85.760 189.385 86.015 190.110 ;
        RECT 80.170 189.200 85.575 189.215 ;
        RECT 86.185 189.200 86.475 189.940 ;
        RECT 86.645 189.370 86.915 190.115 ;
        RECT 80.170 188.975 86.915 189.200 ;
        RECT 76.075 188.555 76.405 188.765 ;
        RECT 75.095 188.265 75.365 188.385 ;
        RECT 75.095 188.220 75.940 188.265 ;
        RECT 75.185 188.095 75.940 188.220 ;
        RECT 76.195 188.155 76.405 188.555 ;
        RECT 76.650 188.555 77.125 188.765 ;
        RECT 77.315 188.555 77.805 188.755 ;
        RECT 76.650 188.155 76.870 188.555 ;
        RECT 74.755 187.735 75.015 188.065 ;
        RECT 75.770 187.945 75.940 188.095 ;
        RECT 75.185 187.565 75.515 187.925 ;
        RECT 75.770 187.735 77.070 187.945 ;
        RECT 77.345 187.565 77.800 188.330 ;
        RECT 77.975 188.245 78.290 188.805 ;
        RECT 78.460 188.555 85.580 188.805 ;
        RECT 77.975 187.565 78.280 188.075 ;
        RECT 78.460 187.745 78.710 188.555 ;
        RECT 78.880 187.565 79.140 188.090 ;
        RECT 79.320 187.745 79.570 188.555 ;
        RECT 85.750 188.385 86.915 188.975 ;
        RECT 87.175 188.950 87.465 190.115 ;
        RECT 87.635 188.975 88.020 189.945 ;
        RECT 88.190 189.655 88.515 190.115 ;
        RECT 89.035 189.485 89.315 189.945 ;
        RECT 88.190 189.265 89.315 189.485 ;
        RECT 80.170 188.215 86.915 188.385 ;
        RECT 87.635 188.305 87.915 188.975 ;
        RECT 88.190 188.805 88.640 189.265 ;
        RECT 89.505 189.095 89.905 189.945 ;
        RECT 90.305 189.655 90.575 190.115 ;
        RECT 90.745 189.485 91.030 189.945 ;
        RECT 88.085 188.475 88.640 188.805 ;
        RECT 88.810 188.535 89.905 189.095 ;
        RECT 88.190 188.365 88.640 188.475 ;
        RECT 79.740 187.565 80.000 188.125 ;
        RECT 80.170 187.760 80.430 188.215 ;
        RECT 80.600 187.565 80.860 188.045 ;
        RECT 81.030 187.760 81.290 188.215 ;
        RECT 81.460 187.565 81.720 188.045 ;
        RECT 81.890 187.760 82.150 188.215 ;
        RECT 82.320 187.565 82.565 188.045 ;
        RECT 82.735 187.760 83.010 188.215 ;
        RECT 83.180 187.565 83.425 188.045 ;
        RECT 83.595 187.760 83.855 188.215 ;
        RECT 84.035 187.565 84.285 188.045 ;
        RECT 84.455 187.760 84.715 188.215 ;
        RECT 84.895 187.565 85.145 188.045 ;
        RECT 85.315 187.760 85.575 188.215 ;
        RECT 85.755 187.565 86.015 188.045 ;
        RECT 86.185 187.760 86.445 188.215 ;
        RECT 86.615 187.565 86.915 188.045 ;
        RECT 87.175 187.565 87.465 188.290 ;
        RECT 87.635 187.735 88.020 188.305 ;
        RECT 88.190 188.195 89.315 188.365 ;
        RECT 88.190 187.565 88.515 188.025 ;
        RECT 89.035 187.735 89.315 188.195 ;
        RECT 89.505 187.735 89.905 188.535 ;
        RECT 90.075 189.265 91.030 189.485 ;
        RECT 90.075 188.365 90.285 189.265 ;
        RECT 90.455 188.535 91.145 189.095 ;
        RECT 91.315 189.025 94.825 190.115 ;
        RECT 95.460 189.735 95.795 190.115 ;
        RECT 90.075 188.195 91.030 188.365 ;
        RECT 90.305 187.565 90.575 188.025 ;
        RECT 90.745 187.735 91.030 188.195 ;
        RECT 91.315 188.335 92.965 188.855 ;
        RECT 93.135 188.505 94.825 189.025 ;
        RECT 91.315 187.565 94.825 188.335 ;
        RECT 95.455 188.245 95.695 189.555 ;
        RECT 95.965 189.145 96.215 189.945 ;
        RECT 96.435 189.395 96.765 190.115 ;
        RECT 96.950 189.145 97.200 189.945 ;
        RECT 97.665 189.315 97.995 190.115 ;
        RECT 98.165 189.685 98.505 189.945 ;
        RECT 95.865 188.975 98.055 189.145 ;
        RECT 95.865 188.065 96.035 188.975 ;
        RECT 97.740 188.805 98.055 188.975 ;
        RECT 95.540 187.735 96.035 188.065 ;
        RECT 96.255 187.840 96.605 188.805 ;
        RECT 96.785 187.835 97.085 188.805 ;
        RECT 97.265 187.835 97.545 188.805 ;
        RECT 97.740 188.555 98.070 188.805 ;
        RECT 97.725 187.565 97.995 188.365 ;
        RECT 98.245 188.285 98.505 189.685 ;
        RECT 98.165 187.775 98.505 188.285 ;
        RECT 98.695 189.060 99.000 189.845 ;
        RECT 99.180 189.645 99.865 190.115 ;
        RECT 99.175 189.125 99.870 189.435 ;
        RECT 98.695 188.255 98.870 189.060 ;
        RECT 100.045 188.955 100.330 189.900 ;
        RECT 100.505 189.665 100.835 190.115 ;
        RECT 101.005 189.495 101.175 189.925 ;
        RECT 99.470 188.805 100.330 188.955 ;
        RECT 99.045 188.785 100.330 188.805 ;
        RECT 100.500 189.265 101.175 189.495 ;
        RECT 99.045 188.425 100.030 188.785 ;
        RECT 100.500 188.615 100.735 189.265 ;
        RECT 98.695 187.735 98.935 188.255 ;
        RECT 99.860 188.090 100.030 188.425 ;
        RECT 100.200 188.285 100.735 188.615 ;
        RECT 100.515 188.135 100.735 188.285 ;
        RECT 100.905 188.245 101.205 189.095 ;
        RECT 101.435 189.025 104.945 190.115 ;
        RECT 101.435 188.335 103.085 188.855 ;
        RECT 103.255 188.505 104.945 189.025 ;
        RECT 105.115 188.975 105.395 190.115 ;
        RECT 105.565 188.965 105.895 189.945 ;
        RECT 106.065 188.975 106.325 190.115 ;
        RECT 106.680 189.145 107.070 189.320 ;
        RECT 107.555 189.315 107.885 190.115 ;
        RECT 108.055 189.325 108.590 189.945 ;
        RECT 108.795 189.560 109.400 190.115 ;
        RECT 109.575 189.605 110.055 189.945 ;
        RECT 110.225 189.570 110.480 190.115 ;
        RECT 108.795 189.460 109.410 189.560 ;
        RECT 106.680 188.975 108.105 189.145 ;
        RECT 105.125 188.535 105.460 188.805 ;
        RECT 105.630 188.365 105.800 188.965 ;
        RECT 105.970 188.555 106.305 188.805 ;
        RECT 99.105 187.565 99.500 188.060 ;
        RECT 99.860 187.895 100.235 188.090 ;
        RECT 100.065 187.750 100.235 187.895 ;
        RECT 100.515 187.760 100.755 188.135 ;
        RECT 100.925 187.565 101.260 188.070 ;
        RECT 101.435 187.565 104.945 188.335 ;
        RECT 105.115 187.565 105.425 188.365 ;
        RECT 105.630 187.735 106.325 188.365 ;
        RECT 106.555 188.245 106.910 188.805 ;
        RECT 107.080 188.075 107.250 188.975 ;
        RECT 107.420 188.245 107.685 188.805 ;
        RECT 107.935 188.475 108.105 188.975 ;
        RECT 108.275 188.305 108.590 189.325 ;
        RECT 109.225 189.435 109.410 189.460 ;
        RECT 108.795 188.840 109.055 189.290 ;
        RECT 109.225 189.190 109.555 189.435 ;
        RECT 109.725 189.115 110.480 189.365 ;
        RECT 110.650 189.245 110.925 189.945 ;
        RECT 109.710 189.080 110.480 189.115 ;
        RECT 109.695 189.070 110.480 189.080 ;
        RECT 109.690 189.055 110.585 189.070 ;
        RECT 109.670 189.040 110.585 189.055 ;
        RECT 109.650 189.030 110.585 189.040 ;
        RECT 109.625 189.020 110.585 189.030 ;
        RECT 109.555 188.990 110.585 189.020 ;
        RECT 109.535 188.960 110.585 188.990 ;
        RECT 109.515 188.930 110.585 188.960 ;
        RECT 109.485 188.905 110.585 188.930 ;
        RECT 109.450 188.870 110.585 188.905 ;
        RECT 109.420 188.865 110.585 188.870 ;
        RECT 109.420 188.860 109.810 188.865 ;
        RECT 109.420 188.850 109.785 188.860 ;
        RECT 109.420 188.845 109.770 188.850 ;
        RECT 109.420 188.840 109.755 188.845 ;
        RECT 108.795 188.835 109.755 188.840 ;
        RECT 108.795 188.825 109.745 188.835 ;
        RECT 108.795 188.820 109.735 188.825 ;
        RECT 108.795 188.810 109.725 188.820 ;
        RECT 108.795 188.800 109.720 188.810 ;
        RECT 108.795 188.795 109.715 188.800 ;
        RECT 108.795 188.780 109.705 188.795 ;
        RECT 108.795 188.765 109.700 188.780 ;
        RECT 108.795 188.740 109.690 188.765 ;
        RECT 108.795 188.670 109.685 188.740 ;
        RECT 106.660 187.565 106.900 188.075 ;
        RECT 107.080 187.745 107.360 188.075 ;
        RECT 107.590 187.565 107.805 188.075 ;
        RECT 107.975 187.735 108.590 188.305 ;
        RECT 108.795 188.115 109.345 188.500 ;
        RECT 109.515 187.945 109.685 188.670 ;
        RECT 108.795 187.775 109.685 187.945 ;
        RECT 109.855 188.270 110.185 188.695 ;
        RECT 110.355 188.470 110.585 188.865 ;
        RECT 109.855 187.785 110.075 188.270 ;
        RECT 110.755 188.215 110.925 189.245 ;
        RECT 111.135 188.975 111.365 190.115 ;
        RECT 111.535 188.965 111.865 189.945 ;
        RECT 112.035 188.975 112.245 190.115 ;
        RECT 111.115 188.555 111.445 188.805 ;
        RECT 110.245 187.565 110.495 188.105 ;
        RECT 110.665 187.735 110.925 188.215 ;
        RECT 111.135 187.565 111.365 188.385 ;
        RECT 111.615 188.365 111.865 188.965 ;
        RECT 112.935 188.950 113.225 190.115 ;
        RECT 113.395 188.975 113.655 190.115 ;
        RECT 113.825 188.965 114.155 189.945 ;
        RECT 114.325 188.975 114.605 190.115 ;
        RECT 114.865 189.185 115.035 189.945 ;
        RECT 115.215 189.355 115.545 190.115 ;
        RECT 114.865 189.015 115.530 189.185 ;
        RECT 115.715 189.040 115.985 189.945 ;
        RECT 113.415 188.555 113.750 188.805 ;
        RECT 111.535 187.735 111.865 188.365 ;
        RECT 112.035 187.565 112.245 188.385 ;
        RECT 113.920 188.365 114.090 188.965 ;
        RECT 115.360 188.870 115.530 189.015 ;
        RECT 114.260 188.535 114.595 188.805 ;
        RECT 114.795 188.465 115.125 188.835 ;
        RECT 115.360 188.540 115.645 188.870 ;
        RECT 112.935 187.565 113.225 188.290 ;
        RECT 113.395 187.735 114.090 188.365 ;
        RECT 114.295 187.565 114.605 188.365 ;
        RECT 115.360 188.285 115.530 188.540 ;
        RECT 114.865 188.115 115.530 188.285 ;
        RECT 115.815 188.240 115.985 189.040 ;
        RECT 116.155 189.025 117.365 190.115 ;
        RECT 117.625 189.445 117.795 189.945 ;
        RECT 117.965 189.615 118.295 190.115 ;
        RECT 117.625 189.275 118.290 189.445 ;
        RECT 114.865 187.735 115.035 188.115 ;
        RECT 115.215 187.565 115.545 187.945 ;
        RECT 115.725 187.735 115.985 188.240 ;
        RECT 116.155 188.315 116.675 188.855 ;
        RECT 116.845 188.485 117.365 189.025 ;
        RECT 117.540 188.455 117.890 189.105 ;
        RECT 116.155 187.565 117.365 188.315 ;
        RECT 118.060 188.285 118.290 189.275 ;
        RECT 117.625 188.115 118.290 188.285 ;
        RECT 117.625 187.825 117.795 188.115 ;
        RECT 117.965 187.565 118.295 187.945 ;
        RECT 118.465 187.825 118.650 189.945 ;
        RECT 118.890 189.655 119.155 190.115 ;
        RECT 119.325 189.520 119.575 189.945 ;
        RECT 119.785 189.670 120.890 189.840 ;
        RECT 119.270 189.390 119.575 189.520 ;
        RECT 118.820 188.195 119.100 189.145 ;
        RECT 119.270 188.285 119.440 189.390 ;
        RECT 119.610 188.605 119.850 189.200 ;
        RECT 120.020 189.135 120.550 189.500 ;
        RECT 120.020 188.435 120.190 189.135 ;
        RECT 120.720 189.055 120.890 189.670 ;
        RECT 121.060 189.315 121.230 190.115 ;
        RECT 121.400 189.615 121.650 189.945 ;
        RECT 121.875 189.645 122.760 189.815 ;
        RECT 120.720 188.965 121.230 189.055 ;
        RECT 119.270 188.155 119.495 188.285 ;
        RECT 119.665 188.215 120.190 188.435 ;
        RECT 120.360 188.795 121.230 188.965 ;
        RECT 118.905 187.565 119.155 188.025 ;
        RECT 119.325 188.015 119.495 188.155 ;
        RECT 120.360 188.015 120.530 188.795 ;
        RECT 121.060 188.725 121.230 188.795 ;
        RECT 120.740 188.545 120.940 188.575 ;
        RECT 121.400 188.545 121.570 189.615 ;
        RECT 121.740 188.725 121.930 189.445 ;
        RECT 120.740 188.245 121.570 188.545 ;
        RECT 122.100 188.515 122.420 189.475 ;
        RECT 119.325 187.845 119.660 188.015 ;
        RECT 119.855 187.845 120.530 188.015 ;
        RECT 120.850 187.565 121.220 188.065 ;
        RECT 121.400 188.015 121.570 188.245 ;
        RECT 121.955 188.185 122.420 188.515 ;
        RECT 122.590 188.805 122.760 189.645 ;
        RECT 122.940 189.615 123.255 190.115 ;
        RECT 123.485 189.385 123.825 189.945 ;
        RECT 122.930 189.010 123.825 189.385 ;
        RECT 123.995 189.105 124.165 190.115 ;
        RECT 123.635 188.805 123.825 189.010 ;
        RECT 124.335 189.055 124.665 189.900 ;
        RECT 124.335 188.975 124.725 189.055 ;
        RECT 125.825 188.975 126.155 190.115 ;
        RECT 126.685 189.145 127.015 189.930 ;
        RECT 127.195 189.560 127.800 190.115 ;
        RECT 127.975 189.605 128.455 189.945 ;
        RECT 128.625 189.570 128.880 190.115 ;
        RECT 127.195 189.460 127.810 189.560 ;
        RECT 127.625 189.435 127.810 189.460 ;
        RECT 126.335 188.975 127.015 189.145 ;
        RECT 124.510 188.925 124.725 188.975 ;
        RECT 122.590 188.475 123.465 188.805 ;
        RECT 123.635 188.475 124.385 188.805 ;
        RECT 122.590 188.015 122.760 188.475 ;
        RECT 123.635 188.305 123.835 188.475 ;
        RECT 124.555 188.345 124.725 188.925 ;
        RECT 125.815 188.555 126.165 188.805 ;
        RECT 126.335 188.375 126.505 188.975 ;
        RECT 127.195 188.840 127.455 189.290 ;
        RECT 127.625 189.190 127.955 189.435 ;
        RECT 128.125 189.115 128.880 189.365 ;
        RECT 129.050 189.245 129.325 189.945 ;
        RECT 128.110 189.080 128.880 189.115 ;
        RECT 128.095 189.070 128.880 189.080 ;
        RECT 128.090 189.055 128.985 189.070 ;
        RECT 128.070 189.040 128.985 189.055 ;
        RECT 128.050 189.030 128.985 189.040 ;
        RECT 128.025 189.020 128.985 189.030 ;
        RECT 127.955 188.990 128.985 189.020 ;
        RECT 127.935 188.960 128.985 188.990 ;
        RECT 127.915 188.930 128.985 188.960 ;
        RECT 127.885 188.905 128.985 188.930 ;
        RECT 127.850 188.870 128.985 188.905 ;
        RECT 127.820 188.865 128.985 188.870 ;
        RECT 127.820 188.860 128.210 188.865 ;
        RECT 127.820 188.850 128.185 188.860 ;
        RECT 127.820 188.845 128.170 188.850 ;
        RECT 127.820 188.840 128.155 188.845 ;
        RECT 127.195 188.835 128.155 188.840 ;
        RECT 127.195 188.825 128.145 188.835 ;
        RECT 127.195 188.820 128.135 188.825 ;
        RECT 127.195 188.810 128.125 188.820 ;
        RECT 126.675 188.555 127.025 188.805 ;
        RECT 127.195 188.800 128.120 188.810 ;
        RECT 127.195 188.795 128.115 188.800 ;
        RECT 127.195 188.780 128.105 188.795 ;
        RECT 127.195 188.765 128.100 188.780 ;
        RECT 127.195 188.740 128.090 188.765 ;
        RECT 127.195 188.670 128.085 188.740 ;
        RECT 124.500 188.305 124.725 188.345 ;
        RECT 121.400 187.845 121.805 188.015 ;
        RECT 121.975 187.845 122.760 188.015 ;
        RECT 123.035 187.565 123.245 188.095 ;
        RECT 123.505 187.780 123.835 188.305 ;
        RECT 124.345 188.220 124.725 188.305 ;
        RECT 124.005 187.565 124.175 188.175 ;
        RECT 124.345 187.785 124.675 188.220 ;
        RECT 125.825 187.565 126.095 188.375 ;
        RECT 126.265 187.735 126.595 188.375 ;
        RECT 126.765 187.565 127.005 188.375 ;
        RECT 127.195 188.115 127.745 188.500 ;
        RECT 127.915 187.945 128.085 188.670 ;
        RECT 127.195 187.775 128.085 187.945 ;
        RECT 128.255 188.270 128.585 188.695 ;
        RECT 128.755 188.470 128.985 188.865 ;
        RECT 128.255 188.245 128.505 188.270 ;
        RECT 128.255 187.785 128.475 188.245 ;
        RECT 129.155 188.215 129.325 189.245 ;
        RECT 128.645 187.565 128.895 188.105 ;
        RECT 129.065 187.735 129.325 188.215 ;
        RECT 129.495 189.245 129.770 189.945 ;
        RECT 129.940 189.570 130.195 190.115 ;
        RECT 130.365 189.605 130.845 189.945 ;
        RECT 131.020 189.560 131.625 190.115 ;
        RECT 131.010 189.460 131.625 189.560 ;
        RECT 131.010 189.435 131.195 189.460 ;
        RECT 129.495 188.215 129.665 189.245 ;
        RECT 129.940 189.115 130.695 189.365 ;
        RECT 130.865 189.190 131.195 189.435 ;
        RECT 129.940 189.080 130.710 189.115 ;
        RECT 129.940 189.070 130.725 189.080 ;
        RECT 129.835 189.055 130.730 189.070 ;
        RECT 129.835 189.040 130.750 189.055 ;
        RECT 129.835 189.030 130.770 189.040 ;
        RECT 129.835 189.020 130.795 189.030 ;
        RECT 129.835 188.990 130.865 189.020 ;
        RECT 129.835 188.960 130.885 188.990 ;
        RECT 129.835 188.930 130.905 188.960 ;
        RECT 129.835 188.905 130.935 188.930 ;
        RECT 129.835 188.870 130.970 188.905 ;
        RECT 129.835 188.865 131.000 188.870 ;
        RECT 129.835 188.470 130.065 188.865 ;
        RECT 130.610 188.860 131.000 188.865 ;
        RECT 130.635 188.850 131.000 188.860 ;
        RECT 130.650 188.845 131.000 188.850 ;
        RECT 130.665 188.840 131.000 188.845 ;
        RECT 131.365 188.840 131.625 189.290 ;
        RECT 131.980 189.145 132.370 189.320 ;
        RECT 132.855 189.315 133.185 190.115 ;
        RECT 133.355 189.325 133.890 189.945 ;
        RECT 131.980 188.975 133.405 189.145 ;
        RECT 130.665 188.835 131.625 188.840 ;
        RECT 130.675 188.825 131.625 188.835 ;
        RECT 130.685 188.820 131.625 188.825 ;
        RECT 130.695 188.810 131.625 188.820 ;
        RECT 130.700 188.800 131.625 188.810 ;
        RECT 130.705 188.795 131.625 188.800 ;
        RECT 130.715 188.780 131.625 188.795 ;
        RECT 130.720 188.765 131.625 188.780 ;
        RECT 130.730 188.740 131.625 188.765 ;
        RECT 130.235 188.270 130.565 188.695 ;
        RECT 129.495 187.735 129.755 188.215 ;
        RECT 129.925 187.565 130.175 188.105 ;
        RECT 130.345 187.785 130.565 188.270 ;
        RECT 130.735 188.670 131.625 188.740 ;
        RECT 130.735 187.945 130.905 188.670 ;
        RECT 131.075 188.115 131.625 188.500 ;
        RECT 131.855 188.245 132.210 188.805 ;
        RECT 132.380 188.075 132.550 188.975 ;
        RECT 132.720 188.245 132.985 188.805 ;
        RECT 133.235 188.475 133.405 188.975 ;
        RECT 133.575 188.305 133.890 189.325 ;
        RECT 134.095 189.025 135.765 190.115 ;
        RECT 130.735 187.775 131.625 187.945 ;
        RECT 131.960 187.565 132.200 188.075 ;
        RECT 132.380 187.745 132.660 188.075 ;
        RECT 132.890 187.565 133.105 188.075 ;
        RECT 133.275 187.735 133.890 188.305 ;
        RECT 134.095 188.335 134.845 188.855 ;
        RECT 135.015 188.505 135.765 189.025 ;
        RECT 135.940 188.975 136.195 190.115 ;
        RECT 136.390 189.565 137.585 189.895 ;
        RECT 136.445 188.805 136.615 189.365 ;
        RECT 136.840 189.145 137.260 189.395 ;
        RECT 137.765 189.315 138.045 190.115 ;
        RECT 136.840 188.975 138.085 189.145 ;
        RECT 138.255 188.975 138.525 189.945 ;
        RECT 137.915 188.805 138.085 188.975 ;
        RECT 135.940 188.555 136.275 188.805 ;
        RECT 136.445 188.475 137.185 188.805 ;
        RECT 137.915 188.475 138.145 188.805 ;
        RECT 136.445 188.385 136.695 188.475 ;
        RECT 134.095 187.565 135.765 188.335 ;
        RECT 135.960 188.215 136.695 188.385 ;
        RECT 137.915 188.305 138.085 188.475 ;
        RECT 135.960 187.745 136.270 188.215 ;
        RECT 137.345 188.135 138.085 188.305 ;
        RECT 138.355 188.240 138.525 188.975 ;
        RECT 138.695 188.950 138.985 190.115 ;
        RECT 139.155 189.680 144.500 190.115 ;
        RECT 136.440 187.565 137.175 188.045 ;
        RECT 137.345 187.785 137.515 188.135 ;
        RECT 137.685 187.565 138.065 187.965 ;
        RECT 138.255 187.895 138.525 188.240 ;
        RECT 138.695 187.565 138.985 188.290 ;
        RECT 140.740 188.110 141.080 188.940 ;
        RECT 142.560 188.430 142.910 189.680 ;
        RECT 144.675 189.025 146.345 190.115 ;
        RECT 146.525 189.305 146.820 190.115 ;
        RECT 144.675 188.335 145.425 188.855 ;
        RECT 145.595 188.505 146.345 189.025 ;
        RECT 147.000 188.805 147.245 189.945 ;
        RECT 147.420 189.305 147.680 190.115 ;
        RECT 148.280 190.110 154.555 190.115 ;
        RECT 147.860 188.805 148.110 189.940 ;
        RECT 148.280 189.315 148.540 190.110 ;
        RECT 148.710 189.215 148.970 189.940 ;
        RECT 149.140 189.385 149.400 190.110 ;
        RECT 149.570 189.215 149.830 189.940 ;
        RECT 150.000 189.385 150.260 190.110 ;
        RECT 150.430 189.215 150.690 189.940 ;
        RECT 150.860 189.385 151.120 190.110 ;
        RECT 151.290 189.215 151.550 189.940 ;
        RECT 151.720 189.385 151.965 190.110 ;
        RECT 152.135 189.215 152.395 189.940 ;
        RECT 152.580 189.385 152.825 190.110 ;
        RECT 152.995 189.215 153.255 189.940 ;
        RECT 153.440 189.385 153.685 190.110 ;
        RECT 153.855 189.215 154.115 189.940 ;
        RECT 154.300 189.385 154.555 190.110 ;
        RECT 148.710 189.200 154.115 189.215 ;
        RECT 154.725 189.200 155.015 189.940 ;
        RECT 155.185 189.370 155.455 190.115 ;
        RECT 148.710 188.975 155.455 189.200 ;
        RECT 139.155 187.565 144.500 188.110 ;
        RECT 144.675 187.565 146.345 188.335 ;
        RECT 146.515 188.245 146.830 188.805 ;
        RECT 147.000 188.555 154.120 188.805 ;
        RECT 146.515 187.565 146.820 188.075 ;
        RECT 147.000 187.745 147.250 188.555 ;
        RECT 147.420 187.565 147.680 188.090 ;
        RECT 147.860 187.745 148.110 188.555 ;
        RECT 154.290 188.385 155.455 188.975 ;
        RECT 155.715 189.025 156.925 190.115 ;
        RECT 155.715 188.485 156.235 189.025 ;
        RECT 148.710 188.215 155.455 188.385 ;
        RECT 156.405 188.315 156.925 188.855 ;
        RECT 148.280 187.565 148.540 188.125 ;
        RECT 148.710 187.760 148.970 188.215 ;
        RECT 149.140 187.565 149.400 188.045 ;
        RECT 149.570 187.760 149.830 188.215 ;
        RECT 150.000 187.565 150.260 188.045 ;
        RECT 150.430 187.760 150.690 188.215 ;
        RECT 150.860 187.565 151.105 188.045 ;
        RECT 151.275 187.760 151.550 188.215 ;
        RECT 151.720 187.565 151.965 188.045 ;
        RECT 152.135 187.760 152.395 188.215 ;
        RECT 152.575 187.565 152.825 188.045 ;
        RECT 152.995 187.760 153.255 188.215 ;
        RECT 153.435 187.565 153.685 188.045 ;
        RECT 153.855 187.760 154.115 188.215 ;
        RECT 154.295 187.565 154.555 188.045 ;
        RECT 154.725 187.760 154.985 188.215 ;
        RECT 155.155 187.565 155.455 188.045 ;
        RECT 155.715 187.565 156.925 188.315 ;
        RECT 22.690 187.395 157.010 187.565 ;
        RECT 22.775 186.645 23.985 187.395 ;
        RECT 24.705 186.845 24.875 187.135 ;
        RECT 25.045 187.015 25.375 187.395 ;
        RECT 24.705 186.675 25.370 186.845 ;
        RECT 22.775 186.105 23.295 186.645 ;
        RECT 23.465 185.935 23.985 186.475 ;
        RECT 22.775 184.845 23.985 185.935 ;
        RECT 24.620 185.855 24.970 186.505 ;
        RECT 25.140 185.685 25.370 186.675 ;
        RECT 24.705 185.515 25.370 185.685 ;
        RECT 24.705 185.015 24.875 185.515 ;
        RECT 25.045 184.845 25.375 185.345 ;
        RECT 25.545 185.015 25.730 187.135 ;
        RECT 25.985 186.935 26.235 187.395 ;
        RECT 26.405 186.945 26.740 187.115 ;
        RECT 26.935 186.945 27.610 187.115 ;
        RECT 26.405 186.805 26.575 186.945 ;
        RECT 25.900 185.815 26.180 186.765 ;
        RECT 26.350 186.675 26.575 186.805 ;
        RECT 26.350 185.570 26.520 186.675 ;
        RECT 26.745 186.525 27.270 186.745 ;
        RECT 26.690 185.760 26.930 186.355 ;
        RECT 27.100 185.825 27.270 186.525 ;
        RECT 27.440 186.165 27.610 186.945 ;
        RECT 27.930 186.895 28.300 187.395 ;
        RECT 28.480 186.945 28.885 187.115 ;
        RECT 29.055 186.945 29.840 187.115 ;
        RECT 28.480 186.715 28.650 186.945 ;
        RECT 27.820 186.415 28.650 186.715 ;
        RECT 29.035 186.445 29.500 186.775 ;
        RECT 27.820 186.385 28.020 186.415 ;
        RECT 28.140 186.165 28.310 186.235 ;
        RECT 27.440 185.995 28.310 186.165 ;
        RECT 27.800 185.905 28.310 185.995 ;
        RECT 26.350 185.440 26.655 185.570 ;
        RECT 27.100 185.460 27.630 185.825 ;
        RECT 25.970 184.845 26.235 185.305 ;
        RECT 26.405 185.015 26.655 185.440 ;
        RECT 27.800 185.290 27.970 185.905 ;
        RECT 26.865 185.120 27.970 185.290 ;
        RECT 28.140 184.845 28.310 185.645 ;
        RECT 28.480 185.345 28.650 186.415 ;
        RECT 28.820 185.515 29.010 186.235 ;
        RECT 29.180 185.485 29.500 186.445 ;
        RECT 29.670 186.485 29.840 186.945 ;
        RECT 30.115 186.865 30.325 187.395 ;
        RECT 30.585 186.655 30.915 187.180 ;
        RECT 31.085 186.785 31.255 187.395 ;
        RECT 31.425 186.740 31.755 187.175 ;
        RECT 31.975 186.745 32.235 187.225 ;
        RECT 32.405 186.935 32.735 187.395 ;
        RECT 32.925 186.755 33.125 187.175 ;
        RECT 31.425 186.655 31.805 186.740 ;
        RECT 30.715 186.485 30.915 186.655 ;
        RECT 31.580 186.615 31.805 186.655 ;
        RECT 29.670 186.155 30.545 186.485 ;
        RECT 30.715 186.155 31.465 186.485 ;
        RECT 28.480 185.015 28.730 185.345 ;
        RECT 29.670 185.315 29.840 186.155 ;
        RECT 30.715 185.950 30.905 186.155 ;
        RECT 31.635 186.035 31.805 186.615 ;
        RECT 31.590 185.985 31.805 186.035 ;
        RECT 30.010 185.575 30.905 185.950 ;
        RECT 31.415 185.905 31.805 185.985 ;
        RECT 28.955 185.145 29.840 185.315 ;
        RECT 30.020 184.845 30.335 185.345 ;
        RECT 30.565 185.015 30.905 185.575 ;
        RECT 31.075 184.845 31.245 185.855 ;
        RECT 31.415 185.060 31.745 185.905 ;
        RECT 31.975 185.715 32.145 186.745 ;
        RECT 32.315 186.055 32.545 186.485 ;
        RECT 32.715 186.235 33.125 186.755 ;
        RECT 33.295 186.910 34.085 187.175 ;
        RECT 33.295 186.055 33.550 186.910 ;
        RECT 34.265 186.575 34.595 186.995 ;
        RECT 34.765 186.575 35.025 187.395 ;
        RECT 35.360 186.885 35.600 187.395 ;
        RECT 35.780 186.885 36.060 187.215 ;
        RECT 36.290 186.885 36.505 187.395 ;
        RECT 34.265 186.485 34.515 186.575 ;
        RECT 33.720 186.235 34.515 186.485 ;
        RECT 32.315 185.885 34.105 186.055 ;
        RECT 31.975 185.015 32.250 185.715 ;
        RECT 32.420 185.590 33.135 185.885 ;
        RECT 33.355 185.525 33.685 185.715 ;
        RECT 32.460 184.845 32.675 185.390 ;
        RECT 32.845 185.015 33.320 185.355 ;
        RECT 33.490 185.350 33.685 185.525 ;
        RECT 33.855 185.520 34.105 185.885 ;
        RECT 33.490 184.845 34.105 185.350 ;
        RECT 34.345 185.015 34.515 186.235 ;
        RECT 34.685 185.525 35.025 186.405 ;
        RECT 35.255 186.155 35.610 186.715 ;
        RECT 35.780 185.985 35.950 186.885 ;
        RECT 36.120 186.155 36.385 186.715 ;
        RECT 36.675 186.655 37.290 187.225 ;
        RECT 36.635 185.985 36.805 186.485 ;
        RECT 35.380 185.815 36.805 185.985 ;
        RECT 35.380 185.640 35.770 185.815 ;
        RECT 34.765 184.845 35.025 185.355 ;
        RECT 36.255 184.845 36.585 185.645 ;
        RECT 36.975 185.635 37.290 186.655 ;
        RECT 36.755 185.015 37.290 185.635 ;
        RECT 37.955 186.720 38.215 187.225 ;
        RECT 38.395 187.015 38.725 187.395 ;
        RECT 38.905 186.845 39.075 187.225 ;
        RECT 37.955 185.920 38.125 186.720 ;
        RECT 38.410 186.675 39.075 186.845 ;
        RECT 38.410 186.420 38.580 186.675 ;
        RECT 39.335 186.625 42.845 187.395 ;
        RECT 43.015 186.645 44.225 187.395 ;
        RECT 44.595 186.765 44.925 187.125 ;
        RECT 45.545 186.935 45.795 187.395 ;
        RECT 45.965 186.935 46.525 187.225 ;
        RECT 38.295 186.090 38.580 186.420 ;
        RECT 38.815 186.125 39.145 186.495 ;
        RECT 39.335 186.105 40.985 186.625 ;
        RECT 38.410 185.945 38.580 186.090 ;
        RECT 37.955 185.015 38.225 185.920 ;
        RECT 38.410 185.775 39.075 185.945 ;
        RECT 41.155 185.935 42.845 186.455 ;
        RECT 43.015 186.105 43.535 186.645 ;
        RECT 44.595 186.575 45.985 186.765 ;
        RECT 45.815 186.485 45.985 186.575 ;
        RECT 43.705 185.935 44.225 186.475 ;
        RECT 38.395 184.845 38.725 185.605 ;
        RECT 38.905 185.015 39.075 185.775 ;
        RECT 39.335 184.845 42.845 185.935 ;
        RECT 43.015 184.845 44.225 185.935 ;
        RECT 44.410 186.155 45.085 186.405 ;
        RECT 45.305 186.155 45.645 186.405 ;
        RECT 45.815 186.155 46.105 186.485 ;
        RECT 44.410 185.795 44.675 186.155 ;
        RECT 45.815 185.905 45.985 186.155 ;
        RECT 45.045 185.735 45.985 185.905 ;
        RECT 44.595 184.845 44.875 185.515 ;
        RECT 45.045 185.185 45.345 185.735 ;
        RECT 46.275 185.565 46.525 186.935 ;
        RECT 46.755 186.575 46.965 187.395 ;
        RECT 47.135 186.595 47.465 187.225 ;
        RECT 47.135 185.995 47.385 186.595 ;
        RECT 47.635 186.575 47.865 187.395 ;
        RECT 48.535 186.670 48.825 187.395 ;
        RECT 48.995 186.645 50.205 187.395 ;
        RECT 50.575 186.765 50.905 187.125 ;
        RECT 51.525 186.935 51.775 187.395 ;
        RECT 51.945 186.935 52.505 187.225 ;
        RECT 47.555 186.155 47.885 186.405 ;
        RECT 48.995 186.105 49.515 186.645 ;
        RECT 50.575 186.575 51.965 186.765 ;
        RECT 51.795 186.485 51.965 186.575 ;
        RECT 45.545 184.845 45.875 185.565 ;
        RECT 46.065 185.015 46.525 185.565 ;
        RECT 46.755 184.845 46.965 185.985 ;
        RECT 47.135 185.015 47.465 185.995 ;
        RECT 47.635 184.845 47.865 185.985 ;
        RECT 48.535 184.845 48.825 186.010 ;
        RECT 49.685 185.935 50.205 186.475 ;
        RECT 48.995 184.845 50.205 185.935 ;
        RECT 50.390 186.155 51.065 186.405 ;
        RECT 51.285 186.155 51.625 186.405 ;
        RECT 51.795 186.155 52.085 186.485 ;
        RECT 50.390 185.795 50.655 186.155 ;
        RECT 51.795 185.905 51.965 186.155 ;
        RECT 51.025 185.735 51.965 185.905 ;
        RECT 50.575 184.845 50.855 185.515 ;
        RECT 51.025 185.185 51.325 185.735 ;
        RECT 52.255 185.565 52.505 186.935 ;
        RECT 52.695 185.815 52.925 187.155 ;
        RECT 53.105 186.315 53.335 187.215 ;
        RECT 53.535 186.615 53.780 187.395 ;
        RECT 53.950 186.855 54.380 187.215 ;
        RECT 54.960 187.025 55.690 187.395 ;
        RECT 53.950 186.665 55.690 186.855 ;
        RECT 53.950 186.435 54.170 186.665 ;
        RECT 53.105 185.635 53.445 186.315 ;
        RECT 51.525 184.845 51.855 185.565 ;
        RECT 52.045 185.015 52.505 185.565 ;
        RECT 52.695 185.435 53.445 185.635 ;
        RECT 53.625 186.135 54.170 186.435 ;
        RECT 52.695 185.045 52.935 185.435 ;
        RECT 53.105 184.845 53.455 185.255 ;
        RECT 53.625 185.025 53.955 186.135 ;
        RECT 54.340 185.865 54.765 186.485 ;
        RECT 54.960 185.865 55.220 186.485 ;
        RECT 55.430 186.155 55.690 186.665 ;
        RECT 54.125 185.495 55.150 185.695 ;
        RECT 54.125 185.025 54.305 185.495 ;
        RECT 54.475 184.845 54.805 185.325 ;
        RECT 54.980 185.025 55.150 185.495 ;
        RECT 55.415 184.845 55.700 185.985 ;
        RECT 55.890 185.025 56.170 187.215 ;
        RECT 56.365 186.895 56.695 187.395 ;
        RECT 56.895 186.825 57.065 187.175 ;
        RECT 57.265 186.995 57.595 187.395 ;
        RECT 57.765 186.825 57.935 187.175 ;
        RECT 58.105 186.995 58.485 187.395 ;
        RECT 56.360 186.155 56.710 186.725 ;
        RECT 56.895 186.655 58.505 186.825 ;
        RECT 58.675 186.720 58.945 187.065 ;
        RECT 58.335 186.485 58.505 186.655 ;
        RECT 56.360 185.695 56.680 185.985 ;
        RECT 56.880 185.865 57.590 186.485 ;
        RECT 57.760 186.155 58.165 186.485 ;
        RECT 58.335 186.155 58.605 186.485 ;
        RECT 58.335 185.985 58.505 186.155 ;
        RECT 58.775 185.985 58.945 186.720 ;
        RECT 57.780 185.815 58.505 185.985 ;
        RECT 57.780 185.695 57.950 185.815 ;
        RECT 56.360 185.525 57.950 185.695 ;
        RECT 56.360 185.065 58.015 185.355 ;
        RECT 58.185 184.845 58.465 185.645 ;
        RECT 58.675 185.015 58.945 185.985 ;
        RECT 60.035 186.895 60.295 187.225 ;
        RECT 60.465 187.035 60.795 187.395 ;
        RECT 61.050 187.015 62.350 187.225 ;
        RECT 60.035 185.695 60.205 186.895 ;
        RECT 61.050 186.865 61.220 187.015 ;
        RECT 60.465 186.740 61.220 186.865 ;
        RECT 60.375 186.695 61.220 186.740 ;
        RECT 60.375 186.575 60.645 186.695 ;
        RECT 60.375 186.000 60.545 186.575 ;
        RECT 60.775 186.135 61.185 186.440 ;
        RECT 61.475 186.405 61.685 186.805 ;
        RECT 61.355 186.195 61.685 186.405 ;
        RECT 61.930 186.405 62.150 186.805 ;
        RECT 62.625 186.630 63.080 187.395 ;
        RECT 63.255 186.895 63.515 187.225 ;
        RECT 63.685 187.035 64.015 187.395 ;
        RECT 64.270 187.015 65.570 187.225 ;
        RECT 61.930 186.195 62.405 186.405 ;
        RECT 62.595 186.205 63.085 186.405 ;
        RECT 60.375 185.965 60.575 186.000 ;
        RECT 61.905 185.965 63.080 186.025 ;
        RECT 60.375 185.855 63.080 185.965 ;
        RECT 60.435 185.795 62.235 185.855 ;
        RECT 61.905 185.765 62.235 185.795 ;
        RECT 60.035 185.015 60.295 185.695 ;
        RECT 60.465 184.845 60.715 185.625 ;
        RECT 60.965 185.595 61.800 185.605 ;
        RECT 62.390 185.595 62.575 185.685 ;
        RECT 60.965 185.395 62.575 185.595 ;
        RECT 60.965 185.015 61.215 185.395 ;
        RECT 62.345 185.355 62.575 185.395 ;
        RECT 62.825 185.235 63.080 185.855 ;
        RECT 61.385 184.845 61.740 185.225 ;
        RECT 62.745 185.015 63.080 185.235 ;
        RECT 63.255 185.695 63.425 186.895 ;
        RECT 64.270 186.865 64.440 187.015 ;
        RECT 63.685 186.740 64.440 186.865 ;
        RECT 63.595 186.695 64.440 186.740 ;
        RECT 63.595 186.575 63.865 186.695 ;
        RECT 63.595 186.000 63.765 186.575 ;
        RECT 63.995 186.135 64.405 186.440 ;
        RECT 64.695 186.405 64.905 186.805 ;
        RECT 64.575 186.195 64.905 186.405 ;
        RECT 65.150 186.405 65.370 186.805 ;
        RECT 65.845 186.630 66.300 187.395 ;
        RECT 66.475 186.655 66.860 187.225 ;
        RECT 67.030 186.935 67.355 187.395 ;
        RECT 67.875 186.765 68.155 187.225 ;
        RECT 65.150 186.195 65.625 186.405 ;
        RECT 65.815 186.205 66.305 186.405 ;
        RECT 63.595 185.965 63.795 186.000 ;
        RECT 65.125 185.965 66.300 186.025 ;
        RECT 63.595 185.855 66.300 185.965 ;
        RECT 63.655 185.795 65.455 185.855 ;
        RECT 65.125 185.765 65.455 185.795 ;
        RECT 63.255 185.015 63.515 185.695 ;
        RECT 63.685 184.845 63.935 185.625 ;
        RECT 64.185 185.595 65.020 185.605 ;
        RECT 65.610 185.595 65.795 185.685 ;
        RECT 64.185 185.395 65.795 185.595 ;
        RECT 64.185 185.015 64.435 185.395 ;
        RECT 65.565 185.355 65.795 185.395 ;
        RECT 66.045 185.235 66.300 185.855 ;
        RECT 64.605 184.845 64.960 185.225 ;
        RECT 65.965 185.015 66.300 185.235 ;
        RECT 66.475 185.985 66.755 186.655 ;
        RECT 67.030 186.595 68.155 186.765 ;
        RECT 67.030 186.485 67.480 186.595 ;
        RECT 66.925 186.155 67.480 186.485 ;
        RECT 68.345 186.425 68.745 187.225 ;
        RECT 69.145 186.935 69.415 187.395 ;
        RECT 69.585 186.765 69.870 187.225 ;
        RECT 66.475 185.015 66.860 185.985 ;
        RECT 67.030 185.695 67.480 186.155 ;
        RECT 67.650 185.865 68.745 186.425 ;
        RECT 67.030 185.475 68.155 185.695 ;
        RECT 67.030 184.845 67.355 185.305 ;
        RECT 67.875 185.015 68.155 185.475 ;
        RECT 68.345 185.015 68.745 185.865 ;
        RECT 68.915 186.595 69.870 186.765 ;
        RECT 70.155 186.655 70.540 187.225 ;
        RECT 70.710 186.935 71.035 187.395 ;
        RECT 71.555 186.765 71.835 187.225 ;
        RECT 68.915 185.695 69.125 186.595 ;
        RECT 69.295 185.865 69.985 186.425 ;
        RECT 70.155 185.985 70.435 186.655 ;
        RECT 70.710 186.595 71.835 186.765 ;
        RECT 70.710 186.485 71.160 186.595 ;
        RECT 70.605 186.155 71.160 186.485 ;
        RECT 72.025 186.425 72.425 187.225 ;
        RECT 72.825 186.935 73.095 187.395 ;
        RECT 73.265 186.765 73.550 187.225 ;
        RECT 68.915 185.475 69.870 185.695 ;
        RECT 69.145 184.845 69.415 185.305 ;
        RECT 69.585 185.015 69.870 185.475 ;
        RECT 70.155 185.015 70.540 185.985 ;
        RECT 70.710 185.695 71.160 186.155 ;
        RECT 71.330 185.865 72.425 186.425 ;
        RECT 70.710 185.475 71.835 185.695 ;
        RECT 70.710 184.845 71.035 185.305 ;
        RECT 71.555 185.015 71.835 185.475 ;
        RECT 72.025 185.015 72.425 185.865 ;
        RECT 72.595 186.595 73.550 186.765 ;
        RECT 74.295 186.670 74.585 187.395 ;
        RECT 74.755 186.645 75.965 187.395 ;
        RECT 76.135 186.895 76.395 187.225 ;
        RECT 76.565 187.035 76.895 187.395 ;
        RECT 77.150 187.015 78.450 187.225 ;
        RECT 72.595 185.695 72.805 186.595 ;
        RECT 72.975 185.865 73.665 186.425 ;
        RECT 74.755 186.105 75.275 186.645 ;
        RECT 72.595 185.475 73.550 185.695 ;
        RECT 72.825 184.845 73.095 185.305 ;
        RECT 73.265 185.015 73.550 185.475 ;
        RECT 74.295 184.845 74.585 186.010 ;
        RECT 75.445 185.935 75.965 186.475 ;
        RECT 74.755 184.845 75.965 185.935 ;
        RECT 76.135 185.695 76.305 186.895 ;
        RECT 77.150 186.865 77.320 187.015 ;
        RECT 76.565 186.740 77.320 186.865 ;
        RECT 76.475 186.695 77.320 186.740 ;
        RECT 76.475 186.575 76.745 186.695 ;
        RECT 76.475 186.000 76.645 186.575 ;
        RECT 76.875 186.135 77.285 186.440 ;
        RECT 77.575 186.405 77.785 186.805 ;
        RECT 77.455 186.195 77.785 186.405 ;
        RECT 78.030 186.405 78.250 186.805 ;
        RECT 78.725 186.630 79.180 187.395 ;
        RECT 79.355 186.655 79.740 187.225 ;
        RECT 79.910 186.935 80.235 187.395 ;
        RECT 80.755 186.765 81.035 187.225 ;
        RECT 78.030 186.195 78.505 186.405 ;
        RECT 78.695 186.205 79.185 186.405 ;
        RECT 76.475 185.965 76.675 186.000 ;
        RECT 78.005 185.965 79.180 186.025 ;
        RECT 76.475 185.855 79.180 185.965 ;
        RECT 76.535 185.795 78.335 185.855 ;
        RECT 78.005 185.765 78.335 185.795 ;
        RECT 76.135 185.015 76.395 185.695 ;
        RECT 76.565 184.845 76.815 185.625 ;
        RECT 77.065 185.595 77.900 185.605 ;
        RECT 78.490 185.595 78.675 185.685 ;
        RECT 77.065 185.395 78.675 185.595 ;
        RECT 77.065 185.015 77.315 185.395 ;
        RECT 78.445 185.355 78.675 185.395 ;
        RECT 78.925 185.235 79.180 185.855 ;
        RECT 77.485 184.845 77.840 185.225 ;
        RECT 78.845 185.015 79.180 185.235 ;
        RECT 79.355 185.985 79.635 186.655 ;
        RECT 79.910 186.595 81.035 186.765 ;
        RECT 79.910 186.485 80.360 186.595 ;
        RECT 79.805 186.155 80.360 186.485 ;
        RECT 81.225 186.425 81.625 187.225 ;
        RECT 82.025 186.935 82.295 187.395 ;
        RECT 82.465 186.765 82.750 187.225 ;
        RECT 79.355 185.015 79.740 185.985 ;
        RECT 79.910 185.695 80.360 186.155 ;
        RECT 80.530 185.865 81.625 186.425 ;
        RECT 79.910 185.475 81.035 185.695 ;
        RECT 79.910 184.845 80.235 185.305 ;
        RECT 80.755 185.015 81.035 185.475 ;
        RECT 81.225 185.015 81.625 185.865 ;
        RECT 81.795 186.595 82.750 186.765 ;
        RECT 83.035 186.895 83.295 187.225 ;
        RECT 83.465 187.035 83.795 187.395 ;
        RECT 84.050 187.015 85.350 187.225 ;
        RECT 83.035 186.885 83.265 186.895 ;
        RECT 81.795 185.695 82.005 186.595 ;
        RECT 82.175 185.865 82.865 186.425 ;
        RECT 83.035 185.695 83.205 186.885 ;
        RECT 84.050 186.865 84.220 187.015 ;
        RECT 83.465 186.740 84.220 186.865 ;
        RECT 83.375 186.695 84.220 186.740 ;
        RECT 83.375 186.575 83.645 186.695 ;
        RECT 83.375 186.000 83.545 186.575 ;
        RECT 83.775 186.135 84.185 186.440 ;
        RECT 84.475 186.405 84.685 186.805 ;
        RECT 84.355 186.195 84.685 186.405 ;
        RECT 84.930 186.405 85.150 186.805 ;
        RECT 85.625 186.630 86.080 187.395 ;
        RECT 86.740 186.745 87.050 187.215 ;
        RECT 87.220 186.915 87.955 187.395 ;
        RECT 88.125 186.825 88.295 187.175 ;
        RECT 88.465 186.995 88.845 187.395 ;
        RECT 86.740 186.575 87.475 186.745 ;
        RECT 88.125 186.655 88.865 186.825 ;
        RECT 89.035 186.720 89.305 187.065 ;
        RECT 87.225 186.485 87.475 186.575 ;
        RECT 88.695 186.485 88.865 186.655 ;
        RECT 84.930 186.195 85.405 186.405 ;
        RECT 85.595 186.205 86.085 186.405 ;
        RECT 86.720 186.155 87.055 186.405 ;
        RECT 87.225 186.155 87.965 186.485 ;
        RECT 88.695 186.155 88.925 186.485 ;
        RECT 83.375 185.965 83.575 186.000 ;
        RECT 84.905 185.965 86.080 186.025 ;
        RECT 83.375 185.855 86.080 185.965 ;
        RECT 83.435 185.795 85.235 185.855 ;
        RECT 84.905 185.765 85.235 185.795 ;
        RECT 81.795 185.475 82.750 185.695 ;
        RECT 82.025 184.845 82.295 185.305 ;
        RECT 82.465 185.015 82.750 185.475 ;
        RECT 83.035 185.015 83.295 185.695 ;
        RECT 83.465 184.845 83.715 185.625 ;
        RECT 83.965 185.595 84.800 185.605 ;
        RECT 85.390 185.595 85.575 185.685 ;
        RECT 83.965 185.395 85.575 185.595 ;
        RECT 83.965 185.015 84.215 185.395 ;
        RECT 85.345 185.355 85.575 185.395 ;
        RECT 85.825 185.235 86.080 185.855 ;
        RECT 84.385 184.845 84.740 185.225 ;
        RECT 85.745 185.015 86.080 185.235 ;
        RECT 86.720 184.845 86.975 185.985 ;
        RECT 87.225 185.595 87.395 186.155 ;
        RECT 88.695 185.985 88.865 186.155 ;
        RECT 89.135 185.985 89.305 186.720 ;
        RECT 87.620 185.815 88.865 185.985 ;
        RECT 87.620 185.565 88.040 185.815 ;
        RECT 87.170 185.065 88.365 185.395 ;
        RECT 88.545 184.845 88.825 185.645 ;
        RECT 89.035 185.015 89.305 185.985 ;
        RECT 89.475 186.720 89.745 187.065 ;
        RECT 89.935 186.995 90.315 187.395 ;
        RECT 90.485 186.825 90.655 187.175 ;
        RECT 90.825 186.915 91.560 187.395 ;
        RECT 89.475 185.985 89.645 186.720 ;
        RECT 89.915 186.655 90.655 186.825 ;
        RECT 91.730 186.745 92.040 187.215 ;
        RECT 89.915 186.485 90.085 186.655 ;
        RECT 91.305 186.575 92.040 186.745 ;
        RECT 92.235 186.625 95.745 187.395 ;
        RECT 91.305 186.485 91.555 186.575 ;
        RECT 89.855 186.155 90.085 186.485 ;
        RECT 90.815 186.155 91.555 186.485 ;
        RECT 91.725 186.155 92.060 186.405 ;
        RECT 89.915 185.985 90.085 186.155 ;
        RECT 89.475 185.015 89.745 185.985 ;
        RECT 89.915 185.815 91.160 185.985 ;
        RECT 89.955 184.845 90.235 185.645 ;
        RECT 90.740 185.565 91.160 185.815 ;
        RECT 91.385 185.595 91.555 186.155 ;
        RECT 92.235 186.105 93.885 186.625 ;
        RECT 90.415 185.065 91.610 185.395 ;
        RECT 91.805 184.845 92.060 185.985 ;
        RECT 94.055 185.935 95.745 186.455 ;
        RECT 92.235 184.845 95.745 185.935 ;
        RECT 96.380 185.795 96.715 187.215 ;
        RECT 96.895 187.025 97.640 187.395 ;
        RECT 98.205 186.855 98.460 187.215 ;
        RECT 98.640 187.025 98.970 187.395 ;
        RECT 99.150 186.855 99.375 187.215 ;
        RECT 96.890 186.665 99.375 186.855 ;
        RECT 100.055 186.670 100.345 187.395 ;
        RECT 101.440 186.890 101.775 187.395 ;
        RECT 101.945 186.825 102.185 187.200 ;
        RECT 102.465 187.065 102.635 187.210 ;
        RECT 102.465 186.870 102.840 187.065 ;
        RECT 103.200 186.900 103.595 187.395 ;
        RECT 96.890 185.975 97.115 186.665 ;
        RECT 97.315 186.155 97.595 186.485 ;
        RECT 97.775 186.155 98.350 186.485 ;
        RECT 98.530 186.155 98.965 186.485 ;
        RECT 99.145 186.155 99.415 186.485 ;
        RECT 96.890 185.795 99.385 185.975 ;
        RECT 96.380 185.025 96.645 185.795 ;
        RECT 96.815 184.845 97.145 185.565 ;
        RECT 97.335 185.385 98.525 185.615 ;
        RECT 97.335 185.025 97.595 185.385 ;
        RECT 97.765 184.845 98.095 185.215 ;
        RECT 98.265 185.025 98.525 185.385 ;
        RECT 99.095 185.025 99.385 185.795 ;
        RECT 100.055 184.845 100.345 186.010 ;
        RECT 101.495 185.865 101.795 186.715 ;
        RECT 101.965 186.675 102.185 186.825 ;
        RECT 101.965 186.345 102.500 186.675 ;
        RECT 102.670 186.535 102.840 186.870 ;
        RECT 103.765 186.705 104.005 187.225 ;
        RECT 101.965 185.695 102.200 186.345 ;
        RECT 102.670 186.175 103.655 186.535 ;
        RECT 101.525 185.465 102.200 185.695 ;
        RECT 102.370 186.155 103.655 186.175 ;
        RECT 102.370 186.005 103.230 186.155 ;
        RECT 101.525 185.035 101.695 185.465 ;
        RECT 101.865 184.845 102.195 185.295 ;
        RECT 102.370 185.060 102.655 186.005 ;
        RECT 103.830 185.900 104.005 186.705 ;
        RECT 104.745 186.845 104.915 187.225 ;
        RECT 105.130 187.015 105.460 187.395 ;
        RECT 104.745 186.675 105.460 186.845 ;
        RECT 104.655 186.125 105.010 186.495 ;
        RECT 105.290 186.485 105.460 186.675 ;
        RECT 105.630 186.650 105.885 187.225 ;
        RECT 105.290 186.155 105.545 186.485 ;
        RECT 105.290 185.945 105.460 186.155 ;
        RECT 102.830 185.525 103.525 185.835 ;
        RECT 102.835 184.845 103.520 185.315 ;
        RECT 103.700 185.115 104.005 185.900 ;
        RECT 104.745 185.775 105.460 185.945 ;
        RECT 105.715 185.920 105.885 186.650 ;
        RECT 106.060 186.555 106.320 187.395 ;
        RECT 107.015 186.575 107.225 187.395 ;
        RECT 107.395 186.595 107.725 187.225 ;
        RECT 107.395 185.995 107.645 186.595 ;
        RECT 107.895 186.575 108.125 187.395 ;
        RECT 108.795 187.015 109.685 187.185 ;
        RECT 108.795 186.460 109.345 186.845 ;
        RECT 107.815 186.155 108.145 186.405 ;
        RECT 109.515 186.290 109.685 187.015 ;
        RECT 108.795 186.220 109.685 186.290 ;
        RECT 109.855 186.690 110.075 187.175 ;
        RECT 110.245 186.855 110.495 187.395 ;
        RECT 110.665 186.745 110.925 187.225 ;
        RECT 109.855 186.265 110.185 186.690 ;
        RECT 108.795 186.195 109.690 186.220 ;
        RECT 108.795 186.180 109.700 186.195 ;
        RECT 108.795 186.165 109.705 186.180 ;
        RECT 108.795 186.160 109.715 186.165 ;
        RECT 108.795 186.150 109.720 186.160 ;
        RECT 108.795 186.140 109.725 186.150 ;
        RECT 108.795 186.135 109.735 186.140 ;
        RECT 108.795 186.125 109.745 186.135 ;
        RECT 108.795 186.120 109.755 186.125 ;
        RECT 104.745 185.015 104.915 185.775 ;
        RECT 105.130 184.845 105.460 185.605 ;
        RECT 105.630 185.015 105.885 185.920 ;
        RECT 106.060 184.845 106.320 185.995 ;
        RECT 107.015 184.845 107.225 185.985 ;
        RECT 107.395 185.015 107.725 185.995 ;
        RECT 107.895 184.845 108.125 185.985 ;
        RECT 108.795 185.670 109.055 186.120 ;
        RECT 109.420 186.115 109.755 186.120 ;
        RECT 109.420 186.110 109.770 186.115 ;
        RECT 109.420 186.100 109.785 186.110 ;
        RECT 109.420 186.095 109.810 186.100 ;
        RECT 110.355 186.095 110.585 186.490 ;
        RECT 109.420 186.090 110.585 186.095 ;
        RECT 109.450 186.055 110.585 186.090 ;
        RECT 109.485 186.030 110.585 186.055 ;
        RECT 109.515 186.000 110.585 186.030 ;
        RECT 109.535 185.970 110.585 186.000 ;
        RECT 109.555 185.940 110.585 185.970 ;
        RECT 109.625 185.930 110.585 185.940 ;
        RECT 109.650 185.920 110.585 185.930 ;
        RECT 109.670 185.905 110.585 185.920 ;
        RECT 109.690 185.890 110.585 185.905 ;
        RECT 109.695 185.880 110.480 185.890 ;
        RECT 109.710 185.845 110.480 185.880 ;
        RECT 109.225 185.525 109.555 185.770 ;
        RECT 109.725 185.595 110.480 185.845 ;
        RECT 110.755 185.715 110.925 186.745 ;
        RECT 112.065 186.740 112.395 187.175 ;
        RECT 112.565 186.785 112.735 187.395 ;
        RECT 112.015 186.655 112.395 186.740 ;
        RECT 112.905 186.655 113.235 187.180 ;
        RECT 113.495 186.865 113.705 187.395 ;
        RECT 113.980 186.945 114.765 187.115 ;
        RECT 114.935 186.945 115.340 187.115 ;
        RECT 112.015 186.615 112.240 186.655 ;
        RECT 112.015 186.035 112.185 186.615 ;
        RECT 112.905 186.485 113.105 186.655 ;
        RECT 113.980 186.485 114.150 186.945 ;
        RECT 112.355 186.155 113.105 186.485 ;
        RECT 113.275 186.155 114.150 186.485 ;
        RECT 112.015 185.985 112.230 186.035 ;
        RECT 112.015 185.905 112.405 185.985 ;
        RECT 109.225 185.500 109.410 185.525 ;
        RECT 108.795 185.400 109.410 185.500 ;
        RECT 108.795 184.845 109.400 185.400 ;
        RECT 109.575 185.015 110.055 185.355 ;
        RECT 110.225 184.845 110.480 185.390 ;
        RECT 110.650 185.015 110.925 185.715 ;
        RECT 112.075 185.060 112.405 185.905 ;
        RECT 112.915 185.950 113.105 186.155 ;
        RECT 112.575 184.845 112.745 185.855 ;
        RECT 112.915 185.575 113.810 185.950 ;
        RECT 112.915 185.015 113.255 185.575 ;
        RECT 113.485 184.845 113.800 185.345 ;
        RECT 113.980 185.315 114.150 186.155 ;
        RECT 114.320 186.445 114.785 186.775 ;
        RECT 115.170 186.715 115.340 186.945 ;
        RECT 115.520 186.895 115.890 187.395 ;
        RECT 116.210 186.945 116.885 187.115 ;
        RECT 117.080 186.945 117.415 187.115 ;
        RECT 114.320 185.485 114.640 186.445 ;
        RECT 115.170 186.415 116.000 186.715 ;
        RECT 114.810 185.515 115.000 186.235 ;
        RECT 115.170 185.345 115.340 186.415 ;
        RECT 115.800 186.385 116.000 186.415 ;
        RECT 115.510 186.165 115.680 186.235 ;
        RECT 116.210 186.165 116.380 186.945 ;
        RECT 117.245 186.805 117.415 186.945 ;
        RECT 117.585 186.935 117.835 187.395 ;
        RECT 115.510 185.995 116.380 186.165 ;
        RECT 116.550 186.525 117.075 186.745 ;
        RECT 117.245 186.675 117.470 186.805 ;
        RECT 115.510 185.905 116.020 185.995 ;
        RECT 113.980 185.145 114.865 185.315 ;
        RECT 115.090 185.015 115.340 185.345 ;
        RECT 115.510 184.845 115.680 185.645 ;
        RECT 115.850 185.290 116.020 185.905 ;
        RECT 116.550 185.825 116.720 186.525 ;
        RECT 116.190 185.460 116.720 185.825 ;
        RECT 116.890 185.760 117.130 186.355 ;
        RECT 117.300 185.570 117.470 186.675 ;
        RECT 117.640 185.815 117.920 186.765 ;
        RECT 117.165 185.440 117.470 185.570 ;
        RECT 115.850 185.120 116.955 185.290 ;
        RECT 117.165 185.015 117.415 185.440 ;
        RECT 117.585 184.845 117.850 185.305 ;
        RECT 118.090 185.015 118.275 187.135 ;
        RECT 118.445 187.015 118.775 187.395 ;
        RECT 118.945 186.845 119.115 187.135 ;
        RECT 118.450 186.675 119.115 186.845 ;
        RECT 118.450 185.685 118.680 186.675 ;
        RECT 119.375 186.625 122.885 187.395 ;
        RECT 123.515 186.720 123.775 187.225 ;
        RECT 123.955 187.015 124.285 187.395 ;
        RECT 124.465 186.845 124.635 187.225 ;
        RECT 118.850 185.855 119.200 186.505 ;
        RECT 119.375 186.105 121.025 186.625 ;
        RECT 121.195 185.935 122.885 186.455 ;
        RECT 118.450 185.515 119.115 185.685 ;
        RECT 118.445 184.845 118.775 185.345 ;
        RECT 118.945 185.015 119.115 185.515 ;
        RECT 119.375 184.845 122.885 185.935 ;
        RECT 123.515 185.920 123.685 186.720 ;
        RECT 123.970 186.675 124.635 186.845 ;
        RECT 123.970 186.420 124.140 186.675 ;
        RECT 125.815 186.670 126.105 187.395 ;
        RECT 126.275 186.745 126.535 187.225 ;
        RECT 126.705 186.855 126.955 187.395 ;
        RECT 123.855 186.090 124.140 186.420 ;
        RECT 124.375 186.125 124.705 186.495 ;
        RECT 123.970 185.945 124.140 186.090 ;
        RECT 123.515 185.015 123.785 185.920 ;
        RECT 123.970 185.775 124.635 185.945 ;
        RECT 123.955 184.845 124.285 185.605 ;
        RECT 124.465 185.015 124.635 185.775 ;
        RECT 125.815 184.845 126.105 186.010 ;
        RECT 126.275 185.715 126.445 186.745 ;
        RECT 127.125 186.690 127.345 187.175 ;
        RECT 126.615 186.095 126.845 186.490 ;
        RECT 127.015 186.265 127.345 186.690 ;
        RECT 127.515 187.015 128.405 187.185 ;
        RECT 127.515 186.290 127.685 187.015 ;
        RECT 128.580 186.905 128.835 187.395 ;
        RECT 129.005 186.885 130.235 187.225 ;
        RECT 127.855 186.460 128.405 186.845 ;
        RECT 127.515 186.220 128.405 186.290 ;
        RECT 127.510 186.195 128.405 186.220 ;
        RECT 127.500 186.180 128.405 186.195 ;
        RECT 127.495 186.165 128.405 186.180 ;
        RECT 127.485 186.160 128.405 186.165 ;
        RECT 127.480 186.150 128.405 186.160 ;
        RECT 128.600 186.155 128.820 186.735 ;
        RECT 127.475 186.140 128.405 186.150 ;
        RECT 127.465 186.135 128.405 186.140 ;
        RECT 127.455 186.125 128.405 186.135 ;
        RECT 127.445 186.120 128.405 186.125 ;
        RECT 127.445 186.115 127.780 186.120 ;
        RECT 127.430 186.110 127.780 186.115 ;
        RECT 127.415 186.100 127.780 186.110 ;
        RECT 127.390 186.095 127.780 186.100 ;
        RECT 126.615 186.090 127.780 186.095 ;
        RECT 126.615 186.055 127.750 186.090 ;
        RECT 126.615 186.030 127.715 186.055 ;
        RECT 126.615 186.000 127.685 186.030 ;
        RECT 126.615 185.970 127.665 186.000 ;
        RECT 126.615 185.940 127.645 185.970 ;
        RECT 126.615 185.930 127.575 185.940 ;
        RECT 126.615 185.920 127.550 185.930 ;
        RECT 126.615 185.905 127.530 185.920 ;
        RECT 126.615 185.890 127.510 185.905 ;
        RECT 126.720 185.880 127.505 185.890 ;
        RECT 126.720 185.845 127.490 185.880 ;
        RECT 126.275 185.015 126.550 185.715 ;
        RECT 126.720 185.595 127.475 185.845 ;
        RECT 127.645 185.525 127.975 185.770 ;
        RECT 128.145 185.670 128.405 186.120 ;
        RECT 129.005 185.985 129.185 186.885 ;
        RECT 129.355 186.155 129.730 186.715 ;
        RECT 129.905 186.655 130.235 186.885 ;
        RECT 130.415 186.645 131.625 187.395 ;
        RECT 131.820 186.745 132.130 187.215 ;
        RECT 132.300 186.915 133.035 187.395 ;
        RECT 133.205 186.825 133.375 187.175 ;
        RECT 133.545 186.995 133.925 187.395 ;
        RECT 129.935 186.155 130.245 186.485 ;
        RECT 130.415 186.105 130.935 186.645 ;
        RECT 131.820 186.575 132.555 186.745 ;
        RECT 133.205 186.655 133.945 186.825 ;
        RECT 134.115 186.720 134.385 187.065 ;
        RECT 132.305 186.485 132.555 186.575 ;
        RECT 133.775 186.485 133.945 186.655 ;
        RECT 127.790 185.500 127.975 185.525 ;
        RECT 127.790 185.400 128.405 185.500 ;
        RECT 126.720 184.845 126.975 185.390 ;
        RECT 127.145 185.015 127.625 185.355 ;
        RECT 127.800 184.845 128.405 185.400 ;
        RECT 128.580 184.845 128.835 185.985 ;
        RECT 129.005 185.815 130.235 185.985 ;
        RECT 131.105 185.935 131.625 186.475 ;
        RECT 131.800 186.155 132.135 186.405 ;
        RECT 132.305 186.155 133.045 186.485 ;
        RECT 133.775 186.155 134.005 186.485 ;
        RECT 129.005 185.015 129.335 185.815 ;
        RECT 129.505 184.845 129.735 185.645 ;
        RECT 129.905 185.015 130.235 185.815 ;
        RECT 130.415 184.845 131.625 185.935 ;
        RECT 131.800 184.845 132.055 185.985 ;
        RECT 132.305 185.595 132.475 186.155 ;
        RECT 133.775 185.985 133.945 186.155 ;
        RECT 134.215 185.985 134.385 186.720 ;
        RECT 132.700 185.815 133.945 185.985 ;
        RECT 132.700 185.565 133.120 185.815 ;
        RECT 132.250 185.065 133.445 185.395 ;
        RECT 133.625 184.845 133.905 185.645 ;
        RECT 134.115 185.015 134.385 185.985 ;
        RECT 135.475 186.675 135.815 187.185 ;
        RECT 135.475 185.275 135.735 186.675 ;
        RECT 135.985 186.595 136.255 187.395 ;
        RECT 135.910 186.155 136.240 186.405 ;
        RECT 136.435 186.155 136.715 187.125 ;
        RECT 136.895 186.155 137.195 187.125 ;
        RECT 137.375 186.155 137.725 187.120 ;
        RECT 137.945 186.895 138.440 187.225 ;
        RECT 135.925 185.985 136.240 186.155 ;
        RECT 137.945 185.985 138.115 186.895 ;
        RECT 135.925 185.815 138.115 185.985 ;
        RECT 135.475 185.015 135.815 185.275 ;
        RECT 135.985 184.845 136.315 185.645 ;
        RECT 136.780 185.015 137.030 185.815 ;
        RECT 137.215 184.845 137.545 185.565 ;
        RECT 137.765 185.015 138.015 185.815 ;
        RECT 138.285 185.405 138.525 186.715 ;
        RECT 138.700 186.630 139.155 187.395 ;
        RECT 139.430 187.015 140.730 187.225 ;
        RECT 140.985 187.035 141.315 187.395 ;
        RECT 140.560 186.865 140.730 187.015 ;
        RECT 141.485 186.895 141.745 187.225 ;
        RECT 141.515 186.885 141.745 186.895 ;
        RECT 139.630 186.405 139.850 186.805 ;
        RECT 138.695 186.205 139.185 186.405 ;
        RECT 139.375 186.195 139.850 186.405 ;
        RECT 140.095 186.405 140.305 186.805 ;
        RECT 140.560 186.740 141.315 186.865 ;
        RECT 140.560 186.695 141.405 186.740 ;
        RECT 141.135 186.575 141.405 186.695 ;
        RECT 140.095 186.195 140.425 186.405 ;
        RECT 140.595 186.135 141.005 186.440 ;
        RECT 138.700 185.965 139.875 186.025 ;
        RECT 141.235 186.000 141.405 186.575 ;
        RECT 141.205 185.965 141.405 186.000 ;
        RECT 138.700 185.855 141.405 185.965 ;
        RECT 138.700 185.235 138.955 185.855 ;
        RECT 139.545 185.795 141.345 185.855 ;
        RECT 139.545 185.765 139.875 185.795 ;
        RECT 141.575 185.695 141.745 186.885 ;
        RECT 141.915 186.625 144.505 187.395 ;
        RECT 141.915 186.105 143.125 186.625 ;
        RECT 144.675 186.575 144.935 187.395 ;
        RECT 145.105 186.575 145.435 186.995 ;
        RECT 145.615 186.910 146.405 187.175 ;
        RECT 145.185 186.485 145.435 186.575 ;
        RECT 143.295 185.935 144.505 186.455 ;
        RECT 139.205 185.595 139.390 185.685 ;
        RECT 139.980 185.595 140.815 185.605 ;
        RECT 139.205 185.395 140.815 185.595 ;
        RECT 139.205 185.355 139.435 185.395 ;
        RECT 138.185 184.845 138.520 185.225 ;
        RECT 138.700 185.015 139.035 185.235 ;
        RECT 140.040 184.845 140.395 185.225 ;
        RECT 140.565 185.015 140.815 185.395 ;
        RECT 141.065 184.845 141.315 185.625 ;
        RECT 141.485 185.015 141.745 185.695 ;
        RECT 141.915 184.845 144.505 185.935 ;
        RECT 144.675 185.525 145.015 186.405 ;
        RECT 145.185 186.235 145.980 186.485 ;
        RECT 144.675 184.845 144.935 185.355 ;
        RECT 145.185 185.015 145.355 186.235 ;
        RECT 146.150 186.055 146.405 186.910 ;
        RECT 146.575 186.755 146.775 187.175 ;
        RECT 146.965 186.935 147.295 187.395 ;
        RECT 146.575 186.235 146.985 186.755 ;
        RECT 147.465 186.745 147.725 187.225 ;
        RECT 147.155 186.055 147.385 186.485 ;
        RECT 145.595 185.885 147.385 186.055 ;
        RECT 145.595 185.520 145.845 185.885 ;
        RECT 146.015 185.525 146.345 185.715 ;
        RECT 146.565 185.590 147.280 185.885 ;
        RECT 147.555 185.715 147.725 186.745 ;
        RECT 146.015 185.350 146.210 185.525 ;
        RECT 145.595 184.845 146.210 185.350 ;
        RECT 146.380 185.015 146.855 185.355 ;
        RECT 147.025 184.845 147.240 185.390 ;
        RECT 147.450 185.015 147.725 185.715 ;
        RECT 147.895 186.745 148.155 187.225 ;
        RECT 148.325 186.855 148.575 187.395 ;
        RECT 147.895 185.715 148.065 186.745 ;
        RECT 148.745 186.715 148.965 187.175 ;
        RECT 148.715 186.690 148.965 186.715 ;
        RECT 148.235 186.095 148.465 186.490 ;
        RECT 148.635 186.265 148.965 186.690 ;
        RECT 149.135 187.015 150.025 187.185 ;
        RECT 149.135 186.290 149.305 187.015 ;
        RECT 149.475 186.460 150.025 186.845 ;
        RECT 150.195 186.720 150.455 187.225 ;
        RECT 150.635 187.015 150.965 187.395 ;
        RECT 151.145 186.845 151.315 187.225 ;
        RECT 149.135 186.220 150.025 186.290 ;
        RECT 149.130 186.195 150.025 186.220 ;
        RECT 149.120 186.180 150.025 186.195 ;
        RECT 149.115 186.165 150.025 186.180 ;
        RECT 149.105 186.160 150.025 186.165 ;
        RECT 149.100 186.150 150.025 186.160 ;
        RECT 149.095 186.140 150.025 186.150 ;
        RECT 149.085 186.135 150.025 186.140 ;
        RECT 149.075 186.125 150.025 186.135 ;
        RECT 149.065 186.120 150.025 186.125 ;
        RECT 149.065 186.115 149.400 186.120 ;
        RECT 149.050 186.110 149.400 186.115 ;
        RECT 149.035 186.100 149.400 186.110 ;
        RECT 149.010 186.095 149.400 186.100 ;
        RECT 148.235 186.090 149.400 186.095 ;
        RECT 148.235 186.055 149.370 186.090 ;
        RECT 148.235 186.030 149.335 186.055 ;
        RECT 148.235 186.000 149.305 186.030 ;
        RECT 148.235 185.970 149.285 186.000 ;
        RECT 148.235 185.940 149.265 185.970 ;
        RECT 148.235 185.930 149.195 185.940 ;
        RECT 148.235 185.920 149.170 185.930 ;
        RECT 148.235 185.905 149.150 185.920 ;
        RECT 148.235 185.890 149.130 185.905 ;
        RECT 148.340 185.880 149.125 185.890 ;
        RECT 148.340 185.845 149.110 185.880 ;
        RECT 147.895 185.015 148.170 185.715 ;
        RECT 148.340 185.595 149.095 185.845 ;
        RECT 149.265 185.525 149.595 185.770 ;
        RECT 149.765 185.670 150.025 186.120 ;
        RECT 150.195 185.920 150.365 186.720 ;
        RECT 150.650 186.675 151.315 186.845 ;
        RECT 150.650 186.420 150.820 186.675 ;
        RECT 151.575 186.670 151.865 187.395 ;
        RECT 152.035 186.625 155.545 187.395 ;
        RECT 155.715 186.645 156.925 187.395 ;
        RECT 150.535 186.090 150.820 186.420 ;
        RECT 151.055 186.125 151.385 186.495 ;
        RECT 152.035 186.105 153.685 186.625 ;
        RECT 150.650 185.945 150.820 186.090 ;
        RECT 149.410 185.500 149.595 185.525 ;
        RECT 149.410 185.400 150.025 185.500 ;
        RECT 148.340 184.845 148.595 185.390 ;
        RECT 148.765 185.015 149.245 185.355 ;
        RECT 149.420 184.845 150.025 185.400 ;
        RECT 150.195 185.015 150.465 185.920 ;
        RECT 150.650 185.775 151.315 185.945 ;
        RECT 150.635 184.845 150.965 185.605 ;
        RECT 151.145 185.015 151.315 185.775 ;
        RECT 151.575 184.845 151.865 186.010 ;
        RECT 153.855 185.935 155.545 186.455 ;
        RECT 152.035 184.845 155.545 185.935 ;
        RECT 155.715 185.935 156.235 186.475 ;
        RECT 156.405 186.105 156.925 186.645 ;
        RECT 155.715 184.845 156.925 185.935 ;
        RECT 22.690 184.675 157.010 184.845 ;
        RECT 22.775 183.585 23.985 184.675 ;
        RECT 24.155 183.585 26.745 184.675 ;
        RECT 22.775 182.875 23.295 183.415 ;
        RECT 23.465 183.045 23.985 183.585 ;
        RECT 24.155 182.895 25.365 183.415 ;
        RECT 25.535 183.065 26.745 183.585 ;
        RECT 26.915 183.600 27.185 184.505 ;
        RECT 27.355 183.915 27.685 184.675 ;
        RECT 27.865 183.745 28.035 184.505 ;
        RECT 22.775 182.125 23.985 182.875 ;
        RECT 24.155 182.125 26.745 182.895 ;
        RECT 26.915 182.800 27.085 183.600 ;
        RECT 27.370 183.575 28.035 183.745 ;
        RECT 28.295 183.585 30.885 184.675 ;
        RECT 31.255 184.005 31.535 184.675 ;
        RECT 31.705 183.785 32.005 184.335 ;
        RECT 32.205 183.955 32.535 184.675 ;
        RECT 32.725 183.955 33.185 184.505 ;
        RECT 33.355 184.120 33.960 184.675 ;
        RECT 34.135 184.165 34.615 184.505 ;
        RECT 34.785 184.130 35.040 184.675 ;
        RECT 33.355 184.020 33.970 184.120 ;
        RECT 27.370 183.430 27.540 183.575 ;
        RECT 27.255 183.100 27.540 183.430 ;
        RECT 27.370 182.845 27.540 183.100 ;
        RECT 27.775 183.025 28.105 183.395 ;
        RECT 28.295 182.895 29.505 183.415 ;
        RECT 29.675 183.065 30.885 183.585 ;
        RECT 31.070 183.365 31.335 183.725 ;
        RECT 31.705 183.615 32.645 183.785 ;
        RECT 32.475 183.365 32.645 183.615 ;
        RECT 31.070 183.115 31.745 183.365 ;
        RECT 31.965 183.115 32.305 183.365 ;
        RECT 32.475 183.035 32.765 183.365 ;
        RECT 32.475 182.945 32.645 183.035 ;
        RECT 26.915 182.295 27.175 182.800 ;
        RECT 27.370 182.675 28.035 182.845 ;
        RECT 27.355 182.125 27.685 182.505 ;
        RECT 27.865 182.295 28.035 182.675 ;
        RECT 28.295 182.125 30.885 182.895 ;
        RECT 31.255 182.755 32.645 182.945 ;
        RECT 31.255 182.395 31.585 182.755 ;
        RECT 32.935 182.585 33.185 183.955 ;
        RECT 33.785 183.995 33.970 184.020 ;
        RECT 33.355 183.400 33.615 183.850 ;
        RECT 33.785 183.750 34.115 183.995 ;
        RECT 34.285 183.675 35.040 183.925 ;
        RECT 35.210 183.805 35.485 184.505 ;
        RECT 34.270 183.640 35.040 183.675 ;
        RECT 34.255 183.630 35.040 183.640 ;
        RECT 34.250 183.615 35.145 183.630 ;
        RECT 34.230 183.600 35.145 183.615 ;
        RECT 34.210 183.590 35.145 183.600 ;
        RECT 34.185 183.580 35.145 183.590 ;
        RECT 34.115 183.550 35.145 183.580 ;
        RECT 34.095 183.520 35.145 183.550 ;
        RECT 34.075 183.490 35.145 183.520 ;
        RECT 34.045 183.465 35.145 183.490 ;
        RECT 34.010 183.430 35.145 183.465 ;
        RECT 33.980 183.425 35.145 183.430 ;
        RECT 33.980 183.420 34.370 183.425 ;
        RECT 33.980 183.410 34.345 183.420 ;
        RECT 33.980 183.405 34.330 183.410 ;
        RECT 33.980 183.400 34.315 183.405 ;
        RECT 33.355 183.395 34.315 183.400 ;
        RECT 33.355 183.385 34.305 183.395 ;
        RECT 33.355 183.380 34.295 183.385 ;
        RECT 33.355 183.370 34.285 183.380 ;
        RECT 33.355 183.360 34.280 183.370 ;
        RECT 33.355 183.355 34.275 183.360 ;
        RECT 33.355 183.340 34.265 183.355 ;
        RECT 33.355 183.325 34.260 183.340 ;
        RECT 33.355 183.300 34.250 183.325 ;
        RECT 33.355 183.230 34.245 183.300 ;
        RECT 33.355 182.675 33.905 183.060 ;
        RECT 32.205 182.125 32.455 182.585 ;
        RECT 32.625 182.295 33.185 182.585 ;
        RECT 34.075 182.505 34.245 183.230 ;
        RECT 33.355 182.335 34.245 182.505 ;
        RECT 34.415 182.830 34.745 183.255 ;
        RECT 34.915 183.030 35.145 183.425 ;
        RECT 34.415 182.345 34.635 182.830 ;
        RECT 35.315 182.775 35.485 183.805 ;
        RECT 35.655 183.510 35.945 184.675 ;
        RECT 36.205 184.005 36.375 184.505 ;
        RECT 36.545 184.175 36.875 184.675 ;
        RECT 36.205 183.835 36.870 184.005 ;
        RECT 36.120 183.015 36.470 183.665 ;
        RECT 34.805 182.125 35.055 182.665 ;
        RECT 35.225 182.295 35.485 182.775 ;
        RECT 35.655 182.125 35.945 182.850 ;
        RECT 36.640 182.845 36.870 183.835 ;
        RECT 36.205 182.675 36.870 182.845 ;
        RECT 36.205 182.385 36.375 182.675 ;
        RECT 36.545 182.125 36.875 182.505 ;
        RECT 37.045 182.385 37.230 184.505 ;
        RECT 37.470 184.215 37.735 184.675 ;
        RECT 37.905 184.080 38.155 184.505 ;
        RECT 38.365 184.230 39.470 184.400 ;
        RECT 37.850 183.950 38.155 184.080 ;
        RECT 37.400 182.755 37.680 183.705 ;
        RECT 37.850 182.845 38.020 183.950 ;
        RECT 38.190 183.165 38.430 183.760 ;
        RECT 38.600 183.695 39.130 184.060 ;
        RECT 38.600 182.995 38.770 183.695 ;
        RECT 39.300 183.615 39.470 184.230 ;
        RECT 39.640 183.875 39.810 184.675 ;
        RECT 39.980 184.175 40.230 184.505 ;
        RECT 40.455 184.205 41.340 184.375 ;
        RECT 39.300 183.525 39.810 183.615 ;
        RECT 37.850 182.715 38.075 182.845 ;
        RECT 38.245 182.775 38.770 182.995 ;
        RECT 38.940 183.355 39.810 183.525 ;
        RECT 37.485 182.125 37.735 182.585 ;
        RECT 37.905 182.575 38.075 182.715 ;
        RECT 38.940 182.575 39.110 183.355 ;
        RECT 39.640 183.285 39.810 183.355 ;
        RECT 39.320 183.105 39.520 183.135 ;
        RECT 39.980 183.105 40.150 184.175 ;
        RECT 40.320 183.285 40.510 184.005 ;
        RECT 39.320 182.805 40.150 183.105 ;
        RECT 40.680 183.075 41.000 184.035 ;
        RECT 37.905 182.405 38.240 182.575 ;
        RECT 38.435 182.405 39.110 182.575 ;
        RECT 39.430 182.125 39.800 182.625 ;
        RECT 39.980 182.575 40.150 182.805 ;
        RECT 40.535 182.745 41.000 183.075 ;
        RECT 41.170 183.365 41.340 184.205 ;
        RECT 41.520 184.175 41.835 184.675 ;
        RECT 42.065 183.945 42.405 184.505 ;
        RECT 41.510 183.570 42.405 183.945 ;
        RECT 42.575 183.665 42.745 184.675 ;
        RECT 42.215 183.365 42.405 183.570 ;
        RECT 42.915 183.615 43.245 184.460 ;
        RECT 42.915 183.535 43.305 183.615 ;
        RECT 43.475 183.585 44.685 184.675 ;
        RECT 44.945 184.005 45.115 184.505 ;
        RECT 45.285 184.175 45.615 184.675 ;
        RECT 44.945 183.835 45.610 184.005 ;
        RECT 43.090 183.485 43.305 183.535 ;
        RECT 41.170 183.035 42.045 183.365 ;
        RECT 42.215 183.035 42.965 183.365 ;
        RECT 41.170 182.575 41.340 183.035 ;
        RECT 42.215 182.865 42.415 183.035 ;
        RECT 43.135 182.905 43.305 183.485 ;
        RECT 43.080 182.865 43.305 182.905 ;
        RECT 39.980 182.405 40.385 182.575 ;
        RECT 40.555 182.405 41.340 182.575 ;
        RECT 41.615 182.125 41.825 182.655 ;
        RECT 42.085 182.340 42.415 182.865 ;
        RECT 42.925 182.780 43.305 182.865 ;
        RECT 43.475 182.875 43.995 183.415 ;
        RECT 44.165 183.045 44.685 183.585 ;
        RECT 44.860 183.015 45.210 183.665 ;
        RECT 42.585 182.125 42.755 182.735 ;
        RECT 42.925 182.345 43.255 182.780 ;
        RECT 43.475 182.125 44.685 182.875 ;
        RECT 45.380 182.845 45.610 183.835 ;
        RECT 44.945 182.675 45.610 182.845 ;
        RECT 44.945 182.385 45.115 182.675 ;
        RECT 45.285 182.125 45.615 182.505 ;
        RECT 45.785 182.385 45.970 184.505 ;
        RECT 46.210 184.215 46.475 184.675 ;
        RECT 46.645 184.080 46.895 184.505 ;
        RECT 47.105 184.230 48.210 184.400 ;
        RECT 46.590 183.950 46.895 184.080 ;
        RECT 46.140 182.755 46.420 183.705 ;
        RECT 46.590 182.845 46.760 183.950 ;
        RECT 46.930 183.165 47.170 183.760 ;
        RECT 47.340 183.695 47.870 184.060 ;
        RECT 47.340 182.995 47.510 183.695 ;
        RECT 48.040 183.615 48.210 184.230 ;
        RECT 48.380 183.875 48.550 184.675 ;
        RECT 48.720 184.175 48.970 184.505 ;
        RECT 49.195 184.205 50.080 184.375 ;
        RECT 48.040 183.525 48.550 183.615 ;
        RECT 46.590 182.715 46.815 182.845 ;
        RECT 46.985 182.775 47.510 182.995 ;
        RECT 47.680 183.355 48.550 183.525 ;
        RECT 46.225 182.125 46.475 182.585 ;
        RECT 46.645 182.575 46.815 182.715 ;
        RECT 47.680 182.575 47.850 183.355 ;
        RECT 48.380 183.285 48.550 183.355 ;
        RECT 48.060 183.105 48.260 183.135 ;
        RECT 48.720 183.105 48.890 184.175 ;
        RECT 49.060 183.285 49.250 184.005 ;
        RECT 48.060 182.805 48.890 183.105 ;
        RECT 49.420 183.075 49.740 184.035 ;
        RECT 46.645 182.405 46.980 182.575 ;
        RECT 47.175 182.405 47.850 182.575 ;
        RECT 48.170 182.125 48.540 182.625 ;
        RECT 48.720 182.575 48.890 182.805 ;
        RECT 49.275 182.745 49.740 183.075 ;
        RECT 49.910 183.365 50.080 184.205 ;
        RECT 50.260 184.175 50.575 184.675 ;
        RECT 50.805 183.945 51.145 184.505 ;
        RECT 50.250 183.570 51.145 183.945 ;
        RECT 51.315 183.665 51.485 184.675 ;
        RECT 50.955 183.365 51.145 183.570 ;
        RECT 51.655 183.615 51.985 184.460 ;
        RECT 51.655 183.535 52.045 183.615 ;
        RECT 51.830 183.485 52.045 183.535 ;
        RECT 49.910 183.035 50.785 183.365 ;
        RECT 50.955 183.035 51.705 183.365 ;
        RECT 49.910 182.575 50.080 183.035 ;
        RECT 50.955 182.865 51.155 183.035 ;
        RECT 51.875 182.905 52.045 183.485 ;
        RECT 51.820 182.865 52.045 182.905 ;
        RECT 48.720 182.405 49.125 182.575 ;
        RECT 49.295 182.405 50.080 182.575 ;
        RECT 50.355 182.125 50.565 182.655 ;
        RECT 50.825 182.340 51.155 182.865 ;
        RECT 51.665 182.780 52.045 182.865 ;
        RECT 52.215 183.535 52.600 184.505 ;
        RECT 52.770 184.215 53.095 184.675 ;
        RECT 53.615 184.045 53.895 184.505 ;
        RECT 52.770 183.825 53.895 184.045 ;
        RECT 52.215 182.865 52.495 183.535 ;
        RECT 52.770 183.365 53.220 183.825 ;
        RECT 54.085 183.655 54.485 184.505 ;
        RECT 54.885 184.215 55.155 184.675 ;
        RECT 55.325 184.045 55.610 184.505 ;
        RECT 52.665 183.035 53.220 183.365 ;
        RECT 53.390 183.095 54.485 183.655 ;
        RECT 52.770 182.925 53.220 183.035 ;
        RECT 51.325 182.125 51.495 182.735 ;
        RECT 51.665 182.345 51.995 182.780 ;
        RECT 52.215 182.295 52.600 182.865 ;
        RECT 52.770 182.755 53.895 182.925 ;
        RECT 52.770 182.125 53.095 182.585 ;
        RECT 53.615 182.295 53.895 182.755 ;
        RECT 54.085 182.295 54.485 183.095 ;
        RECT 54.655 183.825 55.610 184.045 ;
        RECT 54.655 182.925 54.865 183.825 ;
        RECT 55.035 183.095 55.725 183.655 ;
        RECT 55.895 183.495 56.215 184.675 ;
        RECT 56.385 183.655 56.585 184.445 ;
        RECT 56.910 183.845 57.295 184.505 ;
        RECT 57.690 183.915 58.475 184.675 ;
        RECT 56.885 183.745 57.295 183.845 ;
        RECT 56.385 183.485 56.715 183.655 ;
        RECT 56.885 183.535 58.495 183.745 ;
        RECT 56.535 183.365 56.715 183.485 ;
        RECT 55.895 183.115 56.360 183.315 ;
        RECT 56.535 183.115 56.865 183.365 ;
        RECT 57.035 183.315 57.500 183.365 ;
        RECT 57.035 183.145 57.505 183.315 ;
        RECT 57.035 183.115 57.500 183.145 ;
        RECT 57.695 183.115 58.050 183.365 ;
        RECT 58.220 182.935 58.495 183.535 ;
        RECT 54.655 182.755 55.610 182.925 ;
        RECT 54.885 182.125 55.155 182.585 ;
        RECT 55.325 182.295 55.610 182.755 ;
        RECT 55.895 182.735 57.075 182.905 ;
        RECT 55.895 182.320 56.235 182.735 ;
        RECT 56.405 182.125 56.575 182.565 ;
        RECT 56.745 182.515 57.075 182.735 ;
        RECT 57.245 182.755 58.495 182.935 ;
        RECT 57.245 182.685 57.610 182.755 ;
        RECT 56.745 182.335 57.995 182.515 ;
        RECT 58.265 182.125 58.435 182.585 ;
        RECT 58.665 182.405 58.945 184.505 ;
        RECT 59.175 183.535 59.385 184.675 ;
        RECT 59.555 183.525 59.885 184.505 ;
        RECT 60.055 183.535 60.285 184.675 ;
        RECT 59.175 182.125 59.385 182.945 ;
        RECT 59.555 182.925 59.805 183.525 ;
        RECT 61.415 183.510 61.705 184.675 ;
        RECT 61.935 183.535 62.145 184.675 ;
        RECT 62.315 183.525 62.645 184.505 ;
        RECT 62.815 183.535 63.045 184.675 ;
        RECT 63.345 184.005 63.515 184.505 ;
        RECT 63.685 184.175 64.015 184.675 ;
        RECT 63.345 183.835 64.010 184.005 ;
        RECT 59.975 183.115 60.305 183.365 ;
        RECT 59.555 182.295 59.885 182.925 ;
        RECT 60.055 182.125 60.285 182.945 ;
        RECT 61.415 182.125 61.705 182.850 ;
        RECT 61.935 182.125 62.145 182.945 ;
        RECT 62.315 182.925 62.565 183.525 ;
        RECT 62.735 183.115 63.065 183.365 ;
        RECT 63.260 183.015 63.610 183.665 ;
        RECT 62.315 182.295 62.645 182.925 ;
        RECT 62.815 182.125 63.045 182.945 ;
        RECT 63.780 182.845 64.010 183.835 ;
        RECT 63.345 182.675 64.010 182.845 ;
        RECT 63.345 182.385 63.515 182.675 ;
        RECT 63.685 182.125 64.015 182.505 ;
        RECT 64.185 182.385 64.370 184.505 ;
        RECT 64.610 184.215 64.875 184.675 ;
        RECT 65.045 184.080 65.295 184.505 ;
        RECT 65.505 184.230 66.610 184.400 ;
        RECT 64.990 183.950 65.295 184.080 ;
        RECT 64.540 182.755 64.820 183.705 ;
        RECT 64.990 182.845 65.160 183.950 ;
        RECT 65.330 183.165 65.570 183.760 ;
        RECT 65.740 183.695 66.270 184.060 ;
        RECT 65.740 182.995 65.910 183.695 ;
        RECT 66.440 183.615 66.610 184.230 ;
        RECT 66.780 183.875 66.950 184.675 ;
        RECT 67.120 184.175 67.370 184.505 ;
        RECT 67.595 184.205 68.480 184.375 ;
        RECT 66.440 183.525 66.950 183.615 ;
        RECT 64.990 182.715 65.215 182.845 ;
        RECT 65.385 182.775 65.910 182.995 ;
        RECT 66.080 183.355 66.950 183.525 ;
        RECT 64.625 182.125 64.875 182.585 ;
        RECT 65.045 182.575 65.215 182.715 ;
        RECT 66.080 182.575 66.250 183.355 ;
        RECT 66.780 183.285 66.950 183.355 ;
        RECT 66.460 183.105 66.660 183.135 ;
        RECT 67.120 183.105 67.290 184.175 ;
        RECT 67.460 183.285 67.650 184.005 ;
        RECT 66.460 182.805 67.290 183.105 ;
        RECT 67.820 183.075 68.140 184.035 ;
        RECT 65.045 182.405 65.380 182.575 ;
        RECT 65.575 182.405 66.250 182.575 ;
        RECT 66.570 182.125 66.940 182.625 ;
        RECT 67.120 182.575 67.290 182.805 ;
        RECT 67.675 182.745 68.140 183.075 ;
        RECT 68.310 183.365 68.480 184.205 ;
        RECT 68.660 184.175 68.975 184.675 ;
        RECT 69.205 183.945 69.545 184.505 ;
        RECT 68.650 183.570 69.545 183.945 ;
        RECT 69.715 183.665 69.885 184.675 ;
        RECT 69.355 183.365 69.545 183.570 ;
        RECT 70.055 183.615 70.385 184.460 ;
        RECT 70.705 184.005 70.875 184.505 ;
        RECT 71.045 184.175 71.375 184.675 ;
        RECT 70.705 183.835 71.370 184.005 ;
        RECT 70.055 183.535 70.445 183.615 ;
        RECT 70.230 183.485 70.445 183.535 ;
        RECT 68.310 183.035 69.185 183.365 ;
        RECT 69.355 183.035 70.105 183.365 ;
        RECT 68.310 182.575 68.480 183.035 ;
        RECT 69.355 182.865 69.555 183.035 ;
        RECT 70.275 182.905 70.445 183.485 ;
        RECT 70.620 183.015 70.970 183.665 ;
        RECT 70.220 182.865 70.445 182.905 ;
        RECT 67.120 182.405 67.525 182.575 ;
        RECT 67.695 182.405 68.480 182.575 ;
        RECT 68.755 182.125 68.965 182.655 ;
        RECT 69.225 182.340 69.555 182.865 ;
        RECT 70.065 182.780 70.445 182.865 ;
        RECT 71.140 182.845 71.370 183.835 ;
        RECT 69.725 182.125 69.895 182.735 ;
        RECT 70.065 182.345 70.395 182.780 ;
        RECT 70.705 182.675 71.370 182.845 ;
        RECT 70.705 182.385 70.875 182.675 ;
        RECT 71.045 182.125 71.375 182.505 ;
        RECT 71.545 182.385 71.730 184.505 ;
        RECT 71.970 184.215 72.235 184.675 ;
        RECT 72.405 184.080 72.655 184.505 ;
        RECT 72.865 184.230 73.970 184.400 ;
        RECT 72.350 183.950 72.655 184.080 ;
        RECT 71.900 182.755 72.180 183.705 ;
        RECT 72.350 182.845 72.520 183.950 ;
        RECT 72.690 183.165 72.930 183.760 ;
        RECT 73.100 183.695 73.630 184.060 ;
        RECT 73.100 182.995 73.270 183.695 ;
        RECT 73.800 183.615 73.970 184.230 ;
        RECT 74.140 183.875 74.310 184.675 ;
        RECT 74.480 184.175 74.730 184.505 ;
        RECT 74.955 184.205 75.840 184.375 ;
        RECT 73.800 183.525 74.310 183.615 ;
        RECT 72.350 182.715 72.575 182.845 ;
        RECT 72.745 182.775 73.270 182.995 ;
        RECT 73.440 183.355 74.310 183.525 ;
        RECT 71.985 182.125 72.235 182.585 ;
        RECT 72.405 182.575 72.575 182.715 ;
        RECT 73.440 182.575 73.610 183.355 ;
        RECT 74.140 183.285 74.310 183.355 ;
        RECT 73.820 183.105 74.020 183.135 ;
        RECT 74.480 183.105 74.650 184.175 ;
        RECT 74.820 183.285 75.010 184.005 ;
        RECT 73.820 182.805 74.650 183.105 ;
        RECT 75.180 183.075 75.500 184.035 ;
        RECT 72.405 182.405 72.740 182.575 ;
        RECT 72.935 182.405 73.610 182.575 ;
        RECT 73.930 182.125 74.300 182.625 ;
        RECT 74.480 182.575 74.650 182.805 ;
        RECT 75.035 182.745 75.500 183.075 ;
        RECT 75.670 183.365 75.840 184.205 ;
        RECT 76.020 184.175 76.335 184.675 ;
        RECT 76.565 183.945 76.905 184.505 ;
        RECT 76.010 183.570 76.905 183.945 ;
        RECT 77.075 183.665 77.245 184.675 ;
        RECT 76.715 183.365 76.905 183.570 ;
        RECT 77.415 183.615 77.745 184.460 ;
        RECT 78.065 184.005 78.235 184.505 ;
        RECT 78.405 184.175 78.735 184.675 ;
        RECT 78.065 183.835 78.730 184.005 ;
        RECT 77.415 183.535 77.805 183.615 ;
        RECT 77.590 183.485 77.805 183.535 ;
        RECT 75.670 183.035 76.545 183.365 ;
        RECT 76.715 183.035 77.465 183.365 ;
        RECT 75.670 182.575 75.840 183.035 ;
        RECT 76.715 182.865 76.915 183.035 ;
        RECT 77.635 182.905 77.805 183.485 ;
        RECT 77.980 183.015 78.330 183.665 ;
        RECT 77.580 182.865 77.805 182.905 ;
        RECT 74.480 182.405 74.885 182.575 ;
        RECT 75.055 182.405 75.840 182.575 ;
        RECT 76.115 182.125 76.325 182.655 ;
        RECT 76.585 182.340 76.915 182.865 ;
        RECT 77.425 182.780 77.805 182.865 ;
        RECT 78.500 182.845 78.730 183.835 ;
        RECT 77.085 182.125 77.255 182.735 ;
        RECT 77.425 182.345 77.755 182.780 ;
        RECT 78.065 182.675 78.730 182.845 ;
        RECT 78.065 182.385 78.235 182.675 ;
        RECT 78.405 182.125 78.735 182.505 ;
        RECT 78.905 182.385 79.090 184.505 ;
        RECT 79.330 184.215 79.595 184.675 ;
        RECT 79.765 184.080 80.015 184.505 ;
        RECT 80.225 184.230 81.330 184.400 ;
        RECT 79.710 183.950 80.015 184.080 ;
        RECT 79.260 182.755 79.540 183.705 ;
        RECT 79.710 182.845 79.880 183.950 ;
        RECT 80.050 183.165 80.290 183.760 ;
        RECT 80.460 183.695 80.990 184.060 ;
        RECT 80.460 182.995 80.630 183.695 ;
        RECT 81.160 183.615 81.330 184.230 ;
        RECT 81.500 183.875 81.670 184.675 ;
        RECT 81.840 184.175 82.090 184.505 ;
        RECT 82.315 184.205 83.200 184.375 ;
        RECT 81.160 183.525 81.670 183.615 ;
        RECT 79.710 182.715 79.935 182.845 ;
        RECT 80.105 182.775 80.630 182.995 ;
        RECT 80.800 183.355 81.670 183.525 ;
        RECT 79.345 182.125 79.595 182.585 ;
        RECT 79.765 182.575 79.935 182.715 ;
        RECT 80.800 182.575 80.970 183.355 ;
        RECT 81.500 183.285 81.670 183.355 ;
        RECT 81.180 183.105 81.380 183.135 ;
        RECT 81.840 183.105 82.010 184.175 ;
        RECT 82.180 183.285 82.370 184.005 ;
        RECT 81.180 182.805 82.010 183.105 ;
        RECT 82.540 183.075 82.860 184.035 ;
        RECT 79.765 182.405 80.100 182.575 ;
        RECT 80.295 182.405 80.970 182.575 ;
        RECT 81.290 182.125 81.660 182.625 ;
        RECT 81.840 182.575 82.010 182.805 ;
        RECT 82.395 182.745 82.860 183.075 ;
        RECT 83.030 183.365 83.200 184.205 ;
        RECT 83.380 184.175 83.695 184.675 ;
        RECT 83.925 183.945 84.265 184.505 ;
        RECT 83.370 183.570 84.265 183.945 ;
        RECT 84.435 183.665 84.605 184.675 ;
        RECT 84.075 183.365 84.265 183.570 ;
        RECT 84.775 183.615 85.105 184.460 ;
        RECT 84.775 183.535 85.165 183.615 ;
        RECT 85.795 183.535 86.075 184.675 ;
        RECT 84.950 183.485 85.165 183.535 ;
        RECT 86.245 183.525 86.575 184.505 ;
        RECT 86.745 183.535 87.005 184.675 ;
        RECT 83.030 183.035 83.905 183.365 ;
        RECT 84.075 183.035 84.825 183.365 ;
        RECT 83.030 182.575 83.200 183.035 ;
        RECT 84.075 182.865 84.275 183.035 ;
        RECT 84.995 182.905 85.165 183.485 ;
        RECT 86.310 183.485 86.485 183.525 ;
        RECT 87.175 183.510 87.465 184.675 ;
        RECT 87.635 183.535 88.020 184.505 ;
        RECT 88.190 184.215 88.515 184.675 ;
        RECT 89.035 184.045 89.315 184.505 ;
        RECT 88.190 183.825 89.315 184.045 ;
        RECT 85.805 183.095 86.140 183.365 ;
        RECT 86.310 182.925 86.480 183.485 ;
        RECT 86.650 183.115 86.985 183.365 ;
        RECT 84.940 182.865 85.165 182.905 ;
        RECT 81.840 182.405 82.245 182.575 ;
        RECT 82.415 182.405 83.200 182.575 ;
        RECT 83.475 182.125 83.685 182.655 ;
        RECT 83.945 182.340 84.275 182.865 ;
        RECT 84.785 182.780 85.165 182.865 ;
        RECT 84.445 182.125 84.615 182.735 ;
        RECT 84.785 182.345 85.115 182.780 ;
        RECT 85.795 182.125 86.105 182.925 ;
        RECT 86.310 182.295 87.005 182.925 ;
        RECT 87.635 182.865 87.915 183.535 ;
        RECT 88.190 183.365 88.640 183.825 ;
        RECT 89.505 183.655 89.905 184.505 ;
        RECT 90.305 184.215 90.575 184.675 ;
        RECT 90.745 184.045 91.030 184.505 ;
        RECT 88.085 183.035 88.640 183.365 ;
        RECT 88.810 183.095 89.905 183.655 ;
        RECT 88.190 182.925 88.640 183.035 ;
        RECT 87.175 182.125 87.465 182.850 ;
        RECT 87.635 182.295 88.020 182.865 ;
        RECT 88.190 182.755 89.315 182.925 ;
        RECT 88.190 182.125 88.515 182.585 ;
        RECT 89.035 182.295 89.315 182.755 ;
        RECT 89.505 182.295 89.905 183.095 ;
        RECT 90.075 183.825 91.030 184.045 ;
        RECT 91.780 184.285 92.115 184.505 ;
        RECT 93.120 184.295 93.475 184.675 ;
        RECT 90.075 182.925 90.285 183.825 ;
        RECT 91.780 183.665 92.035 184.285 ;
        RECT 92.285 184.125 92.515 184.165 ;
        RECT 93.645 184.125 93.895 184.505 ;
        RECT 92.285 183.925 93.895 184.125 ;
        RECT 92.285 183.835 92.470 183.925 ;
        RECT 93.060 183.915 93.895 183.925 ;
        RECT 94.145 183.895 94.395 184.675 ;
        RECT 94.565 183.825 94.825 184.505 ;
        RECT 92.625 183.725 92.955 183.755 ;
        RECT 92.625 183.665 94.425 183.725 ;
        RECT 90.455 183.095 91.145 183.655 ;
        RECT 91.780 183.555 94.485 183.665 ;
        RECT 91.780 183.495 92.955 183.555 ;
        RECT 94.285 183.520 94.485 183.555 ;
        RECT 91.775 183.115 92.265 183.315 ;
        RECT 92.455 183.115 92.930 183.325 ;
        RECT 90.075 182.755 91.030 182.925 ;
        RECT 90.305 182.125 90.575 182.585 ;
        RECT 90.745 182.295 91.030 182.755 ;
        RECT 91.780 182.125 92.235 182.890 ;
        RECT 92.710 182.715 92.930 183.115 ;
        RECT 93.175 183.115 93.505 183.325 ;
        RECT 93.175 182.715 93.385 183.115 ;
        RECT 93.675 183.080 94.085 183.385 ;
        RECT 94.315 182.945 94.485 183.520 ;
        RECT 94.215 182.825 94.485 182.945 ;
        RECT 93.640 182.780 94.485 182.825 ;
        RECT 93.640 182.655 94.395 182.780 ;
        RECT 93.640 182.505 93.810 182.655 ;
        RECT 94.655 182.625 94.825 183.825 ;
        RECT 95.975 183.615 96.305 184.460 ;
        RECT 96.475 183.665 96.645 184.675 ;
        RECT 96.815 183.945 97.155 184.505 ;
        RECT 97.385 184.175 97.700 184.675 ;
        RECT 97.880 184.205 98.765 184.375 ;
        RECT 95.915 183.535 96.305 183.615 ;
        RECT 96.815 183.570 97.710 183.945 ;
        RECT 95.915 183.485 96.130 183.535 ;
        RECT 95.915 182.905 96.085 183.485 ;
        RECT 96.815 183.365 97.005 183.570 ;
        RECT 97.880 183.365 98.050 184.205 ;
        RECT 98.990 184.175 99.240 184.505 ;
        RECT 96.255 183.035 97.005 183.365 ;
        RECT 97.175 183.035 98.050 183.365 ;
        RECT 95.915 182.865 96.140 182.905 ;
        RECT 96.805 182.865 97.005 183.035 ;
        RECT 95.915 182.780 96.295 182.865 ;
        RECT 92.510 182.295 93.810 182.505 ;
        RECT 94.065 182.125 94.395 182.485 ;
        RECT 94.565 182.295 94.825 182.625 ;
        RECT 95.965 182.345 96.295 182.780 ;
        RECT 96.465 182.125 96.635 182.735 ;
        RECT 96.805 182.340 97.135 182.865 ;
        RECT 97.395 182.125 97.605 182.655 ;
        RECT 97.880 182.575 98.050 183.035 ;
        RECT 98.220 183.075 98.540 184.035 ;
        RECT 98.710 183.285 98.900 184.005 ;
        RECT 99.070 183.105 99.240 184.175 ;
        RECT 99.410 183.875 99.580 184.675 ;
        RECT 99.750 184.230 100.855 184.400 ;
        RECT 99.750 183.615 99.920 184.230 ;
        RECT 101.065 184.080 101.315 184.505 ;
        RECT 101.485 184.215 101.750 184.675 ;
        RECT 100.090 183.695 100.620 184.060 ;
        RECT 101.065 183.950 101.370 184.080 ;
        RECT 99.410 183.525 99.920 183.615 ;
        RECT 99.410 183.355 100.280 183.525 ;
        RECT 99.410 183.285 99.580 183.355 ;
        RECT 99.700 183.105 99.900 183.135 ;
        RECT 98.220 182.745 98.685 183.075 ;
        RECT 99.070 182.805 99.900 183.105 ;
        RECT 99.070 182.575 99.240 182.805 ;
        RECT 97.880 182.405 98.665 182.575 ;
        RECT 98.835 182.405 99.240 182.575 ;
        RECT 99.420 182.125 99.790 182.625 ;
        RECT 100.110 182.575 100.280 183.355 ;
        RECT 100.450 182.995 100.620 183.695 ;
        RECT 100.790 183.165 101.030 183.760 ;
        RECT 100.450 182.775 100.975 182.995 ;
        RECT 101.200 182.845 101.370 183.950 ;
        RECT 101.145 182.715 101.370 182.845 ;
        RECT 101.540 182.755 101.820 183.705 ;
        RECT 101.145 182.575 101.315 182.715 ;
        RECT 100.110 182.405 100.785 182.575 ;
        RECT 100.980 182.405 101.315 182.575 ;
        RECT 101.485 182.125 101.735 182.585 ;
        RECT 101.990 182.385 102.175 184.505 ;
        RECT 102.345 184.175 102.675 184.675 ;
        RECT 102.845 184.005 103.015 184.505 ;
        RECT 103.275 184.240 108.620 184.675 ;
        RECT 102.350 183.835 103.015 184.005 ;
        RECT 102.350 182.845 102.580 183.835 ;
        RECT 102.750 183.015 103.100 183.665 ;
        RECT 102.350 182.675 103.015 182.845 ;
        RECT 102.345 182.125 102.675 182.505 ;
        RECT 102.845 182.385 103.015 182.675 ;
        RECT 104.860 182.670 105.200 183.500 ;
        RECT 106.680 182.990 107.030 184.240 ;
        RECT 109.440 183.705 109.830 183.880 ;
        RECT 110.315 183.875 110.645 184.675 ;
        RECT 110.815 183.885 111.350 184.505 ;
        RECT 109.440 183.535 110.865 183.705 ;
        RECT 109.315 182.805 109.670 183.365 ;
        RECT 103.275 182.125 108.620 182.670 ;
        RECT 109.840 182.635 110.010 183.535 ;
        RECT 110.180 182.805 110.445 183.365 ;
        RECT 110.695 183.035 110.865 183.535 ;
        RECT 111.035 182.865 111.350 183.885 ;
        RECT 111.615 183.535 111.825 184.675 ;
        RECT 111.995 183.525 112.325 184.505 ;
        RECT 112.495 183.535 112.725 184.675 ;
        RECT 109.420 182.125 109.660 182.635 ;
        RECT 109.840 182.305 110.120 182.635 ;
        RECT 110.350 182.125 110.565 182.635 ;
        RECT 110.735 182.295 111.350 182.865 ;
        RECT 111.615 182.125 111.825 182.945 ;
        RECT 111.995 182.925 112.245 183.525 ;
        RECT 112.935 183.510 113.225 184.675 ;
        RECT 113.485 183.745 113.655 184.505 ;
        RECT 113.835 183.915 114.165 184.675 ;
        RECT 113.485 183.575 114.150 183.745 ;
        RECT 114.335 183.600 114.605 184.505 ;
        RECT 114.775 184.240 120.120 184.675 ;
        RECT 113.980 183.430 114.150 183.575 ;
        RECT 112.415 183.115 112.745 183.365 ;
        RECT 113.415 183.025 113.745 183.395 ;
        RECT 113.980 183.100 114.265 183.430 ;
        RECT 111.995 182.295 112.325 182.925 ;
        RECT 112.495 182.125 112.725 182.945 ;
        RECT 112.935 182.125 113.225 182.850 ;
        RECT 113.980 182.845 114.150 183.100 ;
        RECT 113.485 182.675 114.150 182.845 ;
        RECT 114.435 182.800 114.605 183.600 ;
        RECT 113.485 182.295 113.655 182.675 ;
        RECT 113.835 182.125 114.165 182.505 ;
        RECT 114.345 182.295 114.605 182.800 ;
        RECT 116.360 182.670 116.700 183.500 ;
        RECT 118.180 182.990 118.530 184.240 ;
        RECT 121.305 184.005 121.475 184.505 ;
        RECT 121.645 184.175 121.975 184.675 ;
        RECT 121.305 183.835 121.970 184.005 ;
        RECT 121.220 183.015 121.570 183.665 ;
        RECT 121.740 182.845 121.970 183.835 ;
        RECT 121.305 182.675 121.970 182.845 ;
        RECT 114.775 182.125 120.120 182.670 ;
        RECT 121.305 182.385 121.475 182.675 ;
        RECT 121.645 182.125 121.975 182.505 ;
        RECT 122.145 182.385 122.330 184.505 ;
        RECT 122.570 184.215 122.835 184.675 ;
        RECT 123.005 184.080 123.255 184.505 ;
        RECT 123.465 184.230 124.570 184.400 ;
        RECT 122.950 183.950 123.255 184.080 ;
        RECT 122.500 182.755 122.780 183.705 ;
        RECT 122.950 182.845 123.120 183.950 ;
        RECT 123.290 183.165 123.530 183.760 ;
        RECT 123.700 183.695 124.230 184.060 ;
        RECT 123.700 182.995 123.870 183.695 ;
        RECT 124.400 183.615 124.570 184.230 ;
        RECT 124.740 183.875 124.910 184.675 ;
        RECT 125.080 184.175 125.330 184.505 ;
        RECT 125.555 184.205 126.440 184.375 ;
        RECT 124.400 183.525 124.910 183.615 ;
        RECT 122.950 182.715 123.175 182.845 ;
        RECT 123.345 182.775 123.870 182.995 ;
        RECT 124.040 183.355 124.910 183.525 ;
        RECT 122.585 182.125 122.835 182.585 ;
        RECT 123.005 182.575 123.175 182.715 ;
        RECT 124.040 182.575 124.210 183.355 ;
        RECT 124.740 183.285 124.910 183.355 ;
        RECT 124.420 183.105 124.620 183.135 ;
        RECT 125.080 183.105 125.250 184.175 ;
        RECT 125.420 183.285 125.610 184.005 ;
        RECT 124.420 182.805 125.250 183.105 ;
        RECT 125.780 183.075 126.100 184.035 ;
        RECT 123.005 182.405 123.340 182.575 ;
        RECT 123.535 182.405 124.210 182.575 ;
        RECT 124.530 182.125 124.900 182.625 ;
        RECT 125.080 182.575 125.250 182.805 ;
        RECT 125.635 182.745 126.100 183.075 ;
        RECT 126.270 183.365 126.440 184.205 ;
        RECT 126.620 184.175 126.935 184.675 ;
        RECT 127.165 183.945 127.505 184.505 ;
        RECT 126.610 183.570 127.505 183.945 ;
        RECT 127.675 183.665 127.845 184.675 ;
        RECT 127.315 183.365 127.505 183.570 ;
        RECT 128.015 183.615 128.345 184.460 ;
        RECT 128.015 183.535 128.405 183.615 ;
        RECT 128.190 183.485 128.405 183.535 ;
        RECT 126.270 183.035 127.145 183.365 ;
        RECT 127.315 183.035 128.065 183.365 ;
        RECT 126.270 182.575 126.440 183.035 ;
        RECT 127.315 182.865 127.515 183.035 ;
        RECT 128.235 182.905 128.405 183.485 ;
        RECT 128.180 182.865 128.405 182.905 ;
        RECT 125.080 182.405 125.485 182.575 ;
        RECT 125.655 182.405 126.440 182.575 ;
        RECT 126.715 182.125 126.925 182.655 ;
        RECT 127.185 182.340 127.515 182.865 ;
        RECT 128.025 182.780 128.405 182.865 ;
        RECT 127.685 182.125 127.855 182.735 ;
        RECT 128.025 182.345 128.355 182.780 ;
        RECT 128.585 182.305 128.845 184.495 ;
        RECT 129.015 183.945 129.355 184.675 ;
        RECT 129.535 183.765 129.805 184.495 ;
        RECT 129.035 183.545 129.805 183.765 ;
        RECT 129.985 183.785 130.215 184.495 ;
        RECT 130.385 183.965 130.715 184.675 ;
        RECT 130.885 183.785 131.145 184.495 ;
        RECT 129.985 183.545 131.145 183.785 ;
        RECT 129.035 182.875 129.325 183.545 ;
        RECT 131.800 183.535 132.055 184.675 ;
        RECT 132.250 184.125 133.445 184.455 ;
        RECT 132.305 183.365 132.475 183.925 ;
        RECT 132.700 183.705 133.120 183.955 ;
        RECT 133.625 183.875 133.905 184.675 ;
        RECT 132.700 183.535 133.945 183.705 ;
        RECT 134.115 183.535 134.385 184.505 ;
        RECT 135.020 183.535 135.275 184.675 ;
        RECT 135.470 184.125 136.665 184.455 ;
        RECT 133.775 183.365 133.945 183.535 ;
        RECT 129.505 183.055 129.970 183.365 ;
        RECT 130.150 183.055 130.675 183.365 ;
        RECT 129.035 182.675 130.265 182.875 ;
        RECT 129.105 182.125 129.775 182.495 ;
        RECT 129.955 182.305 130.265 182.675 ;
        RECT 130.445 182.415 130.675 183.055 ;
        RECT 130.855 183.035 131.155 183.365 ;
        RECT 131.800 183.115 132.135 183.365 ;
        RECT 132.305 183.035 133.045 183.365 ;
        RECT 133.775 183.035 134.005 183.365 ;
        RECT 132.305 182.945 132.555 183.035 ;
        RECT 130.855 182.125 131.145 182.855 ;
        RECT 131.820 182.775 132.555 182.945 ;
        RECT 133.775 182.865 133.945 183.035 ;
        RECT 131.820 182.305 132.130 182.775 ;
        RECT 133.205 182.695 133.945 182.865 ;
        RECT 134.215 182.800 134.385 183.535 ;
        RECT 135.525 183.365 135.695 183.925 ;
        RECT 135.920 183.705 136.340 183.955 ;
        RECT 136.845 183.875 137.125 184.675 ;
        RECT 135.920 183.535 137.165 183.705 ;
        RECT 137.335 183.535 137.605 184.505 ;
        RECT 136.995 183.365 137.165 183.535 ;
        RECT 135.020 183.115 135.355 183.365 ;
        RECT 135.525 183.035 136.265 183.365 ;
        RECT 136.995 183.035 137.225 183.365 ;
        RECT 135.525 182.945 135.775 183.035 ;
        RECT 132.300 182.125 133.035 182.605 ;
        RECT 133.205 182.345 133.375 182.695 ;
        RECT 133.545 182.125 133.925 182.525 ;
        RECT 134.115 182.455 134.385 182.800 ;
        RECT 135.040 182.775 135.775 182.945 ;
        RECT 136.995 182.865 137.165 183.035 ;
        RECT 135.040 182.305 135.350 182.775 ;
        RECT 136.425 182.695 137.165 182.865 ;
        RECT 137.435 182.800 137.605 183.535 ;
        RECT 138.695 183.510 138.985 184.675 ;
        RECT 139.155 183.535 139.435 184.675 ;
        RECT 139.605 183.525 139.935 184.505 ;
        RECT 140.105 183.535 140.365 184.675 ;
        RECT 141.000 183.525 141.260 184.675 ;
        RECT 141.435 183.600 141.690 184.505 ;
        RECT 141.860 183.915 142.190 184.675 ;
        RECT 142.405 183.745 142.575 184.505 ;
        RECT 139.165 183.095 139.500 183.365 ;
        RECT 139.670 182.925 139.840 183.525 ;
        RECT 140.010 183.115 140.345 183.365 ;
        RECT 135.520 182.125 136.255 182.605 ;
        RECT 136.425 182.345 136.595 182.695 ;
        RECT 136.765 182.125 137.145 182.525 ;
        RECT 137.335 182.455 137.605 182.800 ;
        RECT 138.695 182.125 138.985 182.850 ;
        RECT 139.155 182.125 139.465 182.925 ;
        RECT 139.670 182.295 140.365 182.925 ;
        RECT 141.000 182.125 141.260 182.965 ;
        RECT 141.435 182.870 141.605 183.600 ;
        RECT 141.860 183.575 142.575 183.745 ;
        RECT 142.870 183.885 143.405 184.505 ;
        RECT 141.860 183.365 142.030 183.575 ;
        RECT 141.775 183.035 142.030 183.365 ;
        RECT 141.435 182.295 141.690 182.870 ;
        RECT 141.860 182.845 142.030 183.035 ;
        RECT 142.310 183.025 142.665 183.395 ;
        RECT 142.870 182.865 143.185 183.885 ;
        RECT 143.575 183.875 143.905 184.675 ;
        RECT 145.135 184.165 145.395 184.675 ;
        RECT 144.390 183.705 144.780 183.880 ;
        RECT 143.355 183.535 144.780 183.705 ;
        RECT 143.355 183.035 143.525 183.535 ;
        RECT 141.860 182.675 142.575 182.845 ;
        RECT 141.860 182.125 142.190 182.505 ;
        RECT 142.405 182.295 142.575 182.675 ;
        RECT 142.870 182.295 143.485 182.865 ;
        RECT 143.775 182.805 144.040 183.365 ;
        RECT 144.210 182.635 144.380 183.535 ;
        RECT 144.550 182.805 144.905 183.365 ;
        RECT 145.135 183.115 145.475 183.995 ;
        RECT 145.645 183.285 145.815 184.505 ;
        RECT 146.055 184.170 146.670 184.675 ;
        RECT 146.055 183.635 146.305 184.000 ;
        RECT 146.475 183.995 146.670 184.170 ;
        RECT 146.840 184.165 147.315 184.505 ;
        RECT 147.485 184.130 147.700 184.675 ;
        RECT 146.475 183.805 146.805 183.995 ;
        RECT 147.025 183.635 147.740 183.930 ;
        RECT 147.910 183.805 148.185 184.505 ;
        RECT 146.055 183.465 147.845 183.635 ;
        RECT 145.645 183.035 146.440 183.285 ;
        RECT 145.645 182.945 145.895 183.035 ;
        RECT 143.655 182.125 143.870 182.635 ;
        RECT 144.100 182.305 144.380 182.635 ;
        RECT 144.560 182.125 144.800 182.635 ;
        RECT 145.135 182.125 145.395 182.945 ;
        RECT 145.565 182.525 145.895 182.945 ;
        RECT 146.610 182.610 146.865 183.465 ;
        RECT 146.075 182.345 146.865 182.610 ;
        RECT 147.035 182.765 147.445 183.285 ;
        RECT 147.615 183.035 147.845 183.465 ;
        RECT 148.015 182.775 148.185 183.805 ;
        RECT 148.415 183.615 148.745 184.460 ;
        RECT 148.915 183.665 149.085 184.675 ;
        RECT 149.255 183.945 149.595 184.505 ;
        RECT 149.825 184.175 150.140 184.675 ;
        RECT 150.320 184.205 151.205 184.375 ;
        RECT 148.355 183.535 148.745 183.615 ;
        RECT 149.255 183.570 150.150 183.945 ;
        RECT 148.355 183.485 148.570 183.535 ;
        RECT 148.355 182.905 148.525 183.485 ;
        RECT 149.255 183.365 149.445 183.570 ;
        RECT 150.320 183.365 150.490 184.205 ;
        RECT 151.430 184.175 151.680 184.505 ;
        RECT 148.695 183.035 149.445 183.365 ;
        RECT 149.615 183.035 150.490 183.365 ;
        RECT 148.355 182.865 148.580 182.905 ;
        RECT 149.245 182.865 149.445 183.035 ;
        RECT 148.355 182.780 148.735 182.865 ;
        RECT 147.035 182.345 147.235 182.765 ;
        RECT 147.425 182.125 147.755 182.585 ;
        RECT 147.925 182.295 148.185 182.775 ;
        RECT 148.405 182.345 148.735 182.780 ;
        RECT 148.905 182.125 149.075 182.735 ;
        RECT 149.245 182.340 149.575 182.865 ;
        RECT 149.835 182.125 150.045 182.655 ;
        RECT 150.320 182.575 150.490 183.035 ;
        RECT 150.660 183.075 150.980 184.035 ;
        RECT 151.150 183.285 151.340 184.005 ;
        RECT 151.510 183.105 151.680 184.175 ;
        RECT 151.850 183.875 152.020 184.675 ;
        RECT 152.190 184.230 153.295 184.400 ;
        RECT 152.190 183.615 152.360 184.230 ;
        RECT 153.505 184.080 153.755 184.505 ;
        RECT 153.925 184.215 154.190 184.675 ;
        RECT 152.530 183.695 153.060 184.060 ;
        RECT 153.505 183.950 153.810 184.080 ;
        RECT 151.850 183.525 152.360 183.615 ;
        RECT 151.850 183.355 152.720 183.525 ;
        RECT 151.850 183.285 152.020 183.355 ;
        RECT 152.140 183.105 152.340 183.135 ;
        RECT 150.660 182.745 151.125 183.075 ;
        RECT 151.510 182.805 152.340 183.105 ;
        RECT 151.510 182.575 151.680 182.805 ;
        RECT 150.320 182.405 151.105 182.575 ;
        RECT 151.275 182.405 151.680 182.575 ;
        RECT 151.860 182.125 152.230 182.625 ;
        RECT 152.550 182.575 152.720 183.355 ;
        RECT 152.890 182.995 153.060 183.695 ;
        RECT 153.230 183.165 153.470 183.760 ;
        RECT 152.890 182.775 153.415 182.995 ;
        RECT 153.640 182.845 153.810 183.950 ;
        RECT 153.585 182.715 153.810 182.845 ;
        RECT 153.980 182.755 154.260 183.705 ;
        RECT 153.585 182.575 153.755 182.715 ;
        RECT 152.550 182.405 153.225 182.575 ;
        RECT 153.420 182.405 153.755 182.575 ;
        RECT 153.925 182.125 154.175 182.585 ;
        RECT 154.430 182.385 154.615 184.505 ;
        RECT 154.785 184.175 155.115 184.675 ;
        RECT 155.285 184.005 155.455 184.505 ;
        RECT 154.790 183.835 155.455 184.005 ;
        RECT 154.790 182.845 155.020 183.835 ;
        RECT 155.190 183.015 155.540 183.665 ;
        RECT 155.715 183.585 156.925 184.675 ;
        RECT 155.715 183.045 156.235 183.585 ;
        RECT 156.405 182.875 156.925 183.415 ;
        RECT 154.790 182.675 155.455 182.845 ;
        RECT 154.785 182.125 155.115 182.505 ;
        RECT 155.285 182.385 155.455 182.675 ;
        RECT 155.715 182.125 156.925 182.875 ;
        RECT 22.690 181.955 157.010 182.125 ;
        RECT 22.775 181.205 23.985 181.955 ;
        RECT 25.075 181.280 25.335 181.785 ;
        RECT 25.515 181.575 25.845 181.955 ;
        RECT 26.025 181.405 26.195 181.785 ;
        RECT 22.775 180.665 23.295 181.205 ;
        RECT 23.465 180.495 23.985 181.035 ;
        RECT 22.775 179.405 23.985 180.495 ;
        RECT 25.075 180.480 25.245 181.280 ;
        RECT 25.530 181.235 26.195 181.405 ;
        RECT 25.530 180.980 25.700 181.235 ;
        RECT 26.455 181.185 29.965 181.955 ;
        RECT 31.220 181.445 31.460 181.955 ;
        RECT 31.640 181.445 31.920 181.775 ;
        RECT 32.150 181.445 32.365 181.955 ;
        RECT 25.415 180.650 25.700 180.980 ;
        RECT 25.935 180.685 26.265 181.055 ;
        RECT 26.455 180.665 28.105 181.185 ;
        RECT 25.530 180.505 25.700 180.650 ;
        RECT 25.075 179.575 25.345 180.480 ;
        RECT 25.530 180.335 26.195 180.505 ;
        RECT 28.275 180.495 29.965 181.015 ;
        RECT 31.115 180.715 31.470 181.275 ;
        RECT 31.640 180.545 31.810 181.445 ;
        RECT 31.980 180.715 32.245 181.275 ;
        RECT 32.535 181.215 33.150 181.785 ;
        RECT 32.495 180.545 32.665 181.045 ;
        RECT 25.515 179.405 25.845 180.165 ;
        RECT 26.025 179.575 26.195 180.335 ;
        RECT 26.455 179.405 29.965 180.495 ;
        RECT 31.240 180.375 32.665 180.545 ;
        RECT 31.240 180.200 31.630 180.375 ;
        RECT 32.115 179.405 32.445 180.205 ;
        RECT 32.835 180.195 33.150 181.215 ;
        RECT 33.355 181.185 35.945 181.955 ;
        RECT 33.355 180.665 34.565 181.185 ;
        RECT 36.115 181.135 36.375 181.955 ;
        RECT 36.545 181.135 36.875 181.555 ;
        RECT 37.055 181.470 37.845 181.735 ;
        RECT 36.625 181.045 36.875 181.135 ;
        RECT 34.735 180.495 35.945 181.015 ;
        RECT 32.615 179.575 33.150 180.195 ;
        RECT 33.355 179.405 35.945 180.495 ;
        RECT 36.115 180.085 36.455 180.965 ;
        RECT 36.625 180.795 37.420 181.045 ;
        RECT 36.115 179.405 36.375 179.915 ;
        RECT 36.625 179.575 36.795 180.795 ;
        RECT 37.590 180.615 37.845 181.470 ;
        RECT 38.015 181.315 38.215 181.735 ;
        RECT 38.405 181.495 38.735 181.955 ;
        RECT 38.015 180.795 38.425 181.315 ;
        RECT 38.905 181.305 39.165 181.785 ;
        RECT 38.595 180.615 38.825 181.045 ;
        RECT 37.035 180.445 38.825 180.615 ;
        RECT 37.035 180.080 37.285 180.445 ;
        RECT 37.455 180.085 37.785 180.275 ;
        RECT 38.005 180.150 38.720 180.445 ;
        RECT 38.995 180.275 39.165 181.305 ;
        RECT 39.335 181.185 41.925 181.955 ;
        RECT 39.335 180.665 40.545 181.185 ;
        RECT 42.760 181.175 43.260 181.785 ;
        RECT 40.715 180.495 41.925 181.015 ;
        RECT 42.555 180.715 42.905 180.965 ;
        RECT 43.090 180.545 43.260 181.175 ;
        RECT 43.890 181.305 44.220 181.785 ;
        RECT 44.390 181.495 44.615 181.955 ;
        RECT 44.785 181.305 45.115 181.785 ;
        RECT 43.890 181.135 45.115 181.305 ;
        RECT 45.305 181.155 45.555 181.955 ;
        RECT 45.725 181.155 46.065 181.785 ;
        RECT 43.430 180.765 43.760 180.965 ;
        RECT 43.930 180.765 44.260 180.965 ;
        RECT 44.430 180.765 44.850 180.965 ;
        RECT 45.025 180.795 45.720 180.965 ;
        RECT 45.025 180.545 45.195 180.795 ;
        RECT 45.890 180.545 46.065 181.155 ;
        RECT 46.235 181.185 47.905 181.955 ;
        RECT 48.535 181.230 48.825 181.955 ;
        RECT 48.995 181.185 52.505 181.955 ;
        RECT 52.675 181.205 53.885 181.955 ;
        RECT 46.235 180.665 46.985 181.185 ;
        RECT 37.455 179.910 37.650 180.085 ;
        RECT 37.035 179.405 37.650 179.910 ;
        RECT 37.820 179.575 38.295 179.915 ;
        RECT 38.465 179.405 38.680 179.950 ;
        RECT 38.890 179.575 39.165 180.275 ;
        RECT 39.335 179.405 41.925 180.495 ;
        RECT 42.760 180.375 45.195 180.545 ;
        RECT 42.760 179.575 43.090 180.375 ;
        RECT 43.260 179.405 43.590 180.205 ;
        RECT 43.890 179.575 44.220 180.375 ;
        RECT 44.865 179.405 45.115 180.205 ;
        RECT 45.385 179.405 45.555 180.545 ;
        RECT 45.725 179.575 46.065 180.545 ;
        RECT 47.155 180.495 47.905 181.015 ;
        RECT 48.995 180.665 50.645 181.185 ;
        RECT 46.235 179.405 47.905 180.495 ;
        RECT 48.535 179.405 48.825 180.570 ;
        RECT 50.815 180.495 52.505 181.015 ;
        RECT 52.675 180.665 53.195 181.205 ;
        RECT 54.115 181.135 54.325 181.955 ;
        RECT 54.495 181.155 54.825 181.785 ;
        RECT 53.365 180.495 53.885 181.035 ;
        RECT 54.495 180.555 54.745 181.155 ;
        RECT 54.995 181.135 55.225 181.955 ;
        RECT 55.435 181.185 58.945 181.955 ;
        RECT 59.665 181.405 59.835 181.695 ;
        RECT 60.005 181.575 60.335 181.955 ;
        RECT 59.665 181.235 60.330 181.405 ;
        RECT 54.915 180.715 55.245 180.965 ;
        RECT 55.435 180.665 57.085 181.185 ;
        RECT 48.995 179.405 52.505 180.495 ;
        RECT 52.675 179.405 53.885 180.495 ;
        RECT 54.115 179.405 54.325 180.545 ;
        RECT 54.495 179.575 54.825 180.555 ;
        RECT 54.995 179.405 55.225 180.545 ;
        RECT 57.255 180.495 58.945 181.015 ;
        RECT 55.435 179.405 58.945 180.495 ;
        RECT 59.580 180.415 59.930 181.065 ;
        RECT 60.100 180.245 60.330 181.235 ;
        RECT 59.665 180.075 60.330 180.245 ;
        RECT 59.665 179.575 59.835 180.075 ;
        RECT 60.005 179.405 60.335 179.905 ;
        RECT 60.505 179.575 60.690 181.695 ;
        RECT 60.945 181.495 61.195 181.955 ;
        RECT 61.365 181.505 61.700 181.675 ;
        RECT 61.895 181.505 62.570 181.675 ;
        RECT 61.365 181.365 61.535 181.505 ;
        RECT 60.860 180.375 61.140 181.325 ;
        RECT 61.310 181.235 61.535 181.365 ;
        RECT 61.310 180.130 61.480 181.235 ;
        RECT 61.705 181.085 62.230 181.305 ;
        RECT 61.650 180.320 61.890 180.915 ;
        RECT 62.060 180.385 62.230 181.085 ;
        RECT 62.400 180.725 62.570 181.505 ;
        RECT 62.890 181.455 63.260 181.955 ;
        RECT 63.440 181.505 63.845 181.675 ;
        RECT 64.015 181.505 64.800 181.675 ;
        RECT 63.440 181.275 63.610 181.505 ;
        RECT 62.780 180.975 63.610 181.275 ;
        RECT 63.995 181.005 64.460 181.335 ;
        RECT 62.780 180.945 62.980 180.975 ;
        RECT 63.100 180.725 63.270 180.795 ;
        RECT 62.400 180.555 63.270 180.725 ;
        RECT 62.760 180.465 63.270 180.555 ;
        RECT 61.310 180.000 61.615 180.130 ;
        RECT 62.060 180.020 62.590 180.385 ;
        RECT 60.930 179.405 61.195 179.865 ;
        RECT 61.365 179.575 61.615 180.000 ;
        RECT 62.760 179.850 62.930 180.465 ;
        RECT 61.825 179.680 62.930 179.850 ;
        RECT 63.100 179.405 63.270 180.205 ;
        RECT 63.440 179.905 63.610 180.975 ;
        RECT 63.780 180.075 63.970 180.795 ;
        RECT 64.140 180.045 64.460 181.005 ;
        RECT 64.630 181.045 64.800 181.505 ;
        RECT 65.075 181.425 65.285 181.955 ;
        RECT 65.545 181.215 65.875 181.740 ;
        RECT 66.045 181.345 66.215 181.955 ;
        RECT 66.385 181.300 66.715 181.735 ;
        RECT 66.385 181.215 66.765 181.300 ;
        RECT 65.675 181.045 65.875 181.215 ;
        RECT 66.540 181.175 66.765 181.215 ;
        RECT 64.630 180.715 65.505 181.045 ;
        RECT 65.675 180.715 66.425 181.045 ;
        RECT 63.440 179.575 63.690 179.905 ;
        RECT 64.630 179.875 64.800 180.715 ;
        RECT 65.675 180.510 65.865 180.715 ;
        RECT 66.595 180.595 66.765 181.175 ;
        RECT 66.550 180.545 66.765 180.595 ;
        RECT 64.970 180.135 65.865 180.510 ;
        RECT 66.375 180.465 66.765 180.545 ;
        RECT 66.935 181.215 67.320 181.785 ;
        RECT 67.490 181.495 67.815 181.955 ;
        RECT 68.335 181.325 68.615 181.785 ;
        RECT 66.935 180.545 67.215 181.215 ;
        RECT 67.490 181.155 68.615 181.325 ;
        RECT 67.490 181.045 67.940 181.155 ;
        RECT 67.385 180.715 67.940 181.045 ;
        RECT 68.805 180.985 69.205 181.785 ;
        RECT 69.605 181.495 69.875 181.955 ;
        RECT 70.045 181.325 70.330 181.785 ;
        RECT 63.915 179.705 64.800 179.875 ;
        RECT 64.980 179.405 65.295 179.905 ;
        RECT 65.525 179.575 65.865 180.135 ;
        RECT 66.035 179.405 66.205 180.415 ;
        RECT 66.375 179.620 66.705 180.465 ;
        RECT 66.935 179.575 67.320 180.545 ;
        RECT 67.490 180.255 67.940 180.715 ;
        RECT 68.110 180.425 69.205 180.985 ;
        RECT 67.490 180.035 68.615 180.255 ;
        RECT 67.490 179.405 67.815 179.865 ;
        RECT 68.335 179.575 68.615 180.035 ;
        RECT 68.805 179.575 69.205 180.425 ;
        RECT 69.375 181.155 70.330 181.325 ;
        RECT 70.615 181.185 74.125 181.955 ;
        RECT 74.295 181.230 74.585 181.955 ;
        RECT 74.755 181.185 78.265 181.955 ;
        RECT 78.895 181.455 79.155 181.785 ;
        RECT 79.325 181.595 79.655 181.955 ;
        RECT 79.910 181.575 81.210 181.785 ;
        RECT 78.895 181.445 79.125 181.455 ;
        RECT 69.375 180.255 69.585 181.155 ;
        RECT 69.755 180.425 70.445 180.985 ;
        RECT 70.615 180.665 72.265 181.185 ;
        RECT 72.435 180.495 74.125 181.015 ;
        RECT 74.755 180.665 76.405 181.185 ;
        RECT 69.375 180.035 70.330 180.255 ;
        RECT 69.605 179.405 69.875 179.865 ;
        RECT 70.045 179.575 70.330 180.035 ;
        RECT 70.615 179.405 74.125 180.495 ;
        RECT 74.295 179.405 74.585 180.570 ;
        RECT 76.575 180.495 78.265 181.015 ;
        RECT 74.755 179.405 78.265 180.495 ;
        RECT 78.895 180.255 79.065 181.445 ;
        RECT 79.910 181.425 80.080 181.575 ;
        RECT 79.325 181.300 80.080 181.425 ;
        RECT 79.235 181.255 80.080 181.300 ;
        RECT 79.235 181.135 79.505 181.255 ;
        RECT 79.235 180.560 79.405 181.135 ;
        RECT 79.635 180.695 80.045 181.000 ;
        RECT 80.335 180.965 80.545 181.365 ;
        RECT 80.215 180.755 80.545 180.965 ;
        RECT 80.790 180.965 81.010 181.365 ;
        RECT 81.485 181.190 81.940 181.955 ;
        RECT 82.115 181.185 85.625 181.955 ;
        RECT 85.820 181.305 86.130 181.775 ;
        RECT 86.300 181.475 87.035 181.955 ;
        RECT 87.205 181.385 87.375 181.735 ;
        RECT 87.545 181.555 87.925 181.955 ;
        RECT 80.790 180.755 81.265 180.965 ;
        RECT 81.455 180.765 81.945 180.965 ;
        RECT 82.115 180.665 83.765 181.185 ;
        RECT 85.820 181.135 86.555 181.305 ;
        RECT 87.205 181.215 87.945 181.385 ;
        RECT 88.115 181.280 88.385 181.625 ;
        RECT 88.640 181.455 89.135 181.785 ;
        RECT 86.305 181.045 86.555 181.135 ;
        RECT 87.775 181.045 87.945 181.215 ;
        RECT 79.235 180.525 79.435 180.560 ;
        RECT 80.765 180.525 81.940 180.585 ;
        RECT 79.235 180.415 81.940 180.525 ;
        RECT 83.935 180.495 85.625 181.015 ;
        RECT 85.800 180.715 86.135 180.965 ;
        RECT 86.305 180.715 87.045 181.045 ;
        RECT 87.775 180.715 88.005 181.045 ;
        RECT 79.295 180.355 81.095 180.415 ;
        RECT 80.765 180.325 81.095 180.355 ;
        RECT 78.895 179.575 79.155 180.255 ;
        RECT 79.325 179.405 79.575 180.185 ;
        RECT 79.825 180.155 80.660 180.165 ;
        RECT 81.250 180.155 81.435 180.245 ;
        RECT 79.825 179.955 81.435 180.155 ;
        RECT 79.825 179.575 80.075 179.955 ;
        RECT 81.205 179.915 81.435 179.955 ;
        RECT 81.685 179.795 81.940 180.415 ;
        RECT 80.245 179.405 80.600 179.785 ;
        RECT 81.605 179.575 81.940 179.795 ;
        RECT 82.115 179.405 85.625 180.495 ;
        RECT 85.800 179.405 86.055 180.545 ;
        RECT 86.305 180.155 86.475 180.715 ;
        RECT 87.775 180.545 87.945 180.715 ;
        RECT 88.215 180.545 88.385 181.280 ;
        RECT 86.700 180.375 87.945 180.545 ;
        RECT 86.700 180.125 87.120 180.375 ;
        RECT 86.250 179.625 87.445 179.955 ;
        RECT 87.625 179.405 87.905 180.205 ;
        RECT 88.115 179.575 88.385 180.545 ;
        RECT 88.555 179.965 88.795 181.275 ;
        RECT 88.965 180.545 89.135 181.455 ;
        RECT 89.355 180.715 89.705 181.680 ;
        RECT 89.885 180.715 90.185 181.685 ;
        RECT 90.365 180.715 90.645 181.685 ;
        RECT 90.825 181.155 91.095 181.955 ;
        RECT 91.265 181.235 91.605 181.745 ;
        RECT 90.840 180.715 91.170 180.965 ;
        RECT 90.840 180.545 91.155 180.715 ;
        RECT 88.965 180.375 91.155 180.545 ;
        RECT 88.560 179.405 88.895 179.785 ;
        RECT 89.065 179.575 89.315 180.375 ;
        RECT 89.535 179.405 89.865 180.125 ;
        RECT 90.050 179.575 90.300 180.375 ;
        RECT 90.765 179.405 91.095 180.205 ;
        RECT 91.345 179.835 91.605 181.235 ;
        RECT 92.695 181.135 92.955 181.955 ;
        RECT 93.125 181.135 93.455 181.555 ;
        RECT 93.635 181.470 94.425 181.735 ;
        RECT 93.205 181.045 93.455 181.135 ;
        RECT 92.695 180.085 93.035 180.965 ;
        RECT 93.205 180.795 94.000 181.045 ;
        RECT 91.265 179.575 91.605 179.835 ;
        RECT 92.695 179.405 92.955 179.915 ;
        RECT 93.205 179.575 93.375 180.795 ;
        RECT 94.170 180.615 94.425 181.470 ;
        RECT 94.595 181.315 94.795 181.735 ;
        RECT 94.985 181.495 95.315 181.955 ;
        RECT 94.595 180.795 95.005 181.315 ;
        RECT 95.485 181.305 95.745 181.785 ;
        RECT 96.835 181.575 97.725 181.745 ;
        RECT 95.175 180.615 95.405 181.045 ;
        RECT 93.615 180.445 95.405 180.615 ;
        RECT 93.615 180.080 93.865 180.445 ;
        RECT 94.035 180.085 94.365 180.275 ;
        RECT 94.585 180.150 95.300 180.445 ;
        RECT 95.575 180.275 95.745 181.305 ;
        RECT 96.835 181.020 97.385 181.405 ;
        RECT 97.555 180.850 97.725 181.575 ;
        RECT 94.035 179.910 94.230 180.085 ;
        RECT 93.615 179.405 94.230 179.910 ;
        RECT 94.400 179.575 94.875 179.915 ;
        RECT 95.045 179.405 95.260 179.950 ;
        RECT 95.470 179.575 95.745 180.275 ;
        RECT 96.835 180.780 97.725 180.850 ;
        RECT 97.895 181.250 98.115 181.735 ;
        RECT 98.285 181.415 98.535 181.955 ;
        RECT 98.705 181.305 98.965 181.785 ;
        RECT 97.895 180.825 98.225 181.250 ;
        RECT 96.835 180.755 97.730 180.780 ;
        RECT 96.835 180.740 97.740 180.755 ;
        RECT 96.835 180.725 97.745 180.740 ;
        RECT 96.835 180.720 97.755 180.725 ;
        RECT 96.835 180.710 97.760 180.720 ;
        RECT 96.835 180.700 97.765 180.710 ;
        RECT 96.835 180.695 97.775 180.700 ;
        RECT 96.835 180.685 97.785 180.695 ;
        RECT 96.835 180.680 97.795 180.685 ;
        RECT 96.835 180.230 97.095 180.680 ;
        RECT 97.460 180.675 97.795 180.680 ;
        RECT 97.460 180.670 97.810 180.675 ;
        RECT 97.460 180.660 97.825 180.670 ;
        RECT 97.460 180.655 97.850 180.660 ;
        RECT 98.395 180.655 98.625 181.050 ;
        RECT 97.460 180.650 98.625 180.655 ;
        RECT 97.490 180.615 98.625 180.650 ;
        RECT 97.525 180.590 98.625 180.615 ;
        RECT 97.555 180.560 98.625 180.590 ;
        RECT 97.575 180.530 98.625 180.560 ;
        RECT 97.595 180.500 98.625 180.530 ;
        RECT 97.665 180.490 98.625 180.500 ;
        RECT 97.690 180.480 98.625 180.490 ;
        RECT 97.710 180.465 98.625 180.480 ;
        RECT 97.730 180.450 98.625 180.465 ;
        RECT 97.735 180.440 98.520 180.450 ;
        RECT 97.750 180.405 98.520 180.440 ;
        RECT 97.265 180.085 97.595 180.330 ;
        RECT 97.765 180.155 98.520 180.405 ;
        RECT 98.795 180.275 98.965 181.305 ;
        RECT 100.055 181.230 100.345 181.955 ;
        RECT 100.515 181.185 103.105 181.955 ;
        RECT 100.515 180.665 101.725 181.185 ;
        RECT 103.295 181.145 103.535 181.955 ;
        RECT 103.705 181.145 104.035 181.785 ;
        RECT 104.205 181.145 104.475 181.955 ;
        RECT 104.655 181.185 108.165 181.955 ;
        RECT 108.335 181.205 109.545 181.955 ;
        RECT 109.995 181.325 110.375 181.775 ;
        RECT 97.265 180.060 97.450 180.085 ;
        RECT 96.835 179.960 97.450 180.060 ;
        RECT 96.835 179.405 97.440 179.960 ;
        RECT 97.615 179.575 98.095 179.915 ;
        RECT 98.265 179.405 98.520 179.950 ;
        RECT 98.690 179.575 98.965 180.275 ;
        RECT 100.055 179.405 100.345 180.570 ;
        RECT 101.895 180.495 103.105 181.015 ;
        RECT 103.275 180.715 103.625 180.965 ;
        RECT 103.795 180.545 103.965 181.145 ;
        RECT 104.135 180.715 104.485 180.965 ;
        RECT 104.655 180.665 106.305 181.185 ;
        RECT 100.515 179.405 103.105 180.495 ;
        RECT 103.285 180.375 103.965 180.545 ;
        RECT 103.285 179.590 103.615 180.375 ;
        RECT 104.145 179.405 104.475 180.545 ;
        RECT 106.475 180.495 108.165 181.015 ;
        RECT 108.335 180.665 108.855 181.205 ;
        RECT 109.025 180.495 109.545 181.035 ;
        RECT 104.655 179.405 108.165 180.495 ;
        RECT 108.335 179.405 109.545 180.495 ;
        RECT 109.735 180.375 109.965 181.065 ;
        RECT 110.145 180.875 110.375 181.325 ;
        RECT 110.555 181.175 110.785 181.955 ;
        RECT 110.965 181.245 111.395 181.775 ;
        RECT 110.965 180.995 111.210 181.245 ;
        RECT 111.575 181.045 111.785 181.665 ;
        RECT 111.955 181.225 112.285 181.955 ;
        RECT 112.475 181.185 115.065 181.955 ;
        RECT 110.145 180.195 110.485 180.875 ;
        RECT 109.725 179.995 110.485 180.195 ;
        RECT 110.675 180.695 111.210 180.995 ;
        RECT 111.390 180.695 111.785 181.045 ;
        RECT 111.980 180.695 112.270 181.045 ;
        RECT 109.725 179.605 109.985 179.995 ;
        RECT 110.155 179.405 110.485 179.815 ;
        RECT 110.675 179.585 111.005 180.695 ;
        RECT 112.475 180.665 113.685 181.185 ;
        RECT 115.295 181.135 115.505 181.955 ;
        RECT 115.675 181.155 116.005 181.785 ;
        RECT 111.175 180.315 112.215 180.515 ;
        RECT 113.855 180.495 115.065 181.015 ;
        RECT 115.675 180.555 115.925 181.155 ;
        RECT 116.175 181.135 116.405 181.955 ;
        RECT 116.615 181.185 118.285 181.955 ;
        RECT 118.455 181.215 118.840 181.785 ;
        RECT 119.010 181.495 119.335 181.955 ;
        RECT 119.855 181.325 120.135 181.785 ;
        RECT 116.095 180.715 116.425 180.965 ;
        RECT 116.615 180.665 117.365 181.185 ;
        RECT 111.175 179.585 111.365 180.315 ;
        RECT 111.535 179.405 111.865 180.135 ;
        RECT 112.045 179.585 112.215 180.315 ;
        RECT 112.475 179.405 115.065 180.495 ;
        RECT 115.295 179.405 115.505 180.545 ;
        RECT 115.675 179.575 116.005 180.555 ;
        RECT 116.175 179.405 116.405 180.545 ;
        RECT 117.535 180.495 118.285 181.015 ;
        RECT 116.615 179.405 118.285 180.495 ;
        RECT 118.455 180.545 118.735 181.215 ;
        RECT 119.010 181.155 120.135 181.325 ;
        RECT 119.010 181.045 119.460 181.155 ;
        RECT 118.905 180.715 119.460 181.045 ;
        RECT 120.325 180.985 120.725 181.785 ;
        RECT 121.125 181.495 121.395 181.955 ;
        RECT 121.565 181.325 121.850 181.785 ;
        RECT 118.455 179.575 118.840 180.545 ;
        RECT 119.010 180.255 119.460 180.715 ;
        RECT 119.630 180.425 120.725 180.985 ;
        RECT 119.010 180.035 120.135 180.255 ;
        RECT 119.010 179.405 119.335 179.865 ;
        RECT 119.855 179.575 120.135 180.035 ;
        RECT 120.325 179.575 120.725 180.425 ;
        RECT 120.895 181.155 121.850 181.325 ;
        RECT 122.135 181.455 122.395 181.785 ;
        RECT 122.565 181.595 122.895 181.955 ;
        RECT 123.150 181.575 124.450 181.785 ;
        RECT 120.895 180.255 121.105 181.155 ;
        RECT 121.275 180.425 121.965 180.985 ;
        RECT 122.135 180.255 122.305 181.455 ;
        RECT 123.150 181.425 123.320 181.575 ;
        RECT 122.565 181.300 123.320 181.425 ;
        RECT 122.475 181.255 123.320 181.300 ;
        RECT 122.475 181.135 122.745 181.255 ;
        RECT 122.475 180.560 122.645 181.135 ;
        RECT 122.875 180.695 123.285 181.000 ;
        RECT 123.575 180.965 123.785 181.365 ;
        RECT 123.455 180.755 123.785 180.965 ;
        RECT 124.030 180.965 124.250 181.365 ;
        RECT 124.725 181.190 125.180 181.955 ;
        RECT 125.815 181.230 126.105 181.955 ;
        RECT 126.275 181.215 126.660 181.785 ;
        RECT 126.830 181.495 127.155 181.955 ;
        RECT 127.675 181.325 127.955 181.785 ;
        RECT 124.030 180.755 124.505 180.965 ;
        RECT 124.695 180.765 125.185 180.965 ;
        RECT 122.475 180.525 122.675 180.560 ;
        RECT 124.005 180.525 125.180 180.585 ;
        RECT 122.475 180.415 125.180 180.525 ;
        RECT 122.535 180.355 124.335 180.415 ;
        RECT 124.005 180.325 124.335 180.355 ;
        RECT 120.895 180.035 121.850 180.255 ;
        RECT 121.125 179.405 121.395 179.865 ;
        RECT 121.565 179.575 121.850 180.035 ;
        RECT 122.135 179.575 122.395 180.255 ;
        RECT 122.565 179.405 122.815 180.185 ;
        RECT 123.065 180.155 123.900 180.165 ;
        RECT 124.490 180.155 124.675 180.245 ;
        RECT 123.065 179.955 124.675 180.155 ;
        RECT 123.065 179.575 123.315 179.955 ;
        RECT 124.445 179.915 124.675 179.955 ;
        RECT 124.925 179.795 125.180 180.415 ;
        RECT 123.485 179.405 123.840 179.785 ;
        RECT 124.845 179.575 125.180 179.795 ;
        RECT 125.815 179.405 126.105 180.570 ;
        RECT 126.275 180.545 126.555 181.215 ;
        RECT 126.830 181.155 127.955 181.325 ;
        RECT 126.830 181.045 127.280 181.155 ;
        RECT 126.725 180.715 127.280 181.045 ;
        RECT 128.145 180.985 128.545 181.785 ;
        RECT 128.945 181.495 129.215 181.955 ;
        RECT 129.385 181.325 129.670 181.785 ;
        RECT 126.275 179.575 126.660 180.545 ;
        RECT 126.830 180.255 127.280 180.715 ;
        RECT 127.450 180.425 128.545 180.985 ;
        RECT 126.830 180.035 127.955 180.255 ;
        RECT 126.830 179.405 127.155 179.865 ;
        RECT 127.675 179.575 127.955 180.035 ;
        RECT 128.145 179.575 128.545 180.425 ;
        RECT 128.715 181.155 129.670 181.325 ;
        RECT 129.955 181.185 132.545 181.955 ;
        RECT 132.720 181.450 133.055 181.955 ;
        RECT 133.225 181.385 133.465 181.760 ;
        RECT 133.745 181.625 133.915 181.770 ;
        RECT 133.745 181.430 134.120 181.625 ;
        RECT 134.480 181.460 134.875 181.955 ;
        RECT 128.715 180.255 128.925 181.155 ;
        RECT 129.095 180.425 129.785 180.985 ;
        RECT 129.955 180.665 131.165 181.185 ;
        RECT 131.335 180.495 132.545 181.015 ;
        RECT 128.715 180.035 129.670 180.255 ;
        RECT 128.945 179.405 129.215 179.865 ;
        RECT 129.385 179.575 129.670 180.035 ;
        RECT 129.955 179.405 132.545 180.495 ;
        RECT 132.775 180.425 133.075 181.275 ;
        RECT 133.245 181.235 133.465 181.385 ;
        RECT 133.245 180.905 133.780 181.235 ;
        RECT 133.950 181.095 134.120 181.430 ;
        RECT 135.045 181.265 135.285 181.785 ;
        RECT 133.245 180.255 133.480 180.905 ;
        RECT 133.950 180.735 134.935 181.095 ;
        RECT 132.805 180.025 133.480 180.255 ;
        RECT 133.650 180.715 134.935 180.735 ;
        RECT 133.650 180.565 134.510 180.715 ;
        RECT 132.805 179.595 132.975 180.025 ;
        RECT 133.145 179.405 133.475 179.855 ;
        RECT 133.650 179.620 133.935 180.565 ;
        RECT 135.110 180.460 135.285 181.265 ;
        RECT 135.475 181.185 138.985 181.955 ;
        RECT 139.160 181.450 139.495 181.955 ;
        RECT 139.665 181.385 139.905 181.760 ;
        RECT 140.185 181.625 140.355 181.770 ;
        RECT 140.185 181.430 140.560 181.625 ;
        RECT 140.920 181.460 141.315 181.955 ;
        RECT 135.475 180.665 137.125 181.185 ;
        RECT 137.295 180.495 138.985 181.015 ;
        RECT 134.110 180.085 134.805 180.395 ;
        RECT 134.115 179.405 134.800 179.875 ;
        RECT 134.980 179.675 135.285 180.460 ;
        RECT 135.475 179.405 138.985 180.495 ;
        RECT 139.215 180.425 139.515 181.275 ;
        RECT 139.685 181.235 139.905 181.385 ;
        RECT 139.685 180.905 140.220 181.235 ;
        RECT 140.390 181.095 140.560 181.430 ;
        RECT 141.485 181.265 141.725 181.785 ;
        RECT 139.685 180.255 139.920 180.905 ;
        RECT 140.390 180.735 141.375 181.095 ;
        RECT 139.245 180.025 139.920 180.255 ;
        RECT 140.090 180.715 141.375 180.735 ;
        RECT 140.090 180.565 140.950 180.715 ;
        RECT 139.245 179.595 139.415 180.025 ;
        RECT 139.585 179.405 139.915 179.855 ;
        RECT 140.090 179.620 140.375 180.565 ;
        RECT 141.550 180.460 141.725 181.265 ;
        RECT 141.915 181.185 143.585 181.955 ;
        RECT 144.265 181.300 144.595 181.735 ;
        RECT 144.765 181.345 144.935 181.955 ;
        RECT 144.215 181.215 144.595 181.300 ;
        RECT 145.105 181.215 145.435 181.740 ;
        RECT 145.695 181.425 145.905 181.955 ;
        RECT 146.180 181.505 146.965 181.675 ;
        RECT 147.135 181.505 147.540 181.675 ;
        RECT 141.915 180.665 142.665 181.185 ;
        RECT 144.215 181.175 144.440 181.215 ;
        RECT 142.835 180.495 143.585 181.015 ;
        RECT 140.550 180.085 141.245 180.395 ;
        RECT 140.555 179.405 141.240 179.875 ;
        RECT 141.420 179.675 141.725 180.460 ;
        RECT 141.915 179.405 143.585 180.495 ;
        RECT 144.215 180.595 144.385 181.175 ;
        RECT 145.105 181.045 145.305 181.215 ;
        RECT 146.180 181.045 146.350 181.505 ;
        RECT 144.555 180.715 145.305 181.045 ;
        RECT 145.475 180.715 146.350 181.045 ;
        RECT 144.215 180.545 144.430 180.595 ;
        RECT 144.215 180.465 144.605 180.545 ;
        RECT 144.275 179.620 144.605 180.465 ;
        RECT 145.115 180.510 145.305 180.715 ;
        RECT 144.775 179.405 144.945 180.415 ;
        RECT 145.115 180.135 146.010 180.510 ;
        RECT 145.115 179.575 145.455 180.135 ;
        RECT 145.685 179.405 146.000 179.905 ;
        RECT 146.180 179.875 146.350 180.715 ;
        RECT 146.520 181.005 146.985 181.335 ;
        RECT 147.370 181.275 147.540 181.505 ;
        RECT 147.720 181.455 148.090 181.955 ;
        RECT 148.410 181.505 149.085 181.675 ;
        RECT 149.280 181.505 149.615 181.675 ;
        RECT 146.520 180.045 146.840 181.005 ;
        RECT 147.370 180.975 148.200 181.275 ;
        RECT 147.010 180.075 147.200 180.795 ;
        RECT 147.370 179.905 147.540 180.975 ;
        RECT 148.000 180.945 148.200 180.975 ;
        RECT 147.710 180.725 147.880 180.795 ;
        RECT 148.410 180.725 148.580 181.505 ;
        RECT 149.445 181.365 149.615 181.505 ;
        RECT 149.785 181.495 150.035 181.955 ;
        RECT 147.710 180.555 148.580 180.725 ;
        RECT 148.750 181.085 149.275 181.305 ;
        RECT 149.445 181.235 149.670 181.365 ;
        RECT 147.710 180.465 148.220 180.555 ;
        RECT 146.180 179.705 147.065 179.875 ;
        RECT 147.290 179.575 147.540 179.905 ;
        RECT 147.710 179.405 147.880 180.205 ;
        RECT 148.050 179.850 148.220 180.465 ;
        RECT 148.750 180.385 148.920 181.085 ;
        RECT 148.390 180.020 148.920 180.385 ;
        RECT 149.090 180.320 149.330 180.915 ;
        RECT 149.500 180.130 149.670 181.235 ;
        RECT 149.840 180.375 150.120 181.325 ;
        RECT 149.365 180.000 149.670 180.130 ;
        RECT 148.050 179.680 149.155 179.850 ;
        RECT 149.365 179.575 149.615 180.000 ;
        RECT 149.785 179.405 150.050 179.865 ;
        RECT 150.290 179.575 150.475 181.695 ;
        RECT 150.645 181.575 150.975 181.955 ;
        RECT 151.145 181.405 151.315 181.695 ;
        RECT 150.650 181.235 151.315 181.405 ;
        RECT 150.650 180.245 150.880 181.235 ;
        RECT 151.575 181.230 151.865 181.955 ;
        RECT 152.200 181.445 152.440 181.955 ;
        RECT 152.620 181.445 152.900 181.775 ;
        RECT 153.130 181.445 153.345 181.955 ;
        RECT 151.050 180.415 151.400 181.065 ;
        RECT 152.095 180.715 152.450 181.275 ;
        RECT 150.650 180.075 151.315 180.245 ;
        RECT 150.645 179.405 150.975 179.905 ;
        RECT 151.145 179.575 151.315 180.075 ;
        RECT 151.575 179.405 151.865 180.570 ;
        RECT 152.620 180.545 152.790 181.445 ;
        RECT 152.960 180.715 153.225 181.275 ;
        RECT 153.515 181.215 154.130 181.785 ;
        RECT 153.475 180.545 153.645 181.045 ;
        RECT 152.220 180.375 153.645 180.545 ;
        RECT 152.220 180.200 152.610 180.375 ;
        RECT 153.095 179.405 153.425 180.205 ;
        RECT 153.815 180.195 154.130 181.215 ;
        RECT 153.595 179.575 154.130 180.195 ;
        RECT 154.335 181.280 154.595 181.785 ;
        RECT 154.775 181.575 155.105 181.955 ;
        RECT 155.285 181.405 155.455 181.785 ;
        RECT 154.335 180.480 154.505 181.280 ;
        RECT 154.790 181.235 155.455 181.405 ;
        RECT 154.790 180.980 154.960 181.235 ;
        RECT 155.715 181.205 156.925 181.955 ;
        RECT 154.675 180.650 154.960 180.980 ;
        RECT 155.195 180.685 155.525 181.055 ;
        RECT 154.790 180.505 154.960 180.650 ;
        RECT 154.335 179.575 154.605 180.480 ;
        RECT 154.790 180.335 155.455 180.505 ;
        RECT 154.775 179.405 155.105 180.165 ;
        RECT 155.285 179.575 155.455 180.335 ;
        RECT 155.715 180.495 156.235 181.035 ;
        RECT 156.405 180.665 156.925 181.205 ;
        RECT 155.715 179.405 156.925 180.495 ;
        RECT 22.690 179.235 157.010 179.405 ;
        RECT 22.775 178.145 23.985 179.235 ;
        RECT 24.245 178.565 24.415 179.065 ;
        RECT 24.585 178.735 24.915 179.235 ;
        RECT 24.245 178.395 24.910 178.565 ;
        RECT 22.775 177.435 23.295 177.975 ;
        RECT 23.465 177.605 23.985 178.145 ;
        RECT 24.160 177.575 24.510 178.225 ;
        RECT 22.775 176.685 23.985 177.435 ;
        RECT 24.680 177.405 24.910 178.395 ;
        RECT 24.245 177.235 24.910 177.405 ;
        RECT 24.245 176.945 24.415 177.235 ;
        RECT 24.585 176.685 24.915 177.065 ;
        RECT 25.085 176.945 25.270 179.065 ;
        RECT 25.510 178.775 25.775 179.235 ;
        RECT 25.945 178.640 26.195 179.065 ;
        RECT 26.405 178.790 27.510 178.960 ;
        RECT 25.890 178.510 26.195 178.640 ;
        RECT 25.440 177.315 25.720 178.265 ;
        RECT 25.890 177.405 26.060 178.510 ;
        RECT 26.230 177.725 26.470 178.320 ;
        RECT 26.640 178.255 27.170 178.620 ;
        RECT 26.640 177.555 26.810 178.255 ;
        RECT 27.340 178.175 27.510 178.790 ;
        RECT 27.680 178.435 27.850 179.235 ;
        RECT 28.020 178.735 28.270 179.065 ;
        RECT 28.495 178.765 29.380 178.935 ;
        RECT 27.340 178.085 27.850 178.175 ;
        RECT 25.890 177.275 26.115 177.405 ;
        RECT 26.285 177.335 26.810 177.555 ;
        RECT 26.980 177.915 27.850 178.085 ;
        RECT 25.525 176.685 25.775 177.145 ;
        RECT 25.945 177.135 26.115 177.275 ;
        RECT 26.980 177.135 27.150 177.915 ;
        RECT 27.680 177.845 27.850 177.915 ;
        RECT 27.360 177.665 27.560 177.695 ;
        RECT 28.020 177.665 28.190 178.735 ;
        RECT 28.360 177.845 28.550 178.565 ;
        RECT 27.360 177.365 28.190 177.665 ;
        RECT 28.720 177.635 29.040 178.595 ;
        RECT 25.945 176.965 26.280 177.135 ;
        RECT 26.475 176.965 27.150 177.135 ;
        RECT 27.470 176.685 27.840 177.185 ;
        RECT 28.020 177.135 28.190 177.365 ;
        RECT 28.575 177.305 29.040 177.635 ;
        RECT 29.210 177.925 29.380 178.765 ;
        RECT 29.560 178.735 29.875 179.235 ;
        RECT 30.105 178.505 30.445 179.065 ;
        RECT 29.550 178.130 30.445 178.505 ;
        RECT 30.615 178.225 30.785 179.235 ;
        RECT 30.255 177.925 30.445 178.130 ;
        RECT 30.955 178.175 31.285 179.020 ;
        RECT 31.515 178.365 31.790 179.065 ;
        RECT 32.000 178.690 32.215 179.235 ;
        RECT 32.385 178.725 32.860 179.065 ;
        RECT 33.030 178.730 33.645 179.235 ;
        RECT 33.030 178.555 33.225 178.730 ;
        RECT 30.955 178.095 31.345 178.175 ;
        RECT 31.130 178.045 31.345 178.095 ;
        RECT 29.210 177.595 30.085 177.925 ;
        RECT 30.255 177.595 31.005 177.925 ;
        RECT 29.210 177.135 29.380 177.595 ;
        RECT 30.255 177.425 30.455 177.595 ;
        RECT 31.175 177.465 31.345 178.045 ;
        RECT 31.120 177.425 31.345 177.465 ;
        RECT 28.020 176.965 28.425 177.135 ;
        RECT 28.595 176.965 29.380 177.135 ;
        RECT 29.655 176.685 29.865 177.215 ;
        RECT 30.125 176.900 30.455 177.425 ;
        RECT 30.965 177.340 31.345 177.425 ;
        RECT 30.625 176.685 30.795 177.295 ;
        RECT 30.965 176.905 31.295 177.340 ;
        RECT 31.515 177.335 31.685 178.365 ;
        RECT 31.960 178.195 32.675 178.490 ;
        RECT 32.895 178.365 33.225 178.555 ;
        RECT 33.395 178.195 33.645 178.560 ;
        RECT 31.855 178.025 33.645 178.195 ;
        RECT 31.855 177.595 32.085 178.025 ;
        RECT 31.515 176.855 31.775 177.335 ;
        RECT 32.255 177.325 32.665 177.845 ;
        RECT 31.945 176.685 32.275 177.145 ;
        RECT 32.465 176.905 32.665 177.325 ;
        RECT 32.835 177.170 33.090 178.025 ;
        RECT 33.885 177.845 34.055 179.065 ;
        RECT 34.305 178.725 34.565 179.235 ;
        RECT 33.260 177.595 34.055 177.845 ;
        RECT 34.225 177.675 34.565 178.555 ;
        RECT 35.655 178.070 35.945 179.235 ;
        RECT 36.115 178.365 36.390 179.065 ;
        RECT 36.560 178.690 36.815 179.235 ;
        RECT 36.985 178.725 37.465 179.065 ;
        RECT 37.640 178.680 38.245 179.235 ;
        RECT 37.630 178.580 38.245 178.680 ;
        RECT 37.630 178.555 37.815 178.580 ;
        RECT 33.805 177.505 34.055 177.595 ;
        RECT 32.835 176.905 33.625 177.170 ;
        RECT 33.805 177.085 34.135 177.505 ;
        RECT 34.305 176.685 34.565 177.505 ;
        RECT 35.655 176.685 35.945 177.410 ;
        RECT 36.115 177.335 36.285 178.365 ;
        RECT 36.560 178.235 37.315 178.485 ;
        RECT 37.485 178.310 37.815 178.555 ;
        RECT 36.560 178.200 37.330 178.235 ;
        RECT 36.560 178.190 37.345 178.200 ;
        RECT 36.455 178.175 37.350 178.190 ;
        RECT 36.455 178.160 37.370 178.175 ;
        RECT 36.455 178.150 37.390 178.160 ;
        RECT 36.455 178.140 37.415 178.150 ;
        RECT 36.455 178.110 37.485 178.140 ;
        RECT 36.455 178.080 37.505 178.110 ;
        RECT 36.455 178.050 37.525 178.080 ;
        RECT 36.455 178.025 37.555 178.050 ;
        RECT 36.455 177.990 37.590 178.025 ;
        RECT 36.455 177.985 37.620 177.990 ;
        RECT 36.455 177.590 36.685 177.985 ;
        RECT 37.230 177.980 37.620 177.985 ;
        RECT 37.255 177.970 37.620 177.980 ;
        RECT 37.270 177.965 37.620 177.970 ;
        RECT 37.285 177.960 37.620 177.965 ;
        RECT 37.985 177.960 38.245 178.410 ;
        RECT 38.415 178.145 41.925 179.235 ;
        RECT 42.560 178.855 42.895 179.235 ;
        RECT 37.285 177.955 38.245 177.960 ;
        RECT 37.295 177.945 38.245 177.955 ;
        RECT 37.305 177.940 38.245 177.945 ;
        RECT 37.315 177.930 38.245 177.940 ;
        RECT 37.320 177.920 38.245 177.930 ;
        RECT 37.325 177.915 38.245 177.920 ;
        RECT 37.335 177.900 38.245 177.915 ;
        RECT 37.340 177.885 38.245 177.900 ;
        RECT 37.350 177.860 38.245 177.885 ;
        RECT 36.855 177.390 37.185 177.815 ;
        RECT 36.115 176.855 36.375 177.335 ;
        RECT 36.545 176.685 36.795 177.225 ;
        RECT 36.965 176.905 37.185 177.390 ;
        RECT 37.355 177.790 38.245 177.860 ;
        RECT 37.355 177.065 37.525 177.790 ;
        RECT 37.695 177.235 38.245 177.620 ;
        RECT 38.415 177.455 40.065 177.975 ;
        RECT 40.235 177.625 41.925 178.145 ;
        RECT 37.355 176.895 38.245 177.065 ;
        RECT 38.415 176.685 41.925 177.455 ;
        RECT 42.555 177.365 42.795 178.675 ;
        RECT 43.065 178.265 43.315 179.065 ;
        RECT 43.535 178.515 43.865 179.235 ;
        RECT 44.050 178.265 44.300 179.065 ;
        RECT 44.765 178.435 45.095 179.235 ;
        RECT 45.265 178.805 45.605 179.065 ;
        RECT 42.965 178.095 45.155 178.265 ;
        RECT 42.965 177.185 43.135 178.095 ;
        RECT 44.840 177.925 45.155 178.095 ;
        RECT 42.640 176.855 43.135 177.185 ;
        RECT 43.355 176.960 43.705 177.925 ;
        RECT 43.885 176.955 44.185 177.925 ;
        RECT 44.365 176.955 44.645 177.925 ;
        RECT 44.840 177.675 45.170 177.925 ;
        RECT 44.825 176.685 45.095 177.485 ;
        RECT 45.345 177.405 45.605 178.805 ;
        RECT 45.265 176.895 45.605 177.405 ;
        RECT 45.775 178.805 46.115 179.065 ;
        RECT 45.775 177.405 46.035 178.805 ;
        RECT 46.285 178.435 46.615 179.235 ;
        RECT 47.080 178.265 47.330 179.065 ;
        RECT 47.515 178.515 47.845 179.235 ;
        RECT 48.065 178.265 48.315 179.065 ;
        RECT 48.485 178.855 48.820 179.235 ;
        RECT 46.225 178.095 48.415 178.265 ;
        RECT 46.225 177.925 46.540 178.095 ;
        RECT 46.210 177.675 46.540 177.925 ;
        RECT 45.775 176.895 46.115 177.405 ;
        RECT 46.285 176.685 46.555 177.485 ;
        RECT 46.735 176.955 47.015 177.925 ;
        RECT 47.195 176.955 47.495 177.925 ;
        RECT 47.675 176.960 48.025 177.925 ;
        RECT 48.245 177.185 48.415 178.095 ;
        RECT 48.585 177.365 48.825 178.675 ;
        RECT 49.035 178.095 49.265 179.235 ;
        RECT 49.435 178.085 49.765 179.065 ;
        RECT 49.935 178.095 50.145 179.235 ;
        RECT 51.295 178.415 51.640 179.235 ;
        RECT 49.015 177.675 49.345 177.925 ;
        RECT 48.245 176.855 48.740 177.185 ;
        RECT 49.035 176.685 49.265 177.505 ;
        RECT 49.515 177.485 49.765 178.085 ;
        RECT 51.295 177.675 51.640 178.245 ;
        RECT 51.810 177.925 51.985 179.025 ;
        RECT 52.155 178.655 52.485 178.890 ;
        RECT 52.775 178.835 53.175 179.235 ;
        RECT 54.045 178.835 54.375 179.235 ;
        RECT 52.155 178.485 54.235 178.655 ;
        RECT 52.155 178.095 52.710 178.485 ;
        RECT 51.810 177.675 52.370 177.925 ;
        RECT 52.540 177.845 52.710 178.095 ;
        RECT 52.880 178.095 53.895 178.315 ;
        RECT 54.065 178.215 54.235 178.485 ;
        RECT 54.545 178.395 54.805 179.065 ;
        RECT 52.880 177.955 53.155 178.095 ;
        RECT 54.065 178.045 54.460 178.215 ;
        RECT 52.540 177.675 52.735 177.845 ;
        RECT 49.435 176.855 49.765 177.485 ;
        RECT 49.935 176.685 50.145 177.505 ;
        RECT 51.295 177.325 52.395 177.505 ;
        RECT 51.295 176.920 51.635 177.325 ;
        RECT 51.805 176.685 51.975 177.155 ;
        RECT 52.145 176.920 52.395 177.325 ;
        RECT 52.565 177.290 52.735 177.675 ;
        RECT 52.565 176.920 52.815 177.290 ;
        RECT 52.985 177.165 53.155 177.955 ;
        RECT 53.325 177.505 53.500 177.700 ;
        RECT 53.670 177.675 54.120 177.875 ;
        RECT 54.290 177.595 54.460 178.045 ;
        RECT 53.325 177.335 53.820 177.505 ;
        RECT 54.630 177.425 54.805 178.395 ;
        RECT 54.980 178.095 55.235 179.235 ;
        RECT 55.430 178.685 56.625 179.015 ;
        RECT 55.485 177.925 55.655 178.485 ;
        RECT 55.880 178.265 56.300 178.515 ;
        RECT 56.805 178.435 57.085 179.235 ;
        RECT 55.880 178.095 57.125 178.265 ;
        RECT 57.295 178.095 57.565 179.065 ;
        RECT 57.735 178.095 57.995 179.235 ;
        RECT 56.955 177.925 57.125 178.095 ;
        RECT 54.980 177.675 55.315 177.925 ;
        RECT 55.485 177.595 56.225 177.925 ;
        RECT 56.955 177.595 57.185 177.925 ;
        RECT 55.485 177.505 55.735 177.595 ;
        RECT 53.600 177.195 53.820 177.335 ;
        RECT 52.985 176.995 53.430 177.165 ;
        RECT 53.600 177.025 53.825 177.195 ;
        RECT 53.600 176.980 53.820 177.025 ;
        RECT 54.100 176.685 54.270 177.350 ;
        RECT 54.465 176.855 54.805 177.425 ;
        RECT 55.000 177.335 55.735 177.505 ;
        RECT 56.955 177.425 57.125 177.595 ;
        RECT 55.000 176.865 55.310 177.335 ;
        RECT 56.385 177.255 57.125 177.425 ;
        RECT 57.395 177.360 57.565 178.095 ;
        RECT 58.165 178.085 58.495 179.065 ;
        RECT 58.665 178.095 58.945 179.235 ;
        RECT 59.115 178.145 60.785 179.235 ;
        RECT 57.755 177.675 58.090 177.925 ;
        RECT 58.260 177.535 58.430 178.085 ;
        RECT 58.600 177.655 58.935 177.925 ;
        RECT 58.255 177.485 58.430 177.535 ;
        RECT 55.480 176.685 56.215 177.165 ;
        RECT 56.385 176.905 56.555 177.255 ;
        RECT 56.725 176.685 57.105 177.085 ;
        RECT 57.295 177.015 57.565 177.360 ;
        RECT 57.735 176.855 58.430 177.485 ;
        RECT 58.635 176.685 58.945 177.485 ;
        RECT 59.115 177.455 59.865 177.975 ;
        RECT 60.035 177.625 60.785 178.145 ;
        RECT 61.415 178.070 61.705 179.235 ;
        RECT 61.935 178.175 62.265 179.020 ;
        RECT 62.435 178.225 62.605 179.235 ;
        RECT 62.775 178.505 63.115 179.065 ;
        RECT 63.345 178.735 63.660 179.235 ;
        RECT 63.840 178.765 64.725 178.935 ;
        RECT 61.875 178.095 62.265 178.175 ;
        RECT 62.775 178.130 63.670 178.505 ;
        RECT 61.875 178.045 62.090 178.095 ;
        RECT 61.875 177.465 62.045 178.045 ;
        RECT 62.775 177.925 62.965 178.130 ;
        RECT 63.840 177.925 64.010 178.765 ;
        RECT 64.950 178.735 65.200 179.065 ;
        RECT 62.215 177.595 62.965 177.925 ;
        RECT 63.135 177.595 64.010 177.925 ;
        RECT 59.115 176.685 60.785 177.455 ;
        RECT 61.875 177.425 62.100 177.465 ;
        RECT 62.765 177.425 62.965 177.595 ;
        RECT 61.415 176.685 61.705 177.410 ;
        RECT 61.875 177.340 62.255 177.425 ;
        RECT 61.925 176.905 62.255 177.340 ;
        RECT 62.425 176.685 62.595 177.295 ;
        RECT 62.765 176.900 63.095 177.425 ;
        RECT 63.355 176.685 63.565 177.215 ;
        RECT 63.840 177.135 64.010 177.595 ;
        RECT 64.180 177.635 64.500 178.595 ;
        RECT 64.670 177.845 64.860 178.565 ;
        RECT 65.030 177.665 65.200 178.735 ;
        RECT 65.370 178.435 65.540 179.235 ;
        RECT 65.710 178.790 66.815 178.960 ;
        RECT 65.710 178.175 65.880 178.790 ;
        RECT 67.025 178.640 67.275 179.065 ;
        RECT 67.445 178.775 67.710 179.235 ;
        RECT 66.050 178.255 66.580 178.620 ;
        RECT 67.025 178.510 67.330 178.640 ;
        RECT 65.370 178.085 65.880 178.175 ;
        RECT 65.370 177.915 66.240 178.085 ;
        RECT 65.370 177.845 65.540 177.915 ;
        RECT 65.660 177.665 65.860 177.695 ;
        RECT 64.180 177.305 64.645 177.635 ;
        RECT 65.030 177.365 65.860 177.665 ;
        RECT 65.030 177.135 65.200 177.365 ;
        RECT 63.840 176.965 64.625 177.135 ;
        RECT 64.795 176.965 65.200 177.135 ;
        RECT 65.380 176.685 65.750 177.185 ;
        RECT 66.070 177.135 66.240 177.915 ;
        RECT 66.410 177.555 66.580 178.255 ;
        RECT 66.750 177.725 66.990 178.320 ;
        RECT 66.410 177.335 66.935 177.555 ;
        RECT 67.160 177.405 67.330 178.510 ;
        RECT 67.105 177.275 67.330 177.405 ;
        RECT 67.500 177.315 67.780 178.265 ;
        RECT 67.105 177.135 67.275 177.275 ;
        RECT 66.070 176.965 66.745 177.135 ;
        RECT 66.940 176.965 67.275 177.135 ;
        RECT 67.445 176.685 67.695 177.145 ;
        RECT 67.950 176.945 68.135 179.065 ;
        RECT 68.305 178.735 68.635 179.235 ;
        RECT 68.805 178.565 68.975 179.065 ;
        RECT 68.310 178.395 68.975 178.565 ;
        RECT 68.310 177.405 68.540 178.395 ;
        RECT 69.235 178.385 69.495 179.065 ;
        RECT 69.665 178.455 69.915 179.235 ;
        RECT 70.165 178.685 70.415 179.065 ;
        RECT 70.585 178.855 70.940 179.235 ;
        RECT 71.945 178.845 72.280 179.065 ;
        RECT 71.545 178.685 71.775 178.725 ;
        RECT 70.165 178.485 71.775 178.685 ;
        RECT 70.165 178.475 71.000 178.485 ;
        RECT 71.590 178.395 71.775 178.485 ;
        RECT 68.710 177.575 69.060 178.225 ;
        RECT 68.310 177.235 68.975 177.405 ;
        RECT 68.305 176.685 68.635 177.065 ;
        RECT 68.805 176.945 68.975 177.235 ;
        RECT 69.235 177.195 69.405 178.385 ;
        RECT 71.105 178.285 71.435 178.315 ;
        RECT 69.635 178.225 71.435 178.285 ;
        RECT 72.025 178.225 72.280 178.845 ;
        RECT 72.570 178.605 72.855 179.065 ;
        RECT 73.025 178.775 73.295 179.235 ;
        RECT 72.570 178.385 73.525 178.605 ;
        RECT 69.575 178.115 72.280 178.225 ;
        RECT 69.575 178.080 69.775 178.115 ;
        RECT 69.575 177.505 69.745 178.080 ;
        RECT 71.105 178.055 72.280 178.115 ;
        RECT 69.975 177.640 70.385 177.945 ;
        RECT 70.555 177.675 70.885 177.885 ;
        RECT 69.575 177.385 69.845 177.505 ;
        RECT 69.575 177.340 70.420 177.385 ;
        RECT 69.665 177.215 70.420 177.340 ;
        RECT 70.675 177.275 70.885 177.675 ;
        RECT 71.130 177.675 71.605 177.885 ;
        RECT 71.795 177.675 72.285 177.875 ;
        RECT 71.130 177.275 71.350 177.675 ;
        RECT 72.455 177.655 73.145 178.215 ;
        RECT 73.315 177.485 73.525 178.385 ;
        RECT 69.235 177.185 69.465 177.195 ;
        RECT 69.235 176.855 69.495 177.185 ;
        RECT 70.250 177.065 70.420 177.215 ;
        RECT 69.665 176.685 69.995 177.045 ;
        RECT 70.250 176.855 71.550 177.065 ;
        RECT 71.825 176.685 72.280 177.450 ;
        RECT 72.570 177.315 73.525 177.485 ;
        RECT 73.695 178.215 74.095 179.065 ;
        RECT 74.285 178.605 74.565 179.065 ;
        RECT 75.085 178.775 75.410 179.235 ;
        RECT 74.285 178.385 75.410 178.605 ;
        RECT 73.695 177.655 74.790 178.215 ;
        RECT 74.960 177.925 75.410 178.385 ;
        RECT 75.580 178.095 75.965 179.065 ;
        RECT 76.135 178.145 77.805 179.235 ;
        RECT 78.525 178.565 78.695 179.065 ;
        RECT 78.865 178.735 79.195 179.235 ;
        RECT 78.525 178.395 79.190 178.565 ;
        RECT 72.570 176.855 72.855 177.315 ;
        RECT 73.025 176.685 73.295 177.145 ;
        RECT 73.695 176.855 74.095 177.655 ;
        RECT 74.960 177.595 75.515 177.925 ;
        RECT 74.960 177.485 75.410 177.595 ;
        RECT 74.285 177.315 75.410 177.485 ;
        RECT 75.685 177.425 75.965 178.095 ;
        RECT 74.285 176.855 74.565 177.315 ;
        RECT 75.085 176.685 75.410 177.145 ;
        RECT 75.580 176.855 75.965 177.425 ;
        RECT 76.135 177.455 76.885 177.975 ;
        RECT 77.055 177.625 77.805 178.145 ;
        RECT 78.440 177.575 78.790 178.225 ;
        RECT 76.135 176.685 77.805 177.455 ;
        RECT 78.960 177.405 79.190 178.395 ;
        RECT 78.525 177.235 79.190 177.405 ;
        RECT 78.525 176.945 78.695 177.235 ;
        RECT 78.865 176.685 79.195 177.065 ;
        RECT 79.365 176.945 79.550 179.065 ;
        RECT 79.790 178.775 80.055 179.235 ;
        RECT 80.225 178.640 80.475 179.065 ;
        RECT 80.685 178.790 81.790 178.960 ;
        RECT 80.170 178.510 80.475 178.640 ;
        RECT 79.720 177.315 80.000 178.265 ;
        RECT 80.170 177.405 80.340 178.510 ;
        RECT 80.510 177.725 80.750 178.320 ;
        RECT 80.920 178.255 81.450 178.620 ;
        RECT 80.920 177.555 81.090 178.255 ;
        RECT 81.620 178.175 81.790 178.790 ;
        RECT 81.960 178.435 82.130 179.235 ;
        RECT 82.300 178.735 82.550 179.065 ;
        RECT 82.775 178.765 83.660 178.935 ;
        RECT 81.620 178.085 82.130 178.175 ;
        RECT 80.170 177.275 80.395 177.405 ;
        RECT 80.565 177.335 81.090 177.555 ;
        RECT 81.260 177.915 82.130 178.085 ;
        RECT 79.805 176.685 80.055 177.145 ;
        RECT 80.225 177.135 80.395 177.275 ;
        RECT 81.260 177.135 81.430 177.915 ;
        RECT 81.960 177.845 82.130 177.915 ;
        RECT 81.640 177.665 81.840 177.695 ;
        RECT 82.300 177.665 82.470 178.735 ;
        RECT 82.640 177.845 82.830 178.565 ;
        RECT 81.640 177.365 82.470 177.665 ;
        RECT 83.000 177.635 83.320 178.595 ;
        RECT 80.225 176.965 80.560 177.135 ;
        RECT 80.755 176.965 81.430 177.135 ;
        RECT 81.750 176.685 82.120 177.185 ;
        RECT 82.300 177.135 82.470 177.365 ;
        RECT 82.855 177.305 83.320 177.635 ;
        RECT 83.490 177.925 83.660 178.765 ;
        RECT 83.840 178.735 84.155 179.235 ;
        RECT 84.385 178.505 84.725 179.065 ;
        RECT 83.830 178.130 84.725 178.505 ;
        RECT 84.895 178.225 85.065 179.235 ;
        RECT 84.535 177.925 84.725 178.130 ;
        RECT 85.235 178.175 85.565 179.020 ;
        RECT 85.235 178.095 85.625 178.175 ;
        RECT 85.795 178.145 87.005 179.235 ;
        RECT 85.410 178.045 85.625 178.095 ;
        RECT 83.490 177.595 84.365 177.925 ;
        RECT 84.535 177.595 85.285 177.925 ;
        RECT 83.490 177.135 83.660 177.595 ;
        RECT 84.535 177.425 84.735 177.595 ;
        RECT 85.455 177.465 85.625 178.045 ;
        RECT 85.400 177.425 85.625 177.465 ;
        RECT 82.300 176.965 82.705 177.135 ;
        RECT 82.875 176.965 83.660 177.135 ;
        RECT 83.935 176.685 84.145 177.215 ;
        RECT 84.405 176.900 84.735 177.425 ;
        RECT 85.245 177.340 85.625 177.425 ;
        RECT 85.795 177.435 86.315 177.975 ;
        RECT 86.485 177.605 87.005 178.145 ;
        RECT 87.175 178.070 87.465 179.235 ;
        RECT 87.635 178.145 89.305 179.235 ;
        RECT 87.635 177.455 88.385 177.975 ;
        RECT 88.555 177.625 89.305 178.145 ;
        RECT 89.480 178.095 89.735 179.235 ;
        RECT 89.930 178.685 91.125 179.015 ;
        RECT 89.985 177.925 90.155 178.485 ;
        RECT 90.380 178.265 90.800 178.515 ;
        RECT 91.305 178.435 91.585 179.235 ;
        RECT 90.380 178.095 91.625 178.265 ;
        RECT 91.795 178.095 92.065 179.065 ;
        RECT 92.880 178.265 93.270 178.440 ;
        RECT 93.755 178.435 94.085 179.235 ;
        RECT 94.255 178.445 94.790 179.065 ;
        RECT 92.880 178.095 94.305 178.265 ;
        RECT 91.455 177.925 91.625 178.095 ;
        RECT 89.480 177.675 89.815 177.925 ;
        RECT 89.985 177.595 90.725 177.925 ;
        RECT 91.455 177.595 91.685 177.925 ;
        RECT 89.985 177.505 90.235 177.595 ;
        RECT 84.905 176.685 85.075 177.295 ;
        RECT 85.245 176.905 85.575 177.340 ;
        RECT 85.795 176.685 87.005 177.435 ;
        RECT 87.175 176.685 87.465 177.410 ;
        RECT 87.635 176.685 89.305 177.455 ;
        RECT 89.500 177.335 90.235 177.505 ;
        RECT 91.455 177.425 91.625 177.595 ;
        RECT 89.500 176.865 89.810 177.335 ;
        RECT 90.885 177.255 91.625 177.425 ;
        RECT 91.895 177.360 92.065 178.095 ;
        RECT 92.755 177.365 93.110 177.925 ;
        RECT 89.980 176.685 90.715 177.165 ;
        RECT 90.885 176.905 91.055 177.255 ;
        RECT 91.225 176.685 91.605 177.085 ;
        RECT 91.795 177.015 92.065 177.360 ;
        RECT 93.280 177.195 93.450 178.095 ;
        RECT 93.620 177.365 93.885 177.925 ;
        RECT 94.135 177.595 94.305 178.095 ;
        RECT 94.475 177.425 94.790 178.445 ;
        RECT 92.860 176.685 93.100 177.195 ;
        RECT 93.280 176.865 93.560 177.195 ;
        RECT 93.790 176.685 94.005 177.195 ;
        RECT 94.175 176.855 94.790 177.425 ;
        RECT 94.995 178.365 95.270 179.065 ;
        RECT 95.440 178.690 95.695 179.235 ;
        RECT 95.865 178.725 96.345 179.065 ;
        RECT 96.520 178.680 97.125 179.235 ;
        RECT 96.510 178.580 97.125 178.680 ;
        RECT 96.510 178.555 96.695 178.580 ;
        RECT 94.995 177.335 95.165 178.365 ;
        RECT 95.440 178.235 96.195 178.485 ;
        RECT 96.365 178.310 96.695 178.555 ;
        RECT 95.440 178.200 96.210 178.235 ;
        RECT 95.440 178.190 96.225 178.200 ;
        RECT 95.335 178.175 96.230 178.190 ;
        RECT 95.335 178.160 96.250 178.175 ;
        RECT 95.335 178.150 96.270 178.160 ;
        RECT 95.335 178.140 96.295 178.150 ;
        RECT 95.335 178.110 96.365 178.140 ;
        RECT 95.335 178.080 96.385 178.110 ;
        RECT 95.335 178.050 96.405 178.080 ;
        RECT 95.335 178.025 96.435 178.050 ;
        RECT 95.335 177.990 96.470 178.025 ;
        RECT 95.335 177.985 96.500 177.990 ;
        RECT 95.335 177.590 95.565 177.985 ;
        RECT 96.110 177.980 96.500 177.985 ;
        RECT 96.135 177.970 96.500 177.980 ;
        RECT 96.150 177.965 96.500 177.970 ;
        RECT 96.165 177.960 96.500 177.965 ;
        RECT 96.865 177.960 97.125 178.410 ;
        RECT 97.385 178.305 97.555 179.065 ;
        RECT 97.735 178.475 98.065 179.235 ;
        RECT 97.385 178.135 98.050 178.305 ;
        RECT 98.235 178.160 98.505 179.065 ;
        RECT 96.165 177.955 97.125 177.960 ;
        RECT 97.880 177.990 98.050 178.135 ;
        RECT 96.175 177.945 97.125 177.955 ;
        RECT 96.185 177.940 97.125 177.945 ;
        RECT 96.195 177.930 97.125 177.940 ;
        RECT 96.200 177.920 97.125 177.930 ;
        RECT 96.205 177.915 97.125 177.920 ;
        RECT 96.215 177.900 97.125 177.915 ;
        RECT 96.220 177.885 97.125 177.900 ;
        RECT 96.230 177.860 97.125 177.885 ;
        RECT 95.735 177.390 96.065 177.815 ;
        RECT 94.995 176.855 95.255 177.335 ;
        RECT 95.425 176.685 95.675 177.225 ;
        RECT 95.845 176.905 96.065 177.390 ;
        RECT 96.235 177.790 97.125 177.860 ;
        RECT 96.235 177.065 96.405 177.790 ;
        RECT 96.575 177.235 97.125 177.620 ;
        RECT 97.315 177.585 97.645 177.955 ;
        RECT 97.880 177.660 98.165 177.990 ;
        RECT 97.880 177.405 98.050 177.660 ;
        RECT 97.385 177.235 98.050 177.405 ;
        RECT 98.335 177.360 98.505 178.160 ;
        RECT 96.235 176.895 97.125 177.065 ;
        RECT 97.385 176.855 97.555 177.235 ;
        RECT 97.735 176.685 98.065 177.065 ;
        RECT 98.245 176.855 98.505 177.360 ;
        RECT 99.135 177.630 99.415 179.065 ;
        RECT 99.585 178.460 100.295 179.235 ;
        RECT 100.465 178.290 100.795 179.065 ;
        RECT 99.645 178.075 100.795 178.290 ;
        RECT 99.135 176.855 99.475 177.630 ;
        RECT 99.645 177.505 99.930 178.075 ;
        RECT 100.115 177.675 100.585 177.905 ;
        RECT 100.990 177.875 101.205 178.990 ;
        RECT 101.385 178.515 101.715 179.235 ;
        RECT 101.495 177.875 101.725 178.215 ;
        RECT 100.755 177.695 101.205 177.875 ;
        RECT 100.755 177.675 101.085 177.695 ;
        RECT 101.395 177.675 101.725 177.875 ;
        RECT 101.895 178.045 102.355 179.055 ;
        RECT 103.425 178.725 103.755 179.235 ;
        RECT 104.735 178.605 104.915 179.065 ;
        RECT 105.085 178.775 105.335 179.235 ;
        RECT 105.505 178.855 105.835 179.025 ;
        RECT 106.005 178.970 106.260 179.065 ;
        RECT 105.505 178.605 105.675 178.855 ;
        RECT 106.005 178.800 107.145 178.970 ;
        RECT 107.405 178.835 107.735 179.235 ;
        RECT 106.005 178.665 106.260 178.800 ;
        RECT 102.525 178.385 104.485 178.555 ;
        RECT 104.735 178.435 105.675 178.605 ;
        RECT 105.850 178.495 106.260 178.665 ;
        RECT 106.975 178.575 107.145 178.800 ;
        RECT 99.645 177.315 100.355 177.505 ;
        RECT 100.055 177.175 100.355 177.315 ;
        RECT 100.545 177.315 101.725 177.505 ;
        RECT 100.545 177.235 100.875 177.315 ;
        RECT 100.055 177.165 100.370 177.175 ;
        RECT 100.055 177.155 100.380 177.165 ;
        RECT 100.055 177.150 100.390 177.155 ;
        RECT 99.645 176.685 99.815 177.145 ;
        RECT 100.055 177.140 100.395 177.150 ;
        RECT 100.055 177.135 100.400 177.140 ;
        RECT 100.055 177.125 100.405 177.135 ;
        RECT 100.055 177.120 100.410 177.125 ;
        RECT 100.055 176.855 100.415 177.120 ;
        RECT 101.045 176.685 101.215 177.145 ;
        RECT 101.385 176.855 101.725 177.315 ;
        RECT 101.895 177.425 102.065 178.045 ;
        RECT 102.525 177.845 102.695 178.385 ;
        RECT 102.235 177.675 102.695 177.845 ;
        RECT 102.875 177.595 103.115 178.215 ;
        RECT 103.285 177.595 103.625 178.215 ;
        RECT 103.795 177.595 104.145 178.215 ;
        RECT 104.315 177.425 104.485 178.385 ;
        RECT 101.895 177.255 103.255 177.425 ;
        RECT 101.895 176.855 102.415 177.255 ;
        RECT 102.585 176.685 102.915 177.085 ;
        RECT 103.085 176.910 103.255 177.255 ;
        RECT 103.425 176.685 103.755 177.425 ;
        RECT 103.990 177.255 104.485 177.425 ;
        RECT 104.710 177.365 104.970 178.255 ;
        RECT 105.170 177.955 105.650 178.255 ;
        RECT 105.170 177.365 105.430 177.955 ;
        RECT 105.850 177.470 106.020 178.495 ;
        RECT 106.540 178.315 106.710 178.505 ;
        RECT 106.975 178.405 107.735 178.575 ;
        RECT 105.670 177.300 106.020 177.470 ;
        RECT 106.190 178.145 106.710 178.315 ;
        RECT 106.190 177.425 106.360 178.145 ;
        RECT 106.550 177.595 106.840 177.975 ;
        RECT 107.010 177.595 107.340 178.215 ;
        RECT 107.565 177.925 107.735 178.405 ;
        RECT 107.905 178.125 108.165 179.065 ;
        RECT 108.335 178.145 111.845 179.235 ;
        RECT 107.565 177.595 107.820 177.925 ;
        RECT 103.990 177.005 104.160 177.255 ;
        RECT 104.695 176.685 105.095 177.195 ;
        RECT 105.670 176.855 105.840 177.300 ;
        RECT 106.190 177.255 107.070 177.425 ;
        RECT 107.990 177.410 108.165 178.125 ;
        RECT 106.010 176.685 106.730 177.085 ;
        RECT 106.900 176.855 107.070 177.255 ;
        RECT 107.305 176.685 107.735 177.130 ;
        RECT 107.905 176.855 108.165 177.410 ;
        RECT 108.335 177.455 109.985 177.975 ;
        RECT 110.155 177.625 111.845 178.145 ;
        RECT 112.935 178.070 113.225 179.235 ;
        RECT 113.485 178.565 113.655 179.065 ;
        RECT 113.825 178.735 114.155 179.235 ;
        RECT 113.485 178.395 114.150 178.565 ;
        RECT 113.400 177.575 113.750 178.225 ;
        RECT 108.335 176.685 111.845 177.455 ;
        RECT 112.935 176.685 113.225 177.410 ;
        RECT 113.920 177.405 114.150 178.395 ;
        RECT 113.485 177.235 114.150 177.405 ;
        RECT 113.485 176.945 113.655 177.235 ;
        RECT 113.825 176.685 114.155 177.065 ;
        RECT 114.325 176.945 114.510 179.065 ;
        RECT 114.750 178.775 115.015 179.235 ;
        RECT 115.185 178.640 115.435 179.065 ;
        RECT 115.645 178.790 116.750 178.960 ;
        RECT 115.130 178.510 115.435 178.640 ;
        RECT 114.680 177.315 114.960 178.265 ;
        RECT 115.130 177.405 115.300 178.510 ;
        RECT 115.470 177.725 115.710 178.320 ;
        RECT 115.880 178.255 116.410 178.620 ;
        RECT 115.880 177.555 116.050 178.255 ;
        RECT 116.580 178.175 116.750 178.790 ;
        RECT 116.920 178.435 117.090 179.235 ;
        RECT 117.260 178.735 117.510 179.065 ;
        RECT 117.735 178.765 118.620 178.935 ;
        RECT 116.580 178.085 117.090 178.175 ;
        RECT 115.130 177.275 115.355 177.405 ;
        RECT 115.525 177.335 116.050 177.555 ;
        RECT 116.220 177.915 117.090 178.085 ;
        RECT 114.765 176.685 115.015 177.145 ;
        RECT 115.185 177.135 115.355 177.275 ;
        RECT 116.220 177.135 116.390 177.915 ;
        RECT 116.920 177.845 117.090 177.915 ;
        RECT 116.600 177.665 116.800 177.695 ;
        RECT 117.260 177.665 117.430 178.735 ;
        RECT 117.600 177.845 117.790 178.565 ;
        RECT 116.600 177.365 117.430 177.665 ;
        RECT 117.960 177.635 118.280 178.595 ;
        RECT 115.185 176.965 115.520 177.135 ;
        RECT 115.715 176.965 116.390 177.135 ;
        RECT 116.710 176.685 117.080 177.185 ;
        RECT 117.260 177.135 117.430 177.365 ;
        RECT 117.815 177.305 118.280 177.635 ;
        RECT 118.450 177.925 118.620 178.765 ;
        RECT 118.800 178.735 119.115 179.235 ;
        RECT 119.345 178.505 119.685 179.065 ;
        RECT 118.790 178.130 119.685 178.505 ;
        RECT 119.855 178.225 120.025 179.235 ;
        RECT 119.495 177.925 119.685 178.130 ;
        RECT 120.195 178.175 120.525 179.020 ;
        RECT 120.845 178.565 121.015 179.065 ;
        RECT 121.185 178.735 121.515 179.235 ;
        RECT 120.845 178.395 121.510 178.565 ;
        RECT 120.195 178.095 120.585 178.175 ;
        RECT 120.370 178.045 120.585 178.095 ;
        RECT 118.450 177.595 119.325 177.925 ;
        RECT 119.495 177.595 120.245 177.925 ;
        RECT 118.450 177.135 118.620 177.595 ;
        RECT 119.495 177.425 119.695 177.595 ;
        RECT 120.415 177.465 120.585 178.045 ;
        RECT 120.760 177.575 121.110 178.225 ;
        RECT 120.360 177.425 120.585 177.465 ;
        RECT 117.260 176.965 117.665 177.135 ;
        RECT 117.835 176.965 118.620 177.135 ;
        RECT 118.895 176.685 119.105 177.215 ;
        RECT 119.365 176.900 119.695 177.425 ;
        RECT 120.205 177.340 120.585 177.425 ;
        RECT 121.280 177.405 121.510 178.395 ;
        RECT 119.865 176.685 120.035 177.295 ;
        RECT 120.205 176.905 120.535 177.340 ;
        RECT 120.845 177.235 121.510 177.405 ;
        RECT 120.845 176.945 121.015 177.235 ;
        RECT 121.185 176.685 121.515 177.065 ;
        RECT 121.685 176.945 121.870 179.065 ;
        RECT 122.110 178.775 122.375 179.235 ;
        RECT 122.545 178.640 122.795 179.065 ;
        RECT 123.005 178.790 124.110 178.960 ;
        RECT 122.490 178.510 122.795 178.640 ;
        RECT 122.040 177.315 122.320 178.265 ;
        RECT 122.490 177.405 122.660 178.510 ;
        RECT 122.830 177.725 123.070 178.320 ;
        RECT 123.240 178.255 123.770 178.620 ;
        RECT 123.240 177.555 123.410 178.255 ;
        RECT 123.940 178.175 124.110 178.790 ;
        RECT 124.280 178.435 124.450 179.235 ;
        RECT 124.620 178.735 124.870 179.065 ;
        RECT 125.095 178.765 125.980 178.935 ;
        RECT 123.940 178.085 124.450 178.175 ;
        RECT 122.490 177.275 122.715 177.405 ;
        RECT 122.885 177.335 123.410 177.555 ;
        RECT 123.580 177.915 124.450 178.085 ;
        RECT 122.125 176.685 122.375 177.145 ;
        RECT 122.545 177.135 122.715 177.275 ;
        RECT 123.580 177.135 123.750 177.915 ;
        RECT 124.280 177.845 124.450 177.915 ;
        RECT 123.960 177.665 124.160 177.695 ;
        RECT 124.620 177.665 124.790 178.735 ;
        RECT 124.960 177.845 125.150 178.565 ;
        RECT 123.960 177.365 124.790 177.665 ;
        RECT 125.320 177.635 125.640 178.595 ;
        RECT 122.545 176.965 122.880 177.135 ;
        RECT 123.075 176.965 123.750 177.135 ;
        RECT 124.070 176.685 124.440 177.185 ;
        RECT 124.620 177.135 124.790 177.365 ;
        RECT 125.175 177.305 125.640 177.635 ;
        RECT 125.810 177.925 125.980 178.765 ;
        RECT 126.160 178.735 126.475 179.235 ;
        RECT 126.705 178.505 127.045 179.065 ;
        RECT 126.150 178.130 127.045 178.505 ;
        RECT 127.215 178.225 127.385 179.235 ;
        RECT 126.855 177.925 127.045 178.130 ;
        RECT 127.555 178.175 127.885 179.020 ;
        RECT 128.205 178.615 128.375 179.045 ;
        RECT 128.545 178.785 128.875 179.235 ;
        RECT 128.205 178.385 128.880 178.615 ;
        RECT 127.555 178.095 127.945 178.175 ;
        RECT 127.730 178.045 127.945 178.095 ;
        RECT 125.810 177.595 126.685 177.925 ;
        RECT 126.855 177.595 127.605 177.925 ;
        RECT 125.810 177.135 125.980 177.595 ;
        RECT 126.855 177.425 127.055 177.595 ;
        RECT 127.775 177.465 127.945 178.045 ;
        RECT 127.720 177.425 127.945 177.465 ;
        RECT 124.620 176.965 125.025 177.135 ;
        RECT 125.195 176.965 125.980 177.135 ;
        RECT 126.255 176.685 126.465 177.215 ;
        RECT 126.725 176.900 127.055 177.425 ;
        RECT 127.565 177.340 127.945 177.425 ;
        RECT 128.175 177.365 128.475 178.215 ;
        RECT 128.645 177.735 128.880 178.385 ;
        RECT 129.050 178.075 129.335 179.020 ;
        RECT 129.515 178.765 130.200 179.235 ;
        RECT 129.510 178.245 130.205 178.555 ;
        RECT 130.380 178.180 130.685 178.965 ;
        RECT 129.050 177.925 129.910 178.075 ;
        RECT 130.475 178.045 130.685 178.180 ;
        RECT 130.875 178.145 132.545 179.235 ;
        RECT 133.175 178.435 133.500 179.235 ;
        RECT 129.050 177.905 130.335 177.925 ;
        RECT 128.645 177.405 129.180 177.735 ;
        RECT 129.350 177.545 130.335 177.905 ;
        RECT 127.225 176.685 127.395 177.295 ;
        RECT 127.565 176.905 127.895 177.340 ;
        RECT 128.645 177.255 128.865 177.405 ;
        RECT 128.120 176.685 128.455 177.190 ;
        RECT 128.625 176.880 128.865 177.255 ;
        RECT 129.350 177.210 129.520 177.545 ;
        RECT 130.510 177.375 130.685 178.045 ;
        RECT 129.145 177.015 129.520 177.210 ;
        RECT 129.145 176.870 129.315 177.015 ;
        RECT 129.880 176.685 130.275 177.180 ;
        RECT 130.445 176.855 130.685 177.375 ;
        RECT 130.875 177.455 131.625 177.975 ;
        RECT 131.795 177.625 132.545 178.145 ;
        RECT 133.195 177.675 133.525 178.260 ;
        RECT 133.695 177.925 133.880 179.015 ;
        RECT 134.050 178.265 134.300 179.065 ;
        RECT 134.470 178.435 135.210 179.235 ;
        RECT 135.395 178.265 135.725 179.065 ;
        RECT 135.895 178.435 136.705 179.235 ;
        RECT 134.050 178.095 136.535 178.265 ;
        RECT 136.365 177.925 136.535 178.095 ;
        RECT 133.695 177.675 134.180 177.925 ;
        RECT 134.525 177.595 134.785 177.925 ;
        RECT 130.875 176.685 132.545 177.455 ;
        RECT 133.175 177.305 134.360 177.475 ;
        RECT 133.175 176.855 133.440 177.305 ;
        RECT 133.610 176.685 133.900 177.135 ;
        RECT 134.070 176.855 134.360 177.305 ;
        RECT 134.540 176.990 134.785 177.595 ;
        RECT 135.035 176.990 135.305 177.925 ;
        RECT 135.485 177.675 135.965 177.925 ;
        RECT 135.485 176.990 135.695 177.675 ;
        RECT 136.365 177.595 136.705 177.925 ;
        RECT 136.365 177.505 136.535 177.595 ;
        RECT 135.865 177.335 136.535 177.505 ;
        RECT 135.865 176.855 136.205 177.335 ;
        RECT 136.385 176.685 136.695 177.165 ;
        RECT 136.875 176.855 137.135 179.065 ;
        RECT 137.355 178.095 137.585 179.235 ;
        RECT 137.755 178.085 138.085 179.065 ;
        RECT 138.255 178.095 138.465 179.235 ;
        RECT 137.335 177.675 137.665 177.925 ;
        RECT 137.355 176.685 137.585 177.505 ;
        RECT 137.835 177.485 138.085 178.085 ;
        RECT 138.695 178.070 138.985 179.235 ;
        RECT 139.155 177.630 139.435 179.065 ;
        RECT 139.605 178.460 140.315 179.235 ;
        RECT 140.485 178.290 140.815 179.065 ;
        RECT 139.665 178.075 140.815 178.290 ;
        RECT 137.755 176.855 138.085 177.485 ;
        RECT 138.255 176.685 138.465 177.505 ;
        RECT 138.695 176.685 138.985 177.410 ;
        RECT 139.155 176.855 139.495 177.630 ;
        RECT 139.665 177.505 139.950 178.075 ;
        RECT 140.135 177.675 140.605 177.905 ;
        RECT 141.010 177.875 141.225 178.990 ;
        RECT 141.405 178.515 141.735 179.235 ;
        RECT 141.915 178.365 142.190 179.065 ;
        RECT 142.360 178.690 142.615 179.235 ;
        RECT 142.785 178.725 143.265 179.065 ;
        RECT 143.440 178.680 144.045 179.235 ;
        RECT 143.430 178.580 144.045 178.680 ;
        RECT 143.430 178.555 143.615 178.580 ;
        RECT 141.515 177.875 141.745 178.215 ;
        RECT 140.775 177.695 141.225 177.875 ;
        RECT 140.775 177.675 141.105 177.695 ;
        RECT 141.415 177.675 141.745 177.875 ;
        RECT 139.665 177.315 140.375 177.505 ;
        RECT 140.075 177.175 140.375 177.315 ;
        RECT 140.565 177.315 141.745 177.505 ;
        RECT 140.565 177.235 140.895 177.315 ;
        RECT 140.075 177.165 140.390 177.175 ;
        RECT 140.075 177.155 140.400 177.165 ;
        RECT 140.075 177.150 140.410 177.155 ;
        RECT 139.665 176.685 139.835 177.145 ;
        RECT 140.075 177.140 140.415 177.150 ;
        RECT 140.075 177.135 140.420 177.140 ;
        RECT 140.075 177.125 140.425 177.135 ;
        RECT 140.075 177.120 140.430 177.125 ;
        RECT 140.075 176.855 140.435 177.120 ;
        RECT 141.065 176.685 141.235 177.145 ;
        RECT 141.405 176.855 141.745 177.315 ;
        RECT 141.915 177.335 142.085 178.365 ;
        RECT 142.360 178.235 143.115 178.485 ;
        RECT 143.285 178.310 143.615 178.555 ;
        RECT 142.360 178.200 143.130 178.235 ;
        RECT 142.360 178.190 143.145 178.200 ;
        RECT 142.255 178.175 143.150 178.190 ;
        RECT 142.255 178.160 143.170 178.175 ;
        RECT 142.255 178.150 143.190 178.160 ;
        RECT 142.255 178.140 143.215 178.150 ;
        RECT 142.255 178.110 143.285 178.140 ;
        RECT 142.255 178.080 143.305 178.110 ;
        RECT 142.255 178.050 143.325 178.080 ;
        RECT 142.255 178.025 143.355 178.050 ;
        RECT 142.255 177.990 143.390 178.025 ;
        RECT 142.255 177.985 143.420 177.990 ;
        RECT 142.255 177.590 142.485 177.985 ;
        RECT 143.030 177.980 143.420 177.985 ;
        RECT 143.055 177.970 143.420 177.980 ;
        RECT 143.070 177.965 143.420 177.970 ;
        RECT 143.085 177.960 143.420 177.965 ;
        RECT 143.785 177.960 144.045 178.410 ;
        RECT 144.420 178.265 144.750 179.065 ;
        RECT 144.920 178.435 145.250 179.235 ;
        RECT 145.550 178.265 145.880 179.065 ;
        RECT 146.525 178.435 146.775 179.235 ;
        RECT 144.420 178.095 146.855 178.265 ;
        RECT 147.045 178.095 147.215 179.235 ;
        RECT 147.385 178.095 147.725 179.065 ;
        RECT 147.985 178.565 148.155 179.065 ;
        RECT 148.325 178.735 148.655 179.235 ;
        RECT 147.985 178.395 148.650 178.565 ;
        RECT 143.085 177.955 144.045 177.960 ;
        RECT 143.095 177.945 144.045 177.955 ;
        RECT 143.105 177.940 144.045 177.945 ;
        RECT 143.115 177.930 144.045 177.940 ;
        RECT 143.120 177.920 144.045 177.930 ;
        RECT 143.125 177.915 144.045 177.920 ;
        RECT 143.135 177.900 144.045 177.915 ;
        RECT 143.140 177.885 144.045 177.900 ;
        RECT 143.150 177.860 144.045 177.885 ;
        RECT 142.655 177.390 142.985 177.815 ;
        RECT 142.735 177.365 142.985 177.390 ;
        RECT 141.915 176.855 142.175 177.335 ;
        RECT 142.345 176.685 142.595 177.225 ;
        RECT 142.765 176.905 142.985 177.365 ;
        RECT 143.155 177.790 144.045 177.860 ;
        RECT 143.155 177.065 143.325 177.790 ;
        RECT 144.215 177.675 144.565 177.925 ;
        RECT 143.495 177.235 144.045 177.620 ;
        RECT 144.750 177.465 144.920 178.095 ;
        RECT 145.090 177.675 145.420 177.875 ;
        RECT 145.590 177.675 145.920 177.875 ;
        RECT 146.090 177.675 146.510 177.875 ;
        RECT 146.685 177.845 146.855 178.095 ;
        RECT 146.685 177.675 147.380 177.845 ;
        RECT 143.155 176.895 144.045 177.065 ;
        RECT 144.420 176.855 144.920 177.465 ;
        RECT 145.550 177.335 146.775 177.505 ;
        RECT 147.550 177.485 147.725 178.095 ;
        RECT 147.900 177.575 148.250 178.225 ;
        RECT 145.550 176.855 145.880 177.335 ;
        RECT 146.050 176.685 146.275 177.145 ;
        RECT 146.445 176.855 146.775 177.335 ;
        RECT 146.965 176.685 147.215 177.485 ;
        RECT 147.385 176.855 147.725 177.485 ;
        RECT 148.420 177.405 148.650 178.395 ;
        RECT 147.985 177.235 148.650 177.405 ;
        RECT 147.985 176.945 148.155 177.235 ;
        RECT 148.325 176.685 148.655 177.065 ;
        RECT 148.825 176.945 149.010 179.065 ;
        RECT 149.250 178.775 149.515 179.235 ;
        RECT 149.685 178.640 149.935 179.065 ;
        RECT 150.145 178.790 151.250 178.960 ;
        RECT 149.630 178.510 149.935 178.640 ;
        RECT 149.180 177.315 149.460 178.265 ;
        RECT 149.630 177.405 149.800 178.510 ;
        RECT 149.970 177.725 150.210 178.320 ;
        RECT 150.380 178.255 150.910 178.620 ;
        RECT 150.380 177.555 150.550 178.255 ;
        RECT 151.080 178.175 151.250 178.790 ;
        RECT 151.420 178.435 151.590 179.235 ;
        RECT 151.760 178.735 152.010 179.065 ;
        RECT 152.235 178.765 153.120 178.935 ;
        RECT 151.080 178.085 151.590 178.175 ;
        RECT 149.630 177.275 149.855 177.405 ;
        RECT 150.025 177.335 150.550 177.555 ;
        RECT 150.720 177.915 151.590 178.085 ;
        RECT 149.265 176.685 149.515 177.145 ;
        RECT 149.685 177.135 149.855 177.275 ;
        RECT 150.720 177.135 150.890 177.915 ;
        RECT 151.420 177.845 151.590 177.915 ;
        RECT 151.100 177.665 151.300 177.695 ;
        RECT 151.760 177.665 151.930 178.735 ;
        RECT 152.100 177.845 152.290 178.565 ;
        RECT 151.100 177.365 151.930 177.665 ;
        RECT 152.460 177.635 152.780 178.595 ;
        RECT 149.685 176.965 150.020 177.135 ;
        RECT 150.215 176.965 150.890 177.135 ;
        RECT 151.210 176.685 151.580 177.185 ;
        RECT 151.760 177.135 151.930 177.365 ;
        RECT 152.315 177.305 152.780 177.635 ;
        RECT 152.950 177.925 153.120 178.765 ;
        RECT 153.300 178.735 153.615 179.235 ;
        RECT 153.845 178.505 154.185 179.065 ;
        RECT 153.290 178.130 154.185 178.505 ;
        RECT 154.355 178.225 154.525 179.235 ;
        RECT 153.995 177.925 154.185 178.130 ;
        RECT 154.695 178.175 155.025 179.020 ;
        RECT 154.695 178.095 155.085 178.175 ;
        RECT 154.870 178.045 155.085 178.095 ;
        RECT 152.950 177.595 153.825 177.925 ;
        RECT 153.995 177.595 154.745 177.925 ;
        RECT 152.950 177.135 153.120 177.595 ;
        RECT 153.995 177.425 154.195 177.595 ;
        RECT 154.915 177.465 155.085 178.045 ;
        RECT 155.715 178.145 156.925 179.235 ;
        RECT 155.715 177.605 156.235 178.145 ;
        RECT 154.860 177.425 155.085 177.465 ;
        RECT 156.405 177.435 156.925 177.975 ;
        RECT 151.760 176.965 152.165 177.135 ;
        RECT 152.335 176.965 153.120 177.135 ;
        RECT 153.395 176.685 153.605 177.215 ;
        RECT 153.865 176.900 154.195 177.425 ;
        RECT 154.705 177.340 155.085 177.425 ;
        RECT 154.365 176.685 154.535 177.295 ;
        RECT 154.705 176.905 155.035 177.340 ;
        RECT 155.715 176.685 156.925 177.435 ;
        RECT 22.690 176.515 157.010 176.685 ;
        RECT 22.775 175.765 23.985 176.515 ;
        RECT 25.075 175.840 25.335 176.345 ;
        RECT 25.515 176.135 25.845 176.515 ;
        RECT 26.025 175.965 26.195 176.345 ;
        RECT 22.775 175.225 23.295 175.765 ;
        RECT 23.465 175.055 23.985 175.595 ;
        RECT 22.775 173.965 23.985 175.055 ;
        RECT 25.075 175.040 25.245 175.840 ;
        RECT 25.530 175.795 26.195 175.965 ;
        RECT 25.530 175.540 25.700 175.795 ;
        RECT 26.455 175.745 28.125 176.515 ;
        RECT 28.495 175.885 28.825 176.245 ;
        RECT 29.445 176.055 29.695 176.515 ;
        RECT 29.865 176.055 30.425 176.345 ;
        RECT 25.415 175.210 25.700 175.540 ;
        RECT 25.935 175.245 26.265 175.615 ;
        RECT 26.455 175.225 27.205 175.745 ;
        RECT 28.495 175.695 29.885 175.885 ;
        RECT 29.715 175.605 29.885 175.695 ;
        RECT 25.530 175.065 25.700 175.210 ;
        RECT 25.075 174.135 25.345 175.040 ;
        RECT 25.530 174.895 26.195 175.065 ;
        RECT 27.375 175.055 28.125 175.575 ;
        RECT 25.515 173.965 25.845 174.725 ;
        RECT 26.025 174.135 26.195 174.895 ;
        RECT 26.455 173.965 28.125 175.055 ;
        RECT 28.310 175.275 28.985 175.525 ;
        RECT 29.205 175.275 29.545 175.525 ;
        RECT 29.715 175.275 30.005 175.605 ;
        RECT 28.310 174.915 28.575 175.275 ;
        RECT 29.715 175.025 29.885 175.275 ;
        RECT 28.945 174.855 29.885 175.025 ;
        RECT 28.495 173.965 28.775 174.635 ;
        RECT 28.945 174.305 29.245 174.855 ;
        RECT 30.175 174.685 30.425 176.055 ;
        RECT 30.595 175.695 30.855 176.515 ;
        RECT 31.025 175.695 31.355 176.115 ;
        RECT 31.535 176.030 32.325 176.295 ;
        RECT 31.105 175.605 31.355 175.695 ;
        RECT 29.445 173.965 29.775 174.685 ;
        RECT 29.965 174.135 30.425 174.685 ;
        RECT 30.595 174.645 30.935 175.525 ;
        RECT 31.105 175.355 31.900 175.605 ;
        RECT 30.595 173.965 30.855 174.475 ;
        RECT 31.105 174.135 31.275 175.355 ;
        RECT 32.070 175.175 32.325 176.030 ;
        RECT 32.495 175.875 32.695 176.295 ;
        RECT 32.885 176.055 33.215 176.515 ;
        RECT 32.495 175.355 32.905 175.875 ;
        RECT 33.385 175.865 33.645 176.345 ;
        RECT 33.075 175.175 33.305 175.605 ;
        RECT 31.515 175.005 33.305 175.175 ;
        RECT 31.515 174.640 31.765 175.005 ;
        RECT 31.935 174.645 32.265 174.835 ;
        RECT 32.485 174.710 33.200 175.005 ;
        RECT 33.475 174.835 33.645 175.865 ;
        RECT 31.935 174.470 32.130 174.645 ;
        RECT 31.515 173.965 32.130 174.470 ;
        RECT 32.300 174.135 32.775 174.475 ;
        RECT 32.945 173.965 33.160 174.510 ;
        RECT 33.370 174.135 33.645 174.835 ;
        RECT 33.850 175.775 34.465 176.345 ;
        RECT 34.635 176.005 34.850 176.515 ;
        RECT 35.080 176.005 35.360 176.335 ;
        RECT 35.540 176.005 35.780 176.515 ;
        RECT 33.850 174.755 34.165 175.775 ;
        RECT 34.335 175.105 34.505 175.605 ;
        RECT 34.755 175.275 35.020 175.835 ;
        RECT 35.190 175.105 35.360 176.005 ;
        RECT 36.205 175.965 36.375 176.255 ;
        RECT 36.545 176.135 36.875 176.515 ;
        RECT 35.530 175.275 35.885 175.835 ;
        RECT 36.205 175.795 36.870 175.965 ;
        RECT 34.335 174.935 35.760 175.105 ;
        RECT 36.120 174.975 36.470 175.625 ;
        RECT 33.850 174.135 34.385 174.755 ;
        RECT 34.555 173.965 34.885 174.765 ;
        RECT 35.370 174.760 35.760 174.935 ;
        RECT 36.640 174.805 36.870 175.795 ;
        RECT 36.205 174.635 36.870 174.805 ;
        RECT 36.205 174.135 36.375 174.635 ;
        RECT 36.545 173.965 36.875 174.465 ;
        RECT 37.045 174.135 37.230 176.255 ;
        RECT 37.485 176.055 37.735 176.515 ;
        RECT 37.905 176.065 38.240 176.235 ;
        RECT 38.435 176.065 39.110 176.235 ;
        RECT 37.905 175.925 38.075 176.065 ;
        RECT 37.400 174.935 37.680 175.885 ;
        RECT 37.850 175.795 38.075 175.925 ;
        RECT 37.850 174.690 38.020 175.795 ;
        RECT 38.245 175.645 38.770 175.865 ;
        RECT 38.190 174.880 38.430 175.475 ;
        RECT 38.600 174.945 38.770 175.645 ;
        RECT 38.940 175.285 39.110 176.065 ;
        RECT 39.430 176.015 39.800 176.515 ;
        RECT 39.980 176.065 40.385 176.235 ;
        RECT 40.555 176.065 41.340 176.235 ;
        RECT 39.980 175.835 40.150 176.065 ;
        RECT 39.320 175.535 40.150 175.835 ;
        RECT 40.535 175.565 41.000 175.895 ;
        RECT 39.320 175.505 39.520 175.535 ;
        RECT 39.640 175.285 39.810 175.355 ;
        RECT 38.940 175.115 39.810 175.285 ;
        RECT 39.300 175.025 39.810 175.115 ;
        RECT 37.850 174.560 38.155 174.690 ;
        RECT 38.600 174.580 39.130 174.945 ;
        RECT 37.470 173.965 37.735 174.425 ;
        RECT 37.905 174.135 38.155 174.560 ;
        RECT 39.300 174.410 39.470 175.025 ;
        RECT 38.365 174.240 39.470 174.410 ;
        RECT 39.640 173.965 39.810 174.765 ;
        RECT 39.980 174.465 40.150 175.535 ;
        RECT 40.320 174.635 40.510 175.355 ;
        RECT 40.680 174.605 41.000 175.565 ;
        RECT 41.170 175.605 41.340 176.065 ;
        RECT 41.615 175.985 41.825 176.515 ;
        RECT 42.085 175.775 42.415 176.300 ;
        RECT 42.585 175.905 42.755 176.515 ;
        RECT 42.925 175.860 43.255 176.295 ;
        RECT 42.925 175.775 43.305 175.860 ;
        RECT 42.215 175.605 42.415 175.775 ;
        RECT 43.080 175.735 43.305 175.775 ;
        RECT 41.170 175.275 42.045 175.605 ;
        RECT 42.215 175.275 42.965 175.605 ;
        RECT 39.980 174.135 40.230 174.465 ;
        RECT 41.170 174.435 41.340 175.275 ;
        RECT 42.215 175.070 42.405 175.275 ;
        RECT 43.135 175.155 43.305 175.735 ;
        RECT 44.435 175.695 44.665 176.515 ;
        RECT 44.835 175.715 45.165 176.345 ;
        RECT 44.415 175.275 44.745 175.525 ;
        RECT 43.090 175.105 43.305 175.155 ;
        RECT 44.915 175.115 45.165 175.715 ;
        RECT 45.335 175.695 45.545 176.515 ;
        RECT 45.775 176.015 46.075 176.345 ;
        RECT 46.245 176.035 46.520 176.515 ;
        RECT 41.510 174.695 42.405 175.070 ;
        RECT 42.915 175.025 43.305 175.105 ;
        RECT 40.455 174.265 41.340 174.435 ;
        RECT 41.520 173.965 41.835 174.465 ;
        RECT 42.065 174.135 42.405 174.695 ;
        RECT 42.575 173.965 42.745 174.975 ;
        RECT 42.915 174.180 43.245 175.025 ;
        RECT 44.435 173.965 44.665 175.105 ;
        RECT 44.835 174.135 45.165 175.115 ;
        RECT 45.775 175.105 45.945 176.015 ;
        RECT 46.700 175.865 46.995 176.255 ;
        RECT 47.165 176.035 47.420 176.515 ;
        RECT 47.595 175.865 47.855 176.255 ;
        RECT 48.025 176.035 48.305 176.515 ;
        RECT 46.115 175.275 46.465 175.845 ;
        RECT 46.700 175.695 48.350 175.865 ;
        RECT 48.535 175.790 48.825 176.515 ;
        RECT 46.635 175.355 47.775 175.525 ;
        RECT 46.635 175.105 46.805 175.355 ;
        RECT 47.945 175.185 48.350 175.695 ;
        RECT 45.335 173.965 45.545 175.105 ;
        RECT 45.775 174.935 46.805 175.105 ;
        RECT 47.595 175.015 48.350 175.185 ;
        RECT 45.775 174.135 46.085 174.935 ;
        RECT 47.595 174.765 47.855 175.015 ;
        RECT 46.255 173.965 46.565 174.765 ;
        RECT 46.735 174.595 47.855 174.765 ;
        RECT 46.735 174.135 46.995 174.595 ;
        RECT 47.165 173.965 47.420 174.425 ;
        RECT 47.595 174.135 47.855 174.595 ;
        RECT 48.025 173.965 48.310 174.835 ;
        RECT 48.535 173.965 48.825 175.130 ;
        RECT 49.915 174.135 50.195 176.235 ;
        RECT 50.425 176.055 50.595 176.515 ;
        RECT 50.865 176.125 52.115 176.305 ;
        RECT 51.250 175.885 51.615 175.955 ;
        RECT 50.365 175.705 51.615 175.885 ;
        RECT 51.785 175.905 52.115 176.125 ;
        RECT 52.285 176.075 52.455 176.515 ;
        RECT 52.625 175.905 52.965 176.320 ;
        RECT 51.785 175.735 52.965 175.905 ;
        RECT 50.365 175.105 50.640 175.705 ;
        RECT 53.135 175.695 53.820 176.335 ;
        RECT 53.990 175.695 54.160 176.515 ;
        RECT 54.330 175.865 54.660 176.330 ;
        RECT 54.830 176.045 55.000 176.515 ;
        RECT 55.260 176.125 56.445 176.295 ;
        RECT 56.615 175.955 56.945 176.345 ;
        RECT 55.645 175.865 56.030 175.955 ;
        RECT 54.330 175.695 56.030 175.865 ;
        RECT 56.435 175.775 56.945 175.955 ;
        RECT 57.275 175.775 57.615 176.345 ;
        RECT 57.810 175.850 57.980 176.515 ;
        RECT 58.260 176.175 58.480 176.220 ;
        RECT 58.255 176.005 58.480 176.175 ;
        RECT 58.650 176.035 59.095 176.205 ;
        RECT 58.260 175.865 58.480 176.005 ;
        RECT 50.810 175.275 51.165 175.525 ;
        RECT 51.360 175.495 51.825 175.525 ;
        RECT 51.355 175.325 51.825 175.495 ;
        RECT 51.360 175.275 51.825 175.325 ;
        RECT 51.995 175.275 52.325 175.525 ;
        RECT 52.500 175.325 52.965 175.525 ;
        RECT 52.145 175.155 52.325 175.275 ;
        RECT 50.365 174.895 51.975 175.105 ;
        RECT 52.145 174.985 52.475 175.155 ;
        RECT 51.565 174.795 51.975 174.895 ;
        RECT 50.385 173.965 51.170 174.725 ;
        RECT 51.565 174.135 51.950 174.795 ;
        RECT 52.275 174.195 52.475 174.985 ;
        RECT 52.645 173.965 52.965 175.145 ;
        RECT 53.135 174.725 53.385 175.695 ;
        RECT 53.555 175.315 53.890 175.525 ;
        RECT 54.060 175.315 54.510 175.525 ;
        RECT 54.700 175.495 55.185 175.525 ;
        RECT 54.700 175.325 55.205 175.495 ;
        RECT 54.700 175.315 55.185 175.325 ;
        RECT 53.720 175.145 53.890 175.315 ;
        RECT 53.720 174.975 54.640 175.145 ;
        RECT 53.135 174.135 53.800 174.725 ;
        RECT 53.970 173.965 54.300 174.805 ;
        RECT 54.470 174.725 54.640 174.975 ;
        RECT 54.810 174.895 55.185 175.315 ;
        RECT 55.375 175.275 55.755 175.525 ;
        RECT 55.935 175.315 56.265 175.525 ;
        RECT 55.375 174.895 55.695 175.275 ;
        RECT 56.435 175.145 56.605 175.775 ;
        RECT 56.775 175.315 57.105 175.605 ;
        RECT 55.865 174.975 56.950 175.145 ;
        RECT 55.865 174.725 56.035 174.975 ;
        RECT 54.470 174.555 56.035 174.725 ;
        RECT 54.810 174.135 55.615 174.555 ;
        RECT 56.205 173.965 56.455 174.805 ;
        RECT 56.650 174.135 56.950 174.975 ;
        RECT 57.275 174.805 57.450 175.775 ;
        RECT 58.260 175.695 58.755 175.865 ;
        RECT 57.620 175.155 57.790 175.605 ;
        RECT 57.960 175.325 58.410 175.525 ;
        RECT 58.580 175.500 58.755 175.695 ;
        RECT 58.925 175.245 59.095 176.035 ;
        RECT 59.265 175.910 59.515 176.280 ;
        RECT 59.345 175.525 59.515 175.910 ;
        RECT 59.685 175.875 59.935 176.280 ;
        RECT 60.105 176.045 60.275 176.515 ;
        RECT 60.445 175.875 60.785 176.280 ;
        RECT 59.685 175.695 60.785 175.875 ;
        RECT 60.955 175.715 61.650 176.345 ;
        RECT 61.855 175.715 62.165 176.515 ;
        RECT 63.255 176.015 63.515 176.345 ;
        RECT 63.685 176.155 64.015 176.515 ;
        RECT 64.270 176.135 65.570 176.345 ;
        RECT 63.255 176.005 63.485 176.015 ;
        RECT 59.345 175.355 59.540 175.525 ;
        RECT 57.620 174.985 58.015 175.155 ;
        RECT 58.925 175.105 59.200 175.245 ;
        RECT 57.275 174.135 57.535 174.805 ;
        RECT 57.845 174.715 58.015 174.985 ;
        RECT 58.185 174.885 59.200 175.105 ;
        RECT 59.370 175.105 59.540 175.355 ;
        RECT 59.710 175.275 60.270 175.525 ;
        RECT 59.370 174.715 59.925 175.105 ;
        RECT 57.845 174.545 59.925 174.715 ;
        RECT 57.705 173.965 58.035 174.365 ;
        RECT 58.905 173.965 59.305 174.365 ;
        RECT 59.595 174.310 59.925 174.545 ;
        RECT 60.095 174.175 60.270 175.275 ;
        RECT 60.440 174.955 60.785 175.525 ;
        RECT 60.975 175.275 61.310 175.525 ;
        RECT 61.480 175.115 61.650 175.715 ;
        RECT 61.820 175.275 62.155 175.545 ;
        RECT 60.440 173.965 60.785 174.785 ;
        RECT 60.955 173.965 61.215 175.105 ;
        RECT 61.385 174.135 61.715 175.115 ;
        RECT 61.885 173.965 62.165 175.105 ;
        RECT 63.255 174.815 63.425 176.005 ;
        RECT 64.270 175.985 64.440 176.135 ;
        RECT 63.685 175.860 64.440 175.985 ;
        RECT 63.595 175.815 64.440 175.860 ;
        RECT 63.595 175.695 63.865 175.815 ;
        RECT 63.595 175.120 63.765 175.695 ;
        RECT 63.995 175.255 64.405 175.560 ;
        RECT 64.695 175.525 64.905 175.925 ;
        RECT 64.575 175.315 64.905 175.525 ;
        RECT 65.150 175.525 65.370 175.925 ;
        RECT 65.845 175.750 66.300 176.515 ;
        RECT 66.985 175.860 67.315 176.295 ;
        RECT 67.485 175.905 67.655 176.515 ;
        RECT 66.935 175.775 67.315 175.860 ;
        RECT 67.825 175.775 68.155 176.300 ;
        RECT 68.415 175.985 68.625 176.515 ;
        RECT 68.900 176.065 69.685 176.235 ;
        RECT 69.855 176.065 70.260 176.235 ;
        RECT 66.935 175.735 67.160 175.775 ;
        RECT 65.150 175.315 65.625 175.525 ;
        RECT 65.815 175.325 66.305 175.525 ;
        RECT 66.935 175.155 67.105 175.735 ;
        RECT 67.825 175.605 68.025 175.775 ;
        RECT 68.900 175.605 69.070 176.065 ;
        RECT 67.275 175.275 68.025 175.605 ;
        RECT 68.195 175.275 69.070 175.605 ;
        RECT 63.595 175.085 63.795 175.120 ;
        RECT 65.125 175.085 66.300 175.145 ;
        RECT 63.595 174.975 66.300 175.085 ;
        RECT 66.935 175.105 67.150 175.155 ;
        RECT 66.935 175.025 67.325 175.105 ;
        RECT 63.655 174.915 65.455 174.975 ;
        RECT 65.125 174.885 65.455 174.915 ;
        RECT 63.255 174.135 63.515 174.815 ;
        RECT 63.685 173.965 63.935 174.745 ;
        RECT 64.185 174.715 65.020 174.725 ;
        RECT 65.610 174.715 65.795 174.805 ;
        RECT 64.185 174.515 65.795 174.715 ;
        RECT 64.185 174.135 64.435 174.515 ;
        RECT 65.565 174.475 65.795 174.515 ;
        RECT 66.045 174.355 66.300 174.975 ;
        RECT 64.605 173.965 64.960 174.345 ;
        RECT 65.965 174.135 66.300 174.355 ;
        RECT 66.995 174.180 67.325 175.025 ;
        RECT 67.835 175.070 68.025 175.275 ;
        RECT 67.495 173.965 67.665 174.975 ;
        RECT 67.835 174.695 68.730 175.070 ;
        RECT 67.835 174.135 68.175 174.695 ;
        RECT 68.405 173.965 68.720 174.465 ;
        RECT 68.900 174.435 69.070 175.275 ;
        RECT 69.240 175.565 69.705 175.895 ;
        RECT 70.090 175.835 70.260 176.065 ;
        RECT 70.440 176.015 70.810 176.515 ;
        RECT 71.130 176.065 71.805 176.235 ;
        RECT 72.000 176.065 72.335 176.235 ;
        RECT 69.240 174.605 69.560 175.565 ;
        RECT 70.090 175.535 70.920 175.835 ;
        RECT 69.730 174.635 69.920 175.355 ;
        RECT 70.090 174.465 70.260 175.535 ;
        RECT 70.720 175.505 70.920 175.535 ;
        RECT 70.430 175.285 70.600 175.355 ;
        RECT 71.130 175.285 71.300 176.065 ;
        RECT 72.165 175.925 72.335 176.065 ;
        RECT 72.505 176.055 72.755 176.515 ;
        RECT 70.430 175.115 71.300 175.285 ;
        RECT 71.470 175.645 71.995 175.865 ;
        RECT 72.165 175.795 72.390 175.925 ;
        RECT 70.430 175.025 70.940 175.115 ;
        RECT 68.900 174.265 69.785 174.435 ;
        RECT 70.010 174.135 70.260 174.465 ;
        RECT 70.430 173.965 70.600 174.765 ;
        RECT 70.770 174.410 70.940 175.025 ;
        RECT 71.470 174.945 71.640 175.645 ;
        RECT 71.110 174.580 71.640 174.945 ;
        RECT 71.810 174.880 72.050 175.475 ;
        RECT 72.220 174.690 72.390 175.795 ;
        RECT 72.560 174.935 72.840 175.885 ;
        RECT 72.085 174.560 72.390 174.690 ;
        RECT 70.770 174.240 71.875 174.410 ;
        RECT 72.085 174.135 72.335 174.560 ;
        RECT 72.505 173.965 72.770 174.425 ;
        RECT 73.010 174.135 73.195 176.255 ;
        RECT 73.365 176.135 73.695 176.515 ;
        RECT 73.865 175.965 74.035 176.255 ;
        RECT 73.370 175.795 74.035 175.965 ;
        RECT 73.370 174.805 73.600 175.795 ;
        RECT 74.295 175.790 74.585 176.515 ;
        RECT 74.755 175.775 75.140 176.345 ;
        RECT 75.310 176.055 75.635 176.515 ;
        RECT 76.155 175.885 76.435 176.345 ;
        RECT 73.770 174.975 74.120 175.625 ;
        RECT 73.370 174.635 74.035 174.805 ;
        RECT 73.365 173.965 73.695 174.465 ;
        RECT 73.865 174.135 74.035 174.635 ;
        RECT 74.295 173.965 74.585 175.130 ;
        RECT 74.755 175.105 75.035 175.775 ;
        RECT 75.310 175.715 76.435 175.885 ;
        RECT 75.310 175.605 75.760 175.715 ;
        RECT 75.205 175.275 75.760 175.605 ;
        RECT 76.625 175.545 77.025 176.345 ;
        RECT 77.425 176.055 77.695 176.515 ;
        RECT 77.865 175.885 78.150 176.345 ;
        RECT 74.755 174.135 75.140 175.105 ;
        RECT 75.310 174.815 75.760 175.275 ;
        RECT 75.930 174.985 77.025 175.545 ;
        RECT 75.310 174.595 76.435 174.815 ;
        RECT 75.310 173.965 75.635 174.425 ;
        RECT 76.155 174.135 76.435 174.595 ;
        RECT 76.625 174.135 77.025 174.985 ;
        RECT 77.195 175.715 78.150 175.885 ;
        RECT 78.435 176.015 78.695 176.345 ;
        RECT 78.865 176.155 79.195 176.515 ;
        RECT 79.450 176.135 80.750 176.345 ;
        RECT 78.435 176.005 78.665 176.015 ;
        RECT 77.195 174.815 77.405 175.715 ;
        RECT 77.575 174.985 78.265 175.545 ;
        RECT 78.435 174.815 78.605 176.005 ;
        RECT 79.450 175.985 79.620 176.135 ;
        RECT 78.865 175.860 79.620 175.985 ;
        RECT 78.775 175.815 79.620 175.860 ;
        RECT 78.775 175.695 79.045 175.815 ;
        RECT 78.775 175.120 78.945 175.695 ;
        RECT 79.175 175.255 79.585 175.560 ;
        RECT 79.875 175.525 80.085 175.925 ;
        RECT 79.755 175.315 80.085 175.525 ;
        RECT 80.330 175.525 80.550 175.925 ;
        RECT 81.025 175.750 81.480 176.515 ;
        RECT 82.635 175.695 82.845 176.515 ;
        RECT 83.015 175.715 83.345 176.345 ;
        RECT 80.330 175.315 80.805 175.525 ;
        RECT 80.995 175.325 81.485 175.525 ;
        RECT 78.775 175.085 78.975 175.120 ;
        RECT 80.305 175.085 81.480 175.145 ;
        RECT 83.015 175.115 83.265 175.715 ;
        RECT 83.515 175.695 83.745 176.515 ;
        RECT 83.955 175.715 84.650 176.345 ;
        RECT 84.855 175.715 85.165 176.515 ;
        RECT 85.335 175.865 85.595 176.345 ;
        RECT 85.765 176.055 86.095 176.515 ;
        RECT 86.285 175.875 86.485 176.295 ;
        RECT 84.475 175.665 84.650 175.715 ;
        RECT 83.435 175.275 83.765 175.525 ;
        RECT 83.975 175.275 84.310 175.525 ;
        RECT 84.480 175.115 84.650 175.665 ;
        RECT 84.820 175.275 85.155 175.545 ;
        RECT 78.775 174.975 81.480 175.085 ;
        RECT 78.835 174.915 80.635 174.975 ;
        RECT 80.305 174.885 80.635 174.915 ;
        RECT 77.195 174.595 78.150 174.815 ;
        RECT 77.425 173.965 77.695 174.425 ;
        RECT 77.865 174.135 78.150 174.595 ;
        RECT 78.435 174.135 78.695 174.815 ;
        RECT 78.865 173.965 79.115 174.745 ;
        RECT 79.365 174.715 80.200 174.725 ;
        RECT 80.790 174.715 80.975 174.805 ;
        RECT 79.365 174.515 80.975 174.715 ;
        RECT 79.365 174.135 79.615 174.515 ;
        RECT 80.745 174.475 80.975 174.515 ;
        RECT 81.225 174.355 81.480 174.975 ;
        RECT 79.785 173.965 80.140 174.345 ;
        RECT 81.145 174.135 81.480 174.355 ;
        RECT 82.635 173.965 82.845 175.105 ;
        RECT 83.015 174.135 83.345 175.115 ;
        RECT 83.515 173.965 83.745 175.105 ;
        RECT 83.955 173.965 84.215 175.105 ;
        RECT 84.385 174.135 84.715 175.115 ;
        RECT 84.885 173.965 85.165 175.105 ;
        RECT 85.335 174.835 85.505 175.865 ;
        RECT 85.675 175.175 85.905 175.605 ;
        RECT 86.075 175.355 86.485 175.875 ;
        RECT 86.655 176.030 87.445 176.295 ;
        RECT 86.655 175.175 86.910 176.030 ;
        RECT 87.625 175.695 87.955 176.115 ;
        RECT 88.125 175.695 88.385 176.515 ;
        RECT 88.555 176.135 89.445 176.305 ;
        RECT 87.625 175.605 87.875 175.695 ;
        RECT 87.080 175.355 87.875 175.605 ;
        RECT 88.555 175.580 89.105 175.965 ;
        RECT 85.675 175.005 87.465 175.175 ;
        RECT 85.335 174.135 85.610 174.835 ;
        RECT 85.780 174.710 86.495 175.005 ;
        RECT 86.715 174.645 87.045 174.835 ;
        RECT 85.820 173.965 86.035 174.510 ;
        RECT 86.205 174.135 86.680 174.475 ;
        RECT 86.850 174.470 87.045 174.645 ;
        RECT 87.215 174.640 87.465 175.005 ;
        RECT 86.850 173.965 87.465 174.470 ;
        RECT 87.705 174.135 87.875 175.355 ;
        RECT 88.045 174.645 88.385 175.525 ;
        RECT 89.275 175.410 89.445 176.135 ;
        RECT 88.555 175.340 89.445 175.410 ;
        RECT 89.615 175.810 89.835 176.295 ;
        RECT 90.005 175.975 90.255 176.515 ;
        RECT 90.425 175.865 90.685 176.345 ;
        RECT 90.860 176.010 91.195 176.515 ;
        RECT 91.365 175.945 91.605 176.320 ;
        RECT 91.885 176.185 92.055 176.330 ;
        RECT 91.885 175.990 92.260 176.185 ;
        RECT 92.620 176.020 93.015 176.515 ;
        RECT 89.615 175.385 89.945 175.810 ;
        RECT 88.555 175.315 89.450 175.340 ;
        RECT 88.555 175.300 89.460 175.315 ;
        RECT 88.555 175.285 89.465 175.300 ;
        RECT 88.555 175.280 89.475 175.285 ;
        RECT 88.555 175.270 89.480 175.280 ;
        RECT 88.555 175.260 89.485 175.270 ;
        RECT 88.555 175.255 89.495 175.260 ;
        RECT 88.555 175.245 89.505 175.255 ;
        RECT 88.555 175.240 89.515 175.245 ;
        RECT 88.555 174.790 88.815 175.240 ;
        RECT 89.180 175.235 89.515 175.240 ;
        RECT 89.180 175.230 89.530 175.235 ;
        RECT 89.180 175.220 89.545 175.230 ;
        RECT 89.180 175.215 89.570 175.220 ;
        RECT 90.115 175.215 90.345 175.610 ;
        RECT 89.180 175.210 90.345 175.215 ;
        RECT 89.210 175.175 90.345 175.210 ;
        RECT 89.245 175.150 90.345 175.175 ;
        RECT 89.275 175.120 90.345 175.150 ;
        RECT 89.295 175.090 90.345 175.120 ;
        RECT 89.315 175.060 90.345 175.090 ;
        RECT 89.385 175.050 90.345 175.060 ;
        RECT 89.410 175.040 90.345 175.050 ;
        RECT 89.430 175.025 90.345 175.040 ;
        RECT 89.450 175.010 90.345 175.025 ;
        RECT 89.455 175.000 90.240 175.010 ;
        RECT 89.470 174.965 90.240 175.000 ;
        RECT 88.985 174.645 89.315 174.890 ;
        RECT 89.485 174.715 90.240 174.965 ;
        RECT 90.515 174.835 90.685 175.865 ;
        RECT 90.915 174.985 91.215 175.835 ;
        RECT 91.385 175.795 91.605 175.945 ;
        RECT 91.385 175.465 91.920 175.795 ;
        RECT 92.090 175.655 92.260 175.990 ;
        RECT 93.185 175.825 93.425 176.345 ;
        RECT 88.985 174.620 89.170 174.645 ;
        RECT 88.555 174.520 89.170 174.620 ;
        RECT 88.125 173.965 88.385 174.475 ;
        RECT 88.555 173.965 89.160 174.520 ;
        RECT 89.335 174.135 89.815 174.475 ;
        RECT 89.985 173.965 90.240 174.510 ;
        RECT 90.410 174.135 90.685 174.835 ;
        RECT 91.385 174.815 91.620 175.465 ;
        RECT 92.090 175.295 93.075 175.655 ;
        RECT 90.945 174.585 91.620 174.815 ;
        RECT 91.790 175.275 93.075 175.295 ;
        RECT 91.790 175.125 92.650 175.275 ;
        RECT 90.945 174.155 91.115 174.585 ;
        RECT 91.285 173.965 91.615 174.415 ;
        RECT 91.790 174.180 92.075 175.125 ;
        RECT 93.250 175.020 93.425 175.825 ;
        RECT 93.615 175.895 93.880 176.345 ;
        RECT 94.050 176.065 94.340 176.515 ;
        RECT 94.510 175.895 94.800 176.345 ;
        RECT 93.615 175.725 94.800 175.895 ;
        RECT 94.980 175.605 95.225 176.210 ;
        RECT 92.250 174.645 92.945 174.955 ;
        RECT 92.255 173.965 92.940 174.435 ;
        RECT 93.120 174.235 93.425 175.020 ;
        RECT 93.635 174.940 93.965 175.525 ;
        RECT 94.135 175.275 94.620 175.525 ;
        RECT 94.965 175.275 95.225 175.605 ;
        RECT 95.475 175.275 95.745 176.210 ;
        RECT 95.925 175.525 96.135 176.210 ;
        RECT 96.305 175.865 96.645 176.345 ;
        RECT 96.825 176.035 97.135 176.515 ;
        RECT 96.305 175.695 96.975 175.865 ;
        RECT 96.805 175.605 96.975 175.695 ;
        RECT 95.925 175.275 96.405 175.525 ;
        RECT 96.805 175.275 97.145 175.605 ;
        RECT 93.615 173.965 93.940 174.765 ;
        RECT 94.135 174.185 94.320 175.275 ;
        RECT 96.805 175.105 96.975 175.275 ;
        RECT 94.490 174.935 96.975 175.105 ;
        RECT 94.490 174.135 94.740 174.935 ;
        RECT 94.910 173.965 95.650 174.765 ;
        RECT 95.835 174.135 96.165 174.935 ;
        RECT 96.335 173.965 97.145 174.765 ;
        RECT 97.315 174.135 97.575 176.345 ;
        RECT 97.795 175.695 98.025 176.515 ;
        RECT 98.195 175.715 98.525 176.345 ;
        RECT 97.775 175.275 98.105 175.525 ;
        RECT 98.275 175.115 98.525 175.715 ;
        RECT 98.695 175.695 98.905 176.515 ;
        RECT 100.055 175.790 100.345 176.515 ;
        RECT 100.525 175.785 100.825 176.515 ;
        RECT 101.005 175.605 101.235 176.225 ;
        RECT 101.435 175.955 101.660 176.335 ;
        RECT 101.830 176.125 102.160 176.515 ;
        RECT 102.815 176.015 103.075 176.345 ;
        RECT 103.245 176.155 103.575 176.515 ;
        RECT 103.830 176.135 105.130 176.345 ;
        RECT 102.815 176.005 103.045 176.015 ;
        RECT 101.435 175.775 101.765 175.955 ;
        RECT 100.530 175.275 100.825 175.605 ;
        RECT 101.005 175.275 101.420 175.605 ;
        RECT 97.795 173.965 98.025 175.105 ;
        RECT 98.195 174.135 98.525 175.115 ;
        RECT 98.695 173.965 98.905 175.105 ;
        RECT 100.055 173.965 100.345 175.130 ;
        RECT 101.590 175.105 101.765 175.775 ;
        RECT 101.935 175.275 102.175 175.925 ;
        RECT 100.525 174.745 101.420 175.075 ;
        RECT 101.590 174.915 102.175 175.105 ;
        RECT 100.525 174.575 101.730 174.745 ;
        RECT 100.525 174.145 100.855 174.575 ;
        RECT 101.035 173.965 101.230 174.405 ;
        RECT 101.400 174.145 101.730 174.575 ;
        RECT 101.900 174.145 102.175 174.915 ;
        RECT 102.815 174.815 102.985 176.005 ;
        RECT 103.830 175.985 104.000 176.135 ;
        RECT 103.245 175.860 104.000 175.985 ;
        RECT 103.155 175.815 104.000 175.860 ;
        RECT 103.155 175.695 103.425 175.815 ;
        RECT 103.155 175.120 103.325 175.695 ;
        RECT 103.555 175.255 103.965 175.560 ;
        RECT 104.255 175.525 104.465 175.925 ;
        RECT 104.135 175.315 104.465 175.525 ;
        RECT 104.710 175.525 104.930 175.925 ;
        RECT 105.405 175.750 105.860 176.515 ;
        RECT 106.035 175.715 106.375 176.345 ;
        RECT 106.545 175.715 106.795 176.515 ;
        RECT 106.985 175.865 107.315 176.345 ;
        RECT 107.485 176.055 107.710 176.515 ;
        RECT 107.880 175.865 108.210 176.345 ;
        RECT 104.710 175.315 105.185 175.525 ;
        RECT 105.375 175.325 105.865 175.525 ;
        RECT 103.155 175.085 103.355 175.120 ;
        RECT 104.685 175.085 105.860 175.145 ;
        RECT 103.155 174.975 105.860 175.085 ;
        RECT 103.215 174.915 105.015 174.975 ;
        RECT 104.685 174.885 105.015 174.915 ;
        RECT 102.815 174.135 103.075 174.815 ;
        RECT 103.245 173.965 103.495 174.745 ;
        RECT 103.745 174.715 104.580 174.725 ;
        RECT 105.170 174.715 105.355 174.805 ;
        RECT 103.745 174.515 105.355 174.715 ;
        RECT 103.745 174.135 103.995 174.515 ;
        RECT 105.125 174.475 105.355 174.515 ;
        RECT 105.605 174.355 105.860 174.975 ;
        RECT 104.165 173.965 104.520 174.345 ;
        RECT 105.525 174.135 105.860 174.355 ;
        RECT 106.035 175.105 106.210 175.715 ;
        RECT 106.985 175.695 108.210 175.865 ;
        RECT 108.840 175.735 109.340 176.345 ;
        RECT 110.175 175.775 110.515 176.345 ;
        RECT 110.710 175.850 110.880 176.515 ;
        RECT 111.160 176.175 111.380 176.220 ;
        RECT 111.155 176.005 111.380 176.175 ;
        RECT 111.550 176.035 111.995 176.205 ;
        RECT 111.160 175.865 111.380 176.005 ;
        RECT 106.380 175.355 107.075 175.525 ;
        RECT 106.905 175.105 107.075 175.355 ;
        RECT 107.250 175.325 107.670 175.525 ;
        RECT 107.840 175.325 108.170 175.525 ;
        RECT 108.340 175.325 108.670 175.525 ;
        RECT 108.840 175.105 109.010 175.735 ;
        RECT 109.195 175.275 109.545 175.525 ;
        RECT 106.035 174.135 106.375 175.105 ;
        RECT 106.545 173.965 106.715 175.105 ;
        RECT 106.905 174.935 109.340 175.105 ;
        RECT 106.985 173.965 107.235 174.765 ;
        RECT 107.880 174.135 108.210 174.935 ;
        RECT 108.510 173.965 108.840 174.765 ;
        RECT 109.010 174.135 109.340 174.935 ;
        RECT 110.175 174.805 110.350 175.775 ;
        RECT 111.160 175.695 111.655 175.865 ;
        RECT 110.520 175.155 110.690 175.605 ;
        RECT 110.860 175.325 111.310 175.525 ;
        RECT 111.480 175.500 111.655 175.695 ;
        RECT 111.825 175.245 111.995 176.035 ;
        RECT 112.165 175.910 112.415 176.280 ;
        RECT 112.245 175.525 112.415 175.910 ;
        RECT 112.585 175.875 112.835 176.280 ;
        RECT 113.005 176.045 113.175 176.515 ;
        RECT 113.345 175.875 113.685 176.280 ;
        RECT 112.585 175.695 113.685 175.875 ;
        RECT 114.335 175.825 114.575 176.345 ;
        RECT 114.745 176.020 115.140 176.515 ;
        RECT 115.705 176.185 115.875 176.330 ;
        RECT 115.500 175.990 115.875 176.185 ;
        RECT 112.245 175.355 112.440 175.525 ;
        RECT 110.520 174.985 110.915 175.155 ;
        RECT 111.825 175.105 112.100 175.245 ;
        RECT 110.175 174.135 110.435 174.805 ;
        RECT 110.745 174.715 110.915 174.985 ;
        RECT 111.085 174.885 112.100 175.105 ;
        RECT 112.270 175.105 112.440 175.355 ;
        RECT 112.610 175.275 113.170 175.525 ;
        RECT 112.270 174.715 112.825 175.105 ;
        RECT 110.745 174.545 112.825 174.715 ;
        RECT 110.605 173.965 110.935 174.365 ;
        RECT 111.805 173.965 112.205 174.365 ;
        RECT 112.495 174.310 112.825 174.545 ;
        RECT 112.995 174.175 113.170 175.275 ;
        RECT 113.340 174.955 113.685 175.525 ;
        RECT 114.335 175.020 114.510 175.825 ;
        RECT 115.500 175.655 115.670 175.990 ;
        RECT 116.155 175.945 116.395 176.320 ;
        RECT 116.565 176.010 116.900 176.515 ;
        RECT 116.155 175.795 116.375 175.945 ;
        RECT 114.685 175.295 115.670 175.655 ;
        RECT 115.840 175.465 116.375 175.795 ;
        RECT 114.685 175.275 115.970 175.295 ;
        RECT 115.110 175.125 115.970 175.275 ;
        RECT 113.340 173.965 113.685 174.785 ;
        RECT 114.335 174.235 114.640 175.020 ;
        RECT 114.815 174.645 115.510 174.955 ;
        RECT 114.820 173.965 115.505 174.435 ;
        RECT 115.685 174.180 115.970 175.125 ;
        RECT 116.140 174.815 116.375 175.465 ;
        RECT 116.545 174.985 116.845 175.835 ;
        RECT 117.075 175.765 118.285 176.515 ;
        RECT 118.545 175.965 118.715 176.255 ;
        RECT 118.885 176.135 119.215 176.515 ;
        RECT 118.545 175.795 119.210 175.965 ;
        RECT 117.075 175.225 117.595 175.765 ;
        RECT 117.765 175.055 118.285 175.595 ;
        RECT 116.140 174.585 116.815 174.815 ;
        RECT 116.145 173.965 116.475 174.415 ;
        RECT 116.645 174.155 116.815 174.585 ;
        RECT 117.075 173.965 118.285 175.055 ;
        RECT 118.460 174.975 118.810 175.625 ;
        RECT 118.980 174.805 119.210 175.795 ;
        RECT 118.545 174.635 119.210 174.805 ;
        RECT 118.545 174.135 118.715 174.635 ;
        RECT 118.885 173.965 119.215 174.465 ;
        RECT 119.385 174.135 119.570 176.255 ;
        RECT 119.825 176.055 120.075 176.515 ;
        RECT 120.245 176.065 120.580 176.235 ;
        RECT 120.775 176.065 121.450 176.235 ;
        RECT 120.245 175.925 120.415 176.065 ;
        RECT 119.740 174.935 120.020 175.885 ;
        RECT 120.190 175.795 120.415 175.925 ;
        RECT 120.190 174.690 120.360 175.795 ;
        RECT 120.585 175.645 121.110 175.865 ;
        RECT 120.530 174.880 120.770 175.475 ;
        RECT 120.940 174.945 121.110 175.645 ;
        RECT 121.280 175.285 121.450 176.065 ;
        RECT 121.770 176.015 122.140 176.515 ;
        RECT 122.320 176.065 122.725 176.235 ;
        RECT 122.895 176.065 123.680 176.235 ;
        RECT 122.320 175.835 122.490 176.065 ;
        RECT 121.660 175.535 122.490 175.835 ;
        RECT 122.875 175.565 123.340 175.895 ;
        RECT 121.660 175.505 121.860 175.535 ;
        RECT 121.980 175.285 122.150 175.355 ;
        RECT 121.280 175.115 122.150 175.285 ;
        RECT 121.640 175.025 122.150 175.115 ;
        RECT 120.190 174.560 120.495 174.690 ;
        RECT 120.940 174.580 121.470 174.945 ;
        RECT 119.810 173.965 120.075 174.425 ;
        RECT 120.245 174.135 120.495 174.560 ;
        RECT 121.640 174.410 121.810 175.025 ;
        RECT 120.705 174.240 121.810 174.410 ;
        RECT 121.980 173.965 122.150 174.765 ;
        RECT 122.320 174.465 122.490 175.535 ;
        RECT 122.660 174.635 122.850 175.355 ;
        RECT 123.020 174.605 123.340 175.565 ;
        RECT 123.510 175.605 123.680 176.065 ;
        RECT 123.955 175.985 124.165 176.515 ;
        RECT 124.425 175.775 124.755 176.300 ;
        RECT 124.925 175.905 125.095 176.515 ;
        RECT 125.265 175.860 125.595 176.295 ;
        RECT 125.265 175.775 125.645 175.860 ;
        RECT 125.815 175.790 126.105 176.515 ;
        RECT 124.555 175.605 124.755 175.775 ;
        RECT 125.420 175.735 125.645 175.775 ;
        RECT 123.510 175.275 124.385 175.605 ;
        RECT 124.555 175.275 125.305 175.605 ;
        RECT 122.320 174.135 122.570 174.465 ;
        RECT 123.510 174.435 123.680 175.275 ;
        RECT 124.555 175.070 124.745 175.275 ;
        RECT 125.475 175.155 125.645 175.735 ;
        RECT 125.430 175.105 125.645 175.155 ;
        RECT 126.275 175.775 126.660 176.345 ;
        RECT 126.830 176.055 127.155 176.515 ;
        RECT 127.675 175.885 127.955 176.345 ;
        RECT 123.850 174.695 124.745 175.070 ;
        RECT 125.255 175.025 125.645 175.105 ;
        RECT 122.795 174.265 123.680 174.435 ;
        RECT 123.860 173.965 124.175 174.465 ;
        RECT 124.405 174.135 124.745 174.695 ;
        RECT 124.915 173.965 125.085 174.975 ;
        RECT 125.255 174.180 125.585 175.025 ;
        RECT 125.815 173.965 126.105 175.130 ;
        RECT 126.275 175.105 126.555 175.775 ;
        RECT 126.830 175.715 127.955 175.885 ;
        RECT 126.830 175.605 127.280 175.715 ;
        RECT 126.725 175.275 127.280 175.605 ;
        RECT 128.145 175.545 128.545 176.345 ;
        RECT 128.945 176.055 129.215 176.515 ;
        RECT 129.385 175.885 129.670 176.345 ;
        RECT 126.275 174.135 126.660 175.105 ;
        RECT 126.830 174.815 127.280 175.275 ;
        RECT 127.450 174.985 128.545 175.545 ;
        RECT 126.830 174.595 127.955 174.815 ;
        RECT 126.830 173.965 127.155 174.425 ;
        RECT 127.675 174.135 127.955 174.595 ;
        RECT 128.145 174.135 128.545 174.985 ;
        RECT 128.715 175.715 129.670 175.885 ;
        RECT 129.980 175.865 130.290 176.335 ;
        RECT 130.460 176.035 131.195 176.515 ;
        RECT 131.365 175.945 131.535 176.295 ;
        RECT 131.705 176.115 132.085 176.515 ;
        RECT 128.715 174.815 128.925 175.715 ;
        RECT 129.980 175.695 130.715 175.865 ;
        RECT 131.365 175.775 132.105 175.945 ;
        RECT 132.275 175.840 132.545 176.185 ;
        RECT 130.465 175.605 130.715 175.695 ;
        RECT 131.935 175.605 132.105 175.775 ;
        RECT 129.095 174.985 129.785 175.545 ;
        RECT 129.960 175.275 130.295 175.525 ;
        RECT 130.465 175.275 131.205 175.605 ;
        RECT 131.935 175.275 132.165 175.605 ;
        RECT 128.715 174.595 129.670 174.815 ;
        RECT 128.945 173.965 129.215 174.425 ;
        RECT 129.385 174.135 129.670 174.595 ;
        RECT 129.960 173.965 130.215 175.105 ;
        RECT 130.465 174.715 130.635 175.275 ;
        RECT 131.935 175.105 132.105 175.275 ;
        RECT 132.375 175.155 132.545 175.840 ;
        RECT 132.740 175.865 133.050 176.335 ;
        RECT 133.220 176.035 133.955 176.515 ;
        RECT 134.125 175.945 134.295 176.295 ;
        RECT 134.465 176.115 134.845 176.515 ;
        RECT 132.740 175.695 133.475 175.865 ;
        RECT 134.125 175.775 134.865 175.945 ;
        RECT 135.035 175.840 135.305 176.185 ;
        RECT 133.225 175.605 133.475 175.695 ;
        RECT 134.695 175.605 134.865 175.775 ;
        RECT 132.720 175.275 133.055 175.525 ;
        RECT 133.225 175.275 133.965 175.605 ;
        RECT 134.695 175.275 134.925 175.605 ;
        RECT 132.315 175.105 132.545 175.155 ;
        RECT 130.860 174.935 132.105 175.105 ;
        RECT 130.860 174.685 131.280 174.935 ;
        RECT 130.410 174.185 131.605 174.515 ;
        RECT 131.785 173.965 132.065 174.765 ;
        RECT 132.275 174.135 132.545 175.105 ;
        RECT 132.720 173.965 132.975 175.105 ;
        RECT 133.225 174.715 133.395 175.275 ;
        RECT 134.695 175.105 134.865 175.275 ;
        RECT 135.135 175.105 135.305 175.840 ;
        RECT 135.495 175.785 135.785 176.515 ;
        RECT 135.485 175.275 135.785 175.605 ;
        RECT 135.965 175.585 136.195 176.225 ;
        RECT 136.375 175.965 136.685 176.335 ;
        RECT 136.865 176.145 137.535 176.515 ;
        RECT 136.375 175.765 137.605 175.965 ;
        RECT 135.965 175.275 136.490 175.585 ;
        RECT 136.670 175.275 137.135 175.585 ;
        RECT 133.620 174.935 134.865 175.105 ;
        RECT 133.620 174.685 134.040 174.935 ;
        RECT 133.170 174.185 134.365 174.515 ;
        RECT 134.545 173.965 134.825 174.765 ;
        RECT 135.035 174.135 135.305 175.105 ;
        RECT 137.315 175.095 137.605 175.765 ;
        RECT 135.495 174.855 136.655 175.095 ;
        RECT 135.495 174.145 135.755 174.855 ;
        RECT 135.925 173.965 136.255 174.675 ;
        RECT 136.425 174.145 136.655 174.855 ;
        RECT 136.835 174.875 137.605 175.095 ;
        RECT 136.835 174.145 137.105 174.875 ;
        RECT 137.285 173.965 137.625 174.695 ;
        RECT 137.795 174.145 138.055 176.335 ;
        RECT 138.705 175.785 139.005 176.515 ;
        RECT 139.185 175.605 139.415 176.225 ;
        RECT 139.615 175.955 139.840 176.335 ;
        RECT 140.010 176.125 140.340 176.515 ;
        RECT 139.615 175.775 139.945 175.955 ;
        RECT 138.710 175.275 139.005 175.605 ;
        RECT 139.185 175.275 139.600 175.605 ;
        RECT 139.770 175.105 139.945 175.775 ;
        RECT 140.115 175.275 140.355 175.925 ;
        RECT 140.535 175.745 142.205 176.515 ;
        RECT 140.535 175.225 141.285 175.745 ;
        RECT 142.435 175.695 142.645 176.515 ;
        RECT 142.815 175.715 143.145 176.345 ;
        RECT 138.705 174.745 139.600 175.075 ;
        RECT 139.770 174.915 140.355 175.105 ;
        RECT 141.455 175.055 142.205 175.575 ;
        RECT 142.815 175.115 143.065 175.715 ;
        RECT 143.315 175.695 143.545 176.515 ;
        RECT 144.675 176.135 145.565 176.305 ;
        RECT 144.675 175.580 145.225 175.965 ;
        RECT 143.235 175.275 143.565 175.525 ;
        RECT 145.395 175.410 145.565 176.135 ;
        RECT 144.675 175.340 145.565 175.410 ;
        RECT 145.735 175.810 145.955 176.295 ;
        RECT 146.125 175.975 146.375 176.515 ;
        RECT 146.545 175.865 146.805 176.345 ;
        RECT 145.735 175.385 146.065 175.810 ;
        RECT 144.675 175.315 145.570 175.340 ;
        RECT 144.675 175.300 145.580 175.315 ;
        RECT 144.675 175.285 145.585 175.300 ;
        RECT 144.675 175.280 145.595 175.285 ;
        RECT 144.675 175.270 145.600 175.280 ;
        RECT 144.675 175.260 145.605 175.270 ;
        RECT 144.675 175.255 145.615 175.260 ;
        RECT 144.675 175.245 145.625 175.255 ;
        RECT 144.675 175.240 145.635 175.245 ;
        RECT 138.705 174.575 139.910 174.745 ;
        RECT 138.705 174.145 139.035 174.575 ;
        RECT 139.215 173.965 139.410 174.405 ;
        RECT 139.580 174.145 139.910 174.575 ;
        RECT 140.080 174.145 140.355 174.915 ;
        RECT 140.535 173.965 142.205 175.055 ;
        RECT 142.435 173.965 142.645 175.105 ;
        RECT 142.815 174.135 143.145 175.115 ;
        RECT 143.315 173.965 143.545 175.105 ;
        RECT 144.675 174.790 144.935 175.240 ;
        RECT 145.300 175.235 145.635 175.240 ;
        RECT 145.300 175.230 145.650 175.235 ;
        RECT 145.300 175.220 145.665 175.230 ;
        RECT 145.300 175.215 145.690 175.220 ;
        RECT 146.235 175.215 146.465 175.610 ;
        RECT 145.300 175.210 146.465 175.215 ;
        RECT 145.330 175.175 146.465 175.210 ;
        RECT 145.365 175.150 146.465 175.175 ;
        RECT 145.395 175.120 146.465 175.150 ;
        RECT 145.415 175.090 146.465 175.120 ;
        RECT 145.435 175.060 146.465 175.090 ;
        RECT 145.505 175.050 146.465 175.060 ;
        RECT 145.530 175.040 146.465 175.050 ;
        RECT 145.550 175.025 146.465 175.040 ;
        RECT 145.570 175.010 146.465 175.025 ;
        RECT 145.575 175.000 146.360 175.010 ;
        RECT 145.590 174.965 146.360 175.000 ;
        RECT 145.105 174.645 145.435 174.890 ;
        RECT 145.605 174.715 146.360 174.965 ;
        RECT 146.635 174.835 146.805 175.865 ;
        RECT 147.035 175.695 147.245 176.515 ;
        RECT 147.415 175.715 147.745 176.345 ;
        RECT 147.415 175.115 147.665 175.715 ;
        RECT 147.915 175.695 148.145 176.515 ;
        RECT 148.355 175.765 149.565 176.515 ;
        RECT 147.835 175.275 148.165 175.525 ;
        RECT 148.355 175.225 148.875 175.765 ;
        RECT 149.735 175.715 150.045 176.515 ;
        RECT 150.250 175.715 150.945 176.345 ;
        RECT 151.575 175.790 151.865 176.515 ;
        RECT 152.035 175.775 152.420 176.345 ;
        RECT 152.590 176.055 152.915 176.515 ;
        RECT 153.435 175.885 153.715 176.345 ;
        RECT 145.105 174.620 145.290 174.645 ;
        RECT 144.675 174.520 145.290 174.620 ;
        RECT 144.675 173.965 145.280 174.520 ;
        RECT 145.455 174.135 145.935 174.475 ;
        RECT 146.105 173.965 146.360 174.510 ;
        RECT 146.530 174.135 146.805 174.835 ;
        RECT 147.035 173.965 147.245 175.105 ;
        RECT 147.415 174.135 147.745 175.115 ;
        RECT 147.915 173.965 148.145 175.105 ;
        RECT 149.045 175.055 149.565 175.595 ;
        RECT 149.745 175.275 150.080 175.545 ;
        RECT 150.250 175.115 150.420 175.715 ;
        RECT 150.590 175.275 150.925 175.525 ;
        RECT 148.355 173.965 149.565 175.055 ;
        RECT 149.735 173.965 150.015 175.105 ;
        RECT 150.185 174.135 150.515 175.115 ;
        RECT 150.685 173.965 150.945 175.105 ;
        RECT 151.575 173.965 151.865 175.130 ;
        RECT 152.035 175.105 152.315 175.775 ;
        RECT 152.590 175.715 153.715 175.885 ;
        RECT 152.590 175.605 153.040 175.715 ;
        RECT 152.485 175.275 153.040 175.605 ;
        RECT 153.905 175.545 154.305 176.345 ;
        RECT 154.705 176.055 154.975 176.515 ;
        RECT 155.145 175.885 155.430 176.345 ;
        RECT 152.035 174.135 152.420 175.105 ;
        RECT 152.590 174.815 153.040 175.275 ;
        RECT 153.210 174.985 154.305 175.545 ;
        RECT 152.590 174.595 153.715 174.815 ;
        RECT 152.590 173.965 152.915 174.425 ;
        RECT 153.435 174.135 153.715 174.595 ;
        RECT 153.905 174.135 154.305 174.985 ;
        RECT 154.475 175.715 155.430 175.885 ;
        RECT 155.715 175.765 156.925 176.515 ;
        RECT 154.475 174.815 154.685 175.715 ;
        RECT 154.855 174.985 155.545 175.545 ;
        RECT 155.715 175.055 156.235 175.595 ;
        RECT 156.405 175.225 156.925 175.765 ;
        RECT 154.475 174.595 155.430 174.815 ;
        RECT 154.705 173.965 154.975 174.425 ;
        RECT 155.145 174.135 155.430 174.595 ;
        RECT 155.715 173.965 156.925 175.055 ;
        RECT 22.690 173.795 157.010 173.965 ;
        RECT 22.775 172.705 23.985 173.795 ;
        RECT 24.245 173.125 24.415 173.625 ;
        RECT 24.585 173.295 24.915 173.795 ;
        RECT 24.245 172.955 24.910 173.125 ;
        RECT 22.775 171.995 23.295 172.535 ;
        RECT 23.465 172.165 23.985 172.705 ;
        RECT 24.160 172.135 24.510 172.785 ;
        RECT 22.775 171.245 23.985 171.995 ;
        RECT 24.680 171.965 24.910 172.955 ;
        RECT 24.245 171.795 24.910 171.965 ;
        RECT 24.245 171.505 24.415 171.795 ;
        RECT 24.585 171.245 24.915 171.625 ;
        RECT 25.085 171.505 25.270 173.625 ;
        RECT 25.510 173.335 25.775 173.795 ;
        RECT 25.945 173.200 26.195 173.625 ;
        RECT 26.405 173.350 27.510 173.520 ;
        RECT 25.890 173.070 26.195 173.200 ;
        RECT 25.440 171.875 25.720 172.825 ;
        RECT 25.890 171.965 26.060 173.070 ;
        RECT 26.230 172.285 26.470 172.880 ;
        RECT 26.640 172.815 27.170 173.180 ;
        RECT 26.640 172.115 26.810 172.815 ;
        RECT 27.340 172.735 27.510 173.350 ;
        RECT 27.680 172.995 27.850 173.795 ;
        RECT 28.020 173.295 28.270 173.625 ;
        RECT 28.495 173.325 29.380 173.495 ;
        RECT 27.340 172.645 27.850 172.735 ;
        RECT 25.890 171.835 26.115 171.965 ;
        RECT 26.285 171.895 26.810 172.115 ;
        RECT 26.980 172.475 27.850 172.645 ;
        RECT 25.525 171.245 25.775 171.705 ;
        RECT 25.945 171.695 26.115 171.835 ;
        RECT 26.980 171.695 27.150 172.475 ;
        RECT 27.680 172.405 27.850 172.475 ;
        RECT 27.360 172.225 27.560 172.255 ;
        RECT 28.020 172.225 28.190 173.295 ;
        RECT 28.360 172.405 28.550 173.125 ;
        RECT 27.360 171.925 28.190 172.225 ;
        RECT 28.720 172.195 29.040 173.155 ;
        RECT 25.945 171.525 26.280 171.695 ;
        RECT 26.475 171.525 27.150 171.695 ;
        RECT 27.470 171.245 27.840 171.745 ;
        RECT 28.020 171.695 28.190 171.925 ;
        RECT 28.575 171.865 29.040 172.195 ;
        RECT 29.210 172.485 29.380 173.325 ;
        RECT 29.560 173.295 29.875 173.795 ;
        RECT 30.105 173.065 30.445 173.625 ;
        RECT 29.550 172.690 30.445 173.065 ;
        RECT 30.615 172.785 30.785 173.795 ;
        RECT 30.255 172.485 30.445 172.690 ;
        RECT 30.955 172.735 31.285 173.580 ;
        RECT 30.955 172.655 31.345 172.735 ;
        RECT 31.515 172.705 33.185 173.795 ;
        RECT 31.130 172.605 31.345 172.655 ;
        RECT 29.210 172.155 30.085 172.485 ;
        RECT 30.255 172.155 31.005 172.485 ;
        RECT 29.210 171.695 29.380 172.155 ;
        RECT 30.255 171.985 30.455 172.155 ;
        RECT 31.175 172.025 31.345 172.605 ;
        RECT 31.120 171.985 31.345 172.025 ;
        RECT 28.020 171.525 28.425 171.695 ;
        RECT 28.595 171.525 29.380 171.695 ;
        RECT 29.655 171.245 29.865 171.775 ;
        RECT 30.125 171.460 30.455 171.985 ;
        RECT 30.965 171.900 31.345 171.985 ;
        RECT 31.515 172.015 32.265 172.535 ;
        RECT 32.435 172.185 33.185 172.705 ;
        RECT 33.540 172.825 33.930 173.000 ;
        RECT 34.415 172.995 34.745 173.795 ;
        RECT 34.915 173.005 35.450 173.625 ;
        RECT 33.540 172.655 34.965 172.825 ;
        RECT 30.625 171.245 30.795 171.855 ;
        RECT 30.965 171.465 31.295 171.900 ;
        RECT 31.515 171.245 33.185 172.015 ;
        RECT 33.415 171.925 33.770 172.485 ;
        RECT 33.940 171.755 34.110 172.655 ;
        RECT 34.280 171.925 34.545 172.485 ;
        RECT 34.795 172.155 34.965 172.655 ;
        RECT 35.135 171.985 35.450 173.005 ;
        RECT 35.655 172.630 35.945 173.795 ;
        RECT 36.665 172.865 36.835 173.625 ;
        RECT 37.015 173.035 37.345 173.795 ;
        RECT 36.665 172.695 37.330 172.865 ;
        RECT 37.515 172.720 37.785 173.625 ;
        RECT 37.160 172.550 37.330 172.695 ;
        RECT 36.595 172.145 36.925 172.515 ;
        RECT 37.160 172.220 37.445 172.550 ;
        RECT 33.520 171.245 33.760 171.755 ;
        RECT 33.940 171.425 34.220 171.755 ;
        RECT 34.450 171.245 34.665 171.755 ;
        RECT 34.835 171.415 35.450 171.985 ;
        RECT 35.655 171.245 35.945 171.970 ;
        RECT 37.160 171.965 37.330 172.220 ;
        RECT 36.665 171.795 37.330 171.965 ;
        RECT 37.615 171.920 37.785 172.720 ;
        RECT 37.955 172.705 41.465 173.795 ;
        RECT 36.665 171.415 36.835 171.795 ;
        RECT 37.015 171.245 37.345 171.625 ;
        RECT 37.525 171.415 37.785 171.920 ;
        RECT 37.955 172.015 39.605 172.535 ;
        RECT 39.775 172.185 41.465 172.705 ;
        RECT 42.555 173.365 42.895 173.625 ;
        RECT 37.955 171.245 41.465 172.015 ;
        RECT 42.555 171.965 42.815 173.365 ;
        RECT 43.065 172.995 43.395 173.795 ;
        RECT 43.860 172.825 44.110 173.625 ;
        RECT 44.295 173.075 44.625 173.795 ;
        RECT 44.845 172.825 45.095 173.625 ;
        RECT 45.265 173.415 45.600 173.795 ;
        RECT 45.785 173.455 46.955 173.625 ;
        RECT 43.005 172.655 45.195 172.825 ;
        RECT 43.005 172.485 43.320 172.655 ;
        RECT 42.990 172.235 43.320 172.485 ;
        RECT 42.555 171.455 42.895 171.965 ;
        RECT 43.065 171.245 43.335 172.045 ;
        RECT 43.515 171.515 43.795 172.485 ;
        RECT 43.975 171.515 44.275 172.485 ;
        RECT 44.455 171.520 44.805 172.485 ;
        RECT 45.025 171.745 45.195 172.655 ;
        RECT 45.365 171.925 45.605 173.235 ;
        RECT 45.785 172.785 46.115 173.455 ;
        RECT 46.625 173.415 46.955 173.455 ;
        RECT 47.125 173.415 47.500 173.795 ;
        RECT 46.285 173.245 46.515 173.285 ;
        RECT 46.285 173.195 46.900 173.245 ;
        RECT 47.645 173.195 47.815 173.325 ;
        RECT 46.285 172.995 47.815 173.195 ;
        RECT 48.050 173.015 48.315 173.795 ;
        RECT 48.535 173.360 53.880 173.795 ;
        RECT 46.285 172.955 47.165 172.995 ;
        RECT 47.305 172.785 48.365 172.825 ;
        RECT 45.785 172.655 48.365 172.785 ;
        RECT 45.785 172.605 47.530 172.655 ;
        RECT 45.815 171.925 46.265 172.435 ;
        RECT 46.455 172.235 46.930 172.435 ;
        RECT 46.680 171.835 46.930 172.235 ;
        RECT 47.180 172.235 47.530 172.435 ;
        RECT 47.180 171.835 47.390 172.235 ;
        RECT 47.700 172.155 48.025 172.485 ;
        RECT 48.195 171.985 48.365 172.655 ;
        RECT 47.635 171.815 48.365 171.985 ;
        RECT 45.025 171.415 45.520 171.745 ;
        RECT 45.785 171.245 46.235 171.755 ;
        RECT 47.635 171.665 47.815 171.815 ;
        RECT 50.120 171.790 50.460 172.620 ;
        RECT 51.940 172.110 52.290 173.360 ;
        RECT 54.055 172.705 55.265 173.795 ;
        RECT 54.055 171.995 54.575 172.535 ;
        RECT 54.745 172.165 55.265 172.705 ;
        RECT 55.435 173.365 55.775 173.625 ;
        RECT 46.510 171.415 47.815 171.665 ;
        RECT 47.995 171.245 48.325 171.645 ;
        RECT 48.535 171.245 53.880 171.790 ;
        RECT 54.055 171.245 55.265 171.995 ;
        RECT 55.435 171.965 55.695 173.365 ;
        RECT 55.945 172.995 56.275 173.795 ;
        RECT 56.740 172.825 56.990 173.625 ;
        RECT 57.175 173.075 57.505 173.795 ;
        RECT 57.725 172.825 57.975 173.625 ;
        RECT 58.145 173.415 58.480 173.795 ;
        RECT 55.885 172.655 58.075 172.825 ;
        RECT 55.885 172.485 56.200 172.655 ;
        RECT 55.870 172.235 56.200 172.485 ;
        RECT 55.435 171.455 55.775 171.965 ;
        RECT 55.945 171.245 56.215 172.045 ;
        RECT 56.395 171.515 56.675 172.485 ;
        RECT 56.855 171.515 57.155 172.485 ;
        RECT 57.335 171.520 57.685 172.485 ;
        RECT 57.905 171.745 58.075 172.655 ;
        RECT 58.245 171.925 58.485 173.235 ;
        RECT 58.695 172.655 58.925 173.795 ;
        RECT 59.095 172.645 59.425 173.625 ;
        RECT 59.595 172.655 59.805 173.795 ;
        RECT 60.095 172.655 60.305 173.795 ;
        RECT 58.675 172.235 59.005 172.485 ;
        RECT 57.905 171.415 58.400 171.745 ;
        RECT 58.695 171.245 58.925 172.065 ;
        RECT 59.175 172.045 59.425 172.645 ;
        RECT 60.475 172.645 60.805 173.625 ;
        RECT 60.975 172.655 61.205 173.795 ;
        RECT 59.095 171.415 59.425 172.045 ;
        RECT 59.595 171.245 59.805 172.065 ;
        RECT 60.095 171.245 60.305 172.065 ;
        RECT 60.475 172.045 60.725 172.645 ;
        RECT 61.415 172.630 61.705 173.795 ;
        RECT 62.340 173.405 62.675 173.625 ;
        RECT 63.680 173.415 64.035 173.795 ;
        RECT 62.340 172.785 62.595 173.405 ;
        RECT 62.845 173.245 63.075 173.285 ;
        RECT 64.205 173.245 64.455 173.625 ;
        RECT 62.845 173.045 64.455 173.245 ;
        RECT 62.845 172.955 63.030 173.045 ;
        RECT 63.620 173.035 64.455 173.045 ;
        RECT 64.705 173.015 64.955 173.795 ;
        RECT 65.125 172.945 65.385 173.625 ;
        RECT 63.185 172.845 63.515 172.875 ;
        RECT 63.185 172.785 64.985 172.845 ;
        RECT 62.340 172.675 65.045 172.785 ;
        RECT 62.340 172.615 63.515 172.675 ;
        RECT 64.845 172.640 65.045 172.675 ;
        RECT 60.895 172.235 61.225 172.485 ;
        RECT 62.335 172.235 62.825 172.435 ;
        RECT 63.015 172.235 63.490 172.445 ;
        RECT 60.475 171.415 60.805 172.045 ;
        RECT 60.975 171.245 61.205 172.065 ;
        RECT 61.415 171.245 61.705 171.970 ;
        RECT 62.340 171.245 62.795 172.010 ;
        RECT 63.270 171.835 63.490 172.235 ;
        RECT 63.735 172.235 64.065 172.445 ;
        RECT 63.735 171.835 63.945 172.235 ;
        RECT 64.235 172.200 64.645 172.505 ;
        RECT 64.875 172.065 65.045 172.640 ;
        RECT 64.775 171.945 65.045 172.065 ;
        RECT 64.200 171.900 65.045 171.945 ;
        RECT 64.200 171.775 64.955 171.900 ;
        RECT 64.200 171.625 64.370 171.775 ;
        RECT 65.215 171.755 65.385 172.945 ;
        RECT 65.155 171.745 65.385 171.755 ;
        RECT 63.070 171.415 64.370 171.625 ;
        RECT 64.625 171.245 64.955 171.605 ;
        RECT 65.125 171.415 65.385 171.745 ;
        RECT 65.555 172.655 65.940 173.625 ;
        RECT 66.110 173.335 66.435 173.795 ;
        RECT 66.955 173.165 67.235 173.625 ;
        RECT 66.110 172.945 67.235 173.165 ;
        RECT 65.555 171.985 65.835 172.655 ;
        RECT 66.110 172.485 66.560 172.945 ;
        RECT 67.425 172.775 67.825 173.625 ;
        RECT 68.225 173.335 68.495 173.795 ;
        RECT 68.665 173.165 68.950 173.625 ;
        RECT 66.005 172.155 66.560 172.485 ;
        RECT 66.730 172.215 67.825 172.775 ;
        RECT 66.110 172.045 66.560 172.155 ;
        RECT 65.555 171.415 65.940 171.985 ;
        RECT 66.110 171.875 67.235 172.045 ;
        RECT 66.110 171.245 66.435 171.705 ;
        RECT 66.955 171.415 67.235 171.875 ;
        RECT 67.425 171.415 67.825 172.215 ;
        RECT 67.995 172.945 68.950 173.165 ;
        RECT 69.785 173.125 69.955 173.625 ;
        RECT 70.125 173.295 70.455 173.795 ;
        RECT 69.785 172.955 70.450 173.125 ;
        RECT 67.995 172.045 68.205 172.945 ;
        RECT 68.375 172.215 69.065 172.775 ;
        RECT 69.700 172.135 70.050 172.785 ;
        RECT 67.995 171.875 68.950 172.045 ;
        RECT 70.220 171.965 70.450 172.955 ;
        RECT 68.225 171.245 68.495 171.705 ;
        RECT 68.665 171.415 68.950 171.875 ;
        RECT 69.785 171.795 70.450 171.965 ;
        RECT 69.785 171.505 69.955 171.795 ;
        RECT 70.125 171.245 70.455 171.625 ;
        RECT 70.625 171.505 70.810 173.625 ;
        RECT 71.050 173.335 71.315 173.795 ;
        RECT 71.485 173.200 71.735 173.625 ;
        RECT 71.945 173.350 73.050 173.520 ;
        RECT 71.430 173.070 71.735 173.200 ;
        RECT 70.980 171.875 71.260 172.825 ;
        RECT 71.430 171.965 71.600 173.070 ;
        RECT 71.770 172.285 72.010 172.880 ;
        RECT 72.180 172.815 72.710 173.180 ;
        RECT 72.180 172.115 72.350 172.815 ;
        RECT 72.880 172.735 73.050 173.350 ;
        RECT 73.220 172.995 73.390 173.795 ;
        RECT 73.560 173.295 73.810 173.625 ;
        RECT 74.035 173.325 74.920 173.495 ;
        RECT 72.880 172.645 73.390 172.735 ;
        RECT 71.430 171.835 71.655 171.965 ;
        RECT 71.825 171.895 72.350 172.115 ;
        RECT 72.520 172.475 73.390 172.645 ;
        RECT 71.065 171.245 71.315 171.705 ;
        RECT 71.485 171.695 71.655 171.835 ;
        RECT 72.520 171.695 72.690 172.475 ;
        RECT 73.220 172.405 73.390 172.475 ;
        RECT 72.900 172.225 73.100 172.255 ;
        RECT 73.560 172.225 73.730 173.295 ;
        RECT 73.900 172.405 74.090 173.125 ;
        RECT 72.900 171.925 73.730 172.225 ;
        RECT 74.260 172.195 74.580 173.155 ;
        RECT 71.485 171.525 71.820 171.695 ;
        RECT 72.015 171.525 72.690 171.695 ;
        RECT 73.010 171.245 73.380 171.745 ;
        RECT 73.560 171.695 73.730 171.925 ;
        RECT 74.115 171.865 74.580 172.195 ;
        RECT 74.750 172.485 74.920 173.325 ;
        RECT 75.100 173.295 75.415 173.795 ;
        RECT 75.645 173.065 75.985 173.625 ;
        RECT 75.090 172.690 75.985 173.065 ;
        RECT 76.155 172.785 76.325 173.795 ;
        RECT 75.795 172.485 75.985 172.690 ;
        RECT 76.495 172.735 76.825 173.580 ;
        RECT 77.145 173.125 77.315 173.625 ;
        RECT 77.485 173.295 77.815 173.795 ;
        RECT 77.145 172.955 77.810 173.125 ;
        RECT 76.495 172.655 76.885 172.735 ;
        RECT 76.670 172.605 76.885 172.655 ;
        RECT 74.750 172.155 75.625 172.485 ;
        RECT 75.795 172.155 76.545 172.485 ;
        RECT 74.750 171.695 74.920 172.155 ;
        RECT 75.795 171.985 75.995 172.155 ;
        RECT 76.715 172.025 76.885 172.605 ;
        RECT 77.060 172.135 77.410 172.785 ;
        RECT 76.660 171.985 76.885 172.025 ;
        RECT 73.560 171.525 73.965 171.695 ;
        RECT 74.135 171.525 74.920 171.695 ;
        RECT 75.195 171.245 75.405 171.775 ;
        RECT 75.665 171.460 75.995 171.985 ;
        RECT 76.505 171.900 76.885 171.985 ;
        RECT 77.580 171.965 77.810 172.955 ;
        RECT 76.165 171.245 76.335 171.855 ;
        RECT 76.505 171.465 76.835 171.900 ;
        RECT 77.145 171.795 77.810 171.965 ;
        RECT 77.145 171.505 77.315 171.795 ;
        RECT 77.485 171.245 77.815 171.625 ;
        RECT 77.985 171.505 78.170 173.625 ;
        RECT 78.410 173.335 78.675 173.795 ;
        RECT 78.845 173.200 79.095 173.625 ;
        RECT 79.305 173.350 80.410 173.520 ;
        RECT 78.790 173.070 79.095 173.200 ;
        RECT 78.340 171.875 78.620 172.825 ;
        RECT 78.790 171.965 78.960 173.070 ;
        RECT 79.130 172.285 79.370 172.880 ;
        RECT 79.540 172.815 80.070 173.180 ;
        RECT 79.540 172.115 79.710 172.815 ;
        RECT 80.240 172.735 80.410 173.350 ;
        RECT 80.580 172.995 80.750 173.795 ;
        RECT 80.920 173.295 81.170 173.625 ;
        RECT 81.395 173.325 82.280 173.495 ;
        RECT 80.240 172.645 80.750 172.735 ;
        RECT 78.790 171.835 79.015 171.965 ;
        RECT 79.185 171.895 79.710 172.115 ;
        RECT 79.880 172.475 80.750 172.645 ;
        RECT 78.425 171.245 78.675 171.705 ;
        RECT 78.845 171.695 79.015 171.835 ;
        RECT 79.880 171.695 80.050 172.475 ;
        RECT 80.580 172.405 80.750 172.475 ;
        RECT 80.260 172.225 80.460 172.255 ;
        RECT 80.920 172.225 81.090 173.295 ;
        RECT 81.260 172.405 81.450 173.125 ;
        RECT 80.260 171.925 81.090 172.225 ;
        RECT 81.620 172.195 81.940 173.155 ;
        RECT 78.845 171.525 79.180 171.695 ;
        RECT 79.375 171.525 80.050 171.695 ;
        RECT 80.370 171.245 80.740 171.745 ;
        RECT 80.920 171.695 81.090 171.925 ;
        RECT 81.475 171.865 81.940 172.195 ;
        RECT 82.110 172.485 82.280 173.325 ;
        RECT 82.460 173.295 82.775 173.795 ;
        RECT 83.005 173.065 83.345 173.625 ;
        RECT 82.450 172.690 83.345 173.065 ;
        RECT 83.515 172.785 83.685 173.795 ;
        RECT 83.155 172.485 83.345 172.690 ;
        RECT 83.855 172.735 84.185 173.580 ;
        RECT 83.855 172.655 84.245 172.735 ;
        RECT 84.030 172.605 84.245 172.655 ;
        RECT 82.110 172.155 82.985 172.485 ;
        RECT 83.155 172.155 83.905 172.485 ;
        RECT 82.110 171.695 82.280 172.155 ;
        RECT 83.155 171.985 83.355 172.155 ;
        RECT 84.075 172.025 84.245 172.605 ;
        RECT 84.020 171.985 84.245 172.025 ;
        RECT 80.920 171.525 81.325 171.695 ;
        RECT 81.495 171.525 82.280 171.695 ;
        RECT 82.555 171.245 82.765 171.775 ;
        RECT 83.025 171.460 83.355 171.985 ;
        RECT 83.865 171.900 84.245 171.985 ;
        RECT 84.415 172.720 84.685 173.625 ;
        RECT 84.855 173.035 85.185 173.795 ;
        RECT 85.365 172.865 85.535 173.625 ;
        RECT 84.415 171.920 84.585 172.720 ;
        RECT 84.870 172.695 85.535 172.865 ;
        RECT 85.795 172.705 87.005 173.795 ;
        RECT 84.870 172.550 85.040 172.695 ;
        RECT 84.755 172.220 85.040 172.550 ;
        RECT 84.870 171.965 85.040 172.220 ;
        RECT 85.275 172.145 85.605 172.515 ;
        RECT 85.795 171.995 86.315 172.535 ;
        RECT 86.485 172.165 87.005 172.705 ;
        RECT 87.175 172.630 87.465 173.795 ;
        RECT 87.635 172.655 88.020 173.625 ;
        RECT 88.190 173.335 88.515 173.795 ;
        RECT 89.035 173.165 89.315 173.625 ;
        RECT 88.190 172.945 89.315 173.165 ;
        RECT 83.525 171.245 83.695 171.855 ;
        RECT 83.865 171.465 84.195 171.900 ;
        RECT 84.415 171.415 84.675 171.920 ;
        RECT 84.870 171.795 85.535 171.965 ;
        RECT 84.855 171.245 85.185 171.625 ;
        RECT 85.365 171.415 85.535 171.795 ;
        RECT 85.795 171.245 87.005 171.995 ;
        RECT 87.635 171.985 87.915 172.655 ;
        RECT 88.190 172.485 88.640 172.945 ;
        RECT 89.505 172.775 89.905 173.625 ;
        RECT 90.305 173.335 90.575 173.795 ;
        RECT 90.745 173.165 91.030 173.625 ;
        RECT 88.085 172.155 88.640 172.485 ;
        RECT 88.810 172.215 89.905 172.775 ;
        RECT 88.190 172.045 88.640 172.155 ;
        RECT 87.175 171.245 87.465 171.970 ;
        RECT 87.635 171.415 88.020 171.985 ;
        RECT 88.190 171.875 89.315 172.045 ;
        RECT 88.190 171.245 88.515 171.705 ;
        RECT 89.035 171.415 89.315 171.875 ;
        RECT 89.505 171.415 89.905 172.215 ;
        RECT 90.075 172.945 91.030 173.165 ;
        RECT 90.075 172.045 90.285 172.945 ;
        RECT 90.455 172.215 91.145 172.775 ;
        RECT 91.325 172.655 91.655 173.795 ;
        RECT 92.185 172.825 92.515 173.610 ;
        RECT 91.835 172.655 92.515 172.825 ;
        RECT 93.620 172.655 93.875 173.795 ;
        RECT 94.070 173.245 95.265 173.575 ;
        RECT 91.315 172.235 91.665 172.485 ;
        RECT 91.835 172.055 92.005 172.655 ;
        RECT 94.125 172.485 94.295 173.045 ;
        RECT 94.520 172.825 94.940 173.075 ;
        RECT 95.445 172.995 95.725 173.795 ;
        RECT 94.520 172.655 95.765 172.825 ;
        RECT 95.935 172.655 96.205 173.625 ;
        RECT 96.395 172.905 96.655 173.615 ;
        RECT 96.825 173.085 97.155 173.795 ;
        RECT 97.325 172.905 97.555 173.615 ;
        RECT 96.395 172.665 97.555 172.905 ;
        RECT 97.735 172.885 98.005 173.615 ;
        RECT 98.185 173.065 98.525 173.795 ;
        RECT 97.735 172.665 98.505 172.885 ;
        RECT 95.595 172.485 95.765 172.655 ;
        RECT 92.175 172.235 92.525 172.485 ;
        RECT 93.620 172.235 93.955 172.485 ;
        RECT 94.125 172.155 94.865 172.485 ;
        RECT 95.595 172.155 95.825 172.485 ;
        RECT 94.125 172.065 94.375 172.155 ;
        RECT 90.075 171.875 91.030 172.045 ;
        RECT 90.305 171.245 90.575 171.705 ;
        RECT 90.745 171.415 91.030 171.875 ;
        RECT 91.325 171.245 91.595 172.055 ;
        RECT 91.765 171.415 92.095 172.055 ;
        RECT 92.265 171.245 92.505 172.055 ;
        RECT 93.640 171.895 94.375 172.065 ;
        RECT 95.595 171.985 95.765 172.155 ;
        RECT 93.640 171.425 93.950 171.895 ;
        RECT 95.025 171.815 95.765 171.985 ;
        RECT 96.035 171.920 96.205 172.655 ;
        RECT 96.385 172.155 96.685 172.485 ;
        RECT 96.865 172.175 97.390 172.485 ;
        RECT 97.570 172.175 98.035 172.485 ;
        RECT 94.120 171.245 94.855 171.725 ;
        RECT 95.025 171.465 95.195 171.815 ;
        RECT 95.365 171.245 95.745 171.645 ;
        RECT 95.935 171.575 96.205 171.920 ;
        RECT 96.395 171.245 96.685 171.975 ;
        RECT 96.865 171.535 97.095 172.175 ;
        RECT 98.215 171.995 98.505 172.665 ;
        RECT 97.275 171.795 98.505 171.995 ;
        RECT 97.275 171.425 97.585 171.795 ;
        RECT 97.765 171.245 98.435 171.615 ;
        RECT 98.695 171.425 98.955 173.615 ;
        RECT 99.135 173.360 104.480 173.795 ;
        RECT 104.655 173.360 110.000 173.795 ;
        RECT 100.720 171.790 101.060 172.620 ;
        RECT 102.540 172.110 102.890 173.360 ;
        RECT 106.240 171.790 106.580 172.620 ;
        RECT 108.060 172.110 108.410 173.360 ;
        RECT 110.175 172.705 112.765 173.795 ;
        RECT 110.175 172.015 111.385 172.535 ;
        RECT 111.555 172.185 112.765 172.705 ;
        RECT 112.935 172.630 113.225 173.795 ;
        RECT 113.405 173.185 113.735 173.615 ;
        RECT 113.915 173.355 114.110 173.795 ;
        RECT 114.280 173.185 114.610 173.615 ;
        RECT 113.405 173.015 114.610 173.185 ;
        RECT 113.405 172.685 114.300 173.015 ;
        RECT 114.780 172.845 115.055 173.615 ;
        RECT 114.470 172.655 115.055 172.845 ;
        RECT 115.235 172.705 118.745 173.795 ;
        RECT 113.410 172.155 113.705 172.485 ;
        RECT 113.885 172.155 114.300 172.485 ;
        RECT 99.135 171.245 104.480 171.790 ;
        RECT 104.655 171.245 110.000 171.790 ;
        RECT 110.175 171.245 112.765 172.015 ;
        RECT 112.935 171.245 113.225 171.970 ;
        RECT 113.405 171.245 113.705 171.975 ;
        RECT 113.885 171.535 114.115 172.155 ;
        RECT 114.470 171.985 114.645 172.655 ;
        RECT 114.315 171.805 114.645 171.985 ;
        RECT 114.815 171.835 115.055 172.485 ;
        RECT 115.235 172.015 116.885 172.535 ;
        RECT 117.055 172.185 118.745 172.705 ;
        RECT 119.835 172.945 120.095 173.625 ;
        RECT 120.265 173.015 120.515 173.795 ;
        RECT 120.765 173.245 121.015 173.625 ;
        RECT 121.185 173.415 121.540 173.795 ;
        RECT 122.545 173.405 122.880 173.625 ;
        RECT 122.145 173.245 122.375 173.285 ;
        RECT 120.765 173.045 122.375 173.245 ;
        RECT 120.765 173.035 121.600 173.045 ;
        RECT 122.190 172.955 122.375 173.045 ;
        RECT 114.315 171.425 114.540 171.805 ;
        RECT 114.710 171.245 115.040 171.635 ;
        RECT 115.235 171.245 118.745 172.015 ;
        RECT 119.835 171.745 120.005 172.945 ;
        RECT 121.705 172.845 122.035 172.875 ;
        RECT 120.235 172.785 122.035 172.845 ;
        RECT 122.625 172.785 122.880 173.405 ;
        RECT 123.055 173.360 128.400 173.795 ;
        RECT 120.175 172.675 122.880 172.785 ;
        RECT 120.175 172.640 120.375 172.675 ;
        RECT 120.175 172.065 120.345 172.640 ;
        RECT 121.705 172.615 122.880 172.675 ;
        RECT 120.575 172.200 120.985 172.505 ;
        RECT 121.155 172.235 121.485 172.445 ;
        RECT 120.175 171.945 120.445 172.065 ;
        RECT 120.175 171.900 121.020 171.945 ;
        RECT 120.265 171.775 121.020 171.900 ;
        RECT 121.275 171.835 121.485 172.235 ;
        RECT 121.730 172.235 122.205 172.445 ;
        RECT 122.395 172.235 122.885 172.435 ;
        RECT 121.730 171.835 121.950 172.235 ;
        RECT 119.835 171.415 120.095 171.745 ;
        RECT 120.850 171.625 121.020 171.775 ;
        RECT 120.265 171.245 120.595 171.605 ;
        RECT 120.850 171.415 122.150 171.625 ;
        RECT 122.425 171.245 122.880 172.010 ;
        RECT 124.640 171.790 124.980 172.620 ;
        RECT 126.460 172.110 126.810 173.360 ;
        RECT 129.035 172.655 129.295 173.795 ;
        RECT 129.465 172.645 129.795 173.625 ;
        RECT 129.965 172.655 130.245 173.795 ;
        RECT 130.415 172.705 132.085 173.795 ;
        RECT 129.055 172.235 129.390 172.485 ;
        RECT 129.560 172.045 129.730 172.645 ;
        RECT 129.900 172.215 130.235 172.485 ;
        RECT 123.055 171.245 128.400 171.790 ;
        RECT 129.035 171.415 129.730 172.045 ;
        RECT 129.935 171.245 130.245 172.045 ;
        RECT 130.415 172.015 131.165 172.535 ;
        RECT 131.335 172.185 132.085 172.705 ;
        RECT 132.255 172.655 132.640 173.625 ;
        RECT 132.810 173.335 133.135 173.795 ;
        RECT 133.655 173.165 133.935 173.625 ;
        RECT 132.810 172.945 133.935 173.165 ;
        RECT 130.415 171.245 132.085 172.015 ;
        RECT 132.255 171.985 132.535 172.655 ;
        RECT 132.810 172.485 133.260 172.945 ;
        RECT 134.125 172.775 134.525 173.625 ;
        RECT 134.925 173.335 135.195 173.795 ;
        RECT 135.365 173.165 135.650 173.625 ;
        RECT 132.705 172.155 133.260 172.485 ;
        RECT 133.430 172.215 134.525 172.775 ;
        RECT 132.810 172.045 133.260 172.155 ;
        RECT 132.255 171.415 132.640 171.985 ;
        RECT 132.810 171.875 133.935 172.045 ;
        RECT 132.810 171.245 133.135 171.705 ;
        RECT 133.655 171.415 133.935 171.875 ;
        RECT 134.125 171.415 134.525 172.215 ;
        RECT 134.695 172.945 135.650 173.165 ;
        RECT 134.695 172.045 134.905 172.945 ;
        RECT 135.075 172.215 135.765 172.775 ;
        RECT 135.935 172.705 138.525 173.795 ;
        RECT 134.695 171.875 135.650 172.045 ;
        RECT 134.925 171.245 135.195 171.705 ;
        RECT 135.365 171.415 135.650 171.875 ;
        RECT 135.935 172.015 137.145 172.535 ;
        RECT 137.315 172.185 138.525 172.705 ;
        RECT 138.695 172.630 138.985 173.795 ;
        RECT 139.155 172.705 142.665 173.795 ;
        RECT 139.155 172.015 140.805 172.535 ;
        RECT 140.975 172.185 142.665 172.705 ;
        RECT 142.835 172.605 143.295 173.615 ;
        RECT 144.365 173.285 144.695 173.795 ;
        RECT 143.465 172.945 145.425 173.115 ;
        RECT 135.935 171.245 138.525 172.015 ;
        RECT 138.695 171.245 138.985 171.970 ;
        RECT 139.155 171.245 142.665 172.015 ;
        RECT 142.835 171.985 143.005 172.605 ;
        RECT 143.465 172.405 143.635 172.945 ;
        RECT 143.175 172.235 143.635 172.405 ;
        RECT 143.815 172.155 144.055 172.775 ;
        RECT 144.225 172.155 144.565 172.775 ;
        RECT 144.735 172.155 145.085 172.775 ;
        RECT 145.255 171.985 145.425 172.945 ;
        RECT 145.595 172.705 148.185 173.795 ;
        RECT 148.445 173.125 148.615 173.625 ;
        RECT 148.785 173.295 149.115 173.795 ;
        RECT 148.445 172.955 149.110 173.125 ;
        RECT 142.835 171.815 144.195 171.985 ;
        RECT 142.835 171.415 143.355 171.815 ;
        RECT 143.525 171.245 143.855 171.645 ;
        RECT 144.025 171.470 144.195 171.815 ;
        RECT 144.365 171.245 144.695 171.985 ;
        RECT 144.930 171.815 145.425 171.985 ;
        RECT 145.595 172.015 146.805 172.535 ;
        RECT 146.975 172.185 148.185 172.705 ;
        RECT 148.360 172.135 148.710 172.785 ;
        RECT 144.930 171.565 145.100 171.815 ;
        RECT 145.595 171.245 148.185 172.015 ;
        RECT 148.880 171.965 149.110 172.955 ;
        RECT 148.445 171.795 149.110 171.965 ;
        RECT 148.445 171.505 148.615 171.795 ;
        RECT 148.785 171.245 149.115 171.625 ;
        RECT 149.285 171.505 149.470 173.625 ;
        RECT 149.710 173.335 149.975 173.795 ;
        RECT 150.145 173.200 150.395 173.625 ;
        RECT 150.605 173.350 151.710 173.520 ;
        RECT 150.090 173.070 150.395 173.200 ;
        RECT 149.640 171.875 149.920 172.825 ;
        RECT 150.090 171.965 150.260 173.070 ;
        RECT 150.430 172.285 150.670 172.880 ;
        RECT 150.840 172.815 151.370 173.180 ;
        RECT 150.840 172.115 151.010 172.815 ;
        RECT 151.540 172.735 151.710 173.350 ;
        RECT 151.880 172.995 152.050 173.795 ;
        RECT 152.220 173.295 152.470 173.625 ;
        RECT 152.695 173.325 153.580 173.495 ;
        RECT 151.540 172.645 152.050 172.735 ;
        RECT 150.090 171.835 150.315 171.965 ;
        RECT 150.485 171.895 151.010 172.115 ;
        RECT 151.180 172.475 152.050 172.645 ;
        RECT 149.725 171.245 149.975 171.705 ;
        RECT 150.145 171.695 150.315 171.835 ;
        RECT 151.180 171.695 151.350 172.475 ;
        RECT 151.880 172.405 152.050 172.475 ;
        RECT 151.560 172.225 151.760 172.255 ;
        RECT 152.220 172.225 152.390 173.295 ;
        RECT 152.560 172.405 152.750 173.125 ;
        RECT 151.560 171.925 152.390 172.225 ;
        RECT 152.920 172.195 153.240 173.155 ;
        RECT 150.145 171.525 150.480 171.695 ;
        RECT 150.675 171.525 151.350 171.695 ;
        RECT 151.670 171.245 152.040 171.745 ;
        RECT 152.220 171.695 152.390 171.925 ;
        RECT 152.775 171.865 153.240 172.195 ;
        RECT 153.410 172.485 153.580 173.325 ;
        RECT 153.760 173.295 154.075 173.795 ;
        RECT 154.305 173.065 154.645 173.625 ;
        RECT 153.750 172.690 154.645 173.065 ;
        RECT 154.815 172.785 154.985 173.795 ;
        RECT 154.455 172.485 154.645 172.690 ;
        RECT 155.155 172.735 155.485 173.580 ;
        RECT 155.155 172.655 155.545 172.735 ;
        RECT 155.330 172.605 155.545 172.655 ;
        RECT 153.410 172.155 154.285 172.485 ;
        RECT 154.455 172.155 155.205 172.485 ;
        RECT 153.410 171.695 153.580 172.155 ;
        RECT 154.455 171.985 154.655 172.155 ;
        RECT 155.375 172.025 155.545 172.605 ;
        RECT 155.715 172.705 156.925 173.795 ;
        RECT 155.715 172.165 156.235 172.705 ;
        RECT 155.320 171.985 155.545 172.025 ;
        RECT 156.405 171.995 156.925 172.535 ;
        RECT 152.220 171.525 152.625 171.695 ;
        RECT 152.795 171.525 153.580 171.695 ;
        RECT 153.855 171.245 154.065 171.775 ;
        RECT 154.325 171.460 154.655 171.985 ;
        RECT 155.165 171.900 155.545 171.985 ;
        RECT 154.825 171.245 154.995 171.855 ;
        RECT 155.165 171.465 155.495 171.900 ;
        RECT 155.715 171.245 156.925 171.995 ;
        RECT 22.690 171.075 157.010 171.245 ;
        RECT 22.775 170.325 23.985 171.075 ;
        RECT 24.155 170.530 29.500 171.075 ;
        RECT 22.775 169.785 23.295 170.325 ;
        RECT 23.465 169.615 23.985 170.155 ;
        RECT 25.740 169.700 26.080 170.530 ;
        RECT 29.675 170.325 30.885 171.075 ;
        RECT 31.255 170.445 31.585 170.805 ;
        RECT 32.205 170.615 32.455 171.075 ;
        RECT 32.625 170.615 33.185 170.905 ;
        RECT 22.775 168.525 23.985 169.615 ;
        RECT 27.560 168.960 27.910 170.210 ;
        RECT 29.675 169.785 30.195 170.325 ;
        RECT 31.255 170.255 32.645 170.445 ;
        RECT 32.475 170.165 32.645 170.255 ;
        RECT 30.365 169.615 30.885 170.155 ;
        RECT 24.155 168.525 29.500 168.960 ;
        RECT 29.675 168.525 30.885 169.615 ;
        RECT 31.070 169.835 31.745 170.085 ;
        RECT 31.965 169.835 32.305 170.085 ;
        RECT 32.475 169.835 32.765 170.165 ;
        RECT 31.070 169.475 31.335 169.835 ;
        RECT 32.475 169.585 32.645 169.835 ;
        RECT 31.705 169.415 32.645 169.585 ;
        RECT 31.255 168.525 31.535 169.195 ;
        RECT 31.705 168.865 32.005 169.415 ;
        RECT 32.935 169.245 33.185 170.615 ;
        RECT 33.355 170.255 33.615 171.075 ;
        RECT 33.785 170.255 34.115 170.675 ;
        RECT 34.295 170.590 35.085 170.855 ;
        RECT 33.865 170.165 34.115 170.255 ;
        RECT 32.205 168.525 32.535 169.245 ;
        RECT 32.725 168.695 33.185 169.245 ;
        RECT 33.355 169.205 33.695 170.085 ;
        RECT 33.865 169.915 34.660 170.165 ;
        RECT 33.355 168.525 33.615 169.035 ;
        RECT 33.865 168.695 34.035 169.915 ;
        RECT 34.830 169.735 35.085 170.590 ;
        RECT 35.255 170.435 35.455 170.855 ;
        RECT 35.645 170.615 35.975 171.075 ;
        RECT 35.255 169.915 35.665 170.435 ;
        RECT 36.145 170.425 36.405 170.905 ;
        RECT 35.835 169.735 36.065 170.165 ;
        RECT 34.275 169.565 36.065 169.735 ;
        RECT 34.275 169.200 34.525 169.565 ;
        RECT 34.695 169.205 35.025 169.395 ;
        RECT 35.245 169.270 35.960 169.565 ;
        RECT 36.235 169.395 36.405 170.425 ;
        RECT 34.695 169.030 34.890 169.205 ;
        RECT 34.275 168.525 34.890 169.030 ;
        RECT 35.060 168.695 35.535 169.035 ;
        RECT 35.705 168.525 35.920 169.070 ;
        RECT 36.130 168.695 36.405 169.395 ;
        RECT 36.575 170.425 36.835 170.905 ;
        RECT 37.005 170.535 37.255 171.075 ;
        RECT 36.575 169.395 36.745 170.425 ;
        RECT 37.425 170.370 37.645 170.855 ;
        RECT 36.915 169.775 37.145 170.170 ;
        RECT 37.315 169.945 37.645 170.370 ;
        RECT 37.815 170.695 38.705 170.865 ;
        RECT 37.815 169.970 37.985 170.695 ;
        RECT 38.155 170.140 38.705 170.525 ;
        RECT 38.875 170.400 39.135 170.905 ;
        RECT 39.315 170.695 39.645 171.075 ;
        RECT 39.825 170.525 39.995 170.905 ;
        RECT 37.815 169.900 38.705 169.970 ;
        RECT 37.810 169.875 38.705 169.900 ;
        RECT 37.800 169.860 38.705 169.875 ;
        RECT 37.795 169.845 38.705 169.860 ;
        RECT 37.785 169.840 38.705 169.845 ;
        RECT 37.780 169.830 38.705 169.840 ;
        RECT 37.775 169.820 38.705 169.830 ;
        RECT 37.765 169.815 38.705 169.820 ;
        RECT 37.755 169.805 38.705 169.815 ;
        RECT 37.745 169.800 38.705 169.805 ;
        RECT 37.745 169.795 38.080 169.800 ;
        RECT 37.730 169.790 38.080 169.795 ;
        RECT 37.715 169.780 38.080 169.790 ;
        RECT 37.690 169.775 38.080 169.780 ;
        RECT 36.915 169.770 38.080 169.775 ;
        RECT 36.915 169.735 38.050 169.770 ;
        RECT 36.915 169.710 38.015 169.735 ;
        RECT 36.915 169.680 37.985 169.710 ;
        RECT 36.915 169.650 37.965 169.680 ;
        RECT 36.915 169.620 37.945 169.650 ;
        RECT 36.915 169.610 37.875 169.620 ;
        RECT 36.915 169.600 37.850 169.610 ;
        RECT 36.915 169.585 37.830 169.600 ;
        RECT 36.915 169.570 37.810 169.585 ;
        RECT 37.020 169.560 37.805 169.570 ;
        RECT 37.020 169.525 37.790 169.560 ;
        RECT 36.575 168.695 36.850 169.395 ;
        RECT 37.020 169.275 37.775 169.525 ;
        RECT 37.945 169.205 38.275 169.450 ;
        RECT 38.445 169.350 38.705 169.800 ;
        RECT 38.875 169.600 39.045 170.400 ;
        RECT 39.330 170.355 39.995 170.525 ;
        RECT 39.330 170.100 39.500 170.355 ;
        RECT 40.255 170.305 41.925 171.075 ;
        RECT 42.640 170.575 43.135 170.905 ;
        RECT 39.215 169.770 39.500 170.100 ;
        RECT 39.735 169.805 40.065 170.175 ;
        RECT 40.255 169.785 41.005 170.305 ;
        RECT 39.330 169.625 39.500 169.770 ;
        RECT 38.090 169.180 38.275 169.205 ;
        RECT 38.090 169.080 38.705 169.180 ;
        RECT 37.020 168.525 37.275 169.070 ;
        RECT 37.445 168.695 37.925 169.035 ;
        RECT 38.100 168.525 38.705 169.080 ;
        RECT 38.875 168.695 39.145 169.600 ;
        RECT 39.330 169.455 39.995 169.625 ;
        RECT 41.175 169.615 41.925 170.135 ;
        RECT 39.315 168.525 39.645 169.285 ;
        RECT 39.825 168.695 39.995 169.455 ;
        RECT 40.255 168.525 41.925 169.615 ;
        RECT 42.555 169.085 42.795 170.395 ;
        RECT 42.965 169.665 43.135 170.575 ;
        RECT 43.355 169.835 43.705 170.800 ;
        RECT 43.885 169.835 44.185 170.805 ;
        RECT 44.365 169.835 44.645 170.805 ;
        RECT 44.825 170.275 45.095 171.075 ;
        RECT 45.265 170.355 45.605 170.865 ;
        RECT 44.840 169.835 45.170 170.085 ;
        RECT 44.840 169.665 45.155 169.835 ;
        RECT 42.965 169.495 45.155 169.665 ;
        RECT 42.560 168.525 42.895 168.905 ;
        RECT 43.065 168.695 43.315 169.495 ;
        RECT 43.535 168.525 43.865 169.245 ;
        RECT 44.050 168.695 44.300 169.495 ;
        RECT 44.765 168.525 45.095 169.325 ;
        RECT 45.345 168.955 45.605 170.355 ;
        RECT 45.775 170.305 48.365 171.075 ;
        RECT 48.535 170.350 48.825 171.075 ;
        RECT 49.020 170.425 49.330 170.895 ;
        RECT 49.500 170.595 50.235 171.075 ;
        RECT 50.405 170.505 50.575 170.855 ;
        RECT 50.745 170.675 51.125 171.075 ;
        RECT 45.775 169.785 46.985 170.305 ;
        RECT 49.020 170.255 49.755 170.425 ;
        RECT 50.405 170.335 51.145 170.505 ;
        RECT 51.315 170.400 51.585 170.745 ;
        RECT 49.505 170.165 49.755 170.255 ;
        RECT 50.975 170.165 51.145 170.335 ;
        RECT 47.155 169.615 48.365 170.135 ;
        RECT 49.000 169.835 49.335 170.085 ;
        RECT 49.505 169.835 50.245 170.165 ;
        RECT 50.975 169.835 51.205 170.165 ;
        RECT 45.265 168.695 45.605 168.955 ;
        RECT 45.775 168.525 48.365 169.615 ;
        RECT 48.535 168.525 48.825 169.690 ;
        RECT 49.000 168.525 49.255 169.665 ;
        RECT 49.505 169.275 49.675 169.835 ;
        RECT 50.975 169.665 51.145 169.835 ;
        RECT 51.415 169.665 51.585 170.400 ;
        RECT 51.755 170.305 53.425 171.075 ;
        RECT 54.060 170.545 54.350 170.895 ;
        RECT 54.545 170.715 54.875 171.075 ;
        RECT 55.045 170.545 55.275 170.850 ;
        RECT 54.060 170.375 55.275 170.545 ;
        RECT 55.465 170.395 55.635 170.770 ;
        RECT 51.755 169.785 52.505 170.305 ;
        RECT 55.465 170.225 55.665 170.395 ;
        RECT 55.905 170.345 56.205 171.075 ;
        RECT 55.465 170.205 55.635 170.225 ;
        RECT 49.900 169.495 51.145 169.665 ;
        RECT 49.900 169.245 50.320 169.495 ;
        RECT 49.450 168.745 50.645 169.075 ;
        RECT 50.825 168.525 51.105 169.325 ;
        RECT 51.315 168.695 51.585 169.665 ;
        RECT 52.675 169.615 53.425 170.135 ;
        RECT 54.120 170.055 54.380 170.165 ;
        RECT 54.115 169.885 54.380 170.055 ;
        RECT 54.120 169.835 54.380 169.885 ;
        RECT 54.560 169.835 54.945 170.165 ;
        RECT 55.115 170.035 55.635 170.205 ;
        RECT 56.385 170.165 56.615 170.785 ;
        RECT 56.815 170.515 57.040 170.895 ;
        RECT 57.210 170.685 57.540 171.075 ;
        RECT 56.815 170.335 57.145 170.515 ;
        RECT 51.755 168.525 53.425 169.615 ;
        RECT 54.060 168.525 54.380 169.665 ;
        RECT 54.560 168.785 54.755 169.835 ;
        RECT 55.115 169.655 55.285 170.035 ;
        RECT 54.935 169.375 55.285 169.655 ;
        RECT 55.475 169.505 55.720 169.865 ;
        RECT 55.910 169.835 56.205 170.165 ;
        RECT 56.385 169.835 56.800 170.165 ;
        RECT 56.970 169.665 57.145 170.335 ;
        RECT 57.315 169.835 57.555 170.485 ;
        RECT 57.735 170.305 60.325 171.075 ;
        RECT 60.545 170.420 60.875 170.855 ;
        RECT 61.045 170.465 61.215 171.075 ;
        RECT 60.495 170.335 60.875 170.420 ;
        RECT 61.385 170.335 61.715 170.860 ;
        RECT 61.975 170.545 62.185 171.075 ;
        RECT 62.460 170.625 63.245 170.795 ;
        RECT 63.415 170.625 63.820 170.795 ;
        RECT 57.735 169.785 58.945 170.305 ;
        RECT 60.495 170.295 60.720 170.335 ;
        RECT 54.935 168.695 55.265 169.375 ;
        RECT 55.465 168.525 55.720 169.325 ;
        RECT 55.905 169.305 56.800 169.635 ;
        RECT 56.970 169.475 57.555 169.665 ;
        RECT 59.115 169.615 60.325 170.135 ;
        RECT 55.905 169.135 57.110 169.305 ;
        RECT 55.905 168.705 56.235 169.135 ;
        RECT 56.415 168.525 56.610 168.965 ;
        RECT 56.780 168.705 57.110 169.135 ;
        RECT 57.280 168.705 57.555 169.475 ;
        RECT 57.735 168.525 60.325 169.615 ;
        RECT 60.495 169.715 60.665 170.295 ;
        RECT 61.385 170.165 61.585 170.335 ;
        RECT 62.460 170.165 62.630 170.625 ;
        RECT 60.835 169.835 61.585 170.165 ;
        RECT 61.755 169.835 62.630 170.165 ;
        RECT 60.495 169.665 60.710 169.715 ;
        RECT 60.495 169.585 60.885 169.665 ;
        RECT 60.555 168.740 60.885 169.585 ;
        RECT 61.395 169.630 61.585 169.835 ;
        RECT 61.055 168.525 61.225 169.535 ;
        RECT 61.395 169.255 62.290 169.630 ;
        RECT 61.395 168.695 61.735 169.255 ;
        RECT 61.965 168.525 62.280 169.025 ;
        RECT 62.460 168.995 62.630 169.835 ;
        RECT 62.800 170.125 63.265 170.455 ;
        RECT 63.650 170.395 63.820 170.625 ;
        RECT 64.000 170.575 64.370 171.075 ;
        RECT 64.690 170.625 65.365 170.795 ;
        RECT 65.560 170.625 65.895 170.795 ;
        RECT 62.800 169.165 63.120 170.125 ;
        RECT 63.650 170.095 64.480 170.395 ;
        RECT 63.290 169.195 63.480 169.915 ;
        RECT 63.650 169.025 63.820 170.095 ;
        RECT 64.280 170.065 64.480 170.095 ;
        RECT 63.990 169.845 64.160 169.915 ;
        RECT 64.690 169.845 64.860 170.625 ;
        RECT 65.725 170.485 65.895 170.625 ;
        RECT 66.065 170.615 66.315 171.075 ;
        RECT 63.990 169.675 64.860 169.845 ;
        RECT 65.030 170.205 65.555 170.425 ;
        RECT 65.725 170.355 65.950 170.485 ;
        RECT 63.990 169.585 64.500 169.675 ;
        RECT 62.460 168.825 63.345 168.995 ;
        RECT 63.570 168.695 63.820 169.025 ;
        RECT 63.990 168.525 64.160 169.325 ;
        RECT 64.330 168.970 64.500 169.585 ;
        RECT 65.030 169.505 65.200 170.205 ;
        RECT 64.670 169.140 65.200 169.505 ;
        RECT 65.370 169.440 65.610 170.035 ;
        RECT 65.780 169.250 65.950 170.355 ;
        RECT 66.120 169.495 66.400 170.445 ;
        RECT 65.645 169.120 65.950 169.250 ;
        RECT 64.330 168.800 65.435 168.970 ;
        RECT 65.645 168.695 65.895 169.120 ;
        RECT 66.065 168.525 66.330 168.985 ;
        RECT 66.570 168.695 66.755 170.815 ;
        RECT 66.925 170.695 67.255 171.075 ;
        RECT 67.425 170.525 67.595 170.815 ;
        RECT 68.365 170.605 68.655 171.075 ;
        RECT 66.930 170.355 67.595 170.525 ;
        RECT 68.825 170.435 69.155 170.905 ;
        RECT 69.325 170.605 69.495 171.075 ;
        RECT 69.665 170.435 69.995 170.905 ;
        RECT 68.825 170.425 69.995 170.435 ;
        RECT 68.395 170.395 69.995 170.425 ;
        RECT 66.930 169.365 67.160 170.355 ;
        RECT 68.375 170.255 69.995 170.395 ;
        RECT 70.165 170.255 70.440 171.075 ;
        RECT 70.620 170.310 71.075 171.075 ;
        RECT 71.350 170.695 72.650 170.905 ;
        RECT 72.905 170.715 73.235 171.075 ;
        RECT 72.480 170.545 72.650 170.695 ;
        RECT 73.405 170.575 73.665 170.905 ;
        RECT 68.375 170.225 68.610 170.255 ;
        RECT 67.330 169.535 67.680 170.185 ;
        RECT 68.395 169.715 68.610 170.225 ;
        RECT 71.550 170.085 71.770 170.485 ;
        RECT 68.780 169.885 69.550 170.085 ;
        RECT 69.720 169.885 70.440 170.085 ;
        RECT 70.615 169.885 71.105 170.085 ;
        RECT 71.295 169.875 71.770 170.085 ;
        RECT 72.015 170.085 72.225 170.485 ;
        RECT 72.480 170.420 73.235 170.545 ;
        RECT 72.480 170.375 73.325 170.420 ;
        RECT 73.055 170.255 73.325 170.375 ;
        RECT 72.015 169.875 72.345 170.085 ;
        RECT 72.515 169.815 72.925 170.120 ;
        RECT 68.395 169.495 69.155 169.715 ;
        RECT 66.930 169.195 67.595 169.365 ;
        RECT 66.925 168.525 67.255 169.025 ;
        RECT 67.425 168.695 67.595 169.195 ;
        RECT 68.355 168.865 68.655 169.325 ;
        RECT 68.825 169.035 69.155 169.495 ;
        RECT 69.325 169.495 70.440 169.705 ;
        RECT 69.325 168.865 69.495 169.495 ;
        RECT 68.355 168.695 69.495 168.865 ;
        RECT 69.665 168.525 69.995 169.325 ;
        RECT 70.165 168.695 70.440 169.495 ;
        RECT 70.620 169.645 71.795 169.705 ;
        RECT 73.155 169.680 73.325 170.255 ;
        RECT 73.125 169.645 73.325 169.680 ;
        RECT 70.620 169.535 73.325 169.645 ;
        RECT 70.620 168.915 70.875 169.535 ;
        RECT 71.465 169.475 73.265 169.535 ;
        RECT 71.465 169.445 71.795 169.475 ;
        RECT 73.495 169.375 73.665 170.575 ;
        RECT 74.295 170.350 74.585 171.075 ;
        RECT 74.755 170.325 75.965 171.075 ;
        RECT 76.135 170.575 76.395 170.905 ;
        RECT 76.565 170.715 76.895 171.075 ;
        RECT 77.150 170.695 78.450 170.905 ;
        RECT 74.755 169.785 75.275 170.325 ;
        RECT 71.125 169.275 71.310 169.365 ;
        RECT 71.900 169.275 72.735 169.285 ;
        RECT 71.125 169.075 72.735 169.275 ;
        RECT 71.125 169.035 71.355 169.075 ;
        RECT 70.620 168.695 70.955 168.915 ;
        RECT 71.960 168.525 72.315 168.905 ;
        RECT 72.485 168.695 72.735 169.075 ;
        RECT 72.985 168.525 73.235 169.305 ;
        RECT 73.405 168.695 73.665 169.375 ;
        RECT 74.295 168.525 74.585 169.690 ;
        RECT 75.445 169.615 75.965 170.155 ;
        RECT 74.755 168.525 75.965 169.615 ;
        RECT 76.135 169.375 76.305 170.575 ;
        RECT 77.150 170.545 77.320 170.695 ;
        RECT 76.565 170.420 77.320 170.545 ;
        RECT 76.475 170.375 77.320 170.420 ;
        RECT 76.475 170.255 76.745 170.375 ;
        RECT 76.475 169.680 76.645 170.255 ;
        RECT 76.875 169.815 77.285 170.120 ;
        RECT 77.575 170.085 77.785 170.485 ;
        RECT 77.455 169.875 77.785 170.085 ;
        RECT 78.030 170.085 78.250 170.485 ;
        RECT 78.725 170.310 79.180 171.075 ;
        RECT 79.355 170.575 79.615 170.905 ;
        RECT 79.785 170.715 80.115 171.075 ;
        RECT 80.370 170.695 81.670 170.905 ;
        RECT 78.030 169.875 78.505 170.085 ;
        RECT 78.695 169.885 79.185 170.085 ;
        RECT 76.475 169.645 76.675 169.680 ;
        RECT 78.005 169.645 79.180 169.705 ;
        RECT 76.475 169.535 79.180 169.645 ;
        RECT 76.535 169.475 78.335 169.535 ;
        RECT 78.005 169.445 78.335 169.475 ;
        RECT 76.135 168.695 76.395 169.375 ;
        RECT 76.565 168.525 76.815 169.305 ;
        RECT 77.065 169.275 77.900 169.285 ;
        RECT 78.490 169.275 78.675 169.365 ;
        RECT 77.065 169.075 78.675 169.275 ;
        RECT 77.065 168.695 77.315 169.075 ;
        RECT 78.445 169.035 78.675 169.075 ;
        RECT 78.925 168.915 79.180 169.535 ;
        RECT 77.485 168.525 77.840 168.905 ;
        RECT 78.845 168.695 79.180 168.915 ;
        RECT 79.355 169.375 79.525 170.575 ;
        RECT 80.370 170.545 80.540 170.695 ;
        RECT 79.785 170.420 80.540 170.545 ;
        RECT 79.695 170.375 80.540 170.420 ;
        RECT 79.695 170.255 79.965 170.375 ;
        RECT 79.695 169.680 79.865 170.255 ;
        RECT 80.095 169.815 80.505 170.120 ;
        RECT 80.795 170.085 81.005 170.485 ;
        RECT 80.675 169.875 81.005 170.085 ;
        RECT 81.250 170.085 81.470 170.485 ;
        RECT 81.945 170.310 82.400 171.075 ;
        RECT 82.575 170.335 82.960 170.905 ;
        RECT 83.130 170.615 83.455 171.075 ;
        RECT 83.975 170.445 84.255 170.905 ;
        RECT 81.250 169.875 81.725 170.085 ;
        RECT 81.915 169.885 82.405 170.085 ;
        RECT 79.695 169.645 79.895 169.680 ;
        RECT 81.225 169.645 82.400 169.705 ;
        RECT 79.695 169.535 82.400 169.645 ;
        RECT 79.755 169.475 81.555 169.535 ;
        RECT 81.225 169.445 81.555 169.475 ;
        RECT 79.355 168.695 79.615 169.375 ;
        RECT 79.785 168.525 80.035 169.305 ;
        RECT 80.285 169.275 81.120 169.285 ;
        RECT 81.710 169.275 81.895 169.365 ;
        RECT 80.285 169.075 81.895 169.275 ;
        RECT 80.285 168.695 80.535 169.075 ;
        RECT 81.665 169.035 81.895 169.075 ;
        RECT 82.145 168.915 82.400 169.535 ;
        RECT 80.705 168.525 81.060 168.905 ;
        RECT 82.065 168.695 82.400 168.915 ;
        RECT 82.575 169.665 82.855 170.335 ;
        RECT 83.130 170.275 84.255 170.445 ;
        RECT 83.130 170.165 83.580 170.275 ;
        RECT 83.025 169.835 83.580 170.165 ;
        RECT 84.445 170.105 84.845 170.905 ;
        RECT 85.245 170.615 85.515 171.075 ;
        RECT 85.685 170.445 85.970 170.905 ;
        RECT 82.575 168.695 82.960 169.665 ;
        RECT 83.130 169.375 83.580 169.835 ;
        RECT 83.750 169.545 84.845 170.105 ;
        RECT 83.130 169.155 84.255 169.375 ;
        RECT 83.130 168.525 83.455 168.985 ;
        RECT 83.975 168.695 84.255 169.155 ;
        RECT 84.445 168.695 84.845 169.545 ;
        RECT 85.015 170.275 85.970 170.445 ;
        RECT 86.255 170.305 89.765 171.075 ;
        RECT 89.935 170.325 91.145 171.075 ;
        RECT 91.340 170.425 91.650 170.895 ;
        RECT 91.820 170.595 92.555 171.075 ;
        RECT 92.725 170.505 92.895 170.855 ;
        RECT 93.065 170.675 93.445 171.075 ;
        RECT 85.015 169.375 85.225 170.275 ;
        RECT 85.395 169.545 86.085 170.105 ;
        RECT 86.255 169.785 87.905 170.305 ;
        RECT 88.075 169.615 89.765 170.135 ;
        RECT 89.935 169.785 90.455 170.325 ;
        RECT 91.340 170.255 92.075 170.425 ;
        RECT 92.725 170.335 93.465 170.505 ;
        RECT 93.635 170.400 93.905 170.745 ;
        RECT 94.080 170.570 94.415 171.075 ;
        RECT 94.585 170.505 94.825 170.880 ;
        RECT 95.105 170.745 95.275 170.890 ;
        RECT 95.105 170.550 95.480 170.745 ;
        RECT 95.840 170.580 96.235 171.075 ;
        RECT 91.825 170.165 92.075 170.255 ;
        RECT 93.295 170.165 93.465 170.335 ;
        RECT 90.625 169.615 91.145 170.155 ;
        RECT 91.320 169.835 91.655 170.085 ;
        RECT 91.825 169.835 92.565 170.165 ;
        RECT 93.295 169.835 93.525 170.165 ;
        RECT 85.015 169.155 85.970 169.375 ;
        RECT 85.245 168.525 85.515 168.985 ;
        RECT 85.685 168.695 85.970 169.155 ;
        RECT 86.255 168.525 89.765 169.615 ;
        RECT 89.935 168.525 91.145 169.615 ;
        RECT 91.320 168.525 91.575 169.665 ;
        RECT 91.825 169.275 91.995 169.835 ;
        RECT 93.295 169.665 93.465 169.835 ;
        RECT 93.735 169.665 93.905 170.400 ;
        RECT 92.220 169.495 93.465 169.665 ;
        RECT 92.220 169.245 92.640 169.495 ;
        RECT 91.770 168.745 92.965 169.075 ;
        RECT 93.145 168.525 93.425 169.325 ;
        RECT 93.635 168.695 93.905 169.665 ;
        RECT 94.135 169.545 94.435 170.395 ;
        RECT 94.605 170.355 94.825 170.505 ;
        RECT 94.605 170.025 95.140 170.355 ;
        RECT 95.310 170.215 95.480 170.550 ;
        RECT 96.405 170.385 96.645 170.905 ;
        RECT 94.605 169.375 94.840 170.025 ;
        RECT 95.310 169.855 96.295 170.215 ;
        RECT 94.165 169.145 94.840 169.375 ;
        RECT 95.010 169.835 96.295 169.855 ;
        RECT 95.010 169.685 95.870 169.835 ;
        RECT 94.165 168.715 94.335 169.145 ;
        RECT 94.505 168.525 94.835 168.975 ;
        RECT 95.010 168.740 95.295 169.685 ;
        RECT 96.470 169.580 96.645 170.385 ;
        RECT 96.835 170.305 99.425 171.075 ;
        RECT 100.055 170.350 100.345 171.075 ;
        RECT 100.565 170.420 100.895 170.855 ;
        RECT 101.065 170.465 101.235 171.075 ;
        RECT 100.515 170.335 100.895 170.420 ;
        RECT 101.405 170.335 101.735 170.860 ;
        RECT 101.995 170.545 102.205 171.075 ;
        RECT 102.480 170.625 103.265 170.795 ;
        RECT 103.435 170.625 103.840 170.795 ;
        RECT 96.835 169.785 98.045 170.305 ;
        RECT 100.515 170.295 100.740 170.335 ;
        RECT 98.215 169.615 99.425 170.135 ;
        RECT 100.515 169.715 100.685 170.295 ;
        RECT 101.405 170.165 101.605 170.335 ;
        RECT 102.480 170.165 102.650 170.625 ;
        RECT 100.855 169.835 101.605 170.165 ;
        RECT 101.775 169.835 102.650 170.165 ;
        RECT 95.470 169.205 96.165 169.515 ;
        RECT 95.475 168.525 96.160 168.995 ;
        RECT 96.340 168.795 96.645 169.580 ;
        RECT 96.835 168.525 99.425 169.615 ;
        RECT 100.055 168.525 100.345 169.690 ;
        RECT 100.515 169.665 100.730 169.715 ;
        RECT 100.515 169.585 100.905 169.665 ;
        RECT 100.575 168.740 100.905 169.585 ;
        RECT 101.415 169.630 101.605 169.835 ;
        RECT 101.075 168.525 101.245 169.535 ;
        RECT 101.415 169.255 102.310 169.630 ;
        RECT 101.415 168.695 101.755 169.255 ;
        RECT 101.985 168.525 102.300 169.025 ;
        RECT 102.480 168.995 102.650 169.835 ;
        RECT 102.820 170.125 103.285 170.455 ;
        RECT 103.670 170.395 103.840 170.625 ;
        RECT 104.020 170.575 104.390 171.075 ;
        RECT 104.710 170.625 105.385 170.795 ;
        RECT 105.580 170.625 105.915 170.795 ;
        RECT 102.820 169.165 103.140 170.125 ;
        RECT 103.670 170.095 104.500 170.395 ;
        RECT 103.310 169.195 103.500 169.915 ;
        RECT 103.670 169.025 103.840 170.095 ;
        RECT 104.300 170.065 104.500 170.095 ;
        RECT 104.010 169.845 104.180 169.915 ;
        RECT 104.710 169.845 104.880 170.625 ;
        RECT 105.745 170.485 105.915 170.625 ;
        RECT 106.085 170.615 106.335 171.075 ;
        RECT 104.010 169.675 104.880 169.845 ;
        RECT 105.050 170.205 105.575 170.425 ;
        RECT 105.745 170.355 105.970 170.485 ;
        RECT 104.010 169.585 104.520 169.675 ;
        RECT 102.480 168.825 103.365 168.995 ;
        RECT 103.590 168.695 103.840 169.025 ;
        RECT 104.010 168.525 104.180 169.325 ;
        RECT 104.350 168.970 104.520 169.585 ;
        RECT 105.050 169.505 105.220 170.205 ;
        RECT 104.690 169.140 105.220 169.505 ;
        RECT 105.390 169.440 105.630 170.035 ;
        RECT 105.800 169.250 105.970 170.355 ;
        RECT 106.140 169.495 106.420 170.445 ;
        RECT 105.665 169.120 105.970 169.250 ;
        RECT 104.350 168.800 105.455 168.970 ;
        RECT 105.665 168.695 105.915 169.120 ;
        RECT 106.085 168.525 106.350 168.985 ;
        RECT 106.590 168.695 106.775 170.815 ;
        RECT 106.945 170.695 107.275 171.075 ;
        RECT 107.445 170.525 107.615 170.815 ;
        RECT 106.950 170.355 107.615 170.525 ;
        RECT 106.950 169.365 107.180 170.355 ;
        RECT 107.875 170.305 109.545 171.075 ;
        RECT 109.805 170.525 109.975 170.815 ;
        RECT 110.145 170.695 110.475 171.075 ;
        RECT 109.805 170.355 110.470 170.525 ;
        RECT 107.350 169.535 107.700 170.185 ;
        RECT 107.875 169.785 108.625 170.305 ;
        RECT 108.795 169.615 109.545 170.135 ;
        RECT 106.950 169.195 107.615 169.365 ;
        RECT 106.945 168.525 107.275 169.025 ;
        RECT 107.445 168.695 107.615 169.195 ;
        RECT 107.875 168.525 109.545 169.615 ;
        RECT 109.720 169.535 110.070 170.185 ;
        RECT 110.240 169.365 110.470 170.355 ;
        RECT 109.805 169.195 110.470 169.365 ;
        RECT 109.805 168.695 109.975 169.195 ;
        RECT 110.145 168.525 110.475 169.025 ;
        RECT 110.645 168.695 110.830 170.815 ;
        RECT 111.085 170.615 111.335 171.075 ;
        RECT 111.505 170.625 111.840 170.795 ;
        RECT 112.035 170.625 112.710 170.795 ;
        RECT 111.505 170.485 111.675 170.625 ;
        RECT 111.000 169.495 111.280 170.445 ;
        RECT 111.450 170.355 111.675 170.485 ;
        RECT 111.450 169.250 111.620 170.355 ;
        RECT 111.845 170.205 112.370 170.425 ;
        RECT 111.790 169.440 112.030 170.035 ;
        RECT 112.200 169.505 112.370 170.205 ;
        RECT 112.540 169.845 112.710 170.625 ;
        RECT 113.030 170.575 113.400 171.075 ;
        RECT 113.580 170.625 113.985 170.795 ;
        RECT 114.155 170.625 114.940 170.795 ;
        RECT 113.580 170.395 113.750 170.625 ;
        RECT 112.920 170.095 113.750 170.395 ;
        RECT 114.135 170.125 114.600 170.455 ;
        RECT 112.920 170.065 113.120 170.095 ;
        RECT 113.240 169.845 113.410 169.915 ;
        RECT 112.540 169.675 113.410 169.845 ;
        RECT 112.900 169.585 113.410 169.675 ;
        RECT 111.450 169.120 111.755 169.250 ;
        RECT 112.200 169.140 112.730 169.505 ;
        RECT 111.070 168.525 111.335 168.985 ;
        RECT 111.505 168.695 111.755 169.120 ;
        RECT 112.900 168.970 113.070 169.585 ;
        RECT 111.965 168.800 113.070 168.970 ;
        RECT 113.240 168.525 113.410 169.325 ;
        RECT 113.580 169.025 113.750 170.095 ;
        RECT 113.920 169.195 114.110 169.915 ;
        RECT 114.280 169.165 114.600 170.125 ;
        RECT 114.770 170.165 114.940 170.625 ;
        RECT 115.215 170.545 115.425 171.075 ;
        RECT 115.685 170.335 116.015 170.860 ;
        RECT 116.185 170.465 116.355 171.075 ;
        RECT 116.525 170.420 116.855 170.855 ;
        RECT 116.525 170.335 116.905 170.420 ;
        RECT 115.815 170.165 116.015 170.335 ;
        RECT 116.680 170.295 116.905 170.335 ;
        RECT 114.770 169.835 115.645 170.165 ;
        RECT 115.815 169.835 116.565 170.165 ;
        RECT 113.580 168.695 113.830 169.025 ;
        RECT 114.770 168.995 114.940 169.835 ;
        RECT 115.815 169.630 116.005 169.835 ;
        RECT 116.735 169.715 116.905 170.295 ;
        RECT 116.690 169.665 116.905 169.715 ;
        RECT 115.110 169.255 116.005 169.630 ;
        RECT 116.515 169.585 116.905 169.665 ;
        RECT 117.075 170.335 117.460 170.905 ;
        RECT 117.630 170.615 117.955 171.075 ;
        RECT 118.475 170.445 118.755 170.905 ;
        RECT 117.075 169.665 117.355 170.335 ;
        RECT 117.630 170.275 118.755 170.445 ;
        RECT 117.630 170.165 118.080 170.275 ;
        RECT 117.525 169.835 118.080 170.165 ;
        RECT 118.945 170.105 119.345 170.905 ;
        RECT 119.745 170.615 120.015 171.075 ;
        RECT 120.185 170.445 120.470 170.905 ;
        RECT 114.055 168.825 114.940 168.995 ;
        RECT 115.120 168.525 115.435 169.025 ;
        RECT 115.665 168.695 116.005 169.255 ;
        RECT 116.175 168.525 116.345 169.535 ;
        RECT 116.515 168.740 116.845 169.585 ;
        RECT 117.075 168.695 117.460 169.665 ;
        RECT 117.630 169.375 118.080 169.835 ;
        RECT 118.250 169.545 119.345 170.105 ;
        RECT 117.630 169.155 118.755 169.375 ;
        RECT 117.630 168.525 117.955 168.985 ;
        RECT 118.475 168.695 118.755 169.155 ;
        RECT 118.945 168.695 119.345 169.545 ;
        RECT 119.515 170.275 120.470 170.445 ;
        RECT 120.905 170.275 121.235 171.075 ;
        RECT 121.405 170.425 121.575 170.905 ;
        RECT 121.745 170.595 122.075 171.075 ;
        RECT 122.245 170.425 122.415 170.905 ;
        RECT 122.665 170.595 122.905 171.075 ;
        RECT 123.085 170.425 123.255 170.905 ;
        RECT 119.515 169.375 119.725 170.275 ;
        RECT 121.405 170.255 122.415 170.425 ;
        RECT 122.620 170.255 123.255 170.425 ;
        RECT 123.515 170.305 125.185 171.075 ;
        RECT 125.815 170.350 126.105 171.075 ;
        RECT 126.275 170.335 126.740 170.880 ;
        RECT 119.895 169.545 120.585 170.105 ;
        RECT 121.405 169.715 121.900 170.255 ;
        RECT 122.620 170.085 122.790 170.255 ;
        RECT 122.290 169.915 122.790 170.085 ;
        RECT 119.515 169.155 120.470 169.375 ;
        RECT 119.745 168.525 120.015 168.985 ;
        RECT 120.185 168.695 120.470 169.155 ;
        RECT 120.905 168.525 121.235 169.675 ;
        RECT 121.405 169.545 122.415 169.715 ;
        RECT 121.405 168.695 121.575 169.545 ;
        RECT 121.745 168.525 122.075 169.325 ;
        RECT 122.245 168.695 122.415 169.545 ;
        RECT 122.620 169.675 122.790 169.915 ;
        RECT 122.960 169.845 123.340 170.085 ;
        RECT 123.515 169.785 124.265 170.305 ;
        RECT 122.620 169.505 123.335 169.675 ;
        RECT 124.435 169.615 125.185 170.135 ;
        RECT 122.595 168.525 122.835 169.325 ;
        RECT 123.005 168.695 123.335 169.505 ;
        RECT 123.515 168.525 125.185 169.615 ;
        RECT 125.815 168.525 126.105 169.690 ;
        RECT 126.275 169.375 126.445 170.335 ;
        RECT 127.245 170.255 127.415 171.075 ;
        RECT 127.585 170.425 127.915 170.905 ;
        RECT 128.085 170.685 128.435 171.075 ;
        RECT 128.605 170.505 128.835 170.905 ;
        RECT 128.325 170.425 128.835 170.505 ;
        RECT 127.585 170.335 128.835 170.425 ;
        RECT 129.005 170.335 129.325 170.815 ;
        RECT 129.585 170.525 129.755 170.815 ;
        RECT 129.925 170.695 130.255 171.075 ;
        RECT 129.585 170.355 130.250 170.525 ;
        RECT 127.585 170.255 128.495 170.335 ;
        RECT 126.615 169.715 126.860 170.165 ;
        RECT 127.120 169.885 127.815 170.085 ;
        RECT 127.985 169.915 128.585 170.085 ;
        RECT 127.985 169.715 128.155 169.915 ;
        RECT 128.815 169.745 128.985 170.165 ;
        RECT 126.615 169.545 128.155 169.715 ;
        RECT 128.325 169.575 128.985 169.745 ;
        RECT 128.325 169.375 128.495 169.575 ;
        RECT 129.155 169.405 129.325 170.335 ;
        RECT 129.500 169.535 129.850 170.185 ;
        RECT 126.275 169.205 128.495 169.375 ;
        RECT 128.665 169.205 129.325 169.405 ;
        RECT 130.020 169.365 130.250 170.355 ;
        RECT 126.275 168.525 126.575 169.035 ;
        RECT 126.745 168.695 127.075 169.205 ;
        RECT 128.665 169.035 128.835 169.205 ;
        RECT 129.585 169.195 130.250 169.365 ;
        RECT 127.245 168.525 127.875 169.035 ;
        RECT 128.455 168.865 128.835 169.035 ;
        RECT 129.005 168.525 129.305 169.035 ;
        RECT 129.585 168.695 129.755 169.195 ;
        RECT 129.925 168.525 130.255 169.025 ;
        RECT 130.425 168.695 130.610 170.815 ;
        RECT 130.865 170.615 131.115 171.075 ;
        RECT 131.285 170.625 131.620 170.795 ;
        RECT 131.815 170.625 132.490 170.795 ;
        RECT 131.285 170.485 131.455 170.625 ;
        RECT 130.780 169.495 131.060 170.445 ;
        RECT 131.230 170.355 131.455 170.485 ;
        RECT 131.230 169.250 131.400 170.355 ;
        RECT 131.625 170.205 132.150 170.425 ;
        RECT 131.570 169.440 131.810 170.035 ;
        RECT 131.980 169.505 132.150 170.205 ;
        RECT 132.320 169.845 132.490 170.625 ;
        RECT 132.810 170.575 133.180 171.075 ;
        RECT 133.360 170.625 133.765 170.795 ;
        RECT 133.935 170.625 134.720 170.795 ;
        RECT 133.360 170.395 133.530 170.625 ;
        RECT 132.700 170.095 133.530 170.395 ;
        RECT 133.915 170.125 134.380 170.455 ;
        RECT 132.700 170.065 132.900 170.095 ;
        RECT 133.020 169.845 133.190 169.915 ;
        RECT 132.320 169.675 133.190 169.845 ;
        RECT 132.680 169.585 133.190 169.675 ;
        RECT 131.230 169.120 131.535 169.250 ;
        RECT 131.980 169.140 132.510 169.505 ;
        RECT 130.850 168.525 131.115 168.985 ;
        RECT 131.285 168.695 131.535 169.120 ;
        RECT 132.680 168.970 132.850 169.585 ;
        RECT 131.745 168.800 132.850 168.970 ;
        RECT 133.020 168.525 133.190 169.325 ;
        RECT 133.360 169.025 133.530 170.095 ;
        RECT 133.700 169.195 133.890 169.915 ;
        RECT 134.060 169.165 134.380 170.125 ;
        RECT 134.550 170.165 134.720 170.625 ;
        RECT 134.995 170.545 135.205 171.075 ;
        RECT 135.465 170.335 135.795 170.860 ;
        RECT 135.965 170.465 136.135 171.075 ;
        RECT 136.305 170.420 136.635 170.855 ;
        RECT 136.305 170.335 136.685 170.420 ;
        RECT 135.595 170.165 135.795 170.335 ;
        RECT 136.460 170.295 136.685 170.335 ;
        RECT 134.550 169.835 135.425 170.165 ;
        RECT 135.595 169.835 136.345 170.165 ;
        RECT 133.360 168.695 133.610 169.025 ;
        RECT 134.550 168.995 134.720 169.835 ;
        RECT 135.595 169.630 135.785 169.835 ;
        RECT 136.515 169.715 136.685 170.295 ;
        RECT 136.855 170.325 138.065 171.075 ;
        RECT 136.855 169.785 137.375 170.325 ;
        RECT 138.255 170.265 138.495 171.075 ;
        RECT 138.665 170.265 138.995 170.905 ;
        RECT 139.165 170.265 139.435 171.075 ;
        RECT 139.620 170.310 140.075 171.075 ;
        RECT 140.350 170.695 141.650 170.905 ;
        RECT 141.905 170.715 142.235 171.075 ;
        RECT 141.480 170.545 141.650 170.695 ;
        RECT 142.405 170.575 142.665 170.905 ;
        RECT 142.435 170.565 142.665 170.575 ;
        RECT 136.470 169.665 136.685 169.715 ;
        RECT 134.890 169.255 135.785 169.630 ;
        RECT 136.295 169.585 136.685 169.665 ;
        RECT 137.545 169.615 138.065 170.155 ;
        RECT 138.235 169.835 138.585 170.085 ;
        RECT 138.755 169.665 138.925 170.265 ;
        RECT 140.550 170.085 140.770 170.485 ;
        RECT 139.095 169.835 139.445 170.085 ;
        RECT 139.615 169.885 140.105 170.085 ;
        RECT 140.295 169.875 140.770 170.085 ;
        RECT 141.015 170.085 141.225 170.485 ;
        RECT 141.480 170.420 142.235 170.545 ;
        RECT 141.480 170.375 142.325 170.420 ;
        RECT 142.055 170.255 142.325 170.375 ;
        RECT 141.015 169.875 141.345 170.085 ;
        RECT 141.515 169.815 141.925 170.120 ;
        RECT 133.835 168.825 134.720 168.995 ;
        RECT 134.900 168.525 135.215 169.025 ;
        RECT 135.445 168.695 135.785 169.255 ;
        RECT 135.955 168.525 136.125 169.535 ;
        RECT 136.295 168.740 136.625 169.585 ;
        RECT 136.855 168.525 138.065 169.615 ;
        RECT 138.245 169.495 138.925 169.665 ;
        RECT 138.245 168.710 138.575 169.495 ;
        RECT 139.105 168.525 139.435 169.665 ;
        RECT 139.620 169.645 140.795 169.705 ;
        RECT 142.155 169.680 142.325 170.255 ;
        RECT 142.125 169.645 142.325 169.680 ;
        RECT 139.620 169.535 142.325 169.645 ;
        RECT 139.620 168.915 139.875 169.535 ;
        RECT 140.465 169.475 142.265 169.535 ;
        RECT 140.465 169.445 140.795 169.475 ;
        RECT 142.495 169.375 142.665 170.565 ;
        RECT 142.835 170.325 144.045 171.075 ;
        RECT 144.215 170.350 144.475 170.905 ;
        RECT 144.645 170.630 145.075 171.075 ;
        RECT 145.310 170.505 145.480 170.905 ;
        RECT 145.650 170.675 146.370 171.075 ;
        RECT 142.835 169.785 143.355 170.325 ;
        RECT 143.525 169.615 144.045 170.155 ;
        RECT 140.125 169.275 140.310 169.365 ;
        RECT 140.900 169.275 141.735 169.285 ;
        RECT 140.125 169.075 141.735 169.275 ;
        RECT 140.125 169.035 140.355 169.075 ;
        RECT 139.620 168.695 139.955 168.915 ;
        RECT 140.960 168.525 141.315 168.905 ;
        RECT 141.485 168.695 141.735 169.075 ;
        RECT 141.985 168.525 142.235 169.305 ;
        RECT 142.405 168.695 142.665 169.375 ;
        RECT 142.835 168.525 144.045 169.615 ;
        RECT 144.215 169.635 144.390 170.350 ;
        RECT 145.310 170.335 146.190 170.505 ;
        RECT 146.540 170.460 146.710 170.905 ;
        RECT 147.285 170.565 147.685 171.075 ;
        RECT 144.560 169.835 144.815 170.165 ;
        RECT 144.215 168.695 144.475 169.635 ;
        RECT 144.645 169.355 144.815 169.835 ;
        RECT 145.040 169.545 145.370 170.165 ;
        RECT 145.540 169.785 145.830 170.165 ;
        RECT 146.020 169.615 146.190 170.335 ;
        RECT 145.670 169.445 146.190 169.615 ;
        RECT 146.360 170.290 146.710 170.460 ;
        RECT 147.895 170.425 148.155 170.905 ;
        RECT 148.325 170.535 148.575 171.075 ;
        RECT 144.645 169.185 145.405 169.355 ;
        RECT 145.670 169.255 145.840 169.445 ;
        RECT 146.360 169.265 146.530 170.290 ;
        RECT 146.950 169.805 147.210 170.395 ;
        RECT 146.730 169.505 147.210 169.805 ;
        RECT 147.410 169.505 147.670 170.395 ;
        RECT 147.895 169.395 148.065 170.425 ;
        RECT 148.745 170.370 148.965 170.855 ;
        RECT 148.235 169.775 148.465 170.170 ;
        RECT 148.635 169.945 148.965 170.370 ;
        RECT 149.135 170.695 150.025 170.865 ;
        RECT 149.135 169.970 149.305 170.695 ;
        RECT 149.475 170.140 150.025 170.525 ;
        RECT 150.255 170.255 150.465 171.075 ;
        RECT 150.635 170.275 150.965 170.905 ;
        RECT 149.135 169.900 150.025 169.970 ;
        RECT 149.130 169.875 150.025 169.900 ;
        RECT 149.120 169.860 150.025 169.875 ;
        RECT 149.115 169.845 150.025 169.860 ;
        RECT 149.105 169.840 150.025 169.845 ;
        RECT 149.100 169.830 150.025 169.840 ;
        RECT 149.095 169.820 150.025 169.830 ;
        RECT 149.085 169.815 150.025 169.820 ;
        RECT 149.075 169.805 150.025 169.815 ;
        RECT 149.065 169.800 150.025 169.805 ;
        RECT 149.065 169.795 149.400 169.800 ;
        RECT 149.050 169.790 149.400 169.795 ;
        RECT 149.035 169.780 149.400 169.790 ;
        RECT 149.010 169.775 149.400 169.780 ;
        RECT 148.235 169.770 149.400 169.775 ;
        RECT 148.235 169.735 149.370 169.770 ;
        RECT 148.235 169.710 149.335 169.735 ;
        RECT 148.235 169.680 149.305 169.710 ;
        RECT 148.235 169.650 149.285 169.680 ;
        RECT 148.235 169.620 149.265 169.650 ;
        RECT 148.235 169.610 149.195 169.620 ;
        RECT 148.235 169.600 149.170 169.610 ;
        RECT 148.235 169.585 149.150 169.600 ;
        RECT 148.235 169.570 149.130 169.585 ;
        RECT 148.340 169.560 149.125 169.570 ;
        RECT 148.340 169.525 149.110 169.560 ;
        RECT 145.235 168.960 145.405 169.185 ;
        RECT 146.120 169.095 146.530 169.265 ;
        RECT 146.705 169.155 147.645 169.325 ;
        RECT 146.120 168.960 146.375 169.095 ;
        RECT 144.645 168.525 144.975 168.925 ;
        RECT 145.235 168.790 146.375 168.960 ;
        RECT 146.705 168.905 146.875 169.155 ;
        RECT 146.120 168.695 146.375 168.790 ;
        RECT 146.545 168.735 146.875 168.905 ;
        RECT 147.045 168.525 147.295 168.985 ;
        RECT 147.465 168.695 147.645 169.155 ;
        RECT 147.895 168.695 148.170 169.395 ;
        RECT 148.340 169.275 149.095 169.525 ;
        RECT 149.265 169.205 149.595 169.450 ;
        RECT 149.765 169.350 150.025 169.800 ;
        RECT 150.635 169.675 150.885 170.275 ;
        RECT 151.135 170.255 151.365 171.075 ;
        RECT 151.575 170.350 151.865 171.075 ;
        RECT 152.200 170.565 152.440 171.075 ;
        RECT 152.620 170.565 152.900 170.895 ;
        RECT 153.130 170.565 153.345 171.075 ;
        RECT 151.055 169.835 151.385 170.085 ;
        RECT 152.095 169.835 152.450 170.395 ;
        RECT 149.410 169.180 149.595 169.205 ;
        RECT 149.410 169.080 150.025 169.180 ;
        RECT 148.340 168.525 148.595 169.070 ;
        RECT 148.765 168.695 149.245 169.035 ;
        RECT 149.420 168.525 150.025 169.080 ;
        RECT 150.255 168.525 150.465 169.665 ;
        RECT 150.635 168.695 150.965 169.675 ;
        RECT 151.135 168.525 151.365 169.665 ;
        RECT 151.575 168.525 151.865 169.690 ;
        RECT 152.620 169.665 152.790 170.565 ;
        RECT 152.960 169.835 153.225 170.395 ;
        RECT 153.515 170.335 154.130 170.905 ;
        RECT 153.475 169.665 153.645 170.165 ;
        RECT 152.220 169.495 153.645 169.665 ;
        RECT 152.220 169.320 152.610 169.495 ;
        RECT 153.095 168.525 153.425 169.325 ;
        RECT 153.815 169.315 154.130 170.335 ;
        RECT 154.375 170.255 154.605 171.075 ;
        RECT 154.775 170.275 155.105 170.905 ;
        RECT 154.355 169.835 154.685 170.085 ;
        RECT 154.855 169.675 155.105 170.275 ;
        RECT 155.275 170.255 155.485 171.075 ;
        RECT 155.715 170.325 156.925 171.075 ;
        RECT 153.595 168.695 154.130 169.315 ;
        RECT 154.375 168.525 154.605 169.665 ;
        RECT 154.775 168.695 155.105 169.675 ;
        RECT 155.275 168.525 155.485 169.665 ;
        RECT 155.715 169.615 156.235 170.155 ;
        RECT 156.405 169.785 156.925 170.325 ;
        RECT 155.715 168.525 156.925 169.615 ;
        RECT 22.690 168.355 157.010 168.525 ;
        RECT 22.775 167.265 23.985 168.355 ;
        RECT 24.245 167.685 24.415 168.185 ;
        RECT 24.585 167.855 24.915 168.355 ;
        RECT 24.245 167.515 24.910 167.685 ;
        RECT 22.775 166.555 23.295 167.095 ;
        RECT 23.465 166.725 23.985 167.265 ;
        RECT 24.160 166.695 24.510 167.345 ;
        RECT 22.775 165.805 23.985 166.555 ;
        RECT 24.680 166.525 24.910 167.515 ;
        RECT 24.245 166.355 24.910 166.525 ;
        RECT 24.245 166.065 24.415 166.355 ;
        RECT 24.585 165.805 24.915 166.185 ;
        RECT 25.085 166.065 25.270 168.185 ;
        RECT 25.510 167.895 25.775 168.355 ;
        RECT 25.945 167.760 26.195 168.185 ;
        RECT 26.405 167.910 27.510 168.080 ;
        RECT 25.890 167.630 26.195 167.760 ;
        RECT 25.440 166.435 25.720 167.385 ;
        RECT 25.890 166.525 26.060 167.630 ;
        RECT 26.230 166.845 26.470 167.440 ;
        RECT 26.640 167.375 27.170 167.740 ;
        RECT 26.640 166.675 26.810 167.375 ;
        RECT 27.340 167.295 27.510 167.910 ;
        RECT 27.680 167.555 27.850 168.355 ;
        RECT 28.020 167.855 28.270 168.185 ;
        RECT 28.495 167.885 29.380 168.055 ;
        RECT 27.340 167.205 27.850 167.295 ;
        RECT 25.890 166.395 26.115 166.525 ;
        RECT 26.285 166.455 26.810 166.675 ;
        RECT 26.980 167.035 27.850 167.205 ;
        RECT 25.525 165.805 25.775 166.265 ;
        RECT 25.945 166.255 26.115 166.395 ;
        RECT 26.980 166.255 27.150 167.035 ;
        RECT 27.680 166.965 27.850 167.035 ;
        RECT 27.360 166.785 27.560 166.815 ;
        RECT 28.020 166.785 28.190 167.855 ;
        RECT 28.360 166.965 28.550 167.685 ;
        RECT 27.360 166.485 28.190 166.785 ;
        RECT 28.720 166.755 29.040 167.715 ;
        RECT 25.945 166.085 26.280 166.255 ;
        RECT 26.475 166.085 27.150 166.255 ;
        RECT 27.470 165.805 27.840 166.305 ;
        RECT 28.020 166.255 28.190 166.485 ;
        RECT 28.575 166.425 29.040 166.755 ;
        RECT 29.210 167.045 29.380 167.885 ;
        RECT 29.560 167.855 29.875 168.355 ;
        RECT 30.105 167.625 30.445 168.185 ;
        RECT 29.550 167.250 30.445 167.625 ;
        RECT 30.615 167.345 30.785 168.355 ;
        RECT 30.255 167.045 30.445 167.250 ;
        RECT 30.955 167.295 31.285 168.140 ;
        RECT 31.515 167.485 31.790 168.185 ;
        RECT 32.000 167.810 32.215 168.355 ;
        RECT 32.385 167.845 32.860 168.185 ;
        RECT 33.030 167.850 33.645 168.355 ;
        RECT 33.030 167.675 33.225 167.850 ;
        RECT 30.955 167.215 31.345 167.295 ;
        RECT 31.130 167.165 31.345 167.215 ;
        RECT 29.210 166.715 30.085 167.045 ;
        RECT 30.255 166.715 31.005 167.045 ;
        RECT 29.210 166.255 29.380 166.715 ;
        RECT 30.255 166.545 30.455 166.715 ;
        RECT 31.175 166.585 31.345 167.165 ;
        RECT 31.120 166.545 31.345 166.585 ;
        RECT 28.020 166.085 28.425 166.255 ;
        RECT 28.595 166.085 29.380 166.255 ;
        RECT 29.655 165.805 29.865 166.335 ;
        RECT 30.125 166.020 30.455 166.545 ;
        RECT 30.965 166.460 31.345 166.545 ;
        RECT 30.625 165.805 30.795 166.415 ;
        RECT 30.965 166.025 31.295 166.460 ;
        RECT 31.515 166.455 31.685 167.485 ;
        RECT 31.960 167.315 32.675 167.610 ;
        RECT 32.895 167.485 33.225 167.675 ;
        RECT 33.395 167.315 33.645 167.680 ;
        RECT 31.855 167.145 33.645 167.315 ;
        RECT 31.855 166.715 32.085 167.145 ;
        RECT 31.515 165.975 31.775 166.455 ;
        RECT 32.255 166.445 32.665 166.965 ;
        RECT 31.945 165.805 32.275 166.265 ;
        RECT 32.465 166.025 32.665 166.445 ;
        RECT 32.835 166.290 33.090 167.145 ;
        RECT 33.885 166.965 34.055 168.185 ;
        RECT 34.305 167.845 34.565 168.355 ;
        RECT 33.260 166.715 34.055 166.965 ;
        RECT 34.225 166.795 34.565 167.675 ;
        RECT 35.655 167.190 35.945 168.355 ;
        RECT 37.125 167.685 37.295 168.185 ;
        RECT 37.465 167.855 37.795 168.355 ;
        RECT 37.125 167.515 37.790 167.685 ;
        RECT 33.805 166.625 34.055 166.715 ;
        RECT 37.040 166.695 37.390 167.345 ;
        RECT 32.835 166.025 33.625 166.290 ;
        RECT 33.805 166.205 34.135 166.625 ;
        RECT 34.305 165.805 34.565 166.625 ;
        RECT 35.655 165.805 35.945 166.530 ;
        RECT 37.560 166.525 37.790 167.515 ;
        RECT 37.125 166.355 37.790 166.525 ;
        RECT 37.125 166.065 37.295 166.355 ;
        RECT 37.465 165.805 37.795 166.185 ;
        RECT 37.965 166.065 38.150 168.185 ;
        RECT 38.390 167.895 38.655 168.355 ;
        RECT 38.825 167.760 39.075 168.185 ;
        RECT 39.285 167.910 40.390 168.080 ;
        RECT 38.770 167.630 39.075 167.760 ;
        RECT 38.320 166.435 38.600 167.385 ;
        RECT 38.770 166.525 38.940 167.630 ;
        RECT 39.110 166.845 39.350 167.440 ;
        RECT 39.520 167.375 40.050 167.740 ;
        RECT 39.520 166.675 39.690 167.375 ;
        RECT 40.220 167.295 40.390 167.910 ;
        RECT 40.560 167.555 40.730 168.355 ;
        RECT 40.900 167.855 41.150 168.185 ;
        RECT 41.375 167.885 42.260 168.055 ;
        RECT 40.220 167.205 40.730 167.295 ;
        RECT 38.770 166.395 38.995 166.525 ;
        RECT 39.165 166.455 39.690 166.675 ;
        RECT 39.860 167.035 40.730 167.205 ;
        RECT 38.405 165.805 38.655 166.265 ;
        RECT 38.825 166.255 38.995 166.395 ;
        RECT 39.860 166.255 40.030 167.035 ;
        RECT 40.560 166.965 40.730 167.035 ;
        RECT 40.240 166.785 40.440 166.815 ;
        RECT 40.900 166.785 41.070 167.855 ;
        RECT 41.240 166.965 41.430 167.685 ;
        RECT 40.240 166.485 41.070 166.785 ;
        RECT 41.600 166.755 41.920 167.715 ;
        RECT 38.825 166.085 39.160 166.255 ;
        RECT 39.355 166.085 40.030 166.255 ;
        RECT 40.350 165.805 40.720 166.305 ;
        RECT 40.900 166.255 41.070 166.485 ;
        RECT 41.455 166.425 41.920 166.755 ;
        RECT 42.090 167.045 42.260 167.885 ;
        RECT 42.440 167.855 42.755 168.355 ;
        RECT 42.985 167.625 43.325 168.185 ;
        RECT 42.430 167.250 43.325 167.625 ;
        RECT 43.495 167.345 43.665 168.355 ;
        RECT 43.135 167.045 43.325 167.250 ;
        RECT 43.835 167.295 44.165 168.140 ;
        RECT 44.405 167.295 44.735 168.145 ;
        RECT 43.835 167.215 44.225 167.295 ;
        RECT 44.010 167.165 44.225 167.215 ;
        RECT 42.090 166.715 42.965 167.045 ;
        RECT 43.135 166.715 43.885 167.045 ;
        RECT 42.090 166.255 42.260 166.715 ;
        RECT 43.135 166.545 43.335 166.715 ;
        RECT 44.055 166.585 44.225 167.165 ;
        RECT 44.000 166.545 44.225 166.585 ;
        RECT 40.900 166.085 41.305 166.255 ;
        RECT 41.475 166.085 42.260 166.255 ;
        RECT 42.535 165.805 42.745 166.335 ;
        RECT 43.005 166.020 43.335 166.545 ;
        RECT 43.845 166.460 44.225 166.545 ;
        RECT 44.405 166.530 44.595 167.295 ;
        RECT 44.905 167.215 45.155 168.355 ;
        RECT 45.345 167.715 45.595 168.135 ;
        RECT 45.825 167.885 46.155 168.355 ;
        RECT 46.385 167.715 46.635 168.135 ;
        RECT 45.345 167.545 46.635 167.715 ;
        RECT 46.815 167.715 47.145 168.145 ;
        RECT 46.815 167.545 47.270 167.715 ;
        RECT 45.335 167.045 45.550 167.375 ;
        RECT 44.765 166.715 45.075 167.045 ;
        RECT 45.245 166.715 45.550 167.045 ;
        RECT 45.725 166.715 46.010 167.375 ;
        RECT 46.205 166.715 46.470 167.375 ;
        RECT 46.685 166.715 46.930 167.375 ;
        RECT 44.905 166.545 45.075 166.715 ;
        RECT 47.100 166.545 47.270 167.545 ;
        RECT 47.615 167.265 48.825 168.355 ;
        RECT 49.080 167.735 49.255 168.185 ;
        RECT 49.425 167.915 49.755 168.355 ;
        RECT 50.060 167.765 50.230 168.185 ;
        RECT 50.465 167.945 51.135 168.355 ;
        RECT 51.350 167.765 51.520 168.185 ;
        RECT 51.720 167.945 52.050 168.355 ;
        RECT 49.080 167.565 49.710 167.735 ;
        RECT 43.505 165.805 43.675 166.415 ;
        RECT 43.845 166.025 44.175 166.460 ;
        RECT 44.405 166.020 44.735 166.530 ;
        RECT 44.905 166.375 47.270 166.545 ;
        RECT 47.615 166.555 48.135 167.095 ;
        RECT 48.305 166.725 48.825 167.265 ;
        RECT 48.995 166.715 49.360 167.395 ;
        RECT 49.540 167.045 49.710 167.565 ;
        RECT 50.060 167.595 52.075 167.765 ;
        RECT 49.540 166.715 49.890 167.045 ;
        RECT 44.905 165.805 45.235 166.205 ;
        RECT 46.285 166.035 46.615 166.375 ;
        RECT 46.785 165.805 47.115 166.205 ;
        RECT 47.615 165.805 48.825 166.555 ;
        RECT 49.540 166.545 49.710 166.715 ;
        RECT 49.080 166.375 49.710 166.545 ;
        RECT 49.080 165.975 49.255 166.375 ;
        RECT 50.060 166.305 50.230 167.595 ;
        RECT 49.425 165.805 49.755 166.185 ;
        RECT 50.000 165.975 50.230 166.305 ;
        RECT 50.430 166.140 50.710 167.415 ;
        RECT 50.935 167.335 51.205 167.415 ;
        RECT 50.895 167.165 51.205 167.335 ;
        RECT 50.935 166.140 51.205 167.165 ;
        RECT 51.395 166.385 51.735 167.415 ;
        RECT 51.905 167.045 52.075 167.595 ;
        RECT 52.245 167.215 52.505 168.185 ;
        RECT 51.905 166.715 52.165 167.045 ;
        RECT 52.335 166.525 52.505 167.215 ;
        RECT 51.665 165.805 51.995 166.185 ;
        RECT 52.165 166.060 52.505 166.525 ;
        RECT 52.675 167.215 52.945 168.185 ;
        RECT 53.155 167.555 53.435 168.355 ;
        RECT 53.615 167.805 54.810 168.135 ;
        RECT 53.940 167.385 54.360 167.635 ;
        RECT 53.115 167.215 54.360 167.385 ;
        RECT 52.675 166.480 52.845 167.215 ;
        RECT 53.115 167.045 53.285 167.215 ;
        RECT 54.585 167.045 54.755 167.605 ;
        RECT 55.005 167.215 55.260 168.355 ;
        RECT 55.650 167.555 55.865 168.355 ;
        RECT 56.155 167.385 56.485 168.185 ;
        RECT 56.655 167.555 56.940 168.355 ;
        RECT 57.110 167.385 57.440 168.185 ;
        RECT 55.435 167.215 57.440 167.385 ;
        RECT 57.610 167.215 57.860 168.355 ;
        RECT 58.060 167.315 58.485 167.645 ;
        RECT 53.055 166.715 53.285 167.045 ;
        RECT 54.015 166.715 54.755 167.045 ;
        RECT 54.925 166.795 55.260 167.045 ;
        RECT 53.115 166.545 53.285 166.715 ;
        RECT 54.505 166.625 54.755 166.715 ;
        RECT 52.675 166.135 52.945 166.480 ;
        RECT 53.115 166.375 53.855 166.545 ;
        RECT 54.505 166.455 55.240 166.625 ;
        RECT 52.165 166.015 52.500 166.060 ;
        RECT 53.135 165.805 53.515 166.205 ;
        RECT 53.685 166.025 53.855 166.375 ;
        RECT 54.025 165.805 54.760 166.285 ;
        RECT 54.930 165.985 55.240 166.455 ;
        RECT 55.435 166.545 55.645 167.215 ;
        RECT 55.815 166.715 56.215 167.045 ;
        RECT 55.435 165.975 55.875 166.545 ;
        RECT 56.045 166.315 56.215 166.715 ;
        RECT 56.385 166.485 56.645 167.045 ;
        RECT 56.815 166.485 57.065 167.045 ;
        RECT 57.335 166.715 57.605 167.045 ;
        RECT 57.795 166.715 58.145 167.045 ;
        RECT 58.315 166.545 58.485 167.315 ;
        RECT 58.655 167.265 61.245 168.355 ;
        RECT 57.235 166.375 58.485 166.545 ;
        RECT 57.235 166.315 57.415 166.375 ;
        RECT 56.045 166.145 57.415 166.315 ;
        RECT 57.585 165.805 57.915 166.205 ;
        RECT 58.095 166.165 58.485 166.375 ;
        RECT 58.655 166.575 59.865 167.095 ;
        RECT 60.035 166.745 61.245 167.265 ;
        RECT 61.415 167.190 61.705 168.355 ;
        RECT 61.875 167.265 64.465 168.355 ;
        RECT 65.100 167.355 65.355 168.355 ;
        RECT 61.875 166.575 63.085 167.095 ;
        RECT 63.255 166.745 64.465 167.265 ;
        RECT 58.655 165.805 61.245 166.575 ;
        RECT 61.415 165.805 61.705 166.530 ;
        RECT 61.875 165.805 64.465 166.575 ;
        RECT 65.115 165.805 65.355 166.605 ;
        RECT 65.540 165.975 65.785 168.185 ;
        RECT 65.955 167.905 66.805 168.355 ;
        RECT 66.975 167.725 67.235 168.185 ;
        RECT 66.115 167.505 67.235 167.725 ;
        RECT 66.115 167.050 66.285 167.505 ;
        RECT 67.415 167.335 67.620 167.705 ;
        RECT 67.805 167.370 68.130 168.355 ;
        RECT 65.955 166.560 66.285 167.050 ;
        RECT 66.455 166.730 66.865 167.335 ;
        RECT 67.415 167.165 67.625 167.335 ;
        RECT 68.315 167.215 68.700 168.185 ;
        RECT 68.870 167.895 69.195 168.355 ;
        RECT 69.715 167.725 69.995 168.185 ;
        RECT 68.870 167.505 69.995 167.725 ;
        RECT 67.415 167.120 67.620 167.165 ;
        RECT 67.035 166.745 67.620 167.120 ;
        RECT 67.875 166.715 68.135 167.170 ;
        RECT 65.955 166.355 66.805 166.560 ;
        RECT 68.315 166.545 68.595 167.215 ;
        RECT 68.870 167.045 69.320 167.505 ;
        RECT 70.185 167.335 70.585 168.185 ;
        RECT 70.985 167.895 71.255 168.355 ;
        RECT 71.425 167.725 71.710 168.185 ;
        RECT 68.765 166.715 69.320 167.045 ;
        RECT 69.490 166.775 70.585 167.335 ;
        RECT 68.870 166.605 69.320 166.715 ;
        RECT 65.955 165.805 66.285 166.185 ;
        RECT 66.475 165.975 66.805 166.355 ;
        RECT 66.975 166.355 68.130 166.545 ;
        RECT 66.975 166.185 67.185 166.355 ;
        RECT 67.855 166.215 68.130 166.355 ;
        RECT 67.355 165.805 67.685 166.185 ;
        RECT 68.315 165.975 68.700 166.545 ;
        RECT 68.870 166.435 69.995 166.605 ;
        RECT 68.870 165.805 69.195 166.265 ;
        RECT 69.715 165.975 69.995 166.435 ;
        RECT 70.185 165.975 70.585 166.775 ;
        RECT 70.755 167.505 71.710 167.725 ;
        RECT 70.755 166.605 70.965 167.505 ;
        RECT 71.135 166.775 71.825 167.335 ;
        RECT 71.995 167.265 73.665 168.355 ;
        RECT 73.925 167.610 74.195 168.355 ;
        RECT 74.825 168.350 81.100 168.355 ;
        RECT 74.365 167.440 74.655 168.180 ;
        RECT 74.825 167.625 75.080 168.350 ;
        RECT 75.265 167.455 75.525 168.180 ;
        RECT 75.695 167.625 75.940 168.350 ;
        RECT 76.125 167.455 76.385 168.180 ;
        RECT 76.555 167.625 76.800 168.350 ;
        RECT 76.985 167.455 77.245 168.180 ;
        RECT 77.415 167.625 77.660 168.350 ;
        RECT 77.830 167.455 78.090 168.180 ;
        RECT 78.260 167.625 78.520 168.350 ;
        RECT 78.690 167.455 78.950 168.180 ;
        RECT 79.120 167.625 79.380 168.350 ;
        RECT 79.550 167.455 79.810 168.180 ;
        RECT 79.980 167.625 80.240 168.350 ;
        RECT 80.410 167.455 80.670 168.180 ;
        RECT 80.840 167.555 81.100 168.350 ;
        RECT 75.265 167.440 80.670 167.455 ;
        RECT 70.755 166.435 71.710 166.605 ;
        RECT 70.985 165.805 71.255 166.265 ;
        RECT 71.425 165.975 71.710 166.435 ;
        RECT 71.995 166.575 72.745 167.095 ;
        RECT 72.915 166.745 73.665 167.265 ;
        RECT 73.925 167.215 80.670 167.440 ;
        RECT 73.925 166.625 75.090 167.215 ;
        RECT 81.270 167.045 81.520 168.180 ;
        RECT 81.700 167.545 81.960 168.355 ;
        RECT 82.135 167.045 82.380 168.185 ;
        RECT 82.560 167.545 82.855 168.355 ;
        RECT 83.075 168.015 84.215 168.185 ;
        RECT 83.075 167.555 83.375 168.015 ;
        RECT 83.545 167.385 83.875 167.845 ;
        RECT 83.115 167.335 83.875 167.385 ;
        RECT 83.095 167.165 83.875 167.335 ;
        RECT 84.045 167.385 84.215 168.015 ;
        RECT 84.385 167.555 84.715 168.355 ;
        RECT 84.885 167.385 85.160 168.185 ;
        RECT 84.045 167.175 85.160 167.385 ;
        RECT 85.335 167.265 87.005 168.355 ;
        RECT 75.260 166.795 82.380 167.045 ;
        RECT 71.995 165.805 73.665 166.575 ;
        RECT 73.925 166.455 80.670 166.625 ;
        RECT 73.925 165.805 74.225 166.285 ;
        RECT 74.395 166.000 74.655 166.455 ;
        RECT 74.825 165.805 75.085 166.285 ;
        RECT 75.265 166.000 75.525 166.455 ;
        RECT 75.695 165.805 75.945 166.285 ;
        RECT 76.125 166.000 76.385 166.455 ;
        RECT 76.555 165.805 76.805 166.285 ;
        RECT 76.985 166.000 77.245 166.455 ;
        RECT 77.415 165.805 77.660 166.285 ;
        RECT 77.830 166.000 78.105 166.455 ;
        RECT 78.275 165.805 78.520 166.285 ;
        RECT 78.690 166.000 78.950 166.455 ;
        RECT 79.120 165.805 79.380 166.285 ;
        RECT 79.550 166.000 79.810 166.455 ;
        RECT 79.980 165.805 80.240 166.285 ;
        RECT 80.410 166.000 80.670 166.455 ;
        RECT 80.840 165.805 81.100 166.365 ;
        RECT 81.270 165.985 81.520 166.795 ;
        RECT 81.700 165.805 81.960 166.330 ;
        RECT 82.130 165.985 82.380 166.795 ;
        RECT 82.550 166.485 82.865 167.045 ;
        RECT 83.115 166.625 83.330 167.165 ;
        RECT 83.500 166.795 84.270 166.995 ;
        RECT 84.440 166.795 85.160 166.995 ;
        RECT 83.115 166.455 84.715 166.625 ;
        RECT 83.545 166.445 84.715 166.455 ;
        RECT 82.560 165.805 82.865 166.315 ;
        RECT 83.085 165.805 83.375 166.275 ;
        RECT 83.545 165.975 83.875 166.445 ;
        RECT 84.045 165.805 84.215 166.275 ;
        RECT 84.385 165.975 84.715 166.445 ;
        RECT 84.885 165.805 85.160 166.625 ;
        RECT 85.335 166.575 86.085 167.095 ;
        RECT 86.255 166.745 87.005 167.265 ;
        RECT 87.175 167.190 87.465 168.355 ;
        RECT 87.635 167.800 88.240 168.355 ;
        RECT 88.415 167.845 88.895 168.185 ;
        RECT 89.065 167.810 89.320 168.355 ;
        RECT 87.635 167.700 88.250 167.800 ;
        RECT 88.065 167.675 88.250 167.700 ;
        RECT 87.635 167.080 87.895 167.530 ;
        RECT 88.065 167.430 88.395 167.675 ;
        RECT 88.565 167.355 89.320 167.605 ;
        RECT 89.490 167.485 89.765 168.185 ;
        RECT 88.550 167.320 89.320 167.355 ;
        RECT 88.535 167.310 89.320 167.320 ;
        RECT 88.530 167.295 89.425 167.310 ;
        RECT 88.510 167.280 89.425 167.295 ;
        RECT 88.490 167.270 89.425 167.280 ;
        RECT 88.465 167.260 89.425 167.270 ;
        RECT 88.395 167.230 89.425 167.260 ;
        RECT 88.375 167.200 89.425 167.230 ;
        RECT 88.355 167.170 89.425 167.200 ;
        RECT 88.325 167.145 89.425 167.170 ;
        RECT 88.290 167.110 89.425 167.145 ;
        RECT 88.260 167.105 89.425 167.110 ;
        RECT 88.260 167.100 88.650 167.105 ;
        RECT 88.260 167.090 88.625 167.100 ;
        RECT 88.260 167.085 88.610 167.090 ;
        RECT 88.260 167.080 88.595 167.085 ;
        RECT 87.635 167.075 88.595 167.080 ;
        RECT 87.635 167.065 88.585 167.075 ;
        RECT 87.635 167.060 88.575 167.065 ;
        RECT 87.635 167.050 88.565 167.060 ;
        RECT 87.635 167.040 88.560 167.050 ;
        RECT 87.635 167.035 88.555 167.040 ;
        RECT 87.635 167.020 88.545 167.035 ;
        RECT 87.635 167.005 88.540 167.020 ;
        RECT 87.635 166.980 88.530 167.005 ;
        RECT 87.635 166.910 88.525 166.980 ;
        RECT 85.335 165.805 87.005 166.575 ;
        RECT 87.175 165.805 87.465 166.530 ;
        RECT 87.635 166.355 88.185 166.740 ;
        RECT 88.355 166.185 88.525 166.910 ;
        RECT 87.635 166.015 88.525 166.185 ;
        RECT 88.695 166.510 89.025 166.935 ;
        RECT 89.195 166.710 89.425 167.105 ;
        RECT 88.695 166.025 88.915 166.510 ;
        RECT 89.595 166.455 89.765 167.485 ;
        RECT 89.945 167.385 90.275 168.185 ;
        RECT 90.445 167.555 90.675 168.355 ;
        RECT 90.845 167.385 91.175 168.185 ;
        RECT 89.945 167.215 91.175 167.385 ;
        RECT 91.345 167.215 91.600 168.355 ;
        RECT 91.775 167.920 97.120 168.355 ;
        RECT 89.935 166.715 90.245 167.045 ;
        RECT 89.085 165.805 89.335 166.345 ;
        RECT 89.505 165.975 89.765 166.455 ;
        RECT 89.945 166.315 90.275 166.545 ;
        RECT 90.450 166.485 90.825 167.045 ;
        RECT 90.995 166.315 91.175 167.215 ;
        RECT 91.360 166.465 91.580 167.045 ;
        RECT 93.360 166.350 93.700 167.180 ;
        RECT 95.180 166.670 95.530 167.920 ;
        RECT 97.295 167.265 100.805 168.355 ;
        RECT 100.975 167.265 102.185 168.355 ;
        RECT 102.470 167.725 102.755 168.185 ;
        RECT 102.925 167.895 103.195 168.355 ;
        RECT 102.470 167.505 103.425 167.725 ;
        RECT 97.295 166.575 98.945 167.095 ;
        RECT 99.115 166.745 100.805 167.265 ;
        RECT 89.945 165.975 91.175 166.315 ;
        RECT 91.345 165.805 91.600 166.295 ;
        RECT 91.775 165.805 97.120 166.350 ;
        RECT 97.295 165.805 100.805 166.575 ;
        RECT 100.975 166.555 101.495 167.095 ;
        RECT 101.665 166.725 102.185 167.265 ;
        RECT 102.355 166.775 103.045 167.335 ;
        RECT 103.215 166.605 103.425 167.505 ;
        RECT 100.975 165.805 102.185 166.555 ;
        RECT 102.470 166.435 103.425 166.605 ;
        RECT 103.595 167.335 103.995 168.185 ;
        RECT 104.185 167.725 104.465 168.185 ;
        RECT 104.985 167.895 105.310 168.355 ;
        RECT 104.185 167.505 105.310 167.725 ;
        RECT 103.595 166.775 104.690 167.335 ;
        RECT 104.860 167.045 105.310 167.505 ;
        RECT 105.480 167.215 105.865 168.185 ;
        RECT 102.470 165.975 102.755 166.435 ;
        RECT 102.925 165.805 103.195 166.265 ;
        RECT 103.595 165.975 103.995 166.775 ;
        RECT 104.860 166.715 105.415 167.045 ;
        RECT 104.860 166.605 105.310 166.715 ;
        RECT 104.185 166.435 105.310 166.605 ;
        RECT 105.585 166.545 105.865 167.215 ;
        RECT 104.185 165.975 104.465 166.435 ;
        RECT 104.985 165.805 105.310 166.265 ;
        RECT 105.480 165.975 105.865 166.545 ;
        RECT 106.035 167.505 106.295 168.185 ;
        RECT 106.465 167.575 106.715 168.355 ;
        RECT 106.965 167.805 107.215 168.185 ;
        RECT 107.385 167.975 107.740 168.355 ;
        RECT 108.745 167.965 109.080 168.185 ;
        RECT 108.345 167.805 108.575 167.845 ;
        RECT 106.965 167.605 108.575 167.805 ;
        RECT 106.965 167.595 107.800 167.605 ;
        RECT 108.390 167.515 108.575 167.605 ;
        RECT 106.035 166.305 106.205 167.505 ;
        RECT 107.905 167.405 108.235 167.435 ;
        RECT 106.435 167.345 108.235 167.405 ;
        RECT 108.825 167.345 109.080 167.965 ;
        RECT 106.375 167.235 109.080 167.345 ;
        RECT 106.375 167.200 106.575 167.235 ;
        RECT 106.375 166.625 106.545 167.200 ;
        RECT 107.905 167.175 109.080 167.235 ;
        RECT 109.255 167.505 109.515 168.185 ;
        RECT 109.685 167.575 109.935 168.355 ;
        RECT 110.185 167.805 110.435 168.185 ;
        RECT 110.605 167.975 110.960 168.355 ;
        RECT 111.965 167.965 112.300 168.185 ;
        RECT 111.565 167.805 111.795 167.845 ;
        RECT 110.185 167.605 111.795 167.805 ;
        RECT 110.185 167.595 111.020 167.605 ;
        RECT 111.610 167.515 111.795 167.605 ;
        RECT 106.775 166.760 107.185 167.065 ;
        RECT 107.355 166.795 107.685 167.005 ;
        RECT 106.375 166.505 106.645 166.625 ;
        RECT 106.375 166.460 107.220 166.505 ;
        RECT 106.465 166.335 107.220 166.460 ;
        RECT 107.475 166.395 107.685 166.795 ;
        RECT 107.930 166.795 108.405 167.005 ;
        RECT 108.595 166.795 109.085 166.995 ;
        RECT 107.930 166.395 108.150 166.795 ;
        RECT 106.035 165.975 106.295 166.305 ;
        RECT 107.050 166.185 107.220 166.335 ;
        RECT 106.465 165.805 106.795 166.165 ;
        RECT 107.050 165.975 108.350 166.185 ;
        RECT 108.625 165.805 109.080 166.570 ;
        RECT 109.255 166.305 109.425 167.505 ;
        RECT 111.125 167.405 111.455 167.435 ;
        RECT 109.655 167.345 111.455 167.405 ;
        RECT 112.045 167.345 112.300 167.965 ;
        RECT 109.595 167.235 112.300 167.345 ;
        RECT 109.595 167.200 109.795 167.235 ;
        RECT 109.595 166.625 109.765 167.200 ;
        RECT 111.125 167.175 112.300 167.235 ;
        RECT 112.935 167.190 113.225 168.355 ;
        RECT 113.455 167.215 113.665 168.355 ;
        RECT 113.835 167.205 114.165 168.185 ;
        RECT 114.335 167.215 114.565 168.355 ;
        RECT 115.250 167.370 115.575 168.355 ;
        RECT 116.145 167.725 116.405 168.185 ;
        RECT 116.575 167.905 117.425 168.355 ;
        RECT 109.995 166.760 110.405 167.065 ;
        RECT 110.575 166.795 110.905 167.005 ;
        RECT 109.595 166.505 109.865 166.625 ;
        RECT 109.595 166.460 110.440 166.505 ;
        RECT 109.685 166.335 110.440 166.460 ;
        RECT 110.695 166.395 110.905 166.795 ;
        RECT 111.150 166.795 111.625 167.005 ;
        RECT 111.815 166.795 112.305 166.995 ;
        RECT 111.150 166.395 111.370 166.795 ;
        RECT 109.255 165.975 109.515 166.305 ;
        RECT 110.270 166.185 110.440 166.335 ;
        RECT 109.685 165.805 110.015 166.165 ;
        RECT 110.270 165.975 111.570 166.185 ;
        RECT 111.845 165.805 112.300 166.570 ;
        RECT 112.935 165.805 113.225 166.530 ;
        RECT 113.455 165.805 113.665 166.625 ;
        RECT 113.835 166.605 114.085 167.205 ;
        RECT 114.255 166.795 114.585 167.045 ;
        RECT 115.245 166.715 115.505 167.170 ;
        RECT 115.760 167.120 115.965 167.705 ;
        RECT 116.145 167.505 117.265 167.725 ;
        RECT 115.760 166.995 116.345 167.120 ;
        RECT 115.755 166.825 116.345 166.995 ;
        RECT 115.760 166.745 116.345 166.825 ;
        RECT 116.515 166.730 116.925 167.335 ;
        RECT 117.095 167.050 117.265 167.505 ;
        RECT 113.835 165.975 114.165 166.605 ;
        RECT 114.335 165.805 114.565 166.625 ;
        RECT 117.095 166.560 117.425 167.050 ;
        RECT 115.250 166.355 116.405 166.545 ;
        RECT 115.250 166.215 115.525 166.355 ;
        RECT 116.195 166.185 116.405 166.355 ;
        RECT 116.575 166.355 117.425 166.560 ;
        RECT 115.695 165.805 116.025 166.185 ;
        RECT 116.575 165.975 116.905 166.355 ;
        RECT 117.095 165.805 117.425 166.185 ;
        RECT 117.595 165.975 117.840 168.185 ;
        RECT 118.025 167.355 118.280 168.355 ;
        RECT 119.005 167.685 119.175 168.185 ;
        RECT 119.345 167.855 119.675 168.355 ;
        RECT 119.005 167.515 119.670 167.685 ;
        RECT 118.920 166.695 119.270 167.345 ;
        RECT 118.025 165.805 118.265 166.605 ;
        RECT 119.440 166.525 119.670 167.515 ;
        RECT 119.005 166.355 119.670 166.525 ;
        RECT 119.005 166.065 119.175 166.355 ;
        RECT 119.345 165.805 119.675 166.185 ;
        RECT 119.845 166.065 120.030 168.185 ;
        RECT 120.270 167.895 120.535 168.355 ;
        RECT 120.705 167.760 120.955 168.185 ;
        RECT 121.165 167.910 122.270 168.080 ;
        RECT 120.650 167.630 120.955 167.760 ;
        RECT 120.200 166.435 120.480 167.385 ;
        RECT 120.650 166.525 120.820 167.630 ;
        RECT 120.990 166.845 121.230 167.440 ;
        RECT 121.400 167.375 121.930 167.740 ;
        RECT 121.400 166.675 121.570 167.375 ;
        RECT 122.100 167.295 122.270 167.910 ;
        RECT 122.440 167.555 122.610 168.355 ;
        RECT 122.780 167.855 123.030 168.185 ;
        RECT 123.255 167.885 124.140 168.055 ;
        RECT 122.100 167.205 122.610 167.295 ;
        RECT 120.650 166.395 120.875 166.525 ;
        RECT 121.045 166.455 121.570 166.675 ;
        RECT 121.740 167.035 122.610 167.205 ;
        RECT 120.285 165.805 120.535 166.265 ;
        RECT 120.705 166.255 120.875 166.395 ;
        RECT 121.740 166.255 121.910 167.035 ;
        RECT 122.440 166.965 122.610 167.035 ;
        RECT 122.120 166.785 122.320 166.815 ;
        RECT 122.780 166.785 122.950 167.855 ;
        RECT 123.120 166.965 123.310 167.685 ;
        RECT 122.120 166.485 122.950 166.785 ;
        RECT 123.480 166.755 123.800 167.715 ;
        RECT 120.705 166.085 121.040 166.255 ;
        RECT 121.235 166.085 121.910 166.255 ;
        RECT 122.230 165.805 122.600 166.305 ;
        RECT 122.780 166.255 122.950 166.485 ;
        RECT 123.335 166.425 123.800 166.755 ;
        RECT 123.970 167.045 124.140 167.885 ;
        RECT 124.320 167.855 124.635 168.355 ;
        RECT 124.865 167.625 125.205 168.185 ;
        RECT 124.310 167.250 125.205 167.625 ;
        RECT 125.375 167.345 125.545 168.355 ;
        RECT 125.015 167.045 125.205 167.250 ;
        RECT 125.715 167.295 126.045 168.140 ;
        RECT 126.280 167.965 126.615 168.185 ;
        RECT 127.620 167.975 127.975 168.355 ;
        RECT 126.280 167.345 126.535 167.965 ;
        RECT 126.785 167.805 127.015 167.845 ;
        RECT 128.145 167.805 128.395 168.185 ;
        RECT 126.785 167.605 128.395 167.805 ;
        RECT 126.785 167.515 126.970 167.605 ;
        RECT 127.560 167.595 128.395 167.605 ;
        RECT 128.645 167.575 128.895 168.355 ;
        RECT 129.065 167.505 129.325 168.185 ;
        RECT 129.585 167.685 129.755 168.185 ;
        RECT 129.925 167.855 130.255 168.355 ;
        RECT 129.585 167.515 130.250 167.685 ;
        RECT 127.125 167.405 127.455 167.435 ;
        RECT 127.125 167.345 128.925 167.405 ;
        RECT 125.715 167.215 126.105 167.295 ;
        RECT 125.890 167.165 126.105 167.215 ;
        RECT 126.280 167.235 128.985 167.345 ;
        RECT 126.280 167.175 127.455 167.235 ;
        RECT 128.785 167.200 128.985 167.235 ;
        RECT 123.970 166.715 124.845 167.045 ;
        RECT 125.015 166.715 125.765 167.045 ;
        RECT 123.970 166.255 124.140 166.715 ;
        RECT 125.015 166.545 125.215 166.715 ;
        RECT 125.935 166.585 126.105 167.165 ;
        RECT 126.275 166.795 126.765 166.995 ;
        RECT 126.955 166.795 127.430 167.005 ;
        RECT 125.880 166.545 126.105 166.585 ;
        RECT 122.780 166.085 123.185 166.255 ;
        RECT 123.355 166.085 124.140 166.255 ;
        RECT 124.415 165.805 124.625 166.335 ;
        RECT 124.885 166.020 125.215 166.545 ;
        RECT 125.725 166.460 126.105 166.545 ;
        RECT 125.385 165.805 125.555 166.415 ;
        RECT 125.725 166.025 126.055 166.460 ;
        RECT 126.280 165.805 126.735 166.570 ;
        RECT 127.210 166.395 127.430 166.795 ;
        RECT 127.675 166.795 128.005 167.005 ;
        RECT 127.675 166.395 127.885 166.795 ;
        RECT 128.175 166.760 128.585 167.065 ;
        RECT 128.815 166.625 128.985 167.200 ;
        RECT 128.715 166.505 128.985 166.625 ;
        RECT 128.140 166.460 128.985 166.505 ;
        RECT 128.140 166.335 128.895 166.460 ;
        RECT 128.140 166.185 128.310 166.335 ;
        RECT 129.155 166.315 129.325 167.505 ;
        RECT 129.500 166.695 129.850 167.345 ;
        RECT 130.020 166.525 130.250 167.515 ;
        RECT 129.095 166.305 129.325 166.315 ;
        RECT 127.010 165.975 128.310 166.185 ;
        RECT 128.565 165.805 128.895 166.165 ;
        RECT 129.065 165.975 129.325 166.305 ;
        RECT 129.585 166.355 130.250 166.525 ;
        RECT 129.585 166.065 129.755 166.355 ;
        RECT 129.925 165.805 130.255 166.185 ;
        RECT 130.425 166.065 130.610 168.185 ;
        RECT 130.850 167.895 131.115 168.355 ;
        RECT 131.285 167.760 131.535 168.185 ;
        RECT 131.745 167.910 132.850 168.080 ;
        RECT 131.230 167.630 131.535 167.760 ;
        RECT 130.780 166.435 131.060 167.385 ;
        RECT 131.230 166.525 131.400 167.630 ;
        RECT 131.570 166.845 131.810 167.440 ;
        RECT 131.980 167.375 132.510 167.740 ;
        RECT 131.980 166.675 132.150 167.375 ;
        RECT 132.680 167.295 132.850 167.910 ;
        RECT 133.020 167.555 133.190 168.355 ;
        RECT 133.360 167.855 133.610 168.185 ;
        RECT 133.835 167.885 134.720 168.055 ;
        RECT 132.680 167.205 133.190 167.295 ;
        RECT 131.230 166.395 131.455 166.525 ;
        RECT 131.625 166.455 132.150 166.675 ;
        RECT 132.320 167.035 133.190 167.205 ;
        RECT 130.865 165.805 131.115 166.265 ;
        RECT 131.285 166.255 131.455 166.395 ;
        RECT 132.320 166.255 132.490 167.035 ;
        RECT 133.020 166.965 133.190 167.035 ;
        RECT 132.700 166.785 132.900 166.815 ;
        RECT 133.360 166.785 133.530 167.855 ;
        RECT 133.700 166.965 133.890 167.685 ;
        RECT 132.700 166.485 133.530 166.785 ;
        RECT 134.060 166.755 134.380 167.715 ;
        RECT 131.285 166.085 131.620 166.255 ;
        RECT 131.815 166.085 132.490 166.255 ;
        RECT 132.810 165.805 133.180 166.305 ;
        RECT 133.360 166.255 133.530 166.485 ;
        RECT 133.915 166.425 134.380 166.755 ;
        RECT 134.550 167.045 134.720 167.885 ;
        RECT 134.900 167.855 135.215 168.355 ;
        RECT 135.445 167.625 135.785 168.185 ;
        RECT 134.890 167.250 135.785 167.625 ;
        RECT 135.955 167.345 136.125 168.355 ;
        RECT 135.595 167.045 135.785 167.250 ;
        RECT 136.295 167.295 136.625 168.140 ;
        RECT 136.295 167.215 136.685 167.295 ;
        RECT 136.855 167.265 138.525 168.355 ;
        RECT 136.470 167.165 136.685 167.215 ;
        RECT 134.550 166.715 135.425 167.045 ;
        RECT 135.595 166.715 136.345 167.045 ;
        RECT 134.550 166.255 134.720 166.715 ;
        RECT 135.595 166.545 135.795 166.715 ;
        RECT 136.515 166.585 136.685 167.165 ;
        RECT 136.460 166.545 136.685 166.585 ;
        RECT 133.360 166.085 133.765 166.255 ;
        RECT 133.935 166.085 134.720 166.255 ;
        RECT 134.995 165.805 135.205 166.335 ;
        RECT 135.465 166.020 135.795 166.545 ;
        RECT 136.305 166.460 136.685 166.545 ;
        RECT 136.855 166.575 137.605 167.095 ;
        RECT 137.775 166.745 138.525 167.265 ;
        RECT 138.695 167.190 138.985 168.355 ;
        RECT 139.155 167.215 139.540 168.185 ;
        RECT 139.710 167.895 140.035 168.355 ;
        RECT 140.555 167.725 140.835 168.185 ;
        RECT 139.710 167.505 140.835 167.725 ;
        RECT 135.965 165.805 136.135 166.415 ;
        RECT 136.305 166.025 136.635 166.460 ;
        RECT 136.855 165.805 138.525 166.575 ;
        RECT 139.155 166.545 139.435 167.215 ;
        RECT 139.710 167.045 140.160 167.505 ;
        RECT 141.025 167.335 141.425 168.185 ;
        RECT 141.825 167.895 142.095 168.355 ;
        RECT 142.265 167.725 142.550 168.185 ;
        RECT 139.605 166.715 140.160 167.045 ;
        RECT 140.330 166.775 141.425 167.335 ;
        RECT 139.710 166.605 140.160 166.715 ;
        RECT 138.695 165.805 138.985 166.530 ;
        RECT 139.155 165.975 139.540 166.545 ;
        RECT 139.710 166.435 140.835 166.605 ;
        RECT 139.710 165.805 140.035 166.265 ;
        RECT 140.555 165.975 140.835 166.435 ;
        RECT 141.025 165.975 141.425 166.775 ;
        RECT 141.595 167.505 142.550 167.725 ;
        RECT 141.595 166.605 141.805 167.505 ;
        RECT 143.040 167.385 143.370 168.185 ;
        RECT 143.540 167.555 143.870 168.355 ;
        RECT 144.170 167.385 144.500 168.185 ;
        RECT 145.145 167.555 145.395 168.355 ;
        RECT 141.975 166.775 142.665 167.335 ;
        RECT 143.040 167.215 145.475 167.385 ;
        RECT 145.665 167.215 145.835 168.355 ;
        RECT 146.005 167.215 146.345 168.185 ;
        RECT 147.065 167.425 147.235 168.185 ;
        RECT 147.415 167.595 147.745 168.355 ;
        RECT 147.065 167.255 147.730 167.425 ;
        RECT 147.915 167.280 148.185 168.185 ;
        RECT 148.415 167.295 148.745 168.140 ;
        RECT 148.915 167.345 149.085 168.355 ;
        RECT 149.255 167.625 149.595 168.185 ;
        RECT 149.825 167.855 150.140 168.355 ;
        RECT 150.320 167.885 151.205 168.055 ;
        RECT 142.835 166.795 143.185 167.045 ;
        RECT 141.595 166.435 142.550 166.605 ;
        RECT 143.370 166.585 143.540 167.215 ;
        RECT 143.710 166.795 144.040 166.995 ;
        RECT 144.210 166.795 144.540 166.995 ;
        RECT 144.710 166.795 145.130 166.995 ;
        RECT 145.305 166.965 145.475 167.215 ;
        RECT 145.305 166.795 146.000 166.965 ;
        RECT 141.825 165.805 142.095 166.265 ;
        RECT 142.265 165.975 142.550 166.435 ;
        RECT 143.040 165.975 143.540 166.585 ;
        RECT 144.170 166.455 145.395 166.625 ;
        RECT 146.170 166.605 146.345 167.215 ;
        RECT 147.560 167.110 147.730 167.255 ;
        RECT 146.995 166.705 147.325 167.075 ;
        RECT 147.560 166.780 147.845 167.110 ;
        RECT 144.170 165.975 144.500 166.455 ;
        RECT 144.670 165.805 144.895 166.265 ;
        RECT 145.065 165.975 145.395 166.455 ;
        RECT 145.585 165.805 145.835 166.605 ;
        RECT 146.005 165.975 146.345 166.605 ;
        RECT 147.560 166.525 147.730 166.780 ;
        RECT 147.065 166.355 147.730 166.525 ;
        RECT 148.015 166.480 148.185 167.280 ;
        RECT 147.065 165.975 147.235 166.355 ;
        RECT 147.415 165.805 147.745 166.185 ;
        RECT 147.925 165.975 148.185 166.480 ;
        RECT 148.355 167.215 148.745 167.295 ;
        RECT 149.255 167.250 150.150 167.625 ;
        RECT 148.355 167.165 148.570 167.215 ;
        RECT 148.355 166.585 148.525 167.165 ;
        RECT 149.255 167.045 149.445 167.250 ;
        RECT 150.320 167.045 150.490 167.885 ;
        RECT 151.430 167.855 151.680 168.185 ;
        RECT 148.695 166.715 149.445 167.045 ;
        RECT 149.615 166.715 150.490 167.045 ;
        RECT 148.355 166.545 148.580 166.585 ;
        RECT 149.245 166.545 149.445 166.715 ;
        RECT 148.355 166.460 148.735 166.545 ;
        RECT 148.405 166.025 148.735 166.460 ;
        RECT 148.905 165.805 149.075 166.415 ;
        RECT 149.245 166.020 149.575 166.545 ;
        RECT 149.835 165.805 150.045 166.335 ;
        RECT 150.320 166.255 150.490 166.715 ;
        RECT 150.660 166.755 150.980 167.715 ;
        RECT 151.150 166.965 151.340 167.685 ;
        RECT 151.510 166.785 151.680 167.855 ;
        RECT 151.850 167.555 152.020 168.355 ;
        RECT 152.190 167.910 153.295 168.080 ;
        RECT 152.190 167.295 152.360 167.910 ;
        RECT 153.505 167.760 153.755 168.185 ;
        RECT 153.925 167.895 154.190 168.355 ;
        RECT 152.530 167.375 153.060 167.740 ;
        RECT 153.505 167.630 153.810 167.760 ;
        RECT 151.850 167.205 152.360 167.295 ;
        RECT 151.850 167.035 152.720 167.205 ;
        RECT 151.850 166.965 152.020 167.035 ;
        RECT 152.140 166.785 152.340 166.815 ;
        RECT 150.660 166.425 151.125 166.755 ;
        RECT 151.510 166.485 152.340 166.785 ;
        RECT 151.510 166.255 151.680 166.485 ;
        RECT 150.320 166.085 151.105 166.255 ;
        RECT 151.275 166.085 151.680 166.255 ;
        RECT 151.860 165.805 152.230 166.305 ;
        RECT 152.550 166.255 152.720 167.035 ;
        RECT 152.890 166.675 153.060 167.375 ;
        RECT 153.230 166.845 153.470 167.440 ;
        RECT 152.890 166.455 153.415 166.675 ;
        RECT 153.640 166.525 153.810 167.630 ;
        RECT 153.585 166.395 153.810 166.525 ;
        RECT 153.980 166.435 154.260 167.385 ;
        RECT 153.585 166.255 153.755 166.395 ;
        RECT 152.550 166.085 153.225 166.255 ;
        RECT 153.420 166.085 153.755 166.255 ;
        RECT 153.925 165.805 154.175 166.265 ;
        RECT 154.430 166.065 154.615 168.185 ;
        RECT 154.785 167.855 155.115 168.355 ;
        RECT 155.285 167.685 155.455 168.185 ;
        RECT 154.790 167.515 155.455 167.685 ;
        RECT 154.790 166.525 155.020 167.515 ;
        RECT 155.190 166.695 155.540 167.345 ;
        RECT 155.715 167.265 156.925 168.355 ;
        RECT 155.715 166.725 156.235 167.265 ;
        RECT 156.405 166.555 156.925 167.095 ;
        RECT 154.790 166.355 155.455 166.525 ;
        RECT 154.785 165.805 155.115 166.185 ;
        RECT 155.285 166.065 155.455 166.355 ;
        RECT 155.715 165.805 156.925 166.555 ;
        RECT 22.690 165.635 157.010 165.805 ;
        RECT 22.775 164.885 23.985 165.635 ;
        RECT 22.775 164.345 23.295 164.885 ;
        RECT 24.155 164.865 25.825 165.635 ;
        RECT 25.995 164.960 26.255 165.465 ;
        RECT 26.435 165.255 26.765 165.635 ;
        RECT 26.945 165.085 27.115 165.465 ;
        RECT 23.465 164.175 23.985 164.715 ;
        RECT 24.155 164.345 24.905 164.865 ;
        RECT 25.075 164.175 25.825 164.695 ;
        RECT 22.775 163.085 23.985 164.175 ;
        RECT 24.155 163.085 25.825 164.175 ;
        RECT 25.995 164.160 26.165 164.960 ;
        RECT 26.450 164.915 27.115 165.085 ;
        RECT 26.450 164.660 26.620 164.915 ;
        RECT 27.375 164.865 30.885 165.635 ;
        RECT 32.010 164.895 32.625 165.465 ;
        RECT 32.795 165.125 33.010 165.635 ;
        RECT 33.240 165.125 33.520 165.455 ;
        RECT 33.700 165.125 33.940 165.635 ;
        RECT 26.335 164.330 26.620 164.660 ;
        RECT 26.855 164.365 27.185 164.735 ;
        RECT 27.375 164.345 29.025 164.865 ;
        RECT 26.450 164.185 26.620 164.330 ;
        RECT 25.995 163.255 26.265 164.160 ;
        RECT 26.450 164.015 27.115 164.185 ;
        RECT 29.195 164.175 30.885 164.695 ;
        RECT 26.435 163.085 26.765 163.845 ;
        RECT 26.945 163.255 27.115 164.015 ;
        RECT 27.375 163.085 30.885 164.175 ;
        RECT 32.010 163.875 32.325 164.895 ;
        RECT 32.495 164.225 32.665 164.725 ;
        RECT 32.915 164.395 33.180 164.955 ;
        RECT 33.350 164.225 33.520 165.125 ;
        RECT 33.690 164.395 34.045 164.955 ;
        RECT 34.275 164.865 36.865 165.635 ;
        RECT 34.275 164.345 35.485 164.865 ;
        RECT 37.495 164.815 37.755 165.635 ;
        RECT 37.925 164.815 38.255 165.235 ;
        RECT 38.435 165.150 39.225 165.415 ;
        RECT 38.005 164.725 38.255 164.815 ;
        RECT 32.495 164.055 33.920 164.225 ;
        RECT 35.655 164.175 36.865 164.695 ;
        RECT 32.010 163.255 32.545 163.875 ;
        RECT 32.715 163.085 33.045 163.885 ;
        RECT 33.530 163.880 33.920 164.055 ;
        RECT 34.275 163.085 36.865 164.175 ;
        RECT 37.495 163.765 37.835 164.645 ;
        RECT 38.005 164.475 38.800 164.725 ;
        RECT 37.495 163.085 37.755 163.595 ;
        RECT 38.005 163.255 38.175 164.475 ;
        RECT 38.970 164.295 39.225 165.150 ;
        RECT 39.395 164.995 39.595 165.415 ;
        RECT 39.785 165.175 40.115 165.635 ;
        RECT 39.395 164.475 39.805 164.995 ;
        RECT 40.285 164.985 40.545 165.465 ;
        RECT 39.975 164.295 40.205 164.725 ;
        RECT 38.415 164.125 40.205 164.295 ;
        RECT 38.415 163.760 38.665 164.125 ;
        RECT 38.835 163.765 39.165 163.955 ;
        RECT 39.385 163.830 40.100 164.125 ;
        RECT 40.375 163.955 40.545 164.985 ;
        RECT 40.715 164.865 44.225 165.635 ;
        RECT 44.395 164.885 45.605 165.635 ;
        RECT 45.780 165.130 46.115 165.635 ;
        RECT 46.285 165.065 46.525 165.440 ;
        RECT 46.805 165.305 46.975 165.450 ;
        RECT 46.805 165.110 47.180 165.305 ;
        RECT 47.540 165.140 47.935 165.635 ;
        RECT 40.715 164.345 42.365 164.865 ;
        RECT 42.535 164.175 44.225 164.695 ;
        RECT 44.395 164.345 44.915 164.885 ;
        RECT 45.085 164.175 45.605 164.715 ;
        RECT 38.835 163.590 39.030 163.765 ;
        RECT 38.415 163.085 39.030 163.590 ;
        RECT 39.200 163.255 39.675 163.595 ;
        RECT 39.845 163.085 40.060 163.630 ;
        RECT 40.270 163.255 40.545 163.955 ;
        RECT 40.715 163.085 44.225 164.175 ;
        RECT 44.395 163.085 45.605 164.175 ;
        RECT 45.835 164.105 46.135 164.955 ;
        RECT 46.305 164.915 46.525 165.065 ;
        RECT 46.305 164.585 46.840 164.915 ;
        RECT 47.010 164.775 47.180 165.110 ;
        RECT 48.105 164.945 48.345 165.465 ;
        RECT 46.305 163.935 46.540 164.585 ;
        RECT 47.010 164.415 47.995 164.775 ;
        RECT 45.865 163.705 46.540 163.935 ;
        RECT 46.710 164.395 47.995 164.415 ;
        RECT 46.710 164.245 47.570 164.395 ;
        RECT 45.865 163.275 46.035 163.705 ;
        RECT 46.205 163.085 46.535 163.535 ;
        RECT 46.710 163.300 46.995 164.245 ;
        RECT 48.170 164.140 48.345 164.945 ;
        RECT 48.535 164.910 48.825 165.635 ;
        RECT 49.020 164.985 49.330 165.455 ;
        RECT 49.500 165.155 50.235 165.635 ;
        RECT 50.405 165.065 50.575 165.415 ;
        RECT 50.745 165.235 51.125 165.635 ;
        RECT 49.020 164.815 49.755 164.985 ;
        RECT 50.405 164.895 51.145 165.065 ;
        RECT 51.315 164.960 51.585 165.305 ;
        RECT 49.505 164.725 49.755 164.815 ;
        RECT 50.975 164.725 51.145 164.895 ;
        RECT 49.000 164.395 49.335 164.645 ;
        RECT 49.505 164.395 50.245 164.725 ;
        RECT 50.975 164.395 51.205 164.725 ;
        RECT 47.170 163.765 47.865 164.075 ;
        RECT 47.175 163.085 47.860 163.555 ;
        RECT 48.040 163.355 48.345 164.140 ;
        RECT 48.535 163.085 48.825 164.250 ;
        RECT 49.000 163.085 49.255 164.225 ;
        RECT 49.505 163.835 49.675 164.395 ;
        RECT 50.975 164.225 51.145 164.395 ;
        RECT 51.415 164.225 51.585 164.960 ;
        RECT 51.765 164.905 52.065 165.635 ;
        RECT 52.245 164.725 52.475 165.345 ;
        RECT 52.675 165.075 52.900 165.455 ;
        RECT 53.070 165.245 53.400 165.635 ;
        RECT 52.675 164.895 53.005 165.075 ;
        RECT 51.770 164.395 52.065 164.725 ;
        RECT 52.245 164.395 52.660 164.725 ;
        RECT 49.900 164.055 51.145 164.225 ;
        RECT 49.900 163.805 50.320 164.055 ;
        RECT 49.450 163.305 50.645 163.635 ;
        RECT 50.825 163.085 51.105 163.885 ;
        RECT 51.315 163.255 51.585 164.225 ;
        RECT 52.830 164.225 53.005 164.895 ;
        RECT 53.175 164.395 53.415 165.045 ;
        RECT 54.535 165.005 54.865 165.465 ;
        RECT 55.045 165.175 55.215 165.635 ;
        RECT 55.395 165.005 55.725 165.465 ;
        RECT 55.955 165.175 56.125 165.635 ;
        RECT 56.365 165.295 57.555 165.465 ;
        RECT 56.365 165.005 56.695 165.295 ;
        RECT 57.245 165.125 57.555 165.295 ;
        RECT 57.735 165.175 58.295 165.465 ;
        RECT 58.465 165.175 58.715 165.635 ;
        RECT 54.535 164.835 56.695 165.005 ;
        RECT 54.550 164.275 54.880 164.665 ;
        RECT 55.050 164.445 55.850 164.645 ;
        RECT 56.030 164.275 56.525 164.645 ;
        RECT 51.765 163.865 52.660 164.195 ;
        RECT 52.830 164.035 53.415 164.225 ;
        RECT 54.550 164.105 56.585 164.275 ;
        RECT 51.765 163.695 52.970 163.865 ;
        RECT 51.765 163.265 52.095 163.695 ;
        RECT 52.275 163.085 52.470 163.525 ;
        RECT 52.640 163.265 52.970 163.695 ;
        RECT 53.140 163.265 53.415 164.035 ;
        RECT 56.865 163.935 57.075 165.125 ;
        RECT 57.245 164.320 57.560 164.955 ;
        RECT 54.535 163.085 54.865 163.935 ;
        RECT 55.035 163.425 55.255 163.935 ;
        RECT 55.425 163.755 57.075 163.935 ;
        RECT 55.425 163.595 55.725 163.755 ;
        RECT 55.955 163.425 56.145 163.585 ;
        RECT 55.035 163.255 56.145 163.425 ;
        RECT 56.340 163.085 56.670 163.545 ;
        RECT 56.840 163.255 57.075 163.755 ;
        RECT 57.245 163.085 57.555 164.150 ;
        RECT 57.735 163.805 57.985 165.175 ;
        RECT 59.335 165.005 59.665 165.365 ;
        RECT 58.275 164.815 59.665 165.005 ;
        RECT 60.035 164.865 62.625 165.635 ;
        RECT 63.345 165.085 63.515 165.375 ;
        RECT 63.685 165.255 64.015 165.635 ;
        RECT 63.345 164.915 64.010 165.085 ;
        RECT 58.275 164.725 58.445 164.815 ;
        RECT 58.155 164.395 58.445 164.725 ;
        RECT 58.615 164.395 58.955 164.645 ;
        RECT 59.175 164.395 59.850 164.645 ;
        RECT 58.275 164.145 58.445 164.395 ;
        RECT 58.275 163.975 59.215 164.145 ;
        RECT 59.585 164.035 59.850 164.395 ;
        RECT 60.035 164.345 61.245 164.865 ;
        RECT 61.415 164.175 62.625 164.695 ;
        RECT 57.735 163.255 58.195 163.805 ;
        RECT 58.385 163.085 58.715 163.805 ;
        RECT 58.915 163.425 59.215 163.975 ;
        RECT 59.385 163.085 59.665 163.755 ;
        RECT 60.035 163.085 62.625 164.175 ;
        RECT 63.260 164.095 63.610 164.745 ;
        RECT 63.780 163.925 64.010 164.915 ;
        RECT 63.345 163.755 64.010 163.925 ;
        RECT 63.345 163.255 63.515 163.755 ;
        RECT 63.685 163.085 64.015 163.585 ;
        RECT 64.185 163.255 64.370 165.375 ;
        RECT 64.625 165.175 64.875 165.635 ;
        RECT 65.045 165.185 65.380 165.355 ;
        RECT 65.575 165.185 66.250 165.355 ;
        RECT 65.045 165.045 65.215 165.185 ;
        RECT 64.540 164.055 64.820 165.005 ;
        RECT 64.990 164.915 65.215 165.045 ;
        RECT 64.990 163.810 65.160 164.915 ;
        RECT 65.385 164.765 65.910 164.985 ;
        RECT 65.330 164.000 65.570 164.595 ;
        RECT 65.740 164.065 65.910 164.765 ;
        RECT 66.080 164.405 66.250 165.185 ;
        RECT 66.570 165.135 66.940 165.635 ;
        RECT 67.120 165.185 67.525 165.355 ;
        RECT 67.695 165.185 68.480 165.355 ;
        RECT 67.120 164.955 67.290 165.185 ;
        RECT 66.460 164.655 67.290 164.955 ;
        RECT 67.675 164.685 68.140 165.015 ;
        RECT 66.460 164.625 66.660 164.655 ;
        RECT 66.780 164.405 66.950 164.475 ;
        RECT 66.080 164.235 66.950 164.405 ;
        RECT 66.440 164.145 66.950 164.235 ;
        RECT 64.990 163.680 65.295 163.810 ;
        RECT 65.740 163.700 66.270 164.065 ;
        RECT 64.610 163.085 64.875 163.545 ;
        RECT 65.045 163.255 65.295 163.680 ;
        RECT 66.440 163.530 66.610 164.145 ;
        RECT 65.505 163.360 66.610 163.530 ;
        RECT 66.780 163.085 66.950 163.885 ;
        RECT 67.120 163.585 67.290 164.655 ;
        RECT 67.460 163.755 67.650 164.475 ;
        RECT 67.820 163.725 68.140 164.685 ;
        RECT 68.310 164.725 68.480 165.185 ;
        RECT 68.755 165.105 68.965 165.635 ;
        RECT 69.225 164.895 69.555 165.420 ;
        RECT 69.725 165.025 69.895 165.635 ;
        RECT 70.065 164.980 70.395 165.415 ;
        RECT 70.065 164.895 70.445 164.980 ;
        RECT 69.355 164.725 69.555 164.895 ;
        RECT 70.220 164.855 70.445 164.895 ;
        RECT 68.310 164.395 69.185 164.725 ;
        RECT 69.355 164.395 70.105 164.725 ;
        RECT 67.120 163.255 67.370 163.585 ;
        RECT 68.310 163.555 68.480 164.395 ;
        RECT 69.355 164.190 69.545 164.395 ;
        RECT 70.275 164.275 70.445 164.855 ;
        RECT 70.230 164.225 70.445 164.275 ;
        RECT 68.650 163.815 69.545 164.190 ;
        RECT 70.055 164.145 70.445 164.225 ;
        RECT 70.615 164.895 71.000 165.465 ;
        RECT 71.170 165.175 71.495 165.635 ;
        RECT 72.015 165.005 72.295 165.465 ;
        RECT 70.615 164.225 70.895 164.895 ;
        RECT 71.170 164.835 72.295 165.005 ;
        RECT 71.170 164.725 71.620 164.835 ;
        RECT 71.065 164.395 71.620 164.725 ;
        RECT 72.485 164.665 72.885 165.465 ;
        RECT 73.285 165.175 73.555 165.635 ;
        RECT 73.725 165.005 74.010 165.465 ;
        RECT 67.595 163.385 68.480 163.555 ;
        RECT 68.660 163.085 68.975 163.585 ;
        RECT 69.205 163.255 69.545 163.815 ;
        RECT 69.715 163.085 69.885 164.095 ;
        RECT 70.055 163.300 70.385 164.145 ;
        RECT 70.615 163.255 71.000 164.225 ;
        RECT 71.170 163.935 71.620 164.395 ;
        RECT 71.790 164.105 72.885 164.665 ;
        RECT 71.170 163.715 72.295 163.935 ;
        RECT 71.170 163.085 71.495 163.545 ;
        RECT 72.015 163.255 72.295 163.715 ;
        RECT 72.485 163.255 72.885 164.105 ;
        RECT 73.055 164.835 74.010 165.005 ;
        RECT 74.295 164.910 74.585 165.635 ;
        RECT 74.755 164.865 76.425 165.635 ;
        RECT 77.145 165.085 77.315 165.375 ;
        RECT 77.485 165.255 77.815 165.635 ;
        RECT 77.145 164.915 77.810 165.085 ;
        RECT 73.055 163.935 73.265 164.835 ;
        RECT 73.435 164.105 74.125 164.665 ;
        RECT 74.755 164.345 75.505 164.865 ;
        RECT 73.055 163.715 74.010 163.935 ;
        RECT 73.285 163.085 73.555 163.545 ;
        RECT 73.725 163.255 74.010 163.715 ;
        RECT 74.295 163.085 74.585 164.250 ;
        RECT 75.675 164.175 76.425 164.695 ;
        RECT 74.755 163.085 76.425 164.175 ;
        RECT 77.060 164.095 77.410 164.745 ;
        RECT 77.580 163.925 77.810 164.915 ;
        RECT 77.145 163.755 77.810 163.925 ;
        RECT 77.145 163.255 77.315 163.755 ;
        RECT 77.485 163.085 77.815 163.585 ;
        RECT 77.985 163.255 78.170 165.375 ;
        RECT 78.425 165.175 78.675 165.635 ;
        RECT 78.845 165.185 79.180 165.355 ;
        RECT 79.375 165.185 80.050 165.355 ;
        RECT 78.845 165.045 79.015 165.185 ;
        RECT 78.340 164.055 78.620 165.005 ;
        RECT 78.790 164.915 79.015 165.045 ;
        RECT 78.790 163.810 78.960 164.915 ;
        RECT 79.185 164.765 79.710 164.985 ;
        RECT 79.130 164.000 79.370 164.595 ;
        RECT 79.540 164.065 79.710 164.765 ;
        RECT 79.880 164.405 80.050 165.185 ;
        RECT 80.370 165.135 80.740 165.635 ;
        RECT 80.920 165.185 81.325 165.355 ;
        RECT 81.495 165.185 82.280 165.355 ;
        RECT 80.920 164.955 81.090 165.185 ;
        RECT 80.260 164.655 81.090 164.955 ;
        RECT 81.475 164.685 81.940 165.015 ;
        RECT 80.260 164.625 80.460 164.655 ;
        RECT 80.580 164.405 80.750 164.475 ;
        RECT 79.880 164.235 80.750 164.405 ;
        RECT 80.240 164.145 80.750 164.235 ;
        RECT 78.790 163.680 79.095 163.810 ;
        RECT 79.540 163.700 80.070 164.065 ;
        RECT 78.410 163.085 78.675 163.545 ;
        RECT 78.845 163.255 79.095 163.680 ;
        RECT 80.240 163.530 80.410 164.145 ;
        RECT 79.305 163.360 80.410 163.530 ;
        RECT 80.580 163.085 80.750 163.885 ;
        RECT 80.920 163.585 81.090 164.655 ;
        RECT 81.260 163.755 81.450 164.475 ;
        RECT 81.620 163.725 81.940 164.685 ;
        RECT 82.110 164.725 82.280 165.185 ;
        RECT 82.555 165.105 82.765 165.635 ;
        RECT 83.025 164.895 83.355 165.420 ;
        RECT 83.525 165.025 83.695 165.635 ;
        RECT 83.865 164.980 84.195 165.415 ;
        RECT 85.385 164.980 85.715 165.415 ;
        RECT 85.885 165.025 86.055 165.635 ;
        RECT 83.865 164.895 84.245 164.980 ;
        RECT 83.155 164.725 83.355 164.895 ;
        RECT 84.020 164.855 84.245 164.895 ;
        RECT 82.110 164.395 82.985 164.725 ;
        RECT 83.155 164.395 83.905 164.725 ;
        RECT 80.920 163.255 81.170 163.585 ;
        RECT 82.110 163.555 82.280 164.395 ;
        RECT 83.155 164.190 83.345 164.395 ;
        RECT 84.075 164.275 84.245 164.855 ;
        RECT 84.030 164.225 84.245 164.275 ;
        RECT 82.450 163.815 83.345 164.190 ;
        RECT 83.855 164.145 84.245 164.225 ;
        RECT 85.335 164.895 85.715 164.980 ;
        RECT 86.225 164.895 86.555 165.420 ;
        RECT 86.815 165.105 87.025 165.635 ;
        RECT 87.300 165.185 88.085 165.355 ;
        RECT 88.255 165.185 88.660 165.355 ;
        RECT 85.335 164.855 85.560 164.895 ;
        RECT 85.335 164.275 85.505 164.855 ;
        RECT 86.225 164.725 86.425 164.895 ;
        RECT 87.300 164.725 87.470 165.185 ;
        RECT 85.675 164.395 86.425 164.725 ;
        RECT 86.595 164.395 87.470 164.725 ;
        RECT 85.335 164.225 85.550 164.275 ;
        RECT 85.335 164.145 85.725 164.225 ;
        RECT 81.395 163.385 82.280 163.555 ;
        RECT 82.460 163.085 82.775 163.585 ;
        RECT 83.005 163.255 83.345 163.815 ;
        RECT 83.515 163.085 83.685 164.095 ;
        RECT 83.855 163.300 84.185 164.145 ;
        RECT 85.395 163.300 85.725 164.145 ;
        RECT 86.235 164.190 86.425 164.395 ;
        RECT 85.895 163.085 86.065 164.095 ;
        RECT 86.235 163.815 87.130 164.190 ;
        RECT 86.235 163.255 86.575 163.815 ;
        RECT 86.805 163.085 87.120 163.585 ;
        RECT 87.300 163.555 87.470 164.395 ;
        RECT 87.640 164.685 88.105 165.015 ;
        RECT 88.490 164.955 88.660 165.185 ;
        RECT 88.840 165.135 89.210 165.635 ;
        RECT 89.530 165.185 90.205 165.355 ;
        RECT 90.400 165.185 90.735 165.355 ;
        RECT 87.640 163.725 87.960 164.685 ;
        RECT 88.490 164.655 89.320 164.955 ;
        RECT 88.130 163.755 88.320 164.475 ;
        RECT 88.490 163.585 88.660 164.655 ;
        RECT 89.120 164.625 89.320 164.655 ;
        RECT 88.830 164.405 89.000 164.475 ;
        RECT 89.530 164.405 89.700 165.185 ;
        RECT 90.565 165.045 90.735 165.185 ;
        RECT 90.905 165.175 91.155 165.635 ;
        RECT 88.830 164.235 89.700 164.405 ;
        RECT 89.870 164.765 90.395 164.985 ;
        RECT 90.565 164.915 90.790 165.045 ;
        RECT 88.830 164.145 89.340 164.235 ;
        RECT 87.300 163.385 88.185 163.555 ;
        RECT 88.410 163.255 88.660 163.585 ;
        RECT 88.830 163.085 89.000 163.885 ;
        RECT 89.170 163.530 89.340 164.145 ;
        RECT 89.870 164.065 90.040 164.765 ;
        RECT 89.510 163.700 90.040 164.065 ;
        RECT 90.210 164.000 90.450 164.595 ;
        RECT 90.620 163.810 90.790 164.915 ;
        RECT 90.960 164.055 91.240 165.005 ;
        RECT 90.485 163.680 90.790 163.810 ;
        RECT 89.170 163.360 90.275 163.530 ;
        RECT 90.485 163.255 90.735 163.680 ;
        RECT 90.905 163.085 91.170 163.545 ;
        RECT 91.410 163.255 91.595 165.375 ;
        RECT 91.765 165.255 92.095 165.635 ;
        RECT 92.265 165.085 92.435 165.375 ;
        RECT 91.770 164.915 92.435 165.085 ;
        RECT 92.745 164.980 93.075 165.415 ;
        RECT 93.245 165.025 93.415 165.635 ;
        RECT 91.770 163.925 92.000 164.915 ;
        RECT 92.695 164.895 93.075 164.980 ;
        RECT 93.585 164.895 93.915 165.420 ;
        RECT 94.175 165.105 94.385 165.635 ;
        RECT 94.660 165.185 95.445 165.355 ;
        RECT 95.615 165.185 96.020 165.355 ;
        RECT 92.695 164.855 92.920 164.895 ;
        RECT 92.170 164.095 92.520 164.745 ;
        RECT 92.695 164.275 92.865 164.855 ;
        RECT 93.585 164.725 93.785 164.895 ;
        RECT 94.660 164.725 94.830 165.185 ;
        RECT 93.035 164.395 93.785 164.725 ;
        RECT 93.955 164.395 94.830 164.725 ;
        RECT 92.695 164.225 92.910 164.275 ;
        RECT 92.695 164.145 93.085 164.225 ;
        RECT 91.770 163.755 92.435 163.925 ;
        RECT 91.765 163.085 92.095 163.585 ;
        RECT 92.265 163.255 92.435 163.755 ;
        RECT 92.755 163.300 93.085 164.145 ;
        RECT 93.595 164.190 93.785 164.395 ;
        RECT 93.255 163.085 93.425 164.095 ;
        RECT 93.595 163.815 94.490 164.190 ;
        RECT 93.595 163.255 93.935 163.815 ;
        RECT 94.165 163.085 94.480 163.585 ;
        RECT 94.660 163.555 94.830 164.395 ;
        RECT 95.000 164.685 95.465 165.015 ;
        RECT 95.850 164.955 96.020 165.185 ;
        RECT 96.200 165.135 96.570 165.635 ;
        RECT 96.890 165.185 97.565 165.355 ;
        RECT 97.760 165.185 98.095 165.355 ;
        RECT 95.000 163.725 95.320 164.685 ;
        RECT 95.850 164.655 96.680 164.955 ;
        RECT 95.490 163.755 95.680 164.475 ;
        RECT 95.850 163.585 96.020 164.655 ;
        RECT 96.480 164.625 96.680 164.655 ;
        RECT 96.190 164.405 96.360 164.475 ;
        RECT 96.890 164.405 97.060 165.185 ;
        RECT 97.925 165.045 98.095 165.185 ;
        RECT 98.265 165.175 98.515 165.635 ;
        RECT 96.190 164.235 97.060 164.405 ;
        RECT 97.230 164.765 97.755 164.985 ;
        RECT 97.925 164.915 98.150 165.045 ;
        RECT 96.190 164.145 96.700 164.235 ;
        RECT 94.660 163.385 95.545 163.555 ;
        RECT 95.770 163.255 96.020 163.585 ;
        RECT 96.190 163.085 96.360 163.885 ;
        RECT 96.530 163.530 96.700 164.145 ;
        RECT 97.230 164.065 97.400 164.765 ;
        RECT 96.870 163.700 97.400 164.065 ;
        RECT 97.570 164.000 97.810 164.595 ;
        RECT 97.980 163.810 98.150 164.915 ;
        RECT 98.320 164.055 98.600 165.005 ;
        RECT 97.845 163.680 98.150 163.810 ;
        RECT 96.530 163.360 97.635 163.530 ;
        RECT 97.845 163.255 98.095 163.680 ;
        RECT 98.265 163.085 98.530 163.545 ;
        RECT 98.770 163.255 98.955 165.375 ;
        RECT 99.125 165.255 99.455 165.635 ;
        RECT 99.625 165.085 99.795 165.375 ;
        RECT 99.130 164.915 99.795 165.085 ;
        RECT 99.130 163.925 99.360 164.915 ;
        RECT 100.055 164.910 100.345 165.635 ;
        RECT 100.515 165.005 100.855 165.465 ;
        RECT 101.025 165.175 101.195 165.635 ;
        RECT 101.825 165.200 102.185 165.465 ;
        RECT 101.830 165.195 102.185 165.200 ;
        RECT 101.835 165.185 102.185 165.195 ;
        RECT 101.840 165.180 102.185 165.185 ;
        RECT 101.845 165.170 102.185 165.180 ;
        RECT 102.425 165.175 102.595 165.635 ;
        RECT 101.850 165.165 102.185 165.170 ;
        RECT 101.860 165.155 102.185 165.165 ;
        RECT 101.870 165.145 102.185 165.155 ;
        RECT 101.365 165.005 101.695 165.085 ;
        RECT 100.515 164.815 101.695 165.005 ;
        RECT 101.885 165.005 102.185 165.145 ;
        RECT 101.885 164.815 102.595 165.005 ;
        RECT 99.530 164.095 99.880 164.745 ;
        RECT 100.515 164.445 100.845 164.645 ;
        RECT 101.155 164.625 101.485 164.645 ;
        RECT 101.035 164.445 101.485 164.625 ;
        RECT 99.130 163.755 99.795 163.925 ;
        RECT 99.125 163.085 99.455 163.585 ;
        RECT 99.625 163.255 99.795 163.755 ;
        RECT 100.055 163.085 100.345 164.250 ;
        RECT 100.515 164.105 100.745 164.445 ;
        RECT 100.525 163.085 100.855 163.805 ;
        RECT 101.035 163.330 101.250 164.445 ;
        RECT 101.655 164.415 102.125 164.645 ;
        RECT 102.310 164.245 102.595 164.815 ;
        RECT 102.765 164.690 103.105 165.465 ;
        RECT 103.275 164.835 103.970 165.465 ;
        RECT 104.175 164.835 104.485 165.635 ;
        RECT 101.445 164.030 102.595 164.245 ;
        RECT 101.445 163.255 101.775 164.030 ;
        RECT 101.945 163.085 102.655 163.860 ;
        RECT 102.825 163.255 103.105 164.690 ;
        RECT 103.295 164.395 103.630 164.645 ;
        RECT 103.800 164.235 103.970 164.835 ;
        RECT 104.675 164.825 104.915 165.635 ;
        RECT 105.085 164.825 105.415 165.465 ;
        RECT 105.585 164.825 105.855 165.635 ;
        RECT 106.035 164.865 107.705 165.635 ;
        RECT 108.335 165.135 108.595 165.465 ;
        RECT 108.765 165.275 109.095 165.635 ;
        RECT 109.350 165.255 110.650 165.465 ;
        RECT 104.140 164.395 104.475 164.665 ;
        RECT 104.655 164.395 105.005 164.645 ;
        RECT 103.275 163.085 103.535 164.225 ;
        RECT 103.705 163.255 104.035 164.235 ;
        RECT 105.175 164.225 105.345 164.825 ;
        RECT 105.515 164.395 105.865 164.645 ;
        RECT 106.035 164.345 106.785 164.865 ;
        RECT 104.205 163.085 104.485 164.225 ;
        RECT 104.665 164.055 105.345 164.225 ;
        RECT 104.665 163.270 104.995 164.055 ;
        RECT 105.525 163.085 105.855 164.225 ;
        RECT 106.955 164.175 107.705 164.695 ;
        RECT 106.035 163.085 107.705 164.175 ;
        RECT 108.335 163.935 108.505 165.135 ;
        RECT 109.350 165.105 109.520 165.255 ;
        RECT 108.765 164.980 109.520 165.105 ;
        RECT 108.675 164.935 109.520 164.980 ;
        RECT 108.675 164.815 108.945 164.935 ;
        RECT 108.675 164.240 108.845 164.815 ;
        RECT 109.075 164.375 109.485 164.680 ;
        RECT 109.775 164.645 109.985 165.045 ;
        RECT 109.655 164.435 109.985 164.645 ;
        RECT 110.230 164.645 110.450 165.045 ;
        RECT 110.925 164.870 111.380 165.635 ;
        RECT 111.555 164.885 112.765 165.635 ;
        RECT 112.935 164.895 113.320 165.465 ;
        RECT 113.490 165.175 113.815 165.635 ;
        RECT 114.335 165.005 114.615 165.465 ;
        RECT 110.230 164.435 110.705 164.645 ;
        RECT 110.895 164.445 111.385 164.645 ;
        RECT 111.555 164.345 112.075 164.885 ;
        RECT 108.675 164.205 108.875 164.240 ;
        RECT 110.205 164.205 111.380 164.265 ;
        RECT 108.675 164.095 111.380 164.205 ;
        RECT 112.245 164.175 112.765 164.715 ;
        RECT 108.735 164.035 110.535 164.095 ;
        RECT 110.205 164.005 110.535 164.035 ;
        RECT 108.335 163.255 108.595 163.935 ;
        RECT 108.765 163.085 109.015 163.865 ;
        RECT 109.265 163.835 110.100 163.845 ;
        RECT 110.690 163.835 110.875 163.925 ;
        RECT 109.265 163.635 110.875 163.835 ;
        RECT 109.265 163.255 109.515 163.635 ;
        RECT 110.645 163.595 110.875 163.635 ;
        RECT 111.125 163.475 111.380 164.095 ;
        RECT 109.685 163.085 110.040 163.465 ;
        RECT 111.045 163.255 111.380 163.475 ;
        RECT 111.555 163.085 112.765 164.175 ;
        RECT 112.935 164.225 113.215 164.895 ;
        RECT 113.490 164.835 114.615 165.005 ;
        RECT 113.490 164.725 113.940 164.835 ;
        RECT 113.385 164.395 113.940 164.725 ;
        RECT 114.805 164.665 115.205 165.465 ;
        RECT 115.605 165.175 115.875 165.635 ;
        RECT 116.045 165.005 116.330 165.465 ;
        RECT 116.665 165.165 116.955 165.635 ;
        RECT 112.935 163.255 113.320 164.225 ;
        RECT 113.490 163.935 113.940 164.395 ;
        RECT 114.110 164.105 115.205 164.665 ;
        RECT 113.490 163.715 114.615 163.935 ;
        RECT 113.490 163.085 113.815 163.545 ;
        RECT 114.335 163.255 114.615 163.715 ;
        RECT 114.805 163.255 115.205 164.105 ;
        RECT 115.375 164.835 116.330 165.005 ;
        RECT 117.125 164.995 117.455 165.465 ;
        RECT 117.625 165.165 117.795 165.635 ;
        RECT 117.965 164.995 118.295 165.465 ;
        RECT 117.125 164.985 118.295 164.995 ;
        RECT 115.375 163.935 115.585 164.835 ;
        RECT 116.695 164.815 118.295 164.985 ;
        RECT 118.465 164.815 118.740 165.635 ;
        RECT 119.375 165.135 119.635 165.465 ;
        RECT 119.805 165.275 120.135 165.635 ;
        RECT 120.390 165.255 121.690 165.465 ;
        RECT 119.375 165.125 119.605 165.135 ;
        RECT 115.755 164.105 116.445 164.665 ;
        RECT 116.695 164.275 116.910 164.815 ;
        RECT 117.080 164.445 117.850 164.645 ;
        RECT 118.020 164.445 118.740 164.645 ;
        RECT 116.695 164.055 117.455 164.275 ;
        RECT 115.375 163.715 116.330 163.935 ;
        RECT 115.605 163.085 115.875 163.545 ;
        RECT 116.045 163.255 116.330 163.715 ;
        RECT 116.655 163.425 116.955 163.885 ;
        RECT 117.125 163.595 117.455 164.055 ;
        RECT 117.625 164.055 118.740 164.265 ;
        RECT 117.625 163.425 117.795 164.055 ;
        RECT 116.655 163.255 117.795 163.425 ;
        RECT 117.965 163.085 118.295 163.885 ;
        RECT 118.465 163.255 118.740 164.055 ;
        RECT 119.375 163.935 119.545 165.125 ;
        RECT 120.390 165.105 120.560 165.255 ;
        RECT 119.805 164.980 120.560 165.105 ;
        RECT 119.715 164.935 120.560 164.980 ;
        RECT 119.715 164.815 119.985 164.935 ;
        RECT 119.715 164.240 119.885 164.815 ;
        RECT 120.115 164.375 120.525 164.680 ;
        RECT 120.815 164.645 121.025 165.045 ;
        RECT 120.695 164.435 121.025 164.645 ;
        RECT 121.270 164.645 121.490 165.045 ;
        RECT 121.965 164.870 122.420 165.635 ;
        RECT 122.595 164.865 125.185 165.635 ;
        RECT 125.815 164.910 126.105 165.635 ;
        RECT 126.275 164.895 126.660 165.465 ;
        RECT 126.830 165.175 127.155 165.635 ;
        RECT 127.675 165.005 127.955 165.465 ;
        RECT 121.270 164.435 121.745 164.645 ;
        RECT 121.935 164.445 122.425 164.645 ;
        RECT 122.595 164.345 123.805 164.865 ;
        RECT 119.715 164.205 119.915 164.240 ;
        RECT 121.245 164.205 122.420 164.265 ;
        RECT 119.715 164.095 122.420 164.205 ;
        RECT 123.975 164.175 125.185 164.695 ;
        RECT 119.775 164.035 121.575 164.095 ;
        RECT 121.245 164.005 121.575 164.035 ;
        RECT 119.375 163.255 119.635 163.935 ;
        RECT 119.805 163.085 120.055 163.865 ;
        RECT 120.305 163.835 121.140 163.845 ;
        RECT 121.730 163.835 121.915 163.925 ;
        RECT 120.305 163.635 121.915 163.835 ;
        RECT 120.305 163.255 120.555 163.635 ;
        RECT 121.685 163.595 121.915 163.635 ;
        RECT 122.165 163.475 122.420 164.095 ;
        RECT 120.725 163.085 121.080 163.465 ;
        RECT 122.085 163.255 122.420 163.475 ;
        RECT 122.595 163.085 125.185 164.175 ;
        RECT 125.815 163.085 126.105 164.250 ;
        RECT 126.275 164.225 126.555 164.895 ;
        RECT 126.830 164.835 127.955 165.005 ;
        RECT 126.830 164.725 127.280 164.835 ;
        RECT 126.725 164.395 127.280 164.725 ;
        RECT 128.145 164.665 128.545 165.465 ;
        RECT 128.945 165.175 129.215 165.635 ;
        RECT 129.385 165.005 129.670 165.465 ;
        RECT 126.275 163.255 126.660 164.225 ;
        RECT 126.830 163.935 127.280 164.395 ;
        RECT 127.450 164.105 128.545 164.665 ;
        RECT 126.830 163.715 127.955 163.935 ;
        RECT 126.830 163.085 127.155 163.545 ;
        RECT 127.675 163.255 127.955 163.715 ;
        RECT 128.145 163.255 128.545 164.105 ;
        RECT 128.715 164.835 129.670 165.005 ;
        RECT 129.955 164.885 131.165 165.635 ;
        RECT 131.335 164.895 131.720 165.465 ;
        RECT 131.890 165.175 132.215 165.635 ;
        RECT 132.735 165.005 133.015 165.465 ;
        RECT 128.715 163.935 128.925 164.835 ;
        RECT 129.095 164.105 129.785 164.665 ;
        RECT 129.955 164.345 130.475 164.885 ;
        RECT 130.645 164.175 131.165 164.715 ;
        RECT 128.715 163.715 129.670 163.935 ;
        RECT 128.945 163.085 129.215 163.545 ;
        RECT 129.385 163.255 129.670 163.715 ;
        RECT 129.955 163.085 131.165 164.175 ;
        RECT 131.335 164.225 131.615 164.895 ;
        RECT 131.890 164.835 133.015 165.005 ;
        RECT 131.890 164.725 132.340 164.835 ;
        RECT 131.785 164.395 132.340 164.725 ;
        RECT 133.205 164.665 133.605 165.465 ;
        RECT 134.005 165.175 134.275 165.635 ;
        RECT 134.445 165.005 134.730 165.465 ;
        RECT 131.335 163.255 131.720 164.225 ;
        RECT 131.890 163.935 132.340 164.395 ;
        RECT 132.510 164.105 133.605 164.665 ;
        RECT 131.890 163.715 133.015 163.935 ;
        RECT 131.890 163.085 132.215 163.545 ;
        RECT 132.735 163.255 133.015 163.715 ;
        RECT 133.205 163.255 133.605 164.105 ;
        RECT 133.775 164.835 134.730 165.005 ;
        RECT 135.015 164.895 135.400 165.465 ;
        RECT 135.570 165.175 135.895 165.635 ;
        RECT 136.415 165.005 136.695 165.465 ;
        RECT 133.775 163.935 133.985 164.835 ;
        RECT 134.155 164.105 134.845 164.665 ;
        RECT 135.015 164.225 135.295 164.895 ;
        RECT 135.570 164.835 136.695 165.005 ;
        RECT 135.570 164.725 136.020 164.835 ;
        RECT 135.465 164.395 136.020 164.725 ;
        RECT 136.885 164.665 137.285 165.465 ;
        RECT 137.685 165.175 137.955 165.635 ;
        RECT 138.125 165.005 138.410 165.465 ;
        RECT 133.775 163.715 134.730 163.935 ;
        RECT 134.005 163.085 134.275 163.545 ;
        RECT 134.445 163.255 134.730 163.715 ;
        RECT 135.015 163.255 135.400 164.225 ;
        RECT 135.570 163.935 136.020 164.395 ;
        RECT 136.190 164.105 137.285 164.665 ;
        RECT 135.570 163.715 136.695 163.935 ;
        RECT 135.570 163.085 135.895 163.545 ;
        RECT 136.415 163.255 136.695 163.715 ;
        RECT 136.885 163.255 137.285 164.105 ;
        RECT 137.455 164.835 138.410 165.005 ;
        RECT 138.695 164.865 142.205 165.635 ;
        RECT 137.455 163.935 137.665 164.835 ;
        RECT 137.835 164.105 138.525 164.665 ;
        RECT 138.695 164.345 140.345 164.865 ;
        RECT 143.355 164.815 143.565 165.635 ;
        RECT 143.735 164.835 144.065 165.465 ;
        RECT 140.515 164.175 142.205 164.695 ;
        RECT 143.735 164.235 143.985 164.835 ;
        RECT 144.235 164.815 144.465 165.635 ;
        RECT 144.675 164.895 145.060 165.465 ;
        RECT 145.230 165.175 145.555 165.635 ;
        RECT 146.075 165.005 146.355 165.465 ;
        RECT 144.155 164.395 144.485 164.645 ;
        RECT 137.455 163.715 138.410 163.935 ;
        RECT 137.685 163.085 137.955 163.545 ;
        RECT 138.125 163.255 138.410 163.715 ;
        RECT 138.695 163.085 142.205 164.175 ;
        RECT 143.355 163.085 143.565 164.225 ;
        RECT 143.735 163.255 144.065 164.235 ;
        RECT 144.675 164.225 144.955 164.895 ;
        RECT 145.230 164.835 146.355 165.005 ;
        RECT 145.230 164.725 145.680 164.835 ;
        RECT 145.125 164.395 145.680 164.725 ;
        RECT 146.545 164.665 146.945 165.465 ;
        RECT 147.345 165.175 147.615 165.635 ;
        RECT 147.785 165.005 148.070 165.465 ;
        RECT 148.635 165.005 149.015 165.455 ;
        RECT 144.235 163.085 144.465 164.225 ;
        RECT 144.675 163.255 145.060 164.225 ;
        RECT 145.230 163.935 145.680 164.395 ;
        RECT 145.850 164.105 146.945 164.665 ;
        RECT 145.230 163.715 146.355 163.935 ;
        RECT 145.230 163.085 145.555 163.545 ;
        RECT 146.075 163.255 146.355 163.715 ;
        RECT 146.545 163.255 146.945 164.105 ;
        RECT 147.115 164.835 148.070 165.005 ;
        RECT 147.115 163.935 147.325 164.835 ;
        RECT 147.495 164.105 148.185 164.665 ;
        RECT 148.375 164.055 148.605 164.745 ;
        RECT 148.785 164.555 149.015 165.005 ;
        RECT 149.195 164.855 149.425 165.635 ;
        RECT 149.605 164.925 150.035 165.455 ;
        RECT 149.605 164.675 149.850 164.925 ;
        RECT 150.215 164.725 150.425 165.345 ;
        RECT 150.595 164.905 150.925 165.635 ;
        RECT 151.575 164.910 151.865 165.635 ;
        RECT 152.035 165.255 152.925 165.425 ;
        RECT 147.115 163.715 148.070 163.935 ;
        RECT 148.785 163.875 149.125 164.555 ;
        RECT 147.345 163.085 147.615 163.545 ;
        RECT 147.785 163.255 148.070 163.715 ;
        RECT 148.365 163.675 149.125 163.875 ;
        RECT 149.315 164.375 149.850 164.675 ;
        RECT 150.030 164.375 150.425 164.725 ;
        RECT 150.620 164.375 150.910 164.725 ;
        RECT 152.035 164.700 152.585 165.085 ;
        RECT 152.755 164.530 152.925 165.255 ;
        RECT 152.035 164.460 152.925 164.530 ;
        RECT 153.095 164.955 153.315 165.415 ;
        RECT 153.485 165.095 153.735 165.635 ;
        RECT 153.905 164.985 154.165 165.465 ;
        RECT 153.095 164.930 153.345 164.955 ;
        RECT 153.095 164.505 153.425 164.930 ;
        RECT 152.035 164.435 152.930 164.460 ;
        RECT 152.035 164.420 152.940 164.435 ;
        RECT 152.035 164.405 152.945 164.420 ;
        RECT 152.035 164.400 152.955 164.405 ;
        RECT 152.035 164.390 152.960 164.400 ;
        RECT 152.035 164.380 152.965 164.390 ;
        RECT 152.035 164.375 152.975 164.380 ;
        RECT 148.365 163.285 148.625 163.675 ;
        RECT 148.795 163.085 149.125 163.495 ;
        RECT 149.315 163.265 149.645 164.375 ;
        RECT 152.035 164.365 152.985 164.375 ;
        RECT 152.035 164.360 152.995 164.365 ;
        RECT 149.815 163.995 150.855 164.195 ;
        RECT 149.815 163.265 150.005 163.995 ;
        RECT 150.175 163.085 150.505 163.815 ;
        RECT 150.685 163.265 150.855 163.995 ;
        RECT 151.575 163.085 151.865 164.250 ;
        RECT 152.035 163.910 152.295 164.360 ;
        RECT 152.660 164.355 152.995 164.360 ;
        RECT 152.660 164.350 153.010 164.355 ;
        RECT 152.660 164.340 153.025 164.350 ;
        RECT 152.660 164.335 153.050 164.340 ;
        RECT 153.595 164.335 153.825 164.730 ;
        RECT 152.660 164.330 153.825 164.335 ;
        RECT 152.690 164.295 153.825 164.330 ;
        RECT 152.725 164.270 153.825 164.295 ;
        RECT 152.755 164.240 153.825 164.270 ;
        RECT 152.775 164.210 153.825 164.240 ;
        RECT 152.795 164.180 153.825 164.210 ;
        RECT 152.865 164.170 153.825 164.180 ;
        RECT 152.890 164.160 153.825 164.170 ;
        RECT 152.910 164.145 153.825 164.160 ;
        RECT 152.930 164.130 153.825 164.145 ;
        RECT 152.935 164.120 153.720 164.130 ;
        RECT 152.950 164.085 153.720 164.120 ;
        RECT 152.465 163.765 152.795 164.010 ;
        RECT 152.965 163.835 153.720 164.085 ;
        RECT 153.995 163.955 154.165 164.985 ;
        RECT 152.465 163.740 152.650 163.765 ;
        RECT 152.035 163.640 152.650 163.740 ;
        RECT 152.035 163.085 152.640 163.640 ;
        RECT 152.815 163.255 153.295 163.595 ;
        RECT 153.465 163.085 153.720 163.630 ;
        RECT 153.890 163.255 154.165 163.955 ;
        RECT 154.335 164.960 154.595 165.465 ;
        RECT 154.775 165.255 155.105 165.635 ;
        RECT 155.285 165.085 155.455 165.465 ;
        RECT 154.335 164.160 154.505 164.960 ;
        RECT 154.790 164.915 155.455 165.085 ;
        RECT 154.790 164.660 154.960 164.915 ;
        RECT 155.715 164.885 156.925 165.635 ;
        RECT 154.675 164.330 154.960 164.660 ;
        RECT 155.195 164.365 155.525 164.735 ;
        RECT 154.790 164.185 154.960 164.330 ;
        RECT 154.335 163.255 154.605 164.160 ;
        RECT 154.790 164.015 155.455 164.185 ;
        RECT 154.775 163.085 155.105 163.845 ;
        RECT 155.285 163.255 155.455 164.015 ;
        RECT 155.715 164.175 156.235 164.715 ;
        RECT 156.405 164.345 156.925 164.885 ;
        RECT 155.715 163.085 156.925 164.175 ;
        RECT 22.690 162.915 157.010 163.085 ;
        RECT 22.775 161.825 23.985 162.915 ;
        RECT 22.775 161.115 23.295 161.655 ;
        RECT 23.465 161.285 23.985 161.825 ;
        RECT 25.085 162.305 25.415 162.735 ;
        RECT 25.595 162.475 25.790 162.915 ;
        RECT 25.960 162.305 26.290 162.735 ;
        RECT 25.085 162.135 26.290 162.305 ;
        RECT 25.085 161.805 25.980 162.135 ;
        RECT 26.460 161.965 26.735 162.735 ;
        RECT 26.150 161.775 26.735 161.965 ;
        RECT 26.920 161.775 27.240 162.915 ;
        RECT 25.090 161.275 25.385 161.605 ;
        RECT 25.565 161.275 25.980 161.605 ;
        RECT 22.775 160.365 23.985 161.115 ;
        RECT 25.085 160.365 25.385 161.095 ;
        RECT 25.565 160.655 25.795 161.275 ;
        RECT 26.150 161.105 26.325 161.775 ;
        RECT 27.420 161.605 27.615 162.655 ;
        RECT 27.795 162.065 28.125 162.745 ;
        RECT 28.325 162.115 28.580 162.915 ;
        RECT 27.795 161.785 28.145 162.065 ;
        RECT 25.995 160.925 26.325 161.105 ;
        RECT 26.495 160.955 26.735 161.605 ;
        RECT 26.980 161.555 27.240 161.605 ;
        RECT 26.975 161.385 27.240 161.555 ;
        RECT 26.980 161.275 27.240 161.385 ;
        RECT 27.420 161.275 27.805 161.605 ;
        RECT 27.975 161.405 28.145 161.785 ;
        RECT 28.335 161.575 28.580 161.935 ;
        RECT 28.755 161.775 29.140 162.745 ;
        RECT 29.310 162.455 29.635 162.915 ;
        RECT 30.155 162.285 30.435 162.745 ;
        RECT 29.310 162.065 30.435 162.285 ;
        RECT 27.975 161.235 28.495 161.405 ;
        RECT 28.325 161.215 28.495 161.235 ;
        RECT 25.995 160.545 26.220 160.925 ;
        RECT 26.920 160.895 28.135 161.065 ;
        RECT 26.390 160.365 26.720 160.755 ;
        RECT 26.920 160.545 27.210 160.895 ;
        RECT 27.405 160.365 27.735 160.725 ;
        RECT 27.905 160.590 28.135 160.895 ;
        RECT 28.325 161.045 28.525 161.215 ;
        RECT 28.755 161.105 29.035 161.775 ;
        RECT 29.310 161.605 29.760 162.065 ;
        RECT 30.625 161.895 31.025 162.745 ;
        RECT 31.425 162.455 31.695 162.915 ;
        RECT 31.865 162.285 32.150 162.745 ;
        RECT 29.205 161.275 29.760 161.605 ;
        RECT 29.930 161.335 31.025 161.895 ;
        RECT 29.310 161.165 29.760 161.275 ;
        RECT 28.325 160.670 28.495 161.045 ;
        RECT 28.755 160.535 29.140 161.105 ;
        RECT 29.310 160.995 30.435 161.165 ;
        RECT 29.310 160.365 29.635 160.825 ;
        RECT 30.155 160.535 30.435 160.995 ;
        RECT 30.625 160.535 31.025 161.335 ;
        RECT 31.195 162.065 32.150 162.285 ;
        RECT 31.195 161.165 31.405 162.065 ;
        RECT 32.525 161.985 32.695 162.745 ;
        RECT 32.875 162.155 33.205 162.915 ;
        RECT 31.575 161.335 32.265 161.895 ;
        RECT 32.525 161.815 33.190 161.985 ;
        RECT 33.375 161.840 33.645 162.745 ;
        RECT 33.020 161.670 33.190 161.815 ;
        RECT 32.455 161.265 32.785 161.635 ;
        RECT 33.020 161.340 33.305 161.670 ;
        RECT 31.195 160.995 32.150 161.165 ;
        RECT 33.020 161.085 33.190 161.340 ;
        RECT 31.425 160.365 31.695 160.825 ;
        RECT 31.865 160.535 32.150 160.995 ;
        RECT 32.525 160.915 33.190 161.085 ;
        RECT 33.475 161.040 33.645 161.840 ;
        RECT 33.815 161.825 35.485 162.915 ;
        RECT 32.525 160.535 32.695 160.915 ;
        RECT 32.875 160.365 33.205 160.745 ;
        RECT 33.385 160.535 33.645 161.040 ;
        RECT 33.815 161.135 34.565 161.655 ;
        RECT 34.735 161.305 35.485 161.825 ;
        RECT 35.655 161.750 35.945 162.915 ;
        RECT 33.815 160.365 35.485 161.135 ;
        RECT 35.655 160.365 35.945 161.090 ;
        RECT 36.585 160.545 36.845 162.735 ;
        RECT 37.015 162.185 37.355 162.915 ;
        RECT 37.535 162.005 37.805 162.735 ;
        RECT 37.035 161.785 37.805 162.005 ;
        RECT 37.985 162.025 38.215 162.735 ;
        RECT 38.385 162.205 38.715 162.915 ;
        RECT 38.885 162.025 39.145 162.735 ;
        RECT 39.335 162.405 40.525 162.695 ;
        RECT 37.985 161.785 39.145 162.025 ;
        RECT 39.355 162.065 40.525 162.235 ;
        RECT 40.695 162.115 40.975 162.915 ;
        RECT 37.035 161.115 37.325 161.785 ;
        RECT 39.355 161.775 39.680 162.065 ;
        RECT 40.355 161.945 40.525 162.065 ;
        RECT 39.850 161.605 40.045 161.895 ;
        RECT 40.355 161.775 41.015 161.945 ;
        RECT 41.185 161.775 41.460 162.745 ;
        RECT 41.635 161.825 44.225 162.915 ;
        RECT 40.845 161.605 41.015 161.775 ;
        RECT 37.505 161.295 37.970 161.605 ;
        RECT 38.150 161.295 38.675 161.605 ;
        RECT 37.035 160.915 38.265 161.115 ;
        RECT 37.105 160.365 37.775 160.735 ;
        RECT 37.955 160.545 38.265 160.915 ;
        RECT 38.445 160.655 38.675 161.295 ;
        RECT 38.855 161.275 39.155 161.605 ;
        RECT 39.335 161.275 39.680 161.605 ;
        RECT 39.850 161.275 40.675 161.605 ;
        RECT 40.845 161.275 41.120 161.605 ;
        RECT 40.845 161.105 41.015 161.275 ;
        RECT 38.855 160.365 39.145 161.095 ;
        RECT 39.350 160.935 41.015 161.105 ;
        RECT 41.290 161.040 41.460 161.775 ;
        RECT 39.350 160.585 39.605 160.935 ;
        RECT 39.775 160.365 40.105 160.765 ;
        RECT 40.275 160.585 40.445 160.935 ;
        RECT 40.615 160.365 40.995 160.765 ;
        RECT 41.185 160.695 41.460 161.040 ;
        RECT 41.635 161.135 42.845 161.655 ;
        RECT 43.015 161.305 44.225 161.825 ;
        RECT 44.405 161.945 44.735 162.745 ;
        RECT 44.905 162.115 45.135 162.915 ;
        RECT 45.305 161.945 45.635 162.745 ;
        RECT 44.405 161.775 45.635 161.945 ;
        RECT 45.805 161.775 46.060 162.915 ;
        RECT 46.235 162.480 51.580 162.915 ;
        RECT 44.395 161.275 44.705 161.605 ;
        RECT 41.635 160.365 44.225 161.135 ;
        RECT 44.405 160.875 44.735 161.105 ;
        RECT 44.910 161.045 45.285 161.605 ;
        RECT 45.455 160.875 45.635 161.775 ;
        RECT 45.820 161.025 46.040 161.605 ;
        RECT 47.820 160.910 48.160 161.740 ;
        RECT 49.640 161.230 49.990 162.480 ;
        RECT 51.755 161.825 54.345 162.915 ;
        RECT 51.755 161.135 52.965 161.655 ;
        RECT 53.135 161.305 54.345 161.825 ;
        RECT 44.405 160.535 45.635 160.875 ;
        RECT 45.805 160.365 46.060 160.855 ;
        RECT 46.235 160.365 51.580 160.910 ;
        RECT 51.755 160.365 54.345 161.135 ;
        RECT 54.525 160.545 54.785 162.735 ;
        RECT 54.955 162.185 55.295 162.915 ;
        RECT 55.475 162.005 55.745 162.735 ;
        RECT 54.975 161.785 55.745 162.005 ;
        RECT 55.925 162.025 56.155 162.735 ;
        RECT 56.325 162.205 56.655 162.915 ;
        RECT 56.825 162.025 57.085 162.735 ;
        RECT 55.925 161.785 57.085 162.025 ;
        RECT 54.975 161.115 55.265 161.785 ;
        RECT 57.275 161.775 57.545 162.745 ;
        RECT 57.755 162.115 58.035 162.915 ;
        RECT 58.215 162.365 59.410 162.695 ;
        RECT 58.540 161.945 58.960 162.195 ;
        RECT 57.715 161.775 58.960 161.945 ;
        RECT 55.445 161.295 55.910 161.605 ;
        RECT 56.090 161.295 56.615 161.605 ;
        RECT 54.975 160.915 56.205 161.115 ;
        RECT 55.045 160.365 55.715 160.735 ;
        RECT 55.895 160.545 56.205 160.915 ;
        RECT 56.385 160.655 56.615 161.295 ;
        RECT 56.795 161.275 57.095 161.605 ;
        RECT 56.795 160.365 57.085 161.095 ;
        RECT 57.275 161.040 57.445 161.775 ;
        RECT 57.715 161.605 57.885 161.775 ;
        RECT 59.185 161.605 59.355 162.165 ;
        RECT 59.605 161.775 59.860 162.915 ;
        RECT 60.035 161.825 61.245 162.915 ;
        RECT 57.655 161.275 57.885 161.605 ;
        RECT 58.615 161.275 59.355 161.605 ;
        RECT 59.525 161.355 59.860 161.605 ;
        RECT 57.715 161.105 57.885 161.275 ;
        RECT 59.105 161.185 59.355 161.275 ;
        RECT 57.275 160.695 57.545 161.040 ;
        RECT 57.715 160.935 58.455 161.105 ;
        RECT 59.105 161.015 59.840 161.185 ;
        RECT 57.735 160.365 58.115 160.765 ;
        RECT 58.285 160.585 58.455 160.935 ;
        RECT 58.625 160.365 59.360 160.845 ;
        RECT 59.530 160.545 59.840 161.015 ;
        RECT 60.035 161.115 60.555 161.655 ;
        RECT 60.725 161.285 61.245 161.825 ;
        RECT 61.415 161.750 61.705 162.915 ;
        RECT 61.875 161.825 63.545 162.915 ;
        RECT 61.875 161.135 62.625 161.655 ;
        RECT 62.795 161.305 63.545 161.825 ;
        RECT 63.715 162.065 63.975 162.745 ;
        RECT 64.145 162.135 64.395 162.915 ;
        RECT 64.645 162.365 64.895 162.745 ;
        RECT 65.065 162.535 65.420 162.915 ;
        RECT 66.425 162.525 66.760 162.745 ;
        RECT 66.025 162.365 66.255 162.405 ;
        RECT 64.645 162.165 66.255 162.365 ;
        RECT 64.645 162.155 65.480 162.165 ;
        RECT 66.070 162.075 66.255 162.165 ;
        RECT 60.035 160.365 61.245 161.115 ;
        RECT 61.415 160.365 61.705 161.090 ;
        RECT 61.875 160.365 63.545 161.135 ;
        RECT 63.715 160.865 63.885 162.065 ;
        RECT 65.585 161.965 65.915 161.995 ;
        RECT 64.115 161.905 65.915 161.965 ;
        RECT 66.505 161.905 66.760 162.525 ;
        RECT 64.055 161.795 66.760 161.905 ;
        RECT 66.935 161.825 69.525 162.915 ;
        RECT 70.215 161.855 70.545 162.700 ;
        RECT 70.715 161.905 70.885 162.915 ;
        RECT 71.055 162.185 71.395 162.745 ;
        RECT 71.625 162.415 71.940 162.915 ;
        RECT 72.120 162.445 73.005 162.615 ;
        RECT 64.055 161.760 64.255 161.795 ;
        RECT 64.055 161.185 64.225 161.760 ;
        RECT 65.585 161.735 66.760 161.795 ;
        RECT 64.455 161.320 64.865 161.625 ;
        RECT 65.035 161.355 65.365 161.565 ;
        RECT 64.055 161.065 64.325 161.185 ;
        RECT 64.055 161.020 64.900 161.065 ;
        RECT 64.145 160.895 64.900 161.020 ;
        RECT 65.155 160.955 65.365 161.355 ;
        RECT 65.610 161.355 66.085 161.565 ;
        RECT 66.275 161.355 66.765 161.555 ;
        RECT 65.610 160.955 65.830 161.355 ;
        RECT 66.935 161.135 68.145 161.655 ;
        RECT 68.315 161.305 69.525 161.825 ;
        RECT 70.155 161.775 70.545 161.855 ;
        RECT 71.055 161.810 71.950 162.185 ;
        RECT 70.155 161.725 70.370 161.775 ;
        RECT 70.155 161.145 70.325 161.725 ;
        RECT 71.055 161.605 71.245 161.810 ;
        RECT 72.120 161.605 72.290 162.445 ;
        RECT 73.230 162.415 73.480 162.745 ;
        RECT 70.495 161.275 71.245 161.605 ;
        RECT 71.415 161.275 72.290 161.605 ;
        RECT 63.715 160.535 63.975 160.865 ;
        RECT 64.730 160.745 64.900 160.895 ;
        RECT 64.145 160.365 64.475 160.725 ;
        RECT 64.730 160.535 66.030 160.745 ;
        RECT 66.305 160.365 66.760 161.130 ;
        RECT 66.935 160.365 69.525 161.135 ;
        RECT 70.155 161.105 70.380 161.145 ;
        RECT 71.045 161.105 71.245 161.275 ;
        RECT 70.155 161.020 70.535 161.105 ;
        RECT 70.205 160.585 70.535 161.020 ;
        RECT 70.705 160.365 70.875 160.975 ;
        RECT 71.045 160.580 71.375 161.105 ;
        RECT 71.635 160.365 71.845 160.895 ;
        RECT 72.120 160.815 72.290 161.275 ;
        RECT 72.460 161.315 72.780 162.275 ;
        RECT 72.950 161.525 73.140 162.245 ;
        RECT 73.310 161.345 73.480 162.415 ;
        RECT 73.650 162.115 73.820 162.915 ;
        RECT 73.990 162.470 75.095 162.640 ;
        RECT 73.990 161.855 74.160 162.470 ;
        RECT 75.305 162.320 75.555 162.745 ;
        RECT 75.725 162.455 75.990 162.915 ;
        RECT 74.330 161.935 74.860 162.300 ;
        RECT 75.305 162.190 75.610 162.320 ;
        RECT 73.650 161.765 74.160 161.855 ;
        RECT 73.650 161.595 74.520 161.765 ;
        RECT 73.650 161.525 73.820 161.595 ;
        RECT 73.940 161.345 74.140 161.375 ;
        RECT 72.460 160.985 72.925 161.315 ;
        RECT 73.310 161.045 74.140 161.345 ;
        RECT 73.310 160.815 73.480 161.045 ;
        RECT 72.120 160.645 72.905 160.815 ;
        RECT 73.075 160.645 73.480 160.815 ;
        RECT 73.660 160.365 74.030 160.865 ;
        RECT 74.350 160.815 74.520 161.595 ;
        RECT 74.690 161.235 74.860 161.935 ;
        RECT 75.030 161.405 75.270 162.000 ;
        RECT 74.690 161.015 75.215 161.235 ;
        RECT 75.440 161.085 75.610 162.190 ;
        RECT 75.385 160.955 75.610 161.085 ;
        RECT 75.780 160.995 76.060 161.945 ;
        RECT 75.385 160.815 75.555 160.955 ;
        RECT 74.350 160.645 75.025 160.815 ;
        RECT 75.220 160.645 75.555 160.815 ;
        RECT 75.725 160.365 75.975 160.825 ;
        RECT 76.230 160.625 76.415 162.745 ;
        RECT 76.585 162.415 76.915 162.915 ;
        RECT 77.085 162.245 77.255 162.745 ;
        RECT 76.590 162.075 77.255 162.245 ;
        RECT 76.590 161.085 76.820 162.075 ;
        RECT 76.990 161.255 77.340 161.905 ;
        RECT 77.515 161.825 79.185 162.915 ;
        RECT 79.820 161.915 80.075 162.915 ;
        RECT 77.515 161.135 78.265 161.655 ;
        RECT 78.435 161.305 79.185 161.825 ;
        RECT 76.590 160.915 77.255 161.085 ;
        RECT 76.585 160.365 76.915 160.745 ;
        RECT 77.085 160.625 77.255 160.915 ;
        RECT 77.515 160.365 79.185 161.135 ;
        RECT 79.835 160.365 80.075 161.165 ;
        RECT 80.260 160.535 80.505 162.745 ;
        RECT 80.675 162.465 81.525 162.915 ;
        RECT 81.695 162.285 81.955 162.745 ;
        RECT 80.835 162.065 81.955 162.285 ;
        RECT 80.835 161.610 81.005 162.065 ;
        RECT 80.675 161.120 81.005 161.610 ;
        RECT 81.175 161.290 81.585 161.895 ;
        RECT 82.135 161.680 82.340 162.265 ;
        RECT 82.525 161.930 82.850 162.915 ;
        RECT 83.035 161.825 86.545 162.915 ;
        RECT 81.755 161.555 82.340 161.680 ;
        RECT 81.755 161.385 82.345 161.555 ;
        RECT 81.755 161.305 82.340 161.385 ;
        RECT 82.595 161.275 82.855 161.730 ;
        RECT 83.035 161.135 84.685 161.655 ;
        RECT 84.855 161.305 86.545 161.825 ;
        RECT 87.175 161.750 87.465 162.915 ;
        RECT 80.675 160.915 81.525 161.120 ;
        RECT 80.675 160.365 81.005 160.745 ;
        RECT 81.195 160.535 81.525 160.915 ;
        RECT 81.695 160.915 82.850 161.105 ;
        RECT 81.695 160.745 81.905 160.915 ;
        RECT 82.575 160.775 82.850 160.915 ;
        RECT 82.075 160.365 82.405 160.745 ;
        RECT 83.035 160.365 86.545 161.135 ;
        RECT 87.175 160.365 87.465 161.090 ;
        RECT 88.105 160.545 88.365 162.735 ;
        RECT 88.535 162.185 88.875 162.915 ;
        RECT 89.055 162.005 89.325 162.735 ;
        RECT 88.555 161.785 89.325 162.005 ;
        RECT 89.505 162.025 89.735 162.735 ;
        RECT 89.905 162.205 90.235 162.915 ;
        RECT 90.405 162.025 90.665 162.735 ;
        RECT 89.505 161.785 90.665 162.025 ;
        RECT 90.855 161.840 91.125 162.745 ;
        RECT 91.295 162.155 91.625 162.915 ;
        RECT 91.805 161.985 91.975 162.745 ;
        RECT 88.555 161.115 88.845 161.785 ;
        RECT 89.025 161.295 89.490 161.605 ;
        RECT 89.670 161.295 90.195 161.605 ;
        RECT 88.555 160.915 89.785 161.115 ;
        RECT 88.625 160.365 89.295 160.735 ;
        RECT 89.475 160.545 89.785 160.915 ;
        RECT 89.965 160.655 90.195 161.295 ;
        RECT 90.375 161.275 90.675 161.605 ;
        RECT 90.375 160.365 90.665 161.095 ;
        RECT 90.855 161.040 91.025 161.840 ;
        RECT 91.310 161.815 91.975 161.985 ;
        RECT 92.235 161.825 93.905 162.915 ;
        RECT 94.190 162.285 94.475 162.745 ;
        RECT 94.645 162.455 94.915 162.915 ;
        RECT 94.190 162.065 95.145 162.285 ;
        RECT 91.310 161.670 91.480 161.815 ;
        RECT 91.195 161.340 91.480 161.670 ;
        RECT 91.310 161.085 91.480 161.340 ;
        RECT 91.715 161.265 92.045 161.635 ;
        RECT 92.235 161.135 92.985 161.655 ;
        RECT 93.155 161.305 93.905 161.825 ;
        RECT 94.075 161.335 94.765 161.895 ;
        RECT 94.935 161.165 95.145 162.065 ;
        RECT 90.855 160.535 91.115 161.040 ;
        RECT 91.310 160.915 91.975 161.085 ;
        RECT 91.295 160.365 91.625 160.745 ;
        RECT 91.805 160.535 91.975 160.915 ;
        RECT 92.235 160.365 93.905 161.135 ;
        RECT 94.190 160.995 95.145 161.165 ;
        RECT 95.315 161.895 95.715 162.745 ;
        RECT 95.905 162.285 96.185 162.745 ;
        RECT 96.705 162.455 97.030 162.915 ;
        RECT 95.905 162.065 97.030 162.285 ;
        RECT 95.315 161.335 96.410 161.895 ;
        RECT 96.580 161.605 97.030 162.065 ;
        RECT 97.200 161.775 97.585 162.745 ;
        RECT 97.755 162.405 98.055 162.915 ;
        RECT 98.225 162.235 98.555 162.745 ;
        RECT 98.725 162.405 99.355 162.915 ;
        RECT 99.935 162.405 100.315 162.575 ;
        RECT 100.485 162.405 100.785 162.915 ;
        RECT 100.145 162.235 100.315 162.405 ;
        RECT 94.190 160.535 94.475 160.995 ;
        RECT 94.645 160.365 94.915 160.825 ;
        RECT 95.315 160.535 95.715 161.335 ;
        RECT 96.580 161.275 97.135 161.605 ;
        RECT 96.580 161.165 97.030 161.275 ;
        RECT 95.905 160.995 97.030 161.165 ;
        RECT 97.305 161.105 97.585 161.775 ;
        RECT 95.905 160.535 96.185 160.995 ;
        RECT 96.705 160.365 97.030 160.825 ;
        RECT 97.200 160.535 97.585 161.105 ;
        RECT 97.755 162.065 99.975 162.235 ;
        RECT 97.755 161.105 97.925 162.065 ;
        RECT 98.095 161.725 99.635 161.895 ;
        RECT 98.095 161.275 98.340 161.725 ;
        RECT 98.600 161.355 99.295 161.555 ;
        RECT 99.465 161.525 99.635 161.725 ;
        RECT 99.805 161.865 99.975 162.065 ;
        RECT 100.145 162.035 100.805 162.235 ;
        RECT 99.805 161.695 100.465 161.865 ;
        RECT 99.465 161.355 100.065 161.525 ;
        RECT 100.295 161.275 100.465 161.695 ;
        RECT 97.755 160.560 98.220 161.105 ;
        RECT 98.725 160.365 98.895 161.185 ;
        RECT 99.065 161.105 99.975 161.185 ;
        RECT 100.635 161.105 100.805 162.035 ;
        RECT 100.975 161.825 102.645 162.915 ;
        RECT 103.335 161.855 103.665 162.700 ;
        RECT 103.835 161.905 104.005 162.915 ;
        RECT 104.175 162.185 104.515 162.745 ;
        RECT 104.745 162.415 105.060 162.915 ;
        RECT 105.240 162.445 106.125 162.615 ;
        RECT 99.065 161.015 100.315 161.105 ;
        RECT 99.065 160.535 99.395 161.015 ;
        RECT 99.805 160.935 100.315 161.015 ;
        RECT 99.565 160.365 99.915 160.755 ;
        RECT 100.085 160.535 100.315 160.935 ;
        RECT 100.485 160.625 100.805 161.105 ;
        RECT 100.975 161.135 101.725 161.655 ;
        RECT 101.895 161.305 102.645 161.825 ;
        RECT 103.275 161.775 103.665 161.855 ;
        RECT 104.175 161.810 105.070 162.185 ;
        RECT 103.275 161.725 103.490 161.775 ;
        RECT 103.275 161.145 103.445 161.725 ;
        RECT 104.175 161.605 104.365 161.810 ;
        RECT 105.240 161.605 105.410 162.445 ;
        RECT 106.350 162.415 106.600 162.745 ;
        RECT 103.615 161.275 104.365 161.605 ;
        RECT 104.535 161.275 105.410 161.605 ;
        RECT 100.975 160.365 102.645 161.135 ;
        RECT 103.275 161.105 103.500 161.145 ;
        RECT 104.165 161.105 104.365 161.275 ;
        RECT 103.275 161.020 103.655 161.105 ;
        RECT 103.325 160.585 103.655 161.020 ;
        RECT 103.825 160.365 103.995 160.975 ;
        RECT 104.165 160.580 104.495 161.105 ;
        RECT 104.755 160.365 104.965 160.895 ;
        RECT 105.240 160.815 105.410 161.275 ;
        RECT 105.580 161.315 105.900 162.275 ;
        RECT 106.070 161.525 106.260 162.245 ;
        RECT 106.430 161.345 106.600 162.415 ;
        RECT 106.770 162.115 106.940 162.915 ;
        RECT 107.110 162.470 108.215 162.640 ;
        RECT 107.110 161.855 107.280 162.470 ;
        RECT 108.425 162.320 108.675 162.745 ;
        RECT 108.845 162.455 109.110 162.915 ;
        RECT 107.450 161.935 107.980 162.300 ;
        RECT 108.425 162.190 108.730 162.320 ;
        RECT 106.770 161.765 107.280 161.855 ;
        RECT 106.770 161.595 107.640 161.765 ;
        RECT 106.770 161.525 106.940 161.595 ;
        RECT 107.060 161.345 107.260 161.375 ;
        RECT 105.580 160.985 106.045 161.315 ;
        RECT 106.430 161.045 107.260 161.345 ;
        RECT 106.430 160.815 106.600 161.045 ;
        RECT 105.240 160.645 106.025 160.815 ;
        RECT 106.195 160.645 106.600 160.815 ;
        RECT 106.780 160.365 107.150 160.865 ;
        RECT 107.470 160.815 107.640 161.595 ;
        RECT 107.810 161.235 107.980 161.935 ;
        RECT 108.150 161.405 108.390 162.000 ;
        RECT 107.810 161.015 108.335 161.235 ;
        RECT 108.560 161.085 108.730 162.190 ;
        RECT 108.505 160.955 108.730 161.085 ;
        RECT 108.900 160.995 109.180 161.945 ;
        RECT 108.505 160.815 108.675 160.955 ;
        RECT 107.470 160.645 108.145 160.815 ;
        RECT 108.340 160.645 108.675 160.815 ;
        RECT 108.845 160.365 109.095 160.825 ;
        RECT 109.350 160.625 109.535 162.745 ;
        RECT 109.705 162.415 110.035 162.915 ;
        RECT 110.205 162.245 110.375 162.745 ;
        RECT 109.710 162.075 110.375 162.245 ;
        RECT 109.710 161.085 109.940 162.075 ;
        RECT 110.110 161.255 110.460 161.905 ;
        RECT 110.635 161.825 112.305 162.915 ;
        RECT 110.635 161.135 111.385 161.655 ;
        RECT 111.555 161.305 112.305 161.825 ;
        RECT 112.935 161.750 113.225 162.915 ;
        RECT 113.395 161.825 115.065 162.915 ;
        RECT 115.705 162.195 116.035 162.915 ;
        RECT 113.395 161.135 114.145 161.655 ;
        RECT 114.315 161.305 115.065 161.825 ;
        RECT 115.695 161.555 115.925 161.895 ;
        RECT 116.215 161.555 116.430 162.670 ;
        RECT 116.625 161.970 116.955 162.745 ;
        RECT 117.125 162.140 117.835 162.915 ;
        RECT 116.625 161.755 117.775 161.970 ;
        RECT 115.695 161.355 116.025 161.555 ;
        RECT 116.215 161.375 116.665 161.555 ;
        RECT 116.335 161.355 116.665 161.375 ;
        RECT 116.835 161.355 117.305 161.585 ;
        RECT 117.490 161.185 117.775 161.755 ;
        RECT 118.005 161.310 118.285 162.745 ;
        RECT 118.465 161.775 118.795 162.915 ;
        RECT 119.325 161.945 119.655 162.730 ;
        RECT 119.835 162.480 125.180 162.915 ;
        RECT 125.820 162.525 126.155 162.745 ;
        RECT 127.160 162.535 127.515 162.915 ;
        RECT 118.975 161.775 119.655 161.945 ;
        RECT 118.455 161.355 118.805 161.605 ;
        RECT 109.710 160.915 110.375 161.085 ;
        RECT 109.705 160.365 110.035 160.745 ;
        RECT 110.205 160.625 110.375 160.915 ;
        RECT 110.635 160.365 112.305 161.135 ;
        RECT 112.935 160.365 113.225 161.090 ;
        RECT 113.395 160.365 115.065 161.135 ;
        RECT 115.695 160.995 116.875 161.185 ;
        RECT 115.695 160.535 116.035 160.995 ;
        RECT 116.545 160.915 116.875 160.995 ;
        RECT 117.065 160.995 117.775 161.185 ;
        RECT 117.065 160.855 117.365 160.995 ;
        RECT 117.050 160.845 117.365 160.855 ;
        RECT 117.040 160.835 117.365 160.845 ;
        RECT 117.030 160.830 117.365 160.835 ;
        RECT 116.205 160.365 116.375 160.825 ;
        RECT 117.025 160.820 117.365 160.830 ;
        RECT 117.020 160.815 117.365 160.820 ;
        RECT 117.015 160.805 117.365 160.815 ;
        RECT 117.010 160.800 117.365 160.805 ;
        RECT 117.005 160.535 117.365 160.800 ;
        RECT 117.605 160.365 117.775 160.825 ;
        RECT 117.945 160.535 118.285 161.310 ;
        RECT 118.975 161.175 119.145 161.775 ;
        RECT 119.315 161.355 119.665 161.605 ;
        RECT 118.465 160.365 118.735 161.175 ;
        RECT 118.905 160.535 119.235 161.175 ;
        RECT 119.405 160.365 119.645 161.175 ;
        RECT 121.420 160.910 121.760 161.740 ;
        RECT 123.240 161.230 123.590 162.480 ;
        RECT 125.820 161.905 126.075 162.525 ;
        RECT 126.325 162.365 126.555 162.405 ;
        RECT 127.685 162.365 127.935 162.745 ;
        RECT 126.325 162.165 127.935 162.365 ;
        RECT 126.325 162.075 126.510 162.165 ;
        RECT 127.100 162.155 127.935 162.165 ;
        RECT 128.185 162.135 128.435 162.915 ;
        RECT 128.605 162.065 128.865 162.745 ;
        RECT 129.125 162.245 129.295 162.745 ;
        RECT 129.465 162.415 129.795 162.915 ;
        RECT 129.125 162.075 129.790 162.245 ;
        RECT 126.665 161.965 126.995 161.995 ;
        RECT 126.665 161.905 128.465 161.965 ;
        RECT 125.820 161.795 128.525 161.905 ;
        RECT 125.820 161.735 126.995 161.795 ;
        RECT 128.325 161.760 128.525 161.795 ;
        RECT 125.815 161.355 126.305 161.555 ;
        RECT 126.495 161.355 126.970 161.565 ;
        RECT 119.835 160.365 125.180 160.910 ;
        RECT 125.820 160.365 126.275 161.130 ;
        RECT 126.750 160.955 126.970 161.355 ;
        RECT 127.215 161.355 127.545 161.565 ;
        RECT 127.215 160.955 127.425 161.355 ;
        RECT 127.715 161.320 128.125 161.625 ;
        RECT 128.355 161.185 128.525 161.760 ;
        RECT 128.255 161.065 128.525 161.185 ;
        RECT 127.680 161.020 128.525 161.065 ;
        RECT 127.680 160.895 128.435 161.020 ;
        RECT 127.680 160.745 127.850 160.895 ;
        RECT 128.695 160.875 128.865 162.065 ;
        RECT 129.040 161.255 129.390 161.905 ;
        RECT 129.560 161.085 129.790 162.075 ;
        RECT 128.635 160.865 128.865 160.875 ;
        RECT 126.550 160.535 127.850 160.745 ;
        RECT 128.105 160.365 128.435 160.725 ;
        RECT 128.605 160.535 128.865 160.865 ;
        RECT 129.125 160.915 129.790 161.085 ;
        RECT 129.125 160.625 129.295 160.915 ;
        RECT 129.465 160.365 129.795 160.745 ;
        RECT 129.965 160.625 130.150 162.745 ;
        RECT 130.390 162.455 130.655 162.915 ;
        RECT 130.825 162.320 131.075 162.745 ;
        RECT 131.285 162.470 132.390 162.640 ;
        RECT 130.770 162.190 131.075 162.320 ;
        RECT 130.320 160.995 130.600 161.945 ;
        RECT 130.770 161.085 130.940 162.190 ;
        RECT 131.110 161.405 131.350 162.000 ;
        RECT 131.520 161.935 132.050 162.300 ;
        RECT 131.520 161.235 131.690 161.935 ;
        RECT 132.220 161.855 132.390 162.470 ;
        RECT 132.560 162.115 132.730 162.915 ;
        RECT 132.900 162.415 133.150 162.745 ;
        RECT 133.375 162.445 134.260 162.615 ;
        RECT 132.220 161.765 132.730 161.855 ;
        RECT 130.770 160.955 130.995 161.085 ;
        RECT 131.165 161.015 131.690 161.235 ;
        RECT 131.860 161.595 132.730 161.765 ;
        RECT 130.405 160.365 130.655 160.825 ;
        RECT 130.825 160.815 130.995 160.955 ;
        RECT 131.860 160.815 132.030 161.595 ;
        RECT 132.560 161.525 132.730 161.595 ;
        RECT 132.240 161.345 132.440 161.375 ;
        RECT 132.900 161.345 133.070 162.415 ;
        RECT 133.240 161.525 133.430 162.245 ;
        RECT 132.240 161.045 133.070 161.345 ;
        RECT 133.600 161.315 133.920 162.275 ;
        RECT 130.825 160.645 131.160 160.815 ;
        RECT 131.355 160.645 132.030 160.815 ;
        RECT 132.350 160.365 132.720 160.865 ;
        RECT 132.900 160.815 133.070 161.045 ;
        RECT 133.455 160.985 133.920 161.315 ;
        RECT 134.090 161.605 134.260 162.445 ;
        RECT 134.440 162.415 134.755 162.915 ;
        RECT 134.985 162.185 135.325 162.745 ;
        RECT 134.430 161.810 135.325 162.185 ;
        RECT 135.495 161.905 135.665 162.915 ;
        RECT 135.135 161.605 135.325 161.810 ;
        RECT 135.835 161.855 136.165 162.700 ;
        RECT 135.835 161.775 136.225 161.855 ;
        RECT 137.355 161.775 137.585 162.915 ;
        RECT 136.010 161.725 136.225 161.775 ;
        RECT 137.755 161.765 138.085 162.745 ;
        RECT 138.255 161.775 138.465 162.915 ;
        RECT 134.090 161.275 134.965 161.605 ;
        RECT 135.135 161.275 135.885 161.605 ;
        RECT 134.090 160.815 134.260 161.275 ;
        RECT 135.135 161.105 135.335 161.275 ;
        RECT 136.055 161.145 136.225 161.725 ;
        RECT 137.335 161.355 137.665 161.605 ;
        RECT 136.000 161.105 136.225 161.145 ;
        RECT 132.900 160.645 133.305 160.815 ;
        RECT 133.475 160.645 134.260 160.815 ;
        RECT 134.535 160.365 134.745 160.895 ;
        RECT 135.005 160.580 135.335 161.105 ;
        RECT 135.845 161.020 136.225 161.105 ;
        RECT 135.505 160.365 135.675 160.975 ;
        RECT 135.845 160.585 136.175 161.020 ;
        RECT 137.355 160.365 137.585 161.185 ;
        RECT 137.835 161.165 138.085 161.765 ;
        RECT 138.695 161.750 138.985 162.915 ;
        RECT 139.155 162.095 139.500 162.915 ;
        RECT 139.155 161.355 139.500 161.925 ;
        RECT 139.670 161.605 139.845 162.705 ;
        RECT 140.015 162.335 140.345 162.570 ;
        RECT 140.635 162.515 141.035 162.915 ;
        RECT 141.905 162.515 142.235 162.915 ;
        RECT 140.015 162.165 142.095 162.335 ;
        RECT 140.015 161.775 140.570 162.165 ;
        RECT 139.670 161.355 140.230 161.605 ;
        RECT 140.400 161.525 140.570 161.775 ;
        RECT 140.740 161.775 141.755 161.995 ;
        RECT 141.925 161.895 142.095 162.165 ;
        RECT 142.405 162.075 142.665 162.745 ;
        RECT 140.740 161.635 141.015 161.775 ;
        RECT 141.925 161.725 142.320 161.895 ;
        RECT 140.400 161.355 140.595 161.525 ;
        RECT 137.755 160.535 138.085 161.165 ;
        RECT 138.255 160.365 138.465 161.185 ;
        RECT 138.695 160.365 138.985 161.090 ;
        RECT 139.155 161.005 140.255 161.185 ;
        RECT 139.155 160.600 139.495 161.005 ;
        RECT 139.665 160.365 139.835 160.835 ;
        RECT 140.005 160.600 140.255 161.005 ;
        RECT 140.425 160.970 140.595 161.355 ;
        RECT 140.425 160.600 140.675 160.970 ;
        RECT 140.845 160.845 141.015 161.635 ;
        RECT 141.185 161.185 141.360 161.380 ;
        RECT 141.530 161.355 141.980 161.555 ;
        RECT 142.150 161.275 142.320 161.725 ;
        RECT 141.185 161.015 141.680 161.185 ;
        RECT 142.490 161.105 142.665 162.075 ;
        RECT 142.925 162.295 143.095 162.725 ;
        RECT 143.265 162.465 143.595 162.915 ;
        RECT 142.925 162.065 143.600 162.295 ;
        RECT 141.460 160.875 141.680 161.015 ;
        RECT 140.845 160.675 141.290 160.845 ;
        RECT 141.460 160.705 141.685 160.875 ;
        RECT 141.460 160.660 141.680 160.705 ;
        RECT 141.960 160.365 142.130 161.030 ;
        RECT 142.325 160.535 142.665 161.105 ;
        RECT 142.895 161.045 143.195 161.895 ;
        RECT 143.365 161.415 143.600 162.065 ;
        RECT 143.770 161.755 144.055 162.700 ;
        RECT 144.235 162.445 144.920 162.915 ;
        RECT 144.230 161.925 144.925 162.235 ;
        RECT 145.100 161.860 145.405 162.645 ;
        RECT 146.525 162.105 146.820 162.915 ;
        RECT 143.770 161.605 144.630 161.755 ;
        RECT 143.770 161.585 145.055 161.605 ;
        RECT 143.365 161.085 143.900 161.415 ;
        RECT 144.070 161.225 145.055 161.585 ;
        RECT 143.365 160.935 143.585 161.085 ;
        RECT 142.840 160.365 143.175 160.870 ;
        RECT 143.345 160.560 143.585 160.935 ;
        RECT 144.070 160.890 144.240 161.225 ;
        RECT 145.230 161.055 145.405 161.860 ;
        RECT 147.000 161.605 147.245 162.745 ;
        RECT 147.420 162.105 147.680 162.915 ;
        RECT 148.280 162.910 154.555 162.915 ;
        RECT 147.860 161.605 148.110 162.740 ;
        RECT 148.280 162.115 148.540 162.910 ;
        RECT 148.710 162.015 148.970 162.740 ;
        RECT 149.140 162.185 149.400 162.910 ;
        RECT 149.570 162.015 149.830 162.740 ;
        RECT 150.000 162.185 150.260 162.910 ;
        RECT 150.430 162.015 150.690 162.740 ;
        RECT 150.860 162.185 151.120 162.910 ;
        RECT 151.290 162.015 151.550 162.740 ;
        RECT 151.720 162.185 151.965 162.910 ;
        RECT 152.135 162.015 152.395 162.740 ;
        RECT 152.580 162.185 152.825 162.910 ;
        RECT 152.995 162.015 153.255 162.740 ;
        RECT 153.440 162.185 153.685 162.910 ;
        RECT 153.855 162.015 154.115 162.740 ;
        RECT 154.300 162.185 154.555 162.910 ;
        RECT 148.710 162.000 154.115 162.015 ;
        RECT 154.725 162.000 155.015 162.740 ;
        RECT 155.185 162.170 155.455 162.915 ;
        RECT 148.710 161.775 155.455 162.000 ;
        RECT 143.865 160.695 144.240 160.890 ;
        RECT 143.865 160.550 144.035 160.695 ;
        RECT 144.600 160.365 144.995 160.860 ;
        RECT 145.165 160.535 145.405 161.055 ;
        RECT 146.515 161.045 146.830 161.605 ;
        RECT 147.000 161.355 154.120 161.605 ;
        RECT 146.515 160.365 146.820 160.875 ;
        RECT 147.000 160.545 147.250 161.355 ;
        RECT 147.420 160.365 147.680 160.890 ;
        RECT 147.860 160.545 148.110 161.355 ;
        RECT 154.290 161.185 155.455 161.775 ;
        RECT 155.715 161.825 156.925 162.915 ;
        RECT 155.715 161.285 156.235 161.825 ;
        RECT 148.710 161.015 155.455 161.185 ;
        RECT 156.405 161.115 156.925 161.655 ;
        RECT 148.280 160.365 148.540 160.925 ;
        RECT 148.710 160.560 148.970 161.015 ;
        RECT 149.140 160.365 149.400 160.845 ;
        RECT 149.570 160.560 149.830 161.015 ;
        RECT 150.000 160.365 150.260 160.845 ;
        RECT 150.430 160.560 150.690 161.015 ;
        RECT 150.860 160.365 151.105 160.845 ;
        RECT 151.275 160.560 151.550 161.015 ;
        RECT 151.720 160.365 151.965 160.845 ;
        RECT 152.135 160.560 152.395 161.015 ;
        RECT 152.575 160.365 152.825 160.845 ;
        RECT 152.995 160.560 153.255 161.015 ;
        RECT 153.435 160.365 153.685 160.845 ;
        RECT 153.855 160.560 154.115 161.015 ;
        RECT 154.295 160.365 154.555 160.845 ;
        RECT 154.725 160.560 154.985 161.015 ;
        RECT 155.155 160.365 155.455 160.845 ;
        RECT 155.715 160.365 156.925 161.115 ;
        RECT 22.690 160.195 157.010 160.365 ;
        RECT 22.775 159.445 23.985 160.195 ;
        RECT 25.075 159.455 25.460 160.025 ;
        RECT 25.630 159.735 25.955 160.195 ;
        RECT 26.475 159.565 26.755 160.025 ;
        RECT 22.775 158.905 23.295 159.445 ;
        RECT 23.465 158.735 23.985 159.275 ;
        RECT 22.775 157.645 23.985 158.735 ;
        RECT 25.075 158.785 25.355 159.455 ;
        RECT 25.630 159.395 26.755 159.565 ;
        RECT 25.630 159.285 26.080 159.395 ;
        RECT 25.525 158.955 26.080 159.285 ;
        RECT 26.945 159.225 27.345 160.025 ;
        RECT 27.745 159.735 28.015 160.195 ;
        RECT 28.185 159.565 28.470 160.025 ;
        RECT 28.845 159.715 29.145 160.195 ;
        RECT 25.075 157.815 25.460 158.785 ;
        RECT 25.630 158.495 26.080 158.955 ;
        RECT 26.250 158.665 27.345 159.225 ;
        RECT 25.630 158.275 26.755 158.495 ;
        RECT 25.630 157.645 25.955 158.105 ;
        RECT 26.475 157.815 26.755 158.275 ;
        RECT 26.945 157.815 27.345 158.665 ;
        RECT 27.515 159.395 28.470 159.565 ;
        RECT 29.315 159.545 29.575 160.000 ;
        RECT 29.745 159.715 30.005 160.195 ;
        RECT 30.185 159.545 30.445 160.000 ;
        RECT 30.615 159.715 30.865 160.195 ;
        RECT 31.045 159.545 31.305 160.000 ;
        RECT 31.475 159.715 31.725 160.195 ;
        RECT 31.905 159.545 32.165 160.000 ;
        RECT 32.335 159.715 32.580 160.195 ;
        RECT 32.750 159.545 33.025 160.000 ;
        RECT 33.195 159.715 33.440 160.195 ;
        RECT 33.610 159.545 33.870 160.000 ;
        RECT 34.040 159.715 34.300 160.195 ;
        RECT 34.470 159.545 34.730 160.000 ;
        RECT 34.900 159.715 35.160 160.195 ;
        RECT 35.330 159.545 35.590 160.000 ;
        RECT 35.760 159.635 36.020 160.195 ;
        RECT 27.515 158.495 27.725 159.395 ;
        RECT 28.845 159.375 35.590 159.545 ;
        RECT 27.895 158.665 28.585 159.225 ;
        RECT 28.845 159.175 30.010 159.375 ;
        RECT 36.190 159.205 36.440 160.015 ;
        RECT 36.620 159.670 36.880 160.195 ;
        RECT 37.050 159.205 37.300 160.015 ;
        RECT 37.480 159.685 37.785 160.195 ;
        RECT 38.045 159.645 38.215 159.935 ;
        RECT 38.385 159.815 38.715 160.195 ;
        RECT 28.815 159.005 30.010 159.175 ;
        RECT 28.845 158.785 30.010 159.005 ;
        RECT 30.180 158.955 37.300 159.205 ;
        RECT 37.470 158.955 37.785 159.515 ;
        RECT 38.045 159.475 38.710 159.645 ;
        RECT 28.845 158.560 35.590 158.785 ;
        RECT 27.515 158.275 28.470 158.495 ;
        RECT 27.745 157.645 28.015 158.105 ;
        RECT 28.185 157.815 28.470 158.275 ;
        RECT 28.845 157.645 29.115 158.390 ;
        RECT 29.285 157.820 29.575 158.560 ;
        RECT 30.185 158.545 35.590 158.560 ;
        RECT 29.745 157.650 30.000 158.375 ;
        RECT 30.185 157.820 30.445 158.545 ;
        RECT 30.615 157.650 30.860 158.375 ;
        RECT 31.045 157.820 31.305 158.545 ;
        RECT 31.475 157.650 31.720 158.375 ;
        RECT 31.905 157.820 32.165 158.545 ;
        RECT 32.335 157.650 32.580 158.375 ;
        RECT 32.750 157.820 33.010 158.545 ;
        RECT 33.180 157.650 33.440 158.375 ;
        RECT 33.610 157.820 33.870 158.545 ;
        RECT 34.040 157.650 34.300 158.375 ;
        RECT 34.470 157.820 34.730 158.545 ;
        RECT 34.900 157.650 35.160 158.375 ;
        RECT 35.330 157.820 35.590 158.545 ;
        RECT 35.760 157.650 36.020 158.445 ;
        RECT 36.190 157.820 36.440 158.955 ;
        RECT 29.745 157.645 36.020 157.650 ;
        RECT 36.620 157.645 36.880 158.455 ;
        RECT 37.055 157.815 37.300 158.955 ;
        RECT 37.960 158.655 38.310 159.305 ;
        RECT 38.480 158.485 38.710 159.475 ;
        RECT 37.480 157.645 37.775 158.455 ;
        RECT 38.045 158.315 38.710 158.485 ;
        RECT 38.045 157.815 38.215 158.315 ;
        RECT 38.385 157.645 38.715 158.145 ;
        RECT 38.885 157.815 39.070 159.935 ;
        RECT 39.325 159.735 39.575 160.195 ;
        RECT 39.745 159.745 40.080 159.915 ;
        RECT 40.275 159.745 40.950 159.915 ;
        RECT 39.745 159.605 39.915 159.745 ;
        RECT 39.240 158.615 39.520 159.565 ;
        RECT 39.690 159.475 39.915 159.605 ;
        RECT 39.690 158.370 39.860 159.475 ;
        RECT 40.085 159.325 40.610 159.545 ;
        RECT 40.030 158.560 40.270 159.155 ;
        RECT 40.440 158.625 40.610 159.325 ;
        RECT 40.780 158.965 40.950 159.745 ;
        RECT 41.270 159.695 41.640 160.195 ;
        RECT 41.820 159.745 42.225 159.915 ;
        RECT 42.395 159.745 43.180 159.915 ;
        RECT 41.820 159.515 41.990 159.745 ;
        RECT 41.160 159.215 41.990 159.515 ;
        RECT 42.375 159.245 42.840 159.575 ;
        RECT 41.160 159.185 41.360 159.215 ;
        RECT 41.480 158.965 41.650 159.035 ;
        RECT 40.780 158.795 41.650 158.965 ;
        RECT 41.140 158.705 41.650 158.795 ;
        RECT 39.690 158.240 39.995 158.370 ;
        RECT 40.440 158.260 40.970 158.625 ;
        RECT 39.310 157.645 39.575 158.105 ;
        RECT 39.745 157.815 39.995 158.240 ;
        RECT 41.140 158.090 41.310 158.705 ;
        RECT 40.205 157.920 41.310 158.090 ;
        RECT 41.480 157.645 41.650 158.445 ;
        RECT 41.820 158.145 41.990 159.215 ;
        RECT 42.160 158.315 42.350 159.035 ;
        RECT 42.520 158.285 42.840 159.245 ;
        RECT 43.010 159.285 43.180 159.745 ;
        RECT 43.455 159.665 43.665 160.195 ;
        RECT 43.925 159.455 44.255 159.980 ;
        RECT 44.425 159.585 44.595 160.195 ;
        RECT 44.765 159.540 45.095 159.975 ;
        RECT 44.765 159.455 45.145 159.540 ;
        RECT 44.055 159.285 44.255 159.455 ;
        RECT 44.920 159.415 45.145 159.455 ;
        RECT 43.010 158.955 43.885 159.285 ;
        RECT 44.055 158.955 44.805 159.285 ;
        RECT 41.820 157.815 42.070 158.145 ;
        RECT 43.010 158.115 43.180 158.955 ;
        RECT 44.055 158.750 44.245 158.955 ;
        RECT 44.975 158.835 45.145 159.415 ;
        RECT 44.930 158.785 45.145 158.835 ;
        RECT 43.350 158.375 44.245 158.750 ;
        RECT 44.755 158.705 45.145 158.785 ;
        RECT 42.295 157.945 43.180 158.115 ;
        RECT 43.360 157.645 43.675 158.145 ;
        RECT 43.905 157.815 44.245 158.375 ;
        RECT 44.415 157.645 44.585 158.655 ;
        RECT 44.755 157.860 45.085 158.705 ;
        RECT 45.325 157.825 45.585 160.015 ;
        RECT 45.845 159.825 46.515 160.195 ;
        RECT 46.695 159.645 47.005 160.015 ;
        RECT 45.775 159.445 47.005 159.645 ;
        RECT 45.775 158.775 46.065 159.445 ;
        RECT 47.185 159.265 47.415 159.905 ;
        RECT 47.595 159.465 47.885 160.195 ;
        RECT 48.535 159.470 48.825 160.195 ;
        RECT 48.995 159.425 52.505 160.195 ;
        RECT 53.140 159.690 53.475 160.195 ;
        RECT 53.645 159.625 53.885 160.000 ;
        RECT 54.165 159.865 54.335 160.010 ;
        RECT 54.165 159.670 54.540 159.865 ;
        RECT 54.900 159.700 55.295 160.195 ;
        RECT 46.245 158.955 46.710 159.265 ;
        RECT 46.890 158.955 47.415 159.265 ;
        RECT 47.595 158.955 47.895 159.285 ;
        RECT 48.995 158.905 50.645 159.425 ;
        RECT 45.775 158.555 46.545 158.775 ;
        RECT 45.755 157.645 46.095 158.375 ;
        RECT 46.275 157.825 46.545 158.555 ;
        RECT 46.725 158.535 47.885 158.775 ;
        RECT 46.725 157.825 46.955 158.535 ;
        RECT 47.125 157.645 47.455 158.355 ;
        RECT 47.625 157.825 47.885 158.535 ;
        RECT 48.535 157.645 48.825 158.810 ;
        RECT 50.815 158.735 52.505 159.255 ;
        RECT 48.995 157.645 52.505 158.735 ;
        RECT 53.195 158.665 53.495 159.515 ;
        RECT 53.665 159.475 53.885 159.625 ;
        RECT 53.665 159.145 54.200 159.475 ;
        RECT 54.370 159.335 54.540 159.670 ;
        RECT 55.465 159.505 55.705 160.025 ;
        RECT 53.665 158.495 53.900 159.145 ;
        RECT 54.370 158.975 55.355 159.335 ;
        RECT 53.225 158.265 53.900 158.495 ;
        RECT 54.070 158.955 55.355 158.975 ;
        RECT 54.070 158.805 54.930 158.955 ;
        RECT 53.225 157.835 53.395 158.265 ;
        RECT 53.565 157.645 53.895 158.095 ;
        RECT 54.070 157.860 54.355 158.805 ;
        RECT 55.530 158.700 55.705 159.505 ;
        RECT 55.980 159.625 56.155 160.025 ;
        RECT 56.325 159.815 56.655 160.195 ;
        RECT 56.900 159.695 57.130 160.025 ;
        RECT 55.980 159.455 56.610 159.625 ;
        RECT 56.440 159.285 56.610 159.455 ;
        RECT 54.530 158.325 55.225 158.635 ;
        RECT 54.535 157.645 55.220 158.115 ;
        RECT 55.400 157.915 55.705 158.700 ;
        RECT 55.895 158.605 56.260 159.285 ;
        RECT 56.440 158.955 56.790 159.285 ;
        RECT 56.440 158.435 56.610 158.955 ;
        RECT 55.980 158.265 56.610 158.435 ;
        RECT 56.960 158.405 57.130 159.695 ;
        RECT 57.330 158.585 57.610 159.860 ;
        RECT 57.835 158.835 58.105 159.860 ;
        RECT 58.565 159.815 58.895 160.195 ;
        RECT 59.065 159.940 59.400 159.985 ;
        RECT 57.795 158.665 58.105 158.835 ;
        RECT 57.835 158.585 58.105 158.665 ;
        RECT 58.295 158.585 58.635 159.615 ;
        RECT 59.065 159.475 59.405 159.940 ;
        RECT 59.625 159.540 59.955 159.975 ;
        RECT 60.125 159.585 60.295 160.195 ;
        RECT 58.805 158.955 59.065 159.285 ;
        RECT 58.805 158.405 58.975 158.955 ;
        RECT 59.235 158.785 59.405 159.475 ;
        RECT 55.980 157.815 56.155 158.265 ;
        RECT 56.960 158.235 58.975 158.405 ;
        RECT 56.325 157.645 56.655 158.085 ;
        RECT 56.960 157.815 57.130 158.235 ;
        RECT 57.365 157.645 58.035 158.055 ;
        RECT 58.250 157.815 58.420 158.235 ;
        RECT 58.620 157.645 58.950 158.055 ;
        RECT 59.145 157.815 59.405 158.785 ;
        RECT 59.575 159.455 59.955 159.540 ;
        RECT 60.465 159.455 60.795 159.980 ;
        RECT 61.055 159.665 61.265 160.195 ;
        RECT 61.540 159.745 62.325 159.915 ;
        RECT 62.495 159.745 62.900 159.915 ;
        RECT 59.575 159.415 59.800 159.455 ;
        RECT 59.575 158.835 59.745 159.415 ;
        RECT 60.465 159.285 60.665 159.455 ;
        RECT 61.540 159.285 61.710 159.745 ;
        RECT 59.915 158.955 60.665 159.285 ;
        RECT 60.835 158.955 61.710 159.285 ;
        RECT 59.575 158.785 59.790 158.835 ;
        RECT 59.575 158.705 59.965 158.785 ;
        RECT 59.635 157.860 59.965 158.705 ;
        RECT 60.475 158.750 60.665 158.955 ;
        RECT 60.135 157.645 60.305 158.655 ;
        RECT 60.475 158.375 61.370 158.750 ;
        RECT 60.475 157.815 60.815 158.375 ;
        RECT 61.045 157.645 61.360 158.145 ;
        RECT 61.540 158.115 61.710 158.955 ;
        RECT 61.880 159.245 62.345 159.575 ;
        RECT 62.730 159.515 62.900 159.745 ;
        RECT 63.080 159.695 63.450 160.195 ;
        RECT 63.770 159.745 64.445 159.915 ;
        RECT 64.640 159.745 64.975 159.915 ;
        RECT 61.880 158.285 62.200 159.245 ;
        RECT 62.730 159.215 63.560 159.515 ;
        RECT 62.370 158.315 62.560 159.035 ;
        RECT 62.730 158.145 62.900 159.215 ;
        RECT 63.360 159.185 63.560 159.215 ;
        RECT 63.070 158.965 63.240 159.035 ;
        RECT 63.770 158.965 63.940 159.745 ;
        RECT 64.805 159.605 64.975 159.745 ;
        RECT 65.145 159.735 65.395 160.195 ;
        RECT 63.070 158.795 63.940 158.965 ;
        RECT 64.110 159.325 64.635 159.545 ;
        RECT 64.805 159.475 65.030 159.605 ;
        RECT 63.070 158.705 63.580 158.795 ;
        RECT 61.540 157.945 62.425 158.115 ;
        RECT 62.650 157.815 62.900 158.145 ;
        RECT 63.070 157.645 63.240 158.445 ;
        RECT 63.410 158.090 63.580 158.705 ;
        RECT 64.110 158.625 64.280 159.325 ;
        RECT 63.750 158.260 64.280 158.625 ;
        RECT 64.450 158.560 64.690 159.155 ;
        RECT 64.860 158.370 65.030 159.475 ;
        RECT 65.200 158.615 65.480 159.565 ;
        RECT 64.725 158.240 65.030 158.370 ;
        RECT 63.410 157.920 64.515 158.090 ;
        RECT 64.725 157.815 64.975 158.240 ;
        RECT 65.145 157.645 65.410 158.105 ;
        RECT 65.650 157.815 65.835 159.935 ;
        RECT 66.005 159.815 66.335 160.195 ;
        RECT 66.505 159.645 66.675 159.935 ;
        RECT 66.010 159.475 66.675 159.645 ;
        RECT 66.985 159.540 67.315 159.975 ;
        RECT 67.485 159.585 67.655 160.195 ;
        RECT 66.010 158.485 66.240 159.475 ;
        RECT 66.935 159.455 67.315 159.540 ;
        RECT 67.825 159.455 68.155 159.980 ;
        RECT 68.415 159.665 68.625 160.195 ;
        RECT 68.900 159.745 69.685 159.915 ;
        RECT 69.855 159.745 70.260 159.915 ;
        RECT 66.935 159.415 67.160 159.455 ;
        RECT 66.410 158.655 66.760 159.305 ;
        RECT 66.935 158.835 67.105 159.415 ;
        RECT 67.825 159.285 68.025 159.455 ;
        RECT 68.900 159.285 69.070 159.745 ;
        RECT 67.275 158.955 68.025 159.285 ;
        RECT 68.195 158.955 69.070 159.285 ;
        RECT 66.935 158.785 67.150 158.835 ;
        RECT 66.935 158.705 67.325 158.785 ;
        RECT 66.010 158.315 66.675 158.485 ;
        RECT 66.005 157.645 66.335 158.145 ;
        RECT 66.505 157.815 66.675 158.315 ;
        RECT 66.995 157.860 67.325 158.705 ;
        RECT 67.835 158.750 68.025 158.955 ;
        RECT 67.495 157.645 67.665 158.655 ;
        RECT 67.835 158.375 68.730 158.750 ;
        RECT 67.835 157.815 68.175 158.375 ;
        RECT 68.405 157.645 68.720 158.145 ;
        RECT 68.900 158.115 69.070 158.955 ;
        RECT 69.240 159.245 69.705 159.575 ;
        RECT 70.090 159.515 70.260 159.745 ;
        RECT 70.440 159.695 70.810 160.195 ;
        RECT 71.130 159.745 71.805 159.915 ;
        RECT 72.000 159.745 72.335 159.915 ;
        RECT 69.240 158.285 69.560 159.245 ;
        RECT 70.090 159.215 70.920 159.515 ;
        RECT 69.730 158.315 69.920 159.035 ;
        RECT 70.090 158.145 70.260 159.215 ;
        RECT 70.720 159.185 70.920 159.215 ;
        RECT 70.430 158.965 70.600 159.035 ;
        RECT 71.130 158.965 71.300 159.745 ;
        RECT 72.165 159.605 72.335 159.745 ;
        RECT 72.505 159.735 72.755 160.195 ;
        RECT 70.430 158.795 71.300 158.965 ;
        RECT 71.470 159.325 71.995 159.545 ;
        RECT 72.165 159.475 72.390 159.605 ;
        RECT 70.430 158.705 70.940 158.795 ;
        RECT 68.900 157.945 69.785 158.115 ;
        RECT 70.010 157.815 70.260 158.145 ;
        RECT 70.430 157.645 70.600 158.445 ;
        RECT 70.770 158.090 70.940 158.705 ;
        RECT 71.470 158.625 71.640 159.325 ;
        RECT 71.110 158.260 71.640 158.625 ;
        RECT 71.810 158.560 72.050 159.155 ;
        RECT 72.220 158.370 72.390 159.475 ;
        RECT 72.560 158.615 72.840 159.565 ;
        RECT 72.085 158.240 72.390 158.370 ;
        RECT 70.770 157.920 71.875 158.090 ;
        RECT 72.085 157.815 72.335 158.240 ;
        RECT 72.505 157.645 72.770 158.105 ;
        RECT 73.010 157.815 73.195 159.935 ;
        RECT 73.365 159.815 73.695 160.195 ;
        RECT 73.865 159.645 74.035 159.935 ;
        RECT 73.370 159.475 74.035 159.645 ;
        RECT 73.370 158.485 73.600 159.475 ;
        RECT 74.295 159.470 74.585 160.195 ;
        RECT 74.845 159.645 75.015 160.025 ;
        RECT 75.230 159.815 75.560 160.195 ;
        RECT 74.845 159.475 75.560 159.645 ;
        RECT 73.770 158.655 74.120 159.305 ;
        RECT 74.755 158.925 75.110 159.295 ;
        RECT 75.390 159.285 75.560 159.475 ;
        RECT 75.730 159.450 75.985 160.025 ;
        RECT 75.390 158.955 75.645 159.285 ;
        RECT 73.370 158.315 74.035 158.485 ;
        RECT 73.365 157.645 73.695 158.145 ;
        RECT 73.865 157.815 74.035 158.315 ;
        RECT 74.295 157.645 74.585 158.810 ;
        RECT 75.390 158.745 75.560 158.955 ;
        RECT 74.845 158.575 75.560 158.745 ;
        RECT 75.815 158.720 75.985 159.450 ;
        RECT 76.160 159.355 76.420 160.195 ;
        RECT 76.595 159.425 80.105 160.195 ;
        RECT 80.475 159.565 80.805 159.925 ;
        RECT 81.425 159.735 81.675 160.195 ;
        RECT 81.845 159.735 82.405 160.025 ;
        RECT 76.595 158.905 78.245 159.425 ;
        RECT 80.475 159.375 81.865 159.565 ;
        RECT 81.695 159.285 81.865 159.375 ;
        RECT 74.845 157.815 75.015 158.575 ;
        RECT 75.230 157.645 75.560 158.405 ;
        RECT 75.730 157.815 75.985 158.720 ;
        RECT 76.160 157.645 76.420 158.795 ;
        RECT 78.415 158.735 80.105 159.255 ;
        RECT 76.595 157.645 80.105 158.735 ;
        RECT 80.290 158.955 80.965 159.205 ;
        RECT 81.185 158.955 81.525 159.205 ;
        RECT 81.695 158.955 81.985 159.285 ;
        RECT 80.290 158.595 80.555 158.955 ;
        RECT 81.695 158.705 81.865 158.955 ;
        RECT 80.925 158.535 81.865 158.705 ;
        RECT 80.475 157.645 80.755 158.315 ;
        RECT 80.925 157.985 81.225 158.535 ;
        RECT 82.155 158.365 82.405 159.735 ;
        RECT 81.425 157.645 81.755 158.365 ;
        RECT 81.945 157.815 82.405 158.365 ;
        RECT 82.575 159.520 82.835 160.025 ;
        RECT 83.015 159.815 83.345 160.195 ;
        RECT 83.525 159.645 83.695 160.025 ;
        RECT 82.575 158.720 82.745 159.520 ;
        RECT 83.030 159.475 83.695 159.645 ;
        RECT 83.030 159.220 83.200 159.475 ;
        RECT 83.955 159.425 86.545 160.195 ;
        RECT 82.915 158.890 83.200 159.220 ;
        RECT 83.435 158.925 83.765 159.295 ;
        RECT 83.955 158.905 85.165 159.425 ;
        RECT 87.175 159.375 87.435 160.195 ;
        RECT 87.605 159.375 87.935 159.795 ;
        RECT 88.115 159.625 88.375 160.025 ;
        RECT 88.545 159.795 88.875 160.195 ;
        RECT 89.045 159.625 89.215 159.975 ;
        RECT 89.385 159.795 89.760 160.195 ;
        RECT 88.115 159.455 89.780 159.625 ;
        RECT 89.950 159.520 90.225 159.865 ;
        RECT 87.685 159.285 87.935 159.375 ;
        RECT 89.610 159.285 89.780 159.455 ;
        RECT 83.030 158.745 83.200 158.890 ;
        RECT 82.575 157.815 82.845 158.720 ;
        RECT 83.030 158.575 83.695 158.745 ;
        RECT 85.335 158.735 86.545 159.255 ;
        RECT 87.180 158.955 87.515 159.205 ;
        RECT 87.685 158.955 88.400 159.285 ;
        RECT 88.615 158.955 89.440 159.285 ;
        RECT 89.610 158.955 89.885 159.285 ;
        RECT 83.015 157.645 83.345 158.405 ;
        RECT 83.525 157.815 83.695 158.575 ;
        RECT 83.955 157.645 86.545 158.735 ;
        RECT 87.175 157.645 87.435 158.785 ;
        RECT 87.685 158.395 87.855 158.955 ;
        RECT 88.115 158.495 88.445 158.785 ;
        RECT 88.615 158.665 88.860 158.955 ;
        RECT 89.610 158.785 89.780 158.955 ;
        RECT 90.055 158.785 90.225 159.520 ;
        RECT 89.120 158.615 89.780 158.785 ;
        RECT 89.120 158.495 89.290 158.615 ;
        RECT 88.115 158.325 89.290 158.495 ;
        RECT 87.675 157.825 89.290 158.155 ;
        RECT 89.460 157.645 89.740 158.445 ;
        RECT 89.950 157.815 90.225 158.785 ;
        RECT 90.395 159.695 90.695 160.025 ;
        RECT 90.865 159.715 91.140 160.195 ;
        RECT 90.395 158.785 90.565 159.695 ;
        RECT 91.320 159.545 91.615 159.935 ;
        RECT 91.785 159.715 92.040 160.195 ;
        RECT 92.215 159.545 92.475 159.935 ;
        RECT 92.645 159.715 92.925 160.195 ;
        RECT 90.735 158.955 91.085 159.525 ;
        RECT 91.320 159.375 92.970 159.545 ;
        RECT 91.255 159.035 92.395 159.205 ;
        RECT 91.255 158.785 91.425 159.035 ;
        RECT 92.565 158.865 92.970 159.375 ;
        RECT 93.155 159.445 94.365 160.195 ;
        RECT 94.735 159.565 95.065 159.925 ;
        RECT 95.685 159.735 95.935 160.195 ;
        RECT 96.105 159.735 96.665 160.025 ;
        RECT 93.155 158.905 93.675 159.445 ;
        RECT 94.735 159.375 96.125 159.565 ;
        RECT 95.955 159.285 96.125 159.375 ;
        RECT 90.395 158.615 91.425 158.785 ;
        RECT 92.215 158.695 92.970 158.865 ;
        RECT 93.845 158.735 94.365 159.275 ;
        RECT 90.395 157.815 90.705 158.615 ;
        RECT 92.215 158.445 92.475 158.695 ;
        RECT 90.875 157.645 91.185 158.445 ;
        RECT 91.355 158.275 92.475 158.445 ;
        RECT 91.355 157.815 91.615 158.275 ;
        RECT 91.785 157.645 92.040 158.105 ;
        RECT 92.215 157.815 92.475 158.275 ;
        RECT 92.645 157.645 92.930 158.515 ;
        RECT 93.155 157.645 94.365 158.735 ;
        RECT 94.550 158.955 95.225 159.205 ;
        RECT 95.445 158.955 95.785 159.205 ;
        RECT 95.955 158.955 96.245 159.285 ;
        RECT 94.550 158.595 94.815 158.955 ;
        RECT 95.955 158.705 96.125 158.955 ;
        RECT 95.185 158.535 96.125 158.705 ;
        RECT 94.735 157.645 95.015 158.315 ;
        RECT 95.185 157.985 95.485 158.535 ;
        RECT 96.415 158.365 96.665 159.735 ;
        RECT 96.925 159.645 97.095 160.025 ;
        RECT 97.275 159.815 97.605 160.195 ;
        RECT 96.925 159.475 97.590 159.645 ;
        RECT 97.785 159.520 98.045 160.025 ;
        RECT 96.855 158.925 97.185 159.295 ;
        RECT 97.420 159.220 97.590 159.475 ;
        RECT 97.420 158.890 97.705 159.220 ;
        RECT 97.420 158.745 97.590 158.890 ;
        RECT 95.685 157.645 96.015 158.365 ;
        RECT 96.205 157.815 96.665 158.365 ;
        RECT 96.925 158.575 97.590 158.745 ;
        RECT 97.875 158.720 98.045 159.520 ;
        RECT 98.215 159.425 99.885 160.195 ;
        RECT 100.055 159.470 100.345 160.195 ;
        RECT 100.605 159.715 100.905 160.195 ;
        RECT 101.075 159.545 101.335 160.000 ;
        RECT 101.505 159.715 101.765 160.195 ;
        RECT 101.945 159.545 102.205 160.000 ;
        RECT 102.375 159.715 102.625 160.195 ;
        RECT 102.805 159.545 103.065 160.000 ;
        RECT 103.235 159.715 103.485 160.195 ;
        RECT 103.665 159.545 103.925 160.000 ;
        RECT 104.095 159.715 104.340 160.195 ;
        RECT 104.510 159.545 104.785 160.000 ;
        RECT 104.955 159.715 105.200 160.195 ;
        RECT 105.370 159.545 105.630 160.000 ;
        RECT 105.800 159.715 106.060 160.195 ;
        RECT 106.230 159.545 106.490 160.000 ;
        RECT 106.660 159.715 106.920 160.195 ;
        RECT 107.090 159.545 107.350 160.000 ;
        RECT 107.520 159.635 107.780 160.195 ;
        RECT 98.215 158.905 98.965 159.425 ;
        RECT 100.605 159.375 107.350 159.545 ;
        RECT 99.135 158.735 99.885 159.255 ;
        RECT 96.925 157.815 97.095 158.575 ;
        RECT 97.275 157.645 97.605 158.405 ;
        RECT 97.775 157.815 98.045 158.720 ;
        RECT 98.215 157.645 99.885 158.735 ;
        RECT 100.055 157.645 100.345 158.810 ;
        RECT 100.605 158.785 101.770 159.375 ;
        RECT 107.950 159.205 108.200 160.015 ;
        RECT 108.380 159.670 108.640 160.195 ;
        RECT 108.810 159.205 109.060 160.015 ;
        RECT 109.240 159.685 109.545 160.195 ;
        RECT 109.805 159.645 109.975 159.935 ;
        RECT 110.145 159.815 110.475 160.195 ;
        RECT 101.940 158.955 109.060 159.205 ;
        RECT 109.230 158.955 109.545 159.515 ;
        RECT 109.805 159.475 110.470 159.645 ;
        RECT 100.605 158.560 107.350 158.785 ;
        RECT 100.605 157.645 100.875 158.390 ;
        RECT 101.045 157.820 101.335 158.560 ;
        RECT 101.945 158.545 107.350 158.560 ;
        RECT 101.505 157.650 101.760 158.375 ;
        RECT 101.945 157.820 102.205 158.545 ;
        RECT 102.375 157.650 102.620 158.375 ;
        RECT 102.805 157.820 103.065 158.545 ;
        RECT 103.235 157.650 103.480 158.375 ;
        RECT 103.665 157.820 103.925 158.545 ;
        RECT 104.095 157.650 104.340 158.375 ;
        RECT 104.510 157.820 104.770 158.545 ;
        RECT 104.940 157.650 105.200 158.375 ;
        RECT 105.370 157.820 105.630 158.545 ;
        RECT 105.800 157.650 106.060 158.375 ;
        RECT 106.230 157.820 106.490 158.545 ;
        RECT 106.660 157.650 106.920 158.375 ;
        RECT 107.090 157.820 107.350 158.545 ;
        RECT 107.520 157.650 107.780 158.445 ;
        RECT 107.950 157.820 108.200 158.955 ;
        RECT 101.505 157.645 107.780 157.650 ;
        RECT 108.380 157.645 108.640 158.455 ;
        RECT 108.815 157.815 109.060 158.955 ;
        RECT 109.720 158.655 110.070 159.305 ;
        RECT 110.240 158.485 110.470 159.475 ;
        RECT 109.240 157.645 109.535 158.455 ;
        RECT 109.805 158.315 110.470 158.485 ;
        RECT 109.805 157.815 109.975 158.315 ;
        RECT 110.145 157.645 110.475 158.145 ;
        RECT 110.645 157.815 110.830 159.935 ;
        RECT 111.085 159.735 111.335 160.195 ;
        RECT 111.505 159.745 111.840 159.915 ;
        RECT 112.035 159.745 112.710 159.915 ;
        RECT 111.505 159.605 111.675 159.745 ;
        RECT 111.000 158.615 111.280 159.565 ;
        RECT 111.450 159.475 111.675 159.605 ;
        RECT 111.450 158.370 111.620 159.475 ;
        RECT 111.845 159.325 112.370 159.545 ;
        RECT 111.790 158.560 112.030 159.155 ;
        RECT 112.200 158.625 112.370 159.325 ;
        RECT 112.540 158.965 112.710 159.745 ;
        RECT 113.030 159.695 113.400 160.195 ;
        RECT 113.580 159.745 113.985 159.915 ;
        RECT 114.155 159.745 114.940 159.915 ;
        RECT 113.580 159.515 113.750 159.745 ;
        RECT 112.920 159.215 113.750 159.515 ;
        RECT 114.135 159.245 114.600 159.575 ;
        RECT 112.920 159.185 113.120 159.215 ;
        RECT 113.240 158.965 113.410 159.035 ;
        RECT 112.540 158.795 113.410 158.965 ;
        RECT 112.900 158.705 113.410 158.795 ;
        RECT 111.450 158.240 111.755 158.370 ;
        RECT 112.200 158.260 112.730 158.625 ;
        RECT 111.070 157.645 111.335 158.105 ;
        RECT 111.505 157.815 111.755 158.240 ;
        RECT 112.900 158.090 113.070 158.705 ;
        RECT 111.965 157.920 113.070 158.090 ;
        RECT 113.240 157.645 113.410 158.445 ;
        RECT 113.580 158.145 113.750 159.215 ;
        RECT 113.920 158.315 114.110 159.035 ;
        RECT 114.280 158.285 114.600 159.245 ;
        RECT 114.770 159.285 114.940 159.745 ;
        RECT 115.215 159.665 115.425 160.195 ;
        RECT 115.685 159.455 116.015 159.980 ;
        RECT 116.185 159.585 116.355 160.195 ;
        RECT 116.525 159.540 116.855 159.975 ;
        RECT 116.525 159.455 116.905 159.540 ;
        RECT 115.815 159.285 116.015 159.455 ;
        RECT 116.680 159.415 116.905 159.455 ;
        RECT 114.770 158.955 115.645 159.285 ;
        RECT 115.815 158.955 116.565 159.285 ;
        RECT 113.580 157.815 113.830 158.145 ;
        RECT 114.770 158.115 114.940 158.955 ;
        RECT 115.815 158.750 116.005 158.955 ;
        RECT 116.735 158.835 116.905 159.415 ;
        RECT 116.690 158.785 116.905 158.835 ;
        RECT 115.110 158.375 116.005 158.750 ;
        RECT 116.515 158.705 116.905 158.785 ;
        RECT 117.075 159.520 117.335 160.025 ;
        RECT 117.515 159.815 117.845 160.195 ;
        RECT 118.025 159.645 118.195 160.025 ;
        RECT 117.075 158.720 117.245 159.520 ;
        RECT 117.530 159.475 118.195 159.645 ;
        RECT 117.530 159.220 117.700 159.475 ;
        RECT 118.455 159.425 121.965 160.195 ;
        RECT 122.135 159.445 123.345 160.195 ;
        RECT 123.605 159.645 123.775 160.025 ;
        RECT 123.955 159.815 124.285 160.195 ;
        RECT 123.605 159.475 124.270 159.645 ;
        RECT 124.465 159.520 124.725 160.025 ;
        RECT 117.415 158.890 117.700 159.220 ;
        RECT 117.935 158.925 118.265 159.295 ;
        RECT 118.455 158.905 120.105 159.425 ;
        RECT 117.530 158.745 117.700 158.890 ;
        RECT 114.055 157.945 114.940 158.115 ;
        RECT 115.120 157.645 115.435 158.145 ;
        RECT 115.665 157.815 116.005 158.375 ;
        RECT 116.175 157.645 116.345 158.655 ;
        RECT 116.515 157.860 116.845 158.705 ;
        RECT 117.075 157.815 117.345 158.720 ;
        RECT 117.530 158.575 118.195 158.745 ;
        RECT 120.275 158.735 121.965 159.255 ;
        RECT 122.135 158.905 122.655 159.445 ;
        RECT 122.825 158.735 123.345 159.275 ;
        RECT 123.535 158.925 123.865 159.295 ;
        RECT 124.100 159.220 124.270 159.475 ;
        RECT 124.100 158.890 124.385 159.220 ;
        RECT 124.100 158.745 124.270 158.890 ;
        RECT 117.515 157.645 117.845 158.405 ;
        RECT 118.025 157.815 118.195 158.575 ;
        RECT 118.455 157.645 121.965 158.735 ;
        RECT 122.135 157.645 123.345 158.735 ;
        RECT 123.605 158.575 124.270 158.745 ;
        RECT 124.555 158.720 124.725 159.520 ;
        RECT 125.815 159.470 126.105 160.195 ;
        RECT 126.280 159.430 126.735 160.195 ;
        RECT 127.010 159.815 128.310 160.025 ;
        RECT 128.565 159.835 128.895 160.195 ;
        RECT 128.140 159.665 128.310 159.815 ;
        RECT 129.065 159.695 129.325 160.025 ;
        RECT 127.210 159.205 127.430 159.605 ;
        RECT 126.275 159.005 126.765 159.205 ;
        RECT 126.955 158.995 127.430 159.205 ;
        RECT 127.675 159.205 127.885 159.605 ;
        RECT 128.140 159.540 128.895 159.665 ;
        RECT 128.140 159.495 128.985 159.540 ;
        RECT 128.715 159.375 128.985 159.495 ;
        RECT 127.675 158.995 128.005 159.205 ;
        RECT 128.175 158.935 128.585 159.240 ;
        RECT 123.605 157.815 123.775 158.575 ;
        RECT 123.955 157.645 124.285 158.405 ;
        RECT 124.455 157.815 124.725 158.720 ;
        RECT 125.815 157.645 126.105 158.810 ;
        RECT 126.280 158.765 127.455 158.825 ;
        RECT 128.815 158.800 128.985 159.375 ;
        RECT 128.785 158.765 128.985 158.800 ;
        RECT 126.280 158.655 128.985 158.765 ;
        RECT 126.280 158.035 126.535 158.655 ;
        RECT 127.125 158.595 128.925 158.655 ;
        RECT 127.125 158.565 127.455 158.595 ;
        RECT 129.155 158.495 129.325 159.695 ;
        RECT 129.585 159.645 129.755 159.935 ;
        RECT 129.925 159.815 130.255 160.195 ;
        RECT 129.585 159.475 130.250 159.645 ;
        RECT 129.500 158.655 129.850 159.305 ;
        RECT 126.785 158.395 126.970 158.485 ;
        RECT 127.560 158.395 128.395 158.405 ;
        RECT 126.785 158.195 128.395 158.395 ;
        RECT 126.785 158.155 127.015 158.195 ;
        RECT 126.280 157.815 126.615 158.035 ;
        RECT 127.620 157.645 127.975 158.025 ;
        RECT 128.145 157.815 128.395 158.195 ;
        RECT 128.645 157.645 128.895 158.425 ;
        RECT 129.065 157.815 129.325 158.495 ;
        RECT 130.020 158.485 130.250 159.475 ;
        RECT 129.585 158.315 130.250 158.485 ;
        RECT 129.585 157.815 129.755 158.315 ;
        RECT 129.925 157.645 130.255 158.145 ;
        RECT 130.425 157.815 130.610 159.935 ;
        RECT 130.865 159.735 131.115 160.195 ;
        RECT 131.285 159.745 131.620 159.915 ;
        RECT 131.815 159.745 132.490 159.915 ;
        RECT 131.285 159.605 131.455 159.745 ;
        RECT 130.780 158.615 131.060 159.565 ;
        RECT 131.230 159.475 131.455 159.605 ;
        RECT 131.230 158.370 131.400 159.475 ;
        RECT 131.625 159.325 132.150 159.545 ;
        RECT 131.570 158.560 131.810 159.155 ;
        RECT 131.980 158.625 132.150 159.325 ;
        RECT 132.320 158.965 132.490 159.745 ;
        RECT 132.810 159.695 133.180 160.195 ;
        RECT 133.360 159.745 133.765 159.915 ;
        RECT 133.935 159.745 134.720 159.915 ;
        RECT 133.360 159.515 133.530 159.745 ;
        RECT 132.700 159.215 133.530 159.515 ;
        RECT 133.915 159.245 134.380 159.575 ;
        RECT 132.700 159.185 132.900 159.215 ;
        RECT 133.020 158.965 133.190 159.035 ;
        RECT 132.320 158.795 133.190 158.965 ;
        RECT 132.680 158.705 133.190 158.795 ;
        RECT 131.230 158.240 131.535 158.370 ;
        RECT 131.980 158.260 132.510 158.625 ;
        RECT 130.850 157.645 131.115 158.105 ;
        RECT 131.285 157.815 131.535 158.240 ;
        RECT 132.680 158.090 132.850 158.705 ;
        RECT 131.745 157.920 132.850 158.090 ;
        RECT 133.020 157.645 133.190 158.445 ;
        RECT 133.360 158.145 133.530 159.215 ;
        RECT 133.700 158.315 133.890 159.035 ;
        RECT 134.060 158.285 134.380 159.245 ;
        RECT 134.550 159.285 134.720 159.745 ;
        RECT 134.995 159.665 135.205 160.195 ;
        RECT 135.465 159.455 135.795 159.980 ;
        RECT 135.965 159.585 136.135 160.195 ;
        RECT 136.305 159.540 136.635 159.975 ;
        RECT 136.305 159.455 136.685 159.540 ;
        RECT 135.595 159.285 135.795 159.455 ;
        RECT 136.460 159.415 136.685 159.455 ;
        RECT 134.550 158.955 135.425 159.285 ;
        RECT 135.595 158.955 136.345 159.285 ;
        RECT 133.360 157.815 133.610 158.145 ;
        RECT 134.550 158.115 134.720 158.955 ;
        RECT 135.595 158.750 135.785 158.955 ;
        RECT 136.515 158.835 136.685 159.415 ;
        RECT 136.855 159.425 139.445 160.195 ;
        RECT 139.625 159.465 139.925 160.195 ;
        RECT 136.855 158.905 138.065 159.425 ;
        RECT 140.105 159.285 140.335 159.905 ;
        RECT 140.535 159.635 140.760 160.015 ;
        RECT 140.930 159.805 141.260 160.195 ;
        RECT 140.535 159.455 140.865 159.635 ;
        RECT 136.470 158.785 136.685 158.835 ;
        RECT 134.890 158.375 135.785 158.750 ;
        RECT 136.295 158.705 136.685 158.785 ;
        RECT 138.235 158.735 139.445 159.255 ;
        RECT 139.630 158.955 139.925 159.285 ;
        RECT 140.105 158.955 140.520 159.285 ;
        RECT 140.690 158.785 140.865 159.455 ;
        RECT 141.035 158.955 141.275 159.605 ;
        RECT 141.455 159.425 144.045 160.195 ;
        RECT 144.265 159.540 144.595 159.975 ;
        RECT 144.765 159.585 144.935 160.195 ;
        RECT 144.215 159.455 144.595 159.540 ;
        RECT 145.105 159.455 145.435 159.980 ;
        RECT 145.695 159.665 145.905 160.195 ;
        RECT 146.180 159.745 146.965 159.915 ;
        RECT 147.135 159.745 147.540 159.915 ;
        RECT 141.455 158.905 142.665 159.425 ;
        RECT 144.215 159.415 144.440 159.455 ;
        RECT 133.835 157.945 134.720 158.115 ;
        RECT 134.900 157.645 135.215 158.145 ;
        RECT 135.445 157.815 135.785 158.375 ;
        RECT 135.955 157.645 136.125 158.655 ;
        RECT 136.295 157.860 136.625 158.705 ;
        RECT 136.855 157.645 139.445 158.735 ;
        RECT 139.625 158.425 140.520 158.755 ;
        RECT 140.690 158.595 141.275 158.785 ;
        RECT 142.835 158.735 144.045 159.255 ;
        RECT 139.625 158.255 140.830 158.425 ;
        RECT 139.625 157.825 139.955 158.255 ;
        RECT 140.135 157.645 140.330 158.085 ;
        RECT 140.500 157.825 140.830 158.255 ;
        RECT 141.000 157.825 141.275 158.595 ;
        RECT 141.455 157.645 144.045 158.735 ;
        RECT 144.215 158.835 144.385 159.415 ;
        RECT 145.105 159.285 145.305 159.455 ;
        RECT 146.180 159.285 146.350 159.745 ;
        RECT 144.555 158.955 145.305 159.285 ;
        RECT 145.475 158.955 146.350 159.285 ;
        RECT 144.215 158.785 144.430 158.835 ;
        RECT 144.215 158.705 144.605 158.785 ;
        RECT 144.275 157.860 144.605 158.705 ;
        RECT 145.115 158.750 145.305 158.955 ;
        RECT 144.775 157.645 144.945 158.655 ;
        RECT 145.115 158.375 146.010 158.750 ;
        RECT 145.115 157.815 145.455 158.375 ;
        RECT 145.685 157.645 146.000 158.145 ;
        RECT 146.180 158.115 146.350 158.955 ;
        RECT 146.520 159.245 146.985 159.575 ;
        RECT 147.370 159.515 147.540 159.745 ;
        RECT 147.720 159.695 148.090 160.195 ;
        RECT 148.410 159.745 149.085 159.915 ;
        RECT 149.280 159.745 149.615 159.915 ;
        RECT 146.520 158.285 146.840 159.245 ;
        RECT 147.370 159.215 148.200 159.515 ;
        RECT 147.010 158.315 147.200 159.035 ;
        RECT 147.370 158.145 147.540 159.215 ;
        RECT 148.000 159.185 148.200 159.215 ;
        RECT 147.710 158.965 147.880 159.035 ;
        RECT 148.410 158.965 148.580 159.745 ;
        RECT 149.445 159.605 149.615 159.745 ;
        RECT 149.785 159.735 150.035 160.195 ;
        RECT 147.710 158.795 148.580 158.965 ;
        RECT 148.750 159.325 149.275 159.545 ;
        RECT 149.445 159.475 149.670 159.605 ;
        RECT 147.710 158.705 148.220 158.795 ;
        RECT 146.180 157.945 147.065 158.115 ;
        RECT 147.290 157.815 147.540 158.145 ;
        RECT 147.710 157.645 147.880 158.445 ;
        RECT 148.050 158.090 148.220 158.705 ;
        RECT 148.750 158.625 148.920 159.325 ;
        RECT 148.390 158.260 148.920 158.625 ;
        RECT 149.090 158.560 149.330 159.155 ;
        RECT 149.500 158.370 149.670 159.475 ;
        RECT 149.840 158.615 150.120 159.565 ;
        RECT 149.365 158.240 149.670 158.370 ;
        RECT 148.050 157.920 149.155 158.090 ;
        RECT 149.365 157.815 149.615 158.240 ;
        RECT 149.785 157.645 150.050 158.105 ;
        RECT 150.290 157.815 150.475 159.935 ;
        RECT 150.645 159.815 150.975 160.195 ;
        RECT 151.145 159.645 151.315 159.935 ;
        RECT 150.650 159.475 151.315 159.645 ;
        RECT 150.650 158.485 150.880 159.475 ;
        RECT 151.575 159.470 151.865 160.195 ;
        RECT 152.070 159.455 152.685 160.025 ;
        RECT 152.855 159.685 153.070 160.195 ;
        RECT 153.300 159.685 153.580 160.015 ;
        RECT 153.760 159.685 154.000 160.195 ;
        RECT 151.050 158.655 151.400 159.305 ;
        RECT 150.650 158.315 151.315 158.485 ;
        RECT 150.645 157.645 150.975 158.145 ;
        RECT 151.145 157.815 151.315 158.315 ;
        RECT 151.575 157.645 151.865 158.810 ;
        RECT 152.070 158.435 152.385 159.455 ;
        RECT 152.555 158.785 152.725 159.285 ;
        RECT 152.975 158.955 153.240 159.515 ;
        RECT 153.410 158.785 153.580 159.685 ;
        RECT 153.750 158.955 154.105 159.515 ;
        RECT 154.335 159.395 154.645 160.195 ;
        RECT 154.850 159.395 155.545 160.025 ;
        RECT 155.715 159.445 156.925 160.195 ;
        RECT 154.345 158.955 154.680 159.225 ;
        RECT 154.850 158.795 155.020 159.395 ;
        RECT 155.190 158.955 155.525 159.205 ;
        RECT 152.555 158.615 153.980 158.785 ;
        RECT 152.070 157.815 152.605 158.435 ;
        RECT 152.775 157.645 153.105 158.445 ;
        RECT 153.590 158.440 153.980 158.615 ;
        RECT 154.335 157.645 154.615 158.785 ;
        RECT 154.785 157.815 155.115 158.795 ;
        RECT 155.285 157.645 155.545 158.785 ;
        RECT 155.715 158.735 156.235 159.275 ;
        RECT 156.405 158.905 156.925 159.445 ;
        RECT 155.715 157.645 156.925 158.735 ;
        RECT 22.690 157.475 157.010 157.645 ;
        RECT 22.775 156.385 23.985 157.475 ;
        RECT 24.245 156.805 24.415 157.305 ;
        RECT 24.585 156.975 24.915 157.475 ;
        RECT 24.245 156.635 24.910 156.805 ;
        RECT 22.775 155.675 23.295 156.215 ;
        RECT 23.465 155.845 23.985 156.385 ;
        RECT 24.160 155.815 24.510 156.465 ;
        RECT 22.775 154.925 23.985 155.675 ;
        RECT 24.680 155.645 24.910 156.635 ;
        RECT 24.245 155.475 24.910 155.645 ;
        RECT 24.245 155.185 24.415 155.475 ;
        RECT 24.585 154.925 24.915 155.305 ;
        RECT 25.085 155.185 25.270 157.305 ;
        RECT 25.510 157.015 25.775 157.475 ;
        RECT 25.945 156.880 26.195 157.305 ;
        RECT 26.405 157.030 27.510 157.200 ;
        RECT 25.890 156.750 26.195 156.880 ;
        RECT 25.440 155.555 25.720 156.505 ;
        RECT 25.890 155.645 26.060 156.750 ;
        RECT 26.230 155.965 26.470 156.560 ;
        RECT 26.640 156.495 27.170 156.860 ;
        RECT 26.640 155.795 26.810 156.495 ;
        RECT 27.340 156.415 27.510 157.030 ;
        RECT 27.680 156.675 27.850 157.475 ;
        RECT 28.020 156.975 28.270 157.305 ;
        RECT 28.495 157.005 29.380 157.175 ;
        RECT 27.340 156.325 27.850 156.415 ;
        RECT 25.890 155.515 26.115 155.645 ;
        RECT 26.285 155.575 26.810 155.795 ;
        RECT 26.980 156.155 27.850 156.325 ;
        RECT 25.525 154.925 25.775 155.385 ;
        RECT 25.945 155.375 26.115 155.515 ;
        RECT 26.980 155.375 27.150 156.155 ;
        RECT 27.680 156.085 27.850 156.155 ;
        RECT 27.360 155.905 27.560 155.935 ;
        RECT 28.020 155.905 28.190 156.975 ;
        RECT 28.360 156.085 28.550 156.805 ;
        RECT 27.360 155.605 28.190 155.905 ;
        RECT 28.720 155.875 29.040 156.835 ;
        RECT 25.945 155.205 26.280 155.375 ;
        RECT 26.475 155.205 27.150 155.375 ;
        RECT 27.470 154.925 27.840 155.425 ;
        RECT 28.020 155.375 28.190 155.605 ;
        RECT 28.575 155.545 29.040 155.875 ;
        RECT 29.210 156.165 29.380 157.005 ;
        RECT 29.560 156.975 29.875 157.475 ;
        RECT 30.105 156.745 30.445 157.305 ;
        RECT 29.550 156.370 30.445 156.745 ;
        RECT 30.615 156.465 30.785 157.475 ;
        RECT 30.255 156.165 30.445 156.370 ;
        RECT 30.955 156.415 31.285 157.260 ;
        RECT 32.435 156.965 32.695 157.475 ;
        RECT 30.955 156.335 31.345 156.415 ;
        RECT 31.130 156.285 31.345 156.335 ;
        RECT 29.210 155.835 30.085 156.165 ;
        RECT 30.255 155.835 31.005 156.165 ;
        RECT 29.210 155.375 29.380 155.835 ;
        RECT 30.255 155.665 30.455 155.835 ;
        RECT 31.175 155.705 31.345 156.285 ;
        RECT 32.435 155.915 32.775 156.795 ;
        RECT 32.945 156.085 33.115 157.305 ;
        RECT 33.355 156.970 33.970 157.475 ;
        RECT 33.355 156.435 33.605 156.800 ;
        RECT 33.775 156.795 33.970 156.970 ;
        RECT 34.140 156.965 34.615 157.305 ;
        RECT 34.785 156.930 35.000 157.475 ;
        RECT 33.775 156.605 34.105 156.795 ;
        RECT 34.325 156.435 35.040 156.730 ;
        RECT 35.210 156.605 35.485 157.305 ;
        RECT 33.355 156.265 35.145 156.435 ;
        RECT 32.945 155.835 33.740 156.085 ;
        RECT 32.945 155.745 33.195 155.835 ;
        RECT 31.120 155.665 31.345 155.705 ;
        RECT 28.020 155.205 28.425 155.375 ;
        RECT 28.595 155.205 29.380 155.375 ;
        RECT 29.655 154.925 29.865 155.455 ;
        RECT 30.125 155.140 30.455 155.665 ;
        RECT 30.965 155.580 31.345 155.665 ;
        RECT 30.625 154.925 30.795 155.535 ;
        RECT 30.965 155.145 31.295 155.580 ;
        RECT 32.435 154.925 32.695 155.745 ;
        RECT 32.865 155.325 33.195 155.745 ;
        RECT 33.910 155.410 34.165 156.265 ;
        RECT 33.375 155.145 34.165 155.410 ;
        RECT 34.335 155.565 34.745 156.085 ;
        RECT 34.915 155.835 35.145 156.265 ;
        RECT 35.315 155.575 35.485 156.605 ;
        RECT 35.655 156.310 35.945 157.475 ;
        RECT 36.115 156.920 36.720 157.475 ;
        RECT 36.895 156.965 37.375 157.305 ;
        RECT 37.545 156.930 37.800 157.475 ;
        RECT 36.115 156.820 36.730 156.920 ;
        RECT 36.545 156.795 36.730 156.820 ;
        RECT 36.115 156.200 36.375 156.650 ;
        RECT 36.545 156.550 36.875 156.795 ;
        RECT 37.045 156.475 37.800 156.725 ;
        RECT 37.970 156.605 38.245 157.305 ;
        RECT 38.505 156.805 38.675 157.305 ;
        RECT 38.845 156.975 39.175 157.475 ;
        RECT 38.505 156.635 39.170 156.805 ;
        RECT 37.030 156.440 37.800 156.475 ;
        RECT 37.015 156.430 37.800 156.440 ;
        RECT 37.010 156.415 37.905 156.430 ;
        RECT 36.990 156.400 37.905 156.415 ;
        RECT 36.970 156.390 37.905 156.400 ;
        RECT 36.945 156.380 37.905 156.390 ;
        RECT 36.875 156.350 37.905 156.380 ;
        RECT 36.855 156.320 37.905 156.350 ;
        RECT 36.835 156.290 37.905 156.320 ;
        RECT 36.805 156.265 37.905 156.290 ;
        RECT 36.770 156.230 37.905 156.265 ;
        RECT 36.740 156.225 37.905 156.230 ;
        RECT 36.740 156.220 37.130 156.225 ;
        RECT 36.740 156.210 37.105 156.220 ;
        RECT 36.740 156.205 37.090 156.210 ;
        RECT 36.740 156.200 37.075 156.205 ;
        RECT 36.115 156.195 37.075 156.200 ;
        RECT 36.115 156.185 37.065 156.195 ;
        RECT 36.115 156.180 37.055 156.185 ;
        RECT 36.115 156.170 37.045 156.180 ;
        RECT 36.115 156.160 37.040 156.170 ;
        RECT 36.115 156.155 37.035 156.160 ;
        RECT 36.115 156.140 37.025 156.155 ;
        RECT 36.115 156.125 37.020 156.140 ;
        RECT 36.115 156.100 37.010 156.125 ;
        RECT 36.115 156.030 37.005 156.100 ;
        RECT 34.335 155.145 34.535 155.565 ;
        RECT 34.725 154.925 35.055 155.385 ;
        RECT 35.225 155.095 35.485 155.575 ;
        RECT 35.655 154.925 35.945 155.650 ;
        RECT 36.115 155.475 36.665 155.860 ;
        RECT 36.835 155.305 37.005 156.030 ;
        RECT 36.115 155.135 37.005 155.305 ;
        RECT 37.175 155.630 37.505 156.055 ;
        RECT 37.675 155.830 37.905 156.225 ;
        RECT 37.175 155.145 37.395 155.630 ;
        RECT 38.075 155.575 38.245 156.605 ;
        RECT 38.420 155.815 38.770 156.465 ;
        RECT 38.940 155.645 39.170 156.635 ;
        RECT 37.565 154.925 37.815 155.465 ;
        RECT 37.985 155.095 38.245 155.575 ;
        RECT 38.505 155.475 39.170 155.645 ;
        RECT 38.505 155.185 38.675 155.475 ;
        RECT 38.845 154.925 39.175 155.305 ;
        RECT 39.345 155.185 39.530 157.305 ;
        RECT 39.770 157.015 40.035 157.475 ;
        RECT 40.205 156.880 40.455 157.305 ;
        RECT 40.665 157.030 41.770 157.200 ;
        RECT 40.150 156.750 40.455 156.880 ;
        RECT 39.700 155.555 39.980 156.505 ;
        RECT 40.150 155.645 40.320 156.750 ;
        RECT 40.490 155.965 40.730 156.560 ;
        RECT 40.900 156.495 41.430 156.860 ;
        RECT 40.900 155.795 41.070 156.495 ;
        RECT 41.600 156.415 41.770 157.030 ;
        RECT 41.940 156.675 42.110 157.475 ;
        RECT 42.280 156.975 42.530 157.305 ;
        RECT 42.755 157.005 43.640 157.175 ;
        RECT 41.600 156.325 42.110 156.415 ;
        RECT 40.150 155.515 40.375 155.645 ;
        RECT 40.545 155.575 41.070 155.795 ;
        RECT 41.240 156.155 42.110 156.325 ;
        RECT 39.785 154.925 40.035 155.385 ;
        RECT 40.205 155.375 40.375 155.515 ;
        RECT 41.240 155.375 41.410 156.155 ;
        RECT 41.940 156.085 42.110 156.155 ;
        RECT 41.620 155.905 41.820 155.935 ;
        RECT 42.280 155.905 42.450 156.975 ;
        RECT 42.620 156.085 42.810 156.805 ;
        RECT 41.620 155.605 42.450 155.905 ;
        RECT 42.980 155.875 43.300 156.835 ;
        RECT 40.205 155.205 40.540 155.375 ;
        RECT 40.735 155.205 41.410 155.375 ;
        RECT 41.730 154.925 42.100 155.425 ;
        RECT 42.280 155.375 42.450 155.605 ;
        RECT 42.835 155.545 43.300 155.875 ;
        RECT 43.470 156.165 43.640 157.005 ;
        RECT 43.820 156.975 44.135 157.475 ;
        RECT 44.365 156.745 44.705 157.305 ;
        RECT 43.810 156.370 44.705 156.745 ;
        RECT 44.875 156.465 45.045 157.475 ;
        RECT 44.515 156.165 44.705 156.370 ;
        RECT 45.215 156.415 45.545 157.260 ;
        RECT 45.215 156.335 45.605 156.415 ;
        RECT 46.235 156.335 46.515 157.475 ;
        RECT 45.390 156.285 45.605 156.335 ;
        RECT 46.685 156.325 47.015 157.305 ;
        RECT 47.185 156.335 47.445 157.475 ;
        RECT 47.705 156.805 47.875 157.305 ;
        RECT 48.045 156.975 48.375 157.475 ;
        RECT 47.705 156.635 48.370 156.805 ;
        RECT 43.470 155.835 44.345 156.165 ;
        RECT 44.515 155.835 45.265 156.165 ;
        RECT 43.470 155.375 43.640 155.835 ;
        RECT 44.515 155.665 44.715 155.835 ;
        RECT 45.435 155.705 45.605 156.285 ;
        RECT 46.245 155.895 46.580 156.165 ;
        RECT 46.750 155.775 46.920 156.325 ;
        RECT 47.090 155.915 47.425 156.165 ;
        RECT 47.620 155.815 47.970 156.465 ;
        RECT 46.750 155.725 46.925 155.775 ;
        RECT 45.380 155.665 45.605 155.705 ;
        RECT 42.280 155.205 42.685 155.375 ;
        RECT 42.855 155.205 43.640 155.375 ;
        RECT 43.915 154.925 44.125 155.455 ;
        RECT 44.385 155.140 44.715 155.665 ;
        RECT 45.225 155.580 45.605 155.665 ;
        RECT 44.885 154.925 45.055 155.535 ;
        RECT 45.225 155.145 45.555 155.580 ;
        RECT 46.235 154.925 46.545 155.725 ;
        RECT 46.750 155.095 47.445 155.725 ;
        RECT 48.140 155.645 48.370 156.635 ;
        RECT 47.705 155.475 48.370 155.645 ;
        RECT 47.705 155.185 47.875 155.475 ;
        RECT 48.045 154.925 48.375 155.305 ;
        RECT 48.545 155.185 48.730 157.305 ;
        RECT 48.970 157.015 49.235 157.475 ;
        RECT 49.405 156.880 49.655 157.305 ;
        RECT 49.865 157.030 50.970 157.200 ;
        RECT 49.350 156.750 49.655 156.880 ;
        RECT 48.900 155.555 49.180 156.505 ;
        RECT 49.350 155.645 49.520 156.750 ;
        RECT 49.690 155.965 49.930 156.560 ;
        RECT 50.100 156.495 50.630 156.860 ;
        RECT 50.100 155.795 50.270 156.495 ;
        RECT 50.800 156.415 50.970 157.030 ;
        RECT 51.140 156.675 51.310 157.475 ;
        RECT 51.480 156.975 51.730 157.305 ;
        RECT 51.955 157.005 52.840 157.175 ;
        RECT 50.800 156.325 51.310 156.415 ;
        RECT 49.350 155.515 49.575 155.645 ;
        RECT 49.745 155.575 50.270 155.795 ;
        RECT 50.440 156.155 51.310 156.325 ;
        RECT 48.985 154.925 49.235 155.385 ;
        RECT 49.405 155.375 49.575 155.515 ;
        RECT 50.440 155.375 50.610 156.155 ;
        RECT 51.140 156.085 51.310 156.155 ;
        RECT 50.820 155.905 51.020 155.935 ;
        RECT 51.480 155.905 51.650 156.975 ;
        RECT 51.820 156.085 52.010 156.805 ;
        RECT 50.820 155.605 51.650 155.905 ;
        RECT 52.180 155.875 52.500 156.835 ;
        RECT 49.405 155.205 49.740 155.375 ;
        RECT 49.935 155.205 50.610 155.375 ;
        RECT 50.930 154.925 51.300 155.425 ;
        RECT 51.480 155.375 51.650 155.605 ;
        RECT 52.035 155.545 52.500 155.875 ;
        RECT 52.670 156.165 52.840 157.005 ;
        RECT 53.020 156.975 53.335 157.475 ;
        RECT 53.565 156.745 53.905 157.305 ;
        RECT 53.010 156.370 53.905 156.745 ;
        RECT 54.075 156.465 54.245 157.475 ;
        RECT 53.715 156.165 53.905 156.370 ;
        RECT 54.415 156.415 54.745 157.260 ;
        RECT 54.915 156.560 55.085 157.475 ;
        RECT 54.415 156.335 54.805 156.415 ;
        RECT 55.435 156.385 56.645 157.475 ;
        RECT 54.590 156.285 54.805 156.335 ;
        RECT 52.670 155.835 53.545 156.165 ;
        RECT 53.715 155.835 54.465 156.165 ;
        RECT 52.670 155.375 52.840 155.835 ;
        RECT 53.715 155.665 53.915 155.835 ;
        RECT 54.635 155.705 54.805 156.285 ;
        RECT 54.580 155.665 54.805 155.705 ;
        RECT 51.480 155.205 51.885 155.375 ;
        RECT 52.055 155.205 52.840 155.375 ;
        RECT 53.115 154.925 53.325 155.455 ;
        RECT 53.585 155.140 53.915 155.665 ;
        RECT 54.425 155.580 54.805 155.665 ;
        RECT 55.435 155.675 55.955 156.215 ;
        RECT 56.125 155.845 56.645 156.385 ;
        RECT 56.815 156.335 57.085 157.305 ;
        RECT 57.295 156.675 57.575 157.475 ;
        RECT 57.755 156.925 58.950 157.255 ;
        RECT 58.080 156.505 58.500 156.755 ;
        RECT 57.255 156.335 58.500 156.505 ;
        RECT 54.085 154.925 54.255 155.535 ;
        RECT 54.425 155.145 54.755 155.580 ;
        RECT 54.925 154.925 55.095 155.440 ;
        RECT 55.435 154.925 56.645 155.675 ;
        RECT 56.815 155.600 56.985 156.335 ;
        RECT 57.255 156.165 57.425 156.335 ;
        RECT 58.725 156.165 58.895 156.725 ;
        RECT 59.145 156.335 59.400 157.475 ;
        RECT 59.575 156.385 61.245 157.475 ;
        RECT 57.195 155.835 57.425 156.165 ;
        RECT 58.155 155.835 58.895 156.165 ;
        RECT 59.065 155.915 59.400 156.165 ;
        RECT 57.255 155.665 57.425 155.835 ;
        RECT 58.645 155.745 58.895 155.835 ;
        RECT 56.815 155.255 57.085 155.600 ;
        RECT 57.255 155.495 57.995 155.665 ;
        RECT 58.645 155.575 59.380 155.745 ;
        RECT 57.275 154.925 57.655 155.325 ;
        RECT 57.825 155.145 57.995 155.495 ;
        RECT 58.165 154.925 58.900 155.405 ;
        RECT 59.070 155.105 59.380 155.575 ;
        RECT 59.575 155.695 60.325 156.215 ;
        RECT 60.495 155.865 61.245 156.385 ;
        RECT 61.415 156.310 61.705 157.475 ;
        RECT 61.990 156.845 62.275 157.305 ;
        RECT 62.445 157.015 62.715 157.475 ;
        RECT 61.990 156.625 62.945 156.845 ;
        RECT 61.875 155.895 62.565 156.455 ;
        RECT 62.735 155.725 62.945 156.625 ;
        RECT 59.575 154.925 61.245 155.695 ;
        RECT 61.415 154.925 61.705 155.650 ;
        RECT 61.990 155.555 62.945 155.725 ;
        RECT 63.115 156.455 63.515 157.305 ;
        RECT 63.705 156.845 63.985 157.305 ;
        RECT 64.505 157.015 64.830 157.475 ;
        RECT 63.705 156.625 64.830 156.845 ;
        RECT 63.115 155.895 64.210 156.455 ;
        RECT 64.380 156.165 64.830 156.625 ;
        RECT 65.000 156.335 65.385 157.305 ;
        RECT 65.555 156.385 66.765 157.475 ;
        RECT 67.050 156.845 67.335 157.305 ;
        RECT 67.505 157.015 67.775 157.475 ;
        RECT 67.050 156.625 68.005 156.845 ;
        RECT 61.990 155.095 62.275 155.555 ;
        RECT 62.445 154.925 62.715 155.385 ;
        RECT 63.115 155.095 63.515 155.895 ;
        RECT 64.380 155.835 64.935 156.165 ;
        RECT 64.380 155.725 64.830 155.835 ;
        RECT 63.705 155.555 64.830 155.725 ;
        RECT 65.105 155.665 65.385 156.335 ;
        RECT 63.705 155.095 63.985 155.555 ;
        RECT 64.505 154.925 64.830 155.385 ;
        RECT 65.000 155.095 65.385 155.665 ;
        RECT 65.555 155.675 66.075 156.215 ;
        RECT 66.245 155.845 66.765 156.385 ;
        RECT 66.935 155.895 67.625 156.455 ;
        RECT 67.795 155.725 68.005 156.625 ;
        RECT 65.555 154.925 66.765 155.675 ;
        RECT 67.050 155.555 68.005 155.725 ;
        RECT 68.175 156.455 68.575 157.305 ;
        RECT 68.765 156.845 69.045 157.305 ;
        RECT 69.565 157.015 69.890 157.475 ;
        RECT 68.765 156.625 69.890 156.845 ;
        RECT 68.175 155.895 69.270 156.455 ;
        RECT 69.440 156.165 69.890 156.625 ;
        RECT 70.060 156.335 70.445 157.305 ;
        RECT 71.625 156.805 71.795 157.305 ;
        RECT 71.965 156.975 72.295 157.475 ;
        RECT 71.625 156.635 72.290 156.805 ;
        RECT 67.050 155.095 67.335 155.555 ;
        RECT 67.505 154.925 67.775 155.385 ;
        RECT 68.175 155.095 68.575 155.895 ;
        RECT 69.440 155.835 69.995 156.165 ;
        RECT 69.440 155.725 69.890 155.835 ;
        RECT 68.765 155.555 69.890 155.725 ;
        RECT 70.165 155.665 70.445 156.335 ;
        RECT 71.540 155.815 71.890 156.465 ;
        RECT 68.765 155.095 69.045 155.555 ;
        RECT 69.565 154.925 69.890 155.385 ;
        RECT 70.060 155.095 70.445 155.665 ;
        RECT 72.060 155.645 72.290 156.635 ;
        RECT 71.625 155.475 72.290 155.645 ;
        RECT 71.625 155.185 71.795 155.475 ;
        RECT 71.965 154.925 72.295 155.305 ;
        RECT 72.465 155.185 72.650 157.305 ;
        RECT 72.890 157.015 73.155 157.475 ;
        RECT 73.325 156.880 73.575 157.305 ;
        RECT 73.785 157.030 74.890 157.200 ;
        RECT 73.270 156.750 73.575 156.880 ;
        RECT 72.820 155.555 73.100 156.505 ;
        RECT 73.270 155.645 73.440 156.750 ;
        RECT 73.610 155.965 73.850 156.560 ;
        RECT 74.020 156.495 74.550 156.860 ;
        RECT 74.020 155.795 74.190 156.495 ;
        RECT 74.720 156.415 74.890 157.030 ;
        RECT 75.060 156.675 75.230 157.475 ;
        RECT 75.400 156.975 75.650 157.305 ;
        RECT 75.875 157.005 76.760 157.175 ;
        RECT 74.720 156.325 75.230 156.415 ;
        RECT 73.270 155.515 73.495 155.645 ;
        RECT 73.665 155.575 74.190 155.795 ;
        RECT 74.360 156.155 75.230 156.325 ;
        RECT 72.905 154.925 73.155 155.385 ;
        RECT 73.325 155.375 73.495 155.515 ;
        RECT 74.360 155.375 74.530 156.155 ;
        RECT 75.060 156.085 75.230 156.155 ;
        RECT 74.740 155.905 74.940 155.935 ;
        RECT 75.400 155.905 75.570 156.975 ;
        RECT 75.740 156.085 75.930 156.805 ;
        RECT 74.740 155.605 75.570 155.905 ;
        RECT 76.100 155.875 76.420 156.835 ;
        RECT 73.325 155.205 73.660 155.375 ;
        RECT 73.855 155.205 74.530 155.375 ;
        RECT 74.850 154.925 75.220 155.425 ;
        RECT 75.400 155.375 75.570 155.605 ;
        RECT 75.955 155.545 76.420 155.875 ;
        RECT 76.590 156.165 76.760 157.005 ;
        RECT 76.940 156.975 77.255 157.475 ;
        RECT 77.485 156.745 77.825 157.305 ;
        RECT 76.930 156.370 77.825 156.745 ;
        RECT 77.995 156.465 78.165 157.475 ;
        RECT 77.635 156.165 77.825 156.370 ;
        RECT 78.335 156.415 78.665 157.260 ;
        RECT 78.985 156.805 79.155 157.305 ;
        RECT 79.325 156.975 79.655 157.475 ;
        RECT 78.985 156.635 79.650 156.805 ;
        RECT 78.335 156.335 78.725 156.415 ;
        RECT 78.510 156.285 78.725 156.335 ;
        RECT 76.590 155.835 77.465 156.165 ;
        RECT 77.635 155.835 78.385 156.165 ;
        RECT 76.590 155.375 76.760 155.835 ;
        RECT 77.635 155.665 77.835 155.835 ;
        RECT 78.555 155.705 78.725 156.285 ;
        RECT 78.900 155.815 79.250 156.465 ;
        RECT 78.500 155.665 78.725 155.705 ;
        RECT 75.400 155.205 75.805 155.375 ;
        RECT 75.975 155.205 76.760 155.375 ;
        RECT 77.035 154.925 77.245 155.455 ;
        RECT 77.505 155.140 77.835 155.665 ;
        RECT 78.345 155.580 78.725 155.665 ;
        RECT 79.420 155.645 79.650 156.635 ;
        RECT 78.005 154.925 78.175 155.535 ;
        RECT 78.345 155.145 78.675 155.580 ;
        RECT 78.985 155.475 79.650 155.645 ;
        RECT 78.985 155.185 79.155 155.475 ;
        RECT 79.325 154.925 79.655 155.305 ;
        RECT 79.825 155.185 80.010 157.305 ;
        RECT 80.250 157.015 80.515 157.475 ;
        RECT 80.685 156.880 80.935 157.305 ;
        RECT 81.145 157.030 82.250 157.200 ;
        RECT 80.630 156.750 80.935 156.880 ;
        RECT 80.180 155.555 80.460 156.505 ;
        RECT 80.630 155.645 80.800 156.750 ;
        RECT 80.970 155.965 81.210 156.560 ;
        RECT 81.380 156.495 81.910 156.860 ;
        RECT 81.380 155.795 81.550 156.495 ;
        RECT 82.080 156.415 82.250 157.030 ;
        RECT 82.420 156.675 82.590 157.475 ;
        RECT 82.760 156.975 83.010 157.305 ;
        RECT 83.235 157.005 84.120 157.175 ;
        RECT 82.080 156.325 82.590 156.415 ;
        RECT 80.630 155.515 80.855 155.645 ;
        RECT 81.025 155.575 81.550 155.795 ;
        RECT 81.720 156.155 82.590 156.325 ;
        RECT 80.265 154.925 80.515 155.385 ;
        RECT 80.685 155.375 80.855 155.515 ;
        RECT 81.720 155.375 81.890 156.155 ;
        RECT 82.420 156.085 82.590 156.155 ;
        RECT 82.100 155.905 82.300 155.935 ;
        RECT 82.760 155.905 82.930 156.975 ;
        RECT 83.100 156.085 83.290 156.805 ;
        RECT 82.100 155.605 82.930 155.905 ;
        RECT 83.460 155.875 83.780 156.835 ;
        RECT 80.685 155.205 81.020 155.375 ;
        RECT 81.215 155.205 81.890 155.375 ;
        RECT 82.210 154.925 82.580 155.425 ;
        RECT 82.760 155.375 82.930 155.605 ;
        RECT 83.315 155.545 83.780 155.875 ;
        RECT 83.950 156.165 84.120 157.005 ;
        RECT 84.300 156.975 84.615 157.475 ;
        RECT 84.845 156.745 85.185 157.305 ;
        RECT 84.290 156.370 85.185 156.745 ;
        RECT 85.355 156.465 85.525 157.475 ;
        RECT 84.995 156.165 85.185 156.370 ;
        RECT 85.695 156.415 86.025 157.260 ;
        RECT 85.695 156.335 86.085 156.415 ;
        RECT 85.870 156.285 86.085 156.335 ;
        RECT 87.175 156.310 87.465 157.475 ;
        RECT 87.640 156.905 87.960 157.305 ;
        RECT 87.640 156.455 87.810 156.905 ;
        RECT 88.130 156.675 88.440 157.475 ;
        RECT 88.610 156.845 88.940 157.305 ;
        RECT 89.110 157.015 89.280 157.475 ;
        RECT 89.450 156.845 89.780 157.305 ;
        RECT 89.950 157.015 90.200 157.475 ;
        RECT 90.390 157.015 90.640 157.475 ;
        RECT 88.610 156.795 89.780 156.845 ;
        RECT 90.810 156.845 91.060 157.305 ;
        RECT 91.310 157.015 91.600 157.475 ;
        RECT 91.775 156.920 92.380 157.475 ;
        RECT 92.555 156.965 93.035 157.305 ;
        RECT 93.205 156.930 93.460 157.475 ;
        RECT 90.810 156.795 91.600 156.845 ;
        RECT 91.775 156.820 92.390 156.920 ;
        RECT 88.610 156.625 91.600 156.795 ;
        RECT 92.205 156.795 92.390 156.820 ;
        RECT 91.400 156.455 91.600 156.625 ;
        RECT 83.950 155.835 84.825 156.165 ;
        RECT 84.995 155.835 85.745 156.165 ;
        RECT 83.950 155.375 84.120 155.835 ;
        RECT 84.995 155.665 85.195 155.835 ;
        RECT 85.915 155.705 86.085 156.285 ;
        RECT 85.860 155.665 86.085 155.705 ;
        RECT 82.760 155.205 83.165 155.375 ;
        RECT 83.335 155.205 84.120 155.375 ;
        RECT 84.395 154.925 84.605 155.455 ;
        RECT 84.865 155.140 85.195 155.665 ;
        RECT 85.705 155.580 86.085 155.665 ;
        RECT 87.640 156.285 91.200 156.455 ;
        RECT 91.375 156.285 91.600 156.455 ;
        RECT 85.365 154.925 85.535 155.535 ;
        RECT 85.705 155.145 86.035 155.580 ;
        RECT 87.175 154.925 87.465 155.650 ;
        RECT 87.640 155.495 87.810 156.285 ;
        RECT 87.980 155.915 88.330 156.115 ;
        RECT 88.610 155.915 89.290 156.115 ;
        RECT 89.500 155.915 90.690 156.115 ;
        RECT 90.870 155.915 91.200 156.285 ;
        RECT 91.400 155.745 91.600 156.285 ;
        RECT 91.775 156.200 92.035 156.650 ;
        RECT 92.205 156.550 92.535 156.795 ;
        RECT 92.705 156.475 93.460 156.725 ;
        RECT 93.630 156.605 93.905 157.305 ;
        RECT 92.690 156.440 93.460 156.475 ;
        RECT 92.675 156.430 93.460 156.440 ;
        RECT 92.670 156.415 93.565 156.430 ;
        RECT 92.650 156.400 93.565 156.415 ;
        RECT 92.630 156.390 93.565 156.400 ;
        RECT 92.605 156.380 93.565 156.390 ;
        RECT 92.535 156.350 93.565 156.380 ;
        RECT 92.515 156.320 93.565 156.350 ;
        RECT 92.495 156.290 93.565 156.320 ;
        RECT 92.465 156.265 93.565 156.290 ;
        RECT 92.430 156.230 93.565 156.265 ;
        RECT 92.400 156.225 93.565 156.230 ;
        RECT 92.400 156.220 92.790 156.225 ;
        RECT 92.400 156.210 92.765 156.220 ;
        RECT 92.400 156.205 92.750 156.210 ;
        RECT 92.400 156.200 92.735 156.205 ;
        RECT 91.775 156.195 92.735 156.200 ;
        RECT 91.775 156.185 92.725 156.195 ;
        RECT 91.775 156.180 92.715 156.185 ;
        RECT 91.775 156.170 92.705 156.180 ;
        RECT 91.775 156.160 92.700 156.170 ;
        RECT 91.775 156.155 92.695 156.160 ;
        RECT 91.775 156.140 92.685 156.155 ;
        RECT 91.775 156.125 92.680 156.140 ;
        RECT 91.775 156.100 92.670 156.125 ;
        RECT 91.775 156.030 92.665 156.100 ;
        RECT 87.640 155.095 87.960 155.495 ;
        RECT 88.130 154.925 88.440 155.745 ;
        RECT 88.610 155.555 90.300 155.745 ;
        RECT 88.610 155.095 88.940 155.555 ;
        RECT 89.550 155.475 90.300 155.555 ;
        RECT 89.110 154.925 89.360 155.385 ;
        RECT 90.470 155.305 90.640 155.745 ;
        RECT 90.810 155.475 91.600 155.745 ;
        RECT 91.775 155.475 92.325 155.860 ;
        RECT 92.495 155.305 92.665 156.030 ;
        RECT 89.550 155.095 91.600 155.305 ;
        RECT 91.775 155.135 92.665 155.305 ;
        RECT 92.835 155.630 93.165 156.055 ;
        RECT 93.335 155.830 93.565 156.225 ;
        RECT 92.835 155.145 93.055 155.630 ;
        RECT 93.735 155.575 93.905 156.605 ;
        RECT 94.135 156.415 94.465 157.260 ;
        RECT 94.635 156.465 94.805 157.475 ;
        RECT 94.975 156.745 95.315 157.305 ;
        RECT 95.545 156.975 95.860 157.475 ;
        RECT 96.040 157.005 96.925 157.175 ;
        RECT 94.075 156.335 94.465 156.415 ;
        RECT 94.975 156.370 95.870 156.745 ;
        RECT 94.075 156.285 94.290 156.335 ;
        RECT 94.075 155.705 94.245 156.285 ;
        RECT 94.975 156.165 95.165 156.370 ;
        RECT 96.040 156.165 96.210 157.005 ;
        RECT 97.150 156.975 97.400 157.305 ;
        RECT 94.415 155.835 95.165 156.165 ;
        RECT 95.335 155.835 96.210 156.165 ;
        RECT 94.075 155.665 94.300 155.705 ;
        RECT 94.965 155.665 95.165 155.835 ;
        RECT 94.075 155.580 94.455 155.665 ;
        RECT 93.225 154.925 93.475 155.465 ;
        RECT 93.645 155.095 93.905 155.575 ;
        RECT 94.125 155.145 94.455 155.580 ;
        RECT 94.625 154.925 94.795 155.535 ;
        RECT 94.965 155.140 95.295 155.665 ;
        RECT 95.555 154.925 95.765 155.455 ;
        RECT 96.040 155.375 96.210 155.835 ;
        RECT 96.380 155.875 96.700 156.835 ;
        RECT 96.870 156.085 97.060 156.805 ;
        RECT 97.230 155.905 97.400 156.975 ;
        RECT 97.570 156.675 97.740 157.475 ;
        RECT 97.910 157.030 99.015 157.200 ;
        RECT 97.910 156.415 98.080 157.030 ;
        RECT 99.225 156.880 99.475 157.305 ;
        RECT 99.645 157.015 99.910 157.475 ;
        RECT 98.250 156.495 98.780 156.860 ;
        RECT 99.225 156.750 99.530 156.880 ;
        RECT 97.570 156.325 98.080 156.415 ;
        RECT 97.570 156.155 98.440 156.325 ;
        RECT 97.570 156.085 97.740 156.155 ;
        RECT 97.860 155.905 98.060 155.935 ;
        RECT 96.380 155.545 96.845 155.875 ;
        RECT 97.230 155.605 98.060 155.905 ;
        RECT 97.230 155.375 97.400 155.605 ;
        RECT 96.040 155.205 96.825 155.375 ;
        RECT 96.995 155.205 97.400 155.375 ;
        RECT 97.580 154.925 97.950 155.425 ;
        RECT 98.270 155.375 98.440 156.155 ;
        RECT 98.610 155.795 98.780 156.495 ;
        RECT 98.950 155.965 99.190 156.560 ;
        RECT 98.610 155.575 99.135 155.795 ;
        RECT 99.360 155.645 99.530 156.750 ;
        RECT 99.305 155.515 99.530 155.645 ;
        RECT 99.700 155.555 99.980 156.505 ;
        RECT 99.305 155.375 99.475 155.515 ;
        RECT 98.270 155.205 98.945 155.375 ;
        RECT 99.140 155.205 99.475 155.375 ;
        RECT 99.645 154.925 99.895 155.385 ;
        RECT 100.150 155.185 100.335 157.305 ;
        RECT 100.505 156.975 100.835 157.475 ;
        RECT 101.005 156.805 101.175 157.305 ;
        RECT 100.510 156.635 101.175 156.805 ;
        RECT 100.510 155.645 100.740 156.635 ;
        RECT 100.910 155.815 101.260 156.465 ;
        RECT 101.435 156.385 104.025 157.475 ;
        RECT 104.310 156.845 104.595 157.305 ;
        RECT 104.765 157.015 105.035 157.475 ;
        RECT 104.310 156.625 105.265 156.845 ;
        RECT 101.435 155.695 102.645 156.215 ;
        RECT 102.815 155.865 104.025 156.385 ;
        RECT 104.195 155.895 104.885 156.455 ;
        RECT 105.055 155.725 105.265 156.625 ;
        RECT 100.510 155.475 101.175 155.645 ;
        RECT 100.505 154.925 100.835 155.305 ;
        RECT 101.005 155.185 101.175 155.475 ;
        RECT 101.435 154.925 104.025 155.695 ;
        RECT 104.310 155.555 105.265 155.725 ;
        RECT 105.435 156.455 105.835 157.305 ;
        RECT 106.025 156.845 106.305 157.305 ;
        RECT 106.825 157.015 107.150 157.475 ;
        RECT 106.025 156.625 107.150 156.845 ;
        RECT 105.435 155.895 106.530 156.455 ;
        RECT 106.700 156.165 107.150 156.625 ;
        RECT 107.320 156.335 107.705 157.305 ;
        RECT 104.310 155.095 104.595 155.555 ;
        RECT 104.765 154.925 105.035 155.385 ;
        RECT 105.435 155.095 105.835 155.895 ;
        RECT 106.700 155.835 107.255 156.165 ;
        RECT 106.700 155.725 107.150 155.835 ;
        RECT 106.025 155.555 107.150 155.725 ;
        RECT 107.425 155.665 107.705 156.335 ;
        RECT 107.880 157.085 108.215 157.305 ;
        RECT 109.220 157.095 109.575 157.475 ;
        RECT 107.880 156.465 108.135 157.085 ;
        RECT 108.385 156.925 108.615 156.965 ;
        RECT 109.745 156.925 109.995 157.305 ;
        RECT 108.385 156.725 109.995 156.925 ;
        RECT 108.385 156.635 108.570 156.725 ;
        RECT 109.160 156.715 109.995 156.725 ;
        RECT 110.245 156.695 110.495 157.475 ;
        RECT 110.665 156.625 110.925 157.305 ;
        RECT 108.725 156.525 109.055 156.555 ;
        RECT 108.725 156.465 110.525 156.525 ;
        RECT 107.880 156.355 110.585 156.465 ;
        RECT 107.880 156.295 109.055 156.355 ;
        RECT 110.385 156.320 110.585 156.355 ;
        RECT 107.875 155.915 108.365 156.115 ;
        RECT 108.555 155.915 109.030 156.125 ;
        RECT 106.025 155.095 106.305 155.555 ;
        RECT 106.825 154.925 107.150 155.385 ;
        RECT 107.320 155.095 107.705 155.665 ;
        RECT 107.880 154.925 108.335 155.690 ;
        RECT 108.810 155.515 109.030 155.915 ;
        RECT 109.275 155.915 109.605 156.125 ;
        RECT 109.275 155.515 109.485 155.915 ;
        RECT 109.775 155.880 110.185 156.185 ;
        RECT 110.415 155.745 110.585 156.320 ;
        RECT 110.315 155.625 110.585 155.745 ;
        RECT 109.740 155.580 110.585 155.625 ;
        RECT 109.740 155.455 110.495 155.580 ;
        RECT 109.740 155.305 109.910 155.455 ;
        RECT 110.755 155.425 110.925 156.625 ;
        RECT 111.095 156.385 112.765 157.475 ;
        RECT 108.610 155.095 109.910 155.305 ;
        RECT 110.165 154.925 110.495 155.285 ;
        RECT 110.665 155.095 110.925 155.425 ;
        RECT 111.095 155.695 111.845 156.215 ;
        RECT 112.015 155.865 112.765 156.385 ;
        RECT 112.935 156.310 113.225 157.475 ;
        RECT 114.405 156.805 114.575 157.305 ;
        RECT 114.745 156.975 115.075 157.475 ;
        RECT 114.405 156.635 115.070 156.805 ;
        RECT 114.320 155.815 114.670 156.465 ;
        RECT 111.095 154.925 112.765 155.695 ;
        RECT 112.935 154.925 113.225 155.650 ;
        RECT 114.840 155.645 115.070 156.635 ;
        RECT 114.405 155.475 115.070 155.645 ;
        RECT 114.405 155.185 114.575 155.475 ;
        RECT 114.745 154.925 115.075 155.305 ;
        RECT 115.245 155.185 115.430 157.305 ;
        RECT 115.670 157.015 115.935 157.475 ;
        RECT 116.105 156.880 116.355 157.305 ;
        RECT 116.565 157.030 117.670 157.200 ;
        RECT 116.050 156.750 116.355 156.880 ;
        RECT 115.600 155.555 115.880 156.505 ;
        RECT 116.050 155.645 116.220 156.750 ;
        RECT 116.390 155.965 116.630 156.560 ;
        RECT 116.800 156.495 117.330 156.860 ;
        RECT 116.800 155.795 116.970 156.495 ;
        RECT 117.500 156.415 117.670 157.030 ;
        RECT 117.840 156.675 118.010 157.475 ;
        RECT 118.180 156.975 118.430 157.305 ;
        RECT 118.655 157.005 119.540 157.175 ;
        RECT 117.500 156.325 118.010 156.415 ;
        RECT 116.050 155.515 116.275 155.645 ;
        RECT 116.445 155.575 116.970 155.795 ;
        RECT 117.140 156.155 118.010 156.325 ;
        RECT 115.685 154.925 115.935 155.385 ;
        RECT 116.105 155.375 116.275 155.515 ;
        RECT 117.140 155.375 117.310 156.155 ;
        RECT 117.840 156.085 118.010 156.155 ;
        RECT 117.520 155.905 117.720 155.935 ;
        RECT 118.180 155.905 118.350 156.975 ;
        RECT 118.520 156.085 118.710 156.805 ;
        RECT 117.520 155.605 118.350 155.905 ;
        RECT 118.880 155.875 119.200 156.835 ;
        RECT 116.105 155.205 116.440 155.375 ;
        RECT 116.635 155.205 117.310 155.375 ;
        RECT 117.630 154.925 118.000 155.425 ;
        RECT 118.180 155.375 118.350 155.605 ;
        RECT 118.735 155.545 119.200 155.875 ;
        RECT 119.370 156.165 119.540 157.005 ;
        RECT 119.720 156.975 120.035 157.475 ;
        RECT 120.265 156.745 120.605 157.305 ;
        RECT 119.710 156.370 120.605 156.745 ;
        RECT 120.775 156.465 120.945 157.475 ;
        RECT 120.415 156.165 120.605 156.370 ;
        RECT 121.115 156.415 121.445 157.260 ;
        RECT 121.675 156.755 122.135 157.305 ;
        RECT 122.325 156.755 122.655 157.475 ;
        RECT 121.115 156.335 121.505 156.415 ;
        RECT 121.290 156.285 121.505 156.335 ;
        RECT 119.370 155.835 120.245 156.165 ;
        RECT 120.415 155.835 121.165 156.165 ;
        RECT 119.370 155.375 119.540 155.835 ;
        RECT 120.415 155.665 120.615 155.835 ;
        RECT 121.335 155.705 121.505 156.285 ;
        RECT 121.280 155.665 121.505 155.705 ;
        RECT 118.180 155.205 118.585 155.375 ;
        RECT 118.755 155.205 119.540 155.375 ;
        RECT 119.815 154.925 120.025 155.455 ;
        RECT 120.285 155.140 120.615 155.665 ;
        RECT 121.125 155.580 121.505 155.665 ;
        RECT 120.785 154.925 120.955 155.535 ;
        RECT 121.125 155.145 121.455 155.580 ;
        RECT 121.675 155.385 121.925 156.755 ;
        RECT 122.855 156.585 123.155 157.135 ;
        RECT 123.325 156.805 123.605 157.475 ;
        RECT 122.215 156.415 123.155 156.585 ;
        RECT 122.215 156.165 122.385 156.415 ;
        RECT 123.525 156.165 123.790 156.525 ;
        RECT 124.495 156.415 124.825 157.260 ;
        RECT 124.995 156.465 125.165 157.475 ;
        RECT 125.335 156.745 125.675 157.305 ;
        RECT 125.905 156.975 126.220 157.475 ;
        RECT 126.400 157.005 127.285 157.175 ;
        RECT 122.095 155.835 122.385 156.165 ;
        RECT 122.555 155.915 122.895 156.165 ;
        RECT 123.115 155.915 123.790 156.165 ;
        RECT 124.435 156.335 124.825 156.415 ;
        RECT 125.335 156.370 126.230 156.745 ;
        RECT 124.435 156.285 124.650 156.335 ;
        RECT 122.215 155.745 122.385 155.835 ;
        RECT 122.215 155.555 123.605 155.745 ;
        RECT 124.435 155.705 124.605 156.285 ;
        RECT 125.335 156.165 125.525 156.370 ;
        RECT 126.400 156.165 126.570 157.005 ;
        RECT 127.510 156.975 127.760 157.305 ;
        RECT 124.775 155.835 125.525 156.165 ;
        RECT 125.695 155.835 126.570 156.165 ;
        RECT 124.435 155.665 124.660 155.705 ;
        RECT 125.325 155.665 125.525 155.835 ;
        RECT 124.435 155.580 124.815 155.665 ;
        RECT 121.675 155.095 122.235 155.385 ;
        RECT 122.405 154.925 122.655 155.385 ;
        RECT 123.275 155.195 123.605 155.555 ;
        RECT 124.485 155.145 124.815 155.580 ;
        RECT 124.985 154.925 125.155 155.535 ;
        RECT 125.325 155.140 125.655 155.665 ;
        RECT 125.915 154.925 126.125 155.455 ;
        RECT 126.400 155.375 126.570 155.835 ;
        RECT 126.740 155.875 127.060 156.835 ;
        RECT 127.230 156.085 127.420 156.805 ;
        RECT 127.590 155.905 127.760 156.975 ;
        RECT 127.930 156.675 128.100 157.475 ;
        RECT 128.270 157.030 129.375 157.200 ;
        RECT 128.270 156.415 128.440 157.030 ;
        RECT 129.585 156.880 129.835 157.305 ;
        RECT 130.005 157.015 130.270 157.475 ;
        RECT 128.610 156.495 129.140 156.860 ;
        RECT 129.585 156.750 129.890 156.880 ;
        RECT 127.930 156.325 128.440 156.415 ;
        RECT 127.930 156.155 128.800 156.325 ;
        RECT 127.930 156.085 128.100 156.155 ;
        RECT 128.220 155.905 128.420 155.935 ;
        RECT 126.740 155.545 127.205 155.875 ;
        RECT 127.590 155.605 128.420 155.905 ;
        RECT 127.590 155.375 127.760 155.605 ;
        RECT 126.400 155.205 127.185 155.375 ;
        RECT 127.355 155.205 127.760 155.375 ;
        RECT 127.940 154.925 128.310 155.425 ;
        RECT 128.630 155.375 128.800 156.155 ;
        RECT 128.970 155.795 129.140 156.495 ;
        RECT 129.310 155.965 129.550 156.560 ;
        RECT 128.970 155.575 129.495 155.795 ;
        RECT 129.720 155.645 129.890 156.750 ;
        RECT 129.665 155.515 129.890 155.645 ;
        RECT 130.060 155.555 130.340 156.505 ;
        RECT 129.665 155.375 129.835 155.515 ;
        RECT 128.630 155.205 129.305 155.375 ;
        RECT 129.500 155.205 129.835 155.375 ;
        RECT 130.005 154.925 130.255 155.385 ;
        RECT 130.510 155.185 130.695 157.305 ;
        RECT 130.865 156.975 131.195 157.475 ;
        RECT 131.365 156.805 131.535 157.305 ;
        RECT 131.795 157.040 137.140 157.475 ;
        RECT 130.870 156.635 131.535 156.805 ;
        RECT 130.870 155.645 131.100 156.635 ;
        RECT 131.270 155.815 131.620 156.465 ;
        RECT 130.870 155.475 131.535 155.645 ;
        RECT 130.865 154.925 131.195 155.305 ;
        RECT 131.365 155.185 131.535 155.475 ;
        RECT 133.380 155.470 133.720 156.300 ;
        RECT 135.200 155.790 135.550 157.040 ;
        RECT 137.315 156.400 137.585 157.305 ;
        RECT 137.755 156.715 138.085 157.475 ;
        RECT 138.265 156.545 138.435 157.305 ;
        RECT 137.315 155.600 137.485 156.400 ;
        RECT 137.770 156.375 138.435 156.545 ;
        RECT 137.770 156.230 137.940 156.375 ;
        RECT 138.695 156.310 138.985 157.475 ;
        RECT 139.155 157.040 144.500 157.475 ;
        RECT 137.655 155.900 137.940 156.230 ;
        RECT 137.770 155.645 137.940 155.900 ;
        RECT 138.175 155.825 138.505 156.195 ;
        RECT 131.795 154.925 137.140 155.470 ;
        RECT 137.315 155.095 137.575 155.600 ;
        RECT 137.770 155.475 138.435 155.645 ;
        RECT 137.755 154.925 138.085 155.305 ;
        RECT 138.265 155.095 138.435 155.475 ;
        RECT 138.695 154.925 138.985 155.650 ;
        RECT 140.740 155.470 141.080 156.300 ;
        RECT 142.560 155.790 142.910 157.040 ;
        RECT 144.675 156.385 148.185 157.475 ;
        RECT 148.445 156.805 148.615 157.305 ;
        RECT 148.785 156.975 149.115 157.475 ;
        RECT 148.445 156.635 149.110 156.805 ;
        RECT 144.675 155.695 146.325 156.215 ;
        RECT 146.495 155.865 148.185 156.385 ;
        RECT 148.360 155.815 148.710 156.465 ;
        RECT 139.155 154.925 144.500 155.470 ;
        RECT 144.675 154.925 148.185 155.695 ;
        RECT 148.880 155.645 149.110 156.635 ;
        RECT 148.445 155.475 149.110 155.645 ;
        RECT 148.445 155.185 148.615 155.475 ;
        RECT 148.785 154.925 149.115 155.305 ;
        RECT 149.285 155.185 149.470 157.305 ;
        RECT 149.710 157.015 149.975 157.475 ;
        RECT 150.145 156.880 150.395 157.305 ;
        RECT 150.605 157.030 151.710 157.200 ;
        RECT 150.090 156.750 150.395 156.880 ;
        RECT 149.640 155.555 149.920 156.505 ;
        RECT 150.090 155.645 150.260 156.750 ;
        RECT 150.430 155.965 150.670 156.560 ;
        RECT 150.840 156.495 151.370 156.860 ;
        RECT 150.840 155.795 151.010 156.495 ;
        RECT 151.540 156.415 151.710 157.030 ;
        RECT 151.880 156.675 152.050 157.475 ;
        RECT 152.220 156.975 152.470 157.305 ;
        RECT 152.695 157.005 153.580 157.175 ;
        RECT 151.540 156.325 152.050 156.415 ;
        RECT 150.090 155.515 150.315 155.645 ;
        RECT 150.485 155.575 151.010 155.795 ;
        RECT 151.180 156.155 152.050 156.325 ;
        RECT 149.725 154.925 149.975 155.385 ;
        RECT 150.145 155.375 150.315 155.515 ;
        RECT 151.180 155.375 151.350 156.155 ;
        RECT 151.880 156.085 152.050 156.155 ;
        RECT 151.560 155.905 151.760 155.935 ;
        RECT 152.220 155.905 152.390 156.975 ;
        RECT 152.560 156.085 152.750 156.805 ;
        RECT 151.560 155.605 152.390 155.905 ;
        RECT 152.920 155.875 153.240 156.835 ;
        RECT 150.145 155.205 150.480 155.375 ;
        RECT 150.675 155.205 151.350 155.375 ;
        RECT 151.670 154.925 152.040 155.425 ;
        RECT 152.220 155.375 152.390 155.605 ;
        RECT 152.775 155.545 153.240 155.875 ;
        RECT 153.410 156.165 153.580 157.005 ;
        RECT 153.760 156.975 154.075 157.475 ;
        RECT 154.305 156.745 154.645 157.305 ;
        RECT 153.750 156.370 154.645 156.745 ;
        RECT 154.815 156.465 154.985 157.475 ;
        RECT 154.455 156.165 154.645 156.370 ;
        RECT 155.155 156.415 155.485 157.260 ;
        RECT 155.155 156.335 155.545 156.415 ;
        RECT 155.330 156.285 155.545 156.335 ;
        RECT 153.410 155.835 154.285 156.165 ;
        RECT 154.455 155.835 155.205 156.165 ;
        RECT 153.410 155.375 153.580 155.835 ;
        RECT 154.455 155.665 154.655 155.835 ;
        RECT 155.375 155.705 155.545 156.285 ;
        RECT 155.715 156.385 156.925 157.475 ;
        RECT 155.715 155.845 156.235 156.385 ;
        RECT 155.320 155.665 155.545 155.705 ;
        RECT 156.405 155.675 156.925 156.215 ;
        RECT 152.220 155.205 152.625 155.375 ;
        RECT 152.795 155.205 153.580 155.375 ;
        RECT 153.855 154.925 154.065 155.455 ;
        RECT 154.325 155.140 154.655 155.665 ;
        RECT 155.165 155.580 155.545 155.665 ;
        RECT 154.825 154.925 154.995 155.535 ;
        RECT 155.165 155.145 155.495 155.580 ;
        RECT 155.715 154.925 156.925 155.675 ;
        RECT 22.690 154.755 157.010 154.925 ;
        RECT 22.775 154.005 23.985 154.755 ;
        RECT 22.775 153.465 23.295 154.005 ;
        RECT 24.155 153.985 25.825 154.755 ;
        RECT 25.995 154.080 26.255 154.585 ;
        RECT 26.435 154.375 26.765 154.755 ;
        RECT 26.945 154.205 27.115 154.585 ;
        RECT 27.375 154.210 32.720 154.755 ;
        RECT 32.895 154.210 38.240 154.755 ;
        RECT 23.465 153.295 23.985 153.835 ;
        RECT 24.155 153.465 24.905 153.985 ;
        RECT 25.075 153.295 25.825 153.815 ;
        RECT 22.775 152.205 23.985 153.295 ;
        RECT 24.155 152.205 25.825 153.295 ;
        RECT 25.995 153.280 26.165 154.080 ;
        RECT 26.450 154.035 27.115 154.205 ;
        RECT 26.450 153.780 26.620 154.035 ;
        RECT 26.335 153.450 26.620 153.780 ;
        RECT 26.855 153.485 27.185 153.855 ;
        RECT 26.450 153.305 26.620 153.450 ;
        RECT 28.960 153.380 29.300 154.210 ;
        RECT 25.995 152.375 26.265 153.280 ;
        RECT 26.450 153.135 27.115 153.305 ;
        RECT 26.435 152.205 26.765 152.965 ;
        RECT 26.945 152.375 27.115 153.135 ;
        RECT 30.780 152.640 31.130 153.890 ;
        RECT 34.480 153.380 34.820 154.210 ;
        RECT 39.335 154.080 39.595 154.585 ;
        RECT 39.775 154.375 40.105 154.755 ;
        RECT 40.285 154.205 40.455 154.585 ;
        RECT 36.300 152.640 36.650 153.890 ;
        RECT 39.335 153.280 39.505 154.080 ;
        RECT 39.790 154.035 40.455 154.205 ;
        RECT 40.715 154.105 40.975 154.585 ;
        RECT 41.145 154.215 41.395 154.755 ;
        RECT 39.790 153.780 39.960 154.035 ;
        RECT 39.675 153.450 39.960 153.780 ;
        RECT 40.195 153.485 40.525 153.855 ;
        RECT 39.790 153.305 39.960 153.450 ;
        RECT 27.375 152.205 32.720 152.640 ;
        RECT 32.895 152.205 38.240 152.640 ;
        RECT 39.335 152.375 39.605 153.280 ;
        RECT 39.790 153.135 40.455 153.305 ;
        RECT 39.775 152.205 40.105 152.965 ;
        RECT 40.285 152.375 40.455 153.135 ;
        RECT 40.715 153.075 40.885 154.105 ;
        RECT 41.565 154.050 41.785 154.535 ;
        RECT 41.055 153.455 41.285 153.850 ;
        RECT 41.455 153.625 41.785 154.050 ;
        RECT 41.955 154.375 42.845 154.545 ;
        RECT 41.955 153.650 42.125 154.375 ;
        RECT 42.295 153.820 42.845 154.205 ;
        RECT 43.935 154.015 44.400 154.560 ;
        RECT 41.955 153.580 42.845 153.650 ;
        RECT 41.950 153.555 42.845 153.580 ;
        RECT 41.940 153.540 42.845 153.555 ;
        RECT 41.935 153.525 42.845 153.540 ;
        RECT 41.925 153.520 42.845 153.525 ;
        RECT 41.920 153.510 42.845 153.520 ;
        RECT 41.915 153.500 42.845 153.510 ;
        RECT 41.905 153.495 42.845 153.500 ;
        RECT 41.895 153.485 42.845 153.495 ;
        RECT 41.885 153.480 42.845 153.485 ;
        RECT 41.885 153.475 42.220 153.480 ;
        RECT 41.870 153.470 42.220 153.475 ;
        RECT 41.855 153.460 42.220 153.470 ;
        RECT 41.830 153.455 42.220 153.460 ;
        RECT 41.055 153.450 42.220 153.455 ;
        RECT 41.055 153.415 42.190 153.450 ;
        RECT 41.055 153.390 42.155 153.415 ;
        RECT 41.055 153.360 42.125 153.390 ;
        RECT 41.055 153.330 42.105 153.360 ;
        RECT 41.055 153.300 42.085 153.330 ;
        RECT 41.055 153.290 42.015 153.300 ;
        RECT 41.055 153.280 41.990 153.290 ;
        RECT 41.055 153.265 41.970 153.280 ;
        RECT 41.055 153.250 41.950 153.265 ;
        RECT 41.160 153.240 41.945 153.250 ;
        RECT 41.160 153.205 41.930 153.240 ;
        RECT 40.715 152.375 40.990 153.075 ;
        RECT 41.160 152.955 41.915 153.205 ;
        RECT 42.085 152.885 42.415 153.130 ;
        RECT 42.585 153.030 42.845 153.480 ;
        RECT 43.935 153.055 44.105 154.015 ;
        RECT 44.905 153.935 45.075 154.755 ;
        RECT 45.245 154.105 45.575 154.585 ;
        RECT 45.745 154.365 46.095 154.755 ;
        RECT 46.265 154.185 46.495 154.585 ;
        RECT 45.985 154.105 46.495 154.185 ;
        RECT 45.245 154.015 46.495 154.105 ;
        RECT 46.665 154.015 46.985 154.495 ;
        RECT 45.245 153.935 46.155 154.015 ;
        RECT 44.275 153.395 44.520 153.845 ;
        RECT 44.780 153.565 45.475 153.765 ;
        RECT 45.645 153.595 46.245 153.765 ;
        RECT 45.645 153.395 45.815 153.595 ;
        RECT 46.475 153.425 46.645 153.845 ;
        RECT 44.275 153.225 45.815 153.395 ;
        RECT 45.985 153.255 46.645 153.425 ;
        RECT 45.985 153.055 46.155 153.255 ;
        RECT 46.815 153.085 46.985 154.015 ;
        RECT 47.155 154.005 48.365 154.755 ;
        RECT 48.535 154.030 48.825 154.755 ;
        RECT 49.455 154.015 49.920 154.560 ;
        RECT 47.155 153.465 47.675 154.005 ;
        RECT 47.845 153.295 48.365 153.835 ;
        RECT 43.935 152.885 46.155 153.055 ;
        RECT 46.325 152.885 46.985 153.085 ;
        RECT 42.230 152.860 42.415 152.885 ;
        RECT 42.230 152.760 42.845 152.860 ;
        RECT 41.160 152.205 41.415 152.750 ;
        RECT 41.585 152.375 42.065 152.715 ;
        RECT 42.240 152.205 42.845 152.760 ;
        RECT 43.935 152.205 44.235 152.715 ;
        RECT 44.405 152.375 44.735 152.885 ;
        RECT 46.325 152.715 46.495 152.885 ;
        RECT 44.905 152.205 45.535 152.715 ;
        RECT 46.115 152.545 46.495 152.715 ;
        RECT 46.665 152.205 46.965 152.715 ;
        RECT 47.155 152.205 48.365 153.295 ;
        RECT 48.535 152.205 48.825 153.370 ;
        RECT 49.455 153.055 49.625 154.015 ;
        RECT 50.425 153.935 50.595 154.755 ;
        RECT 50.765 154.105 51.095 154.585 ;
        RECT 51.265 154.365 51.615 154.755 ;
        RECT 51.785 154.185 52.015 154.585 ;
        RECT 51.505 154.105 52.015 154.185 ;
        RECT 50.765 154.015 52.015 154.105 ;
        RECT 52.185 154.015 52.505 154.495 ;
        RECT 50.765 153.935 51.675 154.015 ;
        RECT 49.795 153.395 50.040 153.845 ;
        RECT 50.300 153.565 50.995 153.765 ;
        RECT 51.165 153.595 51.765 153.765 ;
        RECT 51.165 153.395 51.335 153.595 ;
        RECT 51.995 153.425 52.165 153.845 ;
        RECT 49.795 153.225 51.335 153.395 ;
        RECT 51.505 153.255 52.165 153.425 ;
        RECT 51.505 153.055 51.675 153.255 ;
        RECT 52.335 153.085 52.505 154.015 ;
        RECT 52.675 153.985 54.345 154.755 ;
        RECT 54.515 154.015 54.900 154.585 ;
        RECT 55.070 154.295 55.395 154.755 ;
        RECT 55.915 154.125 56.195 154.585 ;
        RECT 52.675 153.465 53.425 153.985 ;
        RECT 53.595 153.295 54.345 153.815 ;
        RECT 49.455 152.885 51.675 153.055 ;
        RECT 51.845 152.885 52.505 153.085 ;
        RECT 49.455 152.205 49.755 152.715 ;
        RECT 49.925 152.375 50.255 152.885 ;
        RECT 51.845 152.715 52.015 152.885 ;
        RECT 50.425 152.205 51.055 152.715 ;
        RECT 51.635 152.545 52.015 152.715 ;
        RECT 52.185 152.205 52.485 152.715 ;
        RECT 52.675 152.205 54.345 153.295 ;
        RECT 54.515 153.345 54.795 154.015 ;
        RECT 55.070 153.955 56.195 154.125 ;
        RECT 55.070 153.845 55.520 153.955 ;
        RECT 54.965 153.515 55.520 153.845 ;
        RECT 56.385 153.785 56.785 154.585 ;
        RECT 57.185 154.295 57.455 154.755 ;
        RECT 57.625 154.125 57.910 154.585 ;
        RECT 54.515 152.375 54.900 153.345 ;
        RECT 55.070 153.055 55.520 153.515 ;
        RECT 55.690 153.225 56.785 153.785 ;
        RECT 55.070 152.835 56.195 153.055 ;
        RECT 55.070 152.205 55.395 152.665 ;
        RECT 55.915 152.375 56.195 152.835 ;
        RECT 56.385 152.375 56.785 153.225 ;
        RECT 56.955 153.955 57.910 154.125 ;
        RECT 58.195 154.080 58.465 154.425 ;
        RECT 58.655 154.355 59.035 154.755 ;
        RECT 59.205 154.185 59.375 154.535 ;
        RECT 59.545 154.275 60.280 154.755 ;
        RECT 56.955 153.055 57.165 153.955 ;
        RECT 57.335 153.225 58.025 153.785 ;
        RECT 58.195 153.345 58.365 154.080 ;
        RECT 58.635 154.015 59.375 154.185 ;
        RECT 60.450 154.105 60.760 154.575 ;
        RECT 58.635 153.845 58.805 154.015 ;
        RECT 60.025 153.935 60.760 154.105 ;
        RECT 60.955 153.985 62.625 154.755 ;
        RECT 63.260 153.990 63.715 154.755 ;
        RECT 63.990 154.375 65.290 154.585 ;
        RECT 65.545 154.395 65.875 154.755 ;
        RECT 65.120 154.225 65.290 154.375 ;
        RECT 66.045 154.255 66.305 154.585 ;
        RECT 66.075 154.245 66.305 154.255 ;
        RECT 60.025 153.845 60.275 153.935 ;
        RECT 58.575 153.515 58.805 153.845 ;
        RECT 59.535 153.515 60.275 153.845 ;
        RECT 60.445 153.515 60.780 153.765 ;
        RECT 58.635 153.345 58.805 153.515 ;
        RECT 56.955 152.835 57.910 153.055 ;
        RECT 57.185 152.205 57.455 152.665 ;
        RECT 57.625 152.375 57.910 152.835 ;
        RECT 58.195 152.375 58.465 153.345 ;
        RECT 58.635 153.175 59.880 153.345 ;
        RECT 58.675 152.205 58.955 153.005 ;
        RECT 59.460 152.925 59.880 153.175 ;
        RECT 60.105 152.955 60.275 153.515 ;
        RECT 60.955 153.465 61.705 153.985 ;
        RECT 59.135 152.425 60.330 152.755 ;
        RECT 60.525 152.205 60.780 153.345 ;
        RECT 61.875 153.295 62.625 153.815 ;
        RECT 64.190 153.765 64.410 154.165 ;
        RECT 63.255 153.565 63.745 153.765 ;
        RECT 63.935 153.555 64.410 153.765 ;
        RECT 64.655 153.765 64.865 154.165 ;
        RECT 65.120 154.100 65.875 154.225 ;
        RECT 65.120 154.055 65.965 154.100 ;
        RECT 65.695 153.935 65.965 154.055 ;
        RECT 64.655 153.555 64.985 153.765 ;
        RECT 65.155 153.495 65.565 153.800 ;
        RECT 60.955 152.205 62.625 153.295 ;
        RECT 63.260 153.325 64.435 153.385 ;
        RECT 65.795 153.360 65.965 153.935 ;
        RECT 65.765 153.325 65.965 153.360 ;
        RECT 63.260 153.215 65.965 153.325 ;
        RECT 63.260 152.595 63.515 153.215 ;
        RECT 64.105 153.155 65.905 153.215 ;
        RECT 64.105 153.125 64.435 153.155 ;
        RECT 66.135 153.055 66.305 154.245 ;
        RECT 63.765 152.955 63.950 153.045 ;
        RECT 64.540 152.955 65.375 152.965 ;
        RECT 63.765 152.755 65.375 152.955 ;
        RECT 63.765 152.715 63.995 152.755 ;
        RECT 63.260 152.375 63.595 152.595 ;
        RECT 64.600 152.205 64.955 152.585 ;
        RECT 65.125 152.375 65.375 152.755 ;
        RECT 65.625 152.205 65.875 152.985 ;
        RECT 66.045 152.375 66.305 153.055 ;
        RECT 66.475 154.255 66.735 154.585 ;
        RECT 66.905 154.395 67.235 154.755 ;
        RECT 67.490 154.375 68.790 154.585 ;
        RECT 66.475 154.245 66.705 154.255 ;
        RECT 66.475 153.055 66.645 154.245 ;
        RECT 67.490 154.225 67.660 154.375 ;
        RECT 66.905 154.100 67.660 154.225 ;
        RECT 66.815 154.055 67.660 154.100 ;
        RECT 66.815 153.935 67.085 154.055 ;
        RECT 66.815 153.360 66.985 153.935 ;
        RECT 67.215 153.495 67.625 153.800 ;
        RECT 67.915 153.765 68.125 154.165 ;
        RECT 67.795 153.555 68.125 153.765 ;
        RECT 68.370 153.765 68.590 154.165 ;
        RECT 69.065 153.990 69.520 154.755 ;
        RECT 69.700 154.250 70.035 154.755 ;
        RECT 70.205 154.185 70.445 154.560 ;
        RECT 70.725 154.425 70.895 154.570 ;
        RECT 70.725 154.230 71.100 154.425 ;
        RECT 71.460 154.260 71.855 154.755 ;
        RECT 68.370 153.555 68.845 153.765 ;
        RECT 69.035 153.565 69.525 153.765 ;
        RECT 66.815 153.325 67.015 153.360 ;
        RECT 68.345 153.325 69.520 153.385 ;
        RECT 66.815 153.215 69.520 153.325 ;
        RECT 69.755 153.225 70.055 154.075 ;
        RECT 70.225 154.035 70.445 154.185 ;
        RECT 70.225 153.705 70.760 154.035 ;
        RECT 70.930 153.895 71.100 154.230 ;
        RECT 72.025 154.065 72.265 154.585 ;
        RECT 66.875 153.155 68.675 153.215 ;
        RECT 68.345 153.125 68.675 153.155 ;
        RECT 66.475 152.375 66.735 153.055 ;
        RECT 66.905 152.205 67.155 152.985 ;
        RECT 67.405 152.955 68.240 152.965 ;
        RECT 68.830 152.955 69.015 153.045 ;
        RECT 67.405 152.755 69.015 152.955 ;
        RECT 67.405 152.375 67.655 152.755 ;
        RECT 68.785 152.715 69.015 152.755 ;
        RECT 69.265 152.595 69.520 153.215 ;
        RECT 70.225 153.055 70.460 153.705 ;
        RECT 70.930 153.535 71.915 153.895 ;
        RECT 67.825 152.205 68.180 152.585 ;
        RECT 69.185 152.375 69.520 152.595 ;
        RECT 69.785 152.825 70.460 153.055 ;
        RECT 70.630 153.515 71.915 153.535 ;
        RECT 70.630 153.365 71.490 153.515 ;
        RECT 69.785 152.395 69.955 152.825 ;
        RECT 70.125 152.205 70.455 152.655 ;
        RECT 70.630 152.420 70.915 153.365 ;
        RECT 72.090 153.260 72.265 154.065 ;
        RECT 72.460 153.915 72.720 154.755 ;
        RECT 72.895 154.010 73.150 154.585 ;
        RECT 73.320 154.375 73.650 154.755 ;
        RECT 73.865 154.205 74.035 154.585 ;
        RECT 73.320 154.035 74.035 154.205 ;
        RECT 71.090 152.885 71.785 153.195 ;
        RECT 71.095 152.205 71.780 152.675 ;
        RECT 71.960 152.475 72.265 153.260 ;
        RECT 72.460 152.205 72.720 153.355 ;
        RECT 72.895 153.280 73.065 154.010 ;
        RECT 73.320 153.845 73.490 154.035 ;
        RECT 74.295 154.030 74.585 154.755 ;
        RECT 75.215 154.255 75.475 154.585 ;
        RECT 75.645 154.395 75.975 154.755 ;
        RECT 76.230 154.375 77.530 154.585 ;
        RECT 75.215 154.245 75.445 154.255 ;
        RECT 73.235 153.515 73.490 153.845 ;
        RECT 73.320 153.305 73.490 153.515 ;
        RECT 73.770 153.485 74.125 153.855 ;
        RECT 72.895 152.375 73.150 153.280 ;
        RECT 73.320 153.135 74.035 153.305 ;
        RECT 73.320 152.205 73.650 152.965 ;
        RECT 73.865 152.375 74.035 153.135 ;
        RECT 74.295 152.205 74.585 153.370 ;
        RECT 75.215 153.055 75.385 154.245 ;
        RECT 76.230 154.225 76.400 154.375 ;
        RECT 75.645 154.100 76.400 154.225 ;
        RECT 75.555 154.055 76.400 154.100 ;
        RECT 75.555 153.935 75.825 154.055 ;
        RECT 75.555 153.360 75.725 153.935 ;
        RECT 75.955 153.495 76.365 153.800 ;
        RECT 76.655 153.765 76.865 154.165 ;
        RECT 76.535 153.555 76.865 153.765 ;
        RECT 77.110 153.765 77.330 154.165 ;
        RECT 77.805 153.990 78.260 154.755 ;
        RECT 78.435 154.015 78.820 154.585 ;
        RECT 78.990 154.295 79.315 154.755 ;
        RECT 79.835 154.125 80.115 154.585 ;
        RECT 77.110 153.555 77.585 153.765 ;
        RECT 77.775 153.565 78.265 153.765 ;
        RECT 75.555 153.325 75.755 153.360 ;
        RECT 77.085 153.325 78.260 153.385 ;
        RECT 75.555 153.215 78.260 153.325 ;
        RECT 75.615 153.155 77.415 153.215 ;
        RECT 77.085 153.125 77.415 153.155 ;
        RECT 75.215 152.375 75.475 153.055 ;
        RECT 75.645 152.205 75.895 152.985 ;
        RECT 76.145 152.955 76.980 152.965 ;
        RECT 77.570 152.955 77.755 153.045 ;
        RECT 76.145 152.755 77.755 152.955 ;
        RECT 76.145 152.375 76.395 152.755 ;
        RECT 77.525 152.715 77.755 152.755 ;
        RECT 78.005 152.595 78.260 153.215 ;
        RECT 76.565 152.205 76.920 152.585 ;
        RECT 77.925 152.375 78.260 152.595 ;
        RECT 78.435 153.345 78.715 154.015 ;
        RECT 78.990 153.955 80.115 154.125 ;
        RECT 78.990 153.845 79.440 153.955 ;
        RECT 78.885 153.515 79.440 153.845 ;
        RECT 80.305 153.785 80.705 154.585 ;
        RECT 81.105 154.295 81.375 154.755 ;
        RECT 81.545 154.125 81.830 154.585 ;
        RECT 78.435 152.375 78.820 153.345 ;
        RECT 78.990 153.055 79.440 153.515 ;
        RECT 79.610 153.225 80.705 153.785 ;
        RECT 78.990 152.835 80.115 153.055 ;
        RECT 78.990 152.205 79.315 152.665 ;
        RECT 79.835 152.375 80.115 152.835 ;
        RECT 80.305 152.375 80.705 153.225 ;
        RECT 80.875 153.955 81.830 154.125 ;
        RECT 83.040 154.015 83.295 154.585 ;
        RECT 83.465 154.355 83.795 154.755 ;
        RECT 84.220 154.220 84.750 154.585 ;
        RECT 84.220 154.185 84.395 154.220 ;
        RECT 83.465 154.015 84.395 154.185 ;
        RECT 80.875 153.055 81.085 153.955 ;
        RECT 81.255 153.225 81.945 153.785 ;
        RECT 83.040 153.345 83.210 154.015 ;
        RECT 83.465 153.845 83.635 154.015 ;
        RECT 83.380 153.515 83.635 153.845 ;
        RECT 83.860 153.515 84.055 153.845 ;
        RECT 80.875 152.835 81.830 153.055 ;
        RECT 81.105 152.205 81.375 152.665 ;
        RECT 81.545 152.375 81.830 152.835 ;
        RECT 83.040 152.375 83.375 153.345 ;
        RECT 83.545 152.205 83.715 153.345 ;
        RECT 83.885 152.545 84.055 153.515 ;
        RECT 84.225 152.885 84.395 154.015 ;
        RECT 84.565 153.225 84.735 154.025 ;
        RECT 84.940 153.735 85.215 154.585 ;
        RECT 84.935 153.565 85.215 153.735 ;
        RECT 84.940 153.425 85.215 153.565 ;
        RECT 85.385 153.225 85.575 154.585 ;
        RECT 85.755 154.220 86.265 154.755 ;
        RECT 86.485 153.945 86.730 154.550 ;
        RECT 85.775 153.775 87.005 153.945 ;
        RECT 87.905 153.935 88.235 154.755 ;
        RECT 88.405 154.125 88.735 154.585 ;
        RECT 88.905 154.295 89.075 154.755 ;
        RECT 89.245 154.125 89.575 154.585 ;
        RECT 89.745 154.295 89.995 154.755 ;
        RECT 90.185 154.375 93.875 154.585 ;
        RECT 94.065 154.295 94.315 154.755 ;
        RECT 90.185 154.125 91.775 154.205 ;
        RECT 88.405 153.935 91.775 154.125 ;
        RECT 91.945 153.935 93.455 154.205 ;
        RECT 94.485 154.125 94.825 154.585 ;
        RECT 93.625 153.935 94.825 154.125 ;
        RECT 84.565 153.055 85.575 153.225 ;
        RECT 85.745 153.210 86.495 153.400 ;
        RECT 84.225 152.715 85.350 152.885 ;
        RECT 85.745 152.545 85.915 153.210 ;
        RECT 86.665 152.965 87.005 153.775 ;
        RECT 91.945 153.765 92.115 153.935 ;
        RECT 93.625 153.765 93.905 153.935 ;
        RECT 88.410 153.565 90.120 153.765 ;
        RECT 90.430 153.565 91.640 153.765 ;
        RECT 91.810 153.395 92.115 153.765 ;
        RECT 92.285 153.565 93.905 153.765 ;
        RECT 94.130 153.565 94.480 153.765 ;
        RECT 94.650 153.395 94.825 153.935 ;
        RECT 83.885 152.375 85.915 152.545 ;
        RECT 86.085 152.205 86.255 152.965 ;
        RECT 86.490 152.555 87.005 152.965 ;
        RECT 87.905 152.205 88.235 153.395 ;
        RECT 88.405 153.175 93.455 153.395 ;
        RECT 88.405 152.375 88.735 153.175 ;
        RECT 88.905 152.205 89.075 153.005 ;
        RECT 89.245 152.375 89.575 153.175 ;
        RECT 89.745 152.205 90.435 153.005 ;
        RECT 90.605 152.375 90.935 153.175 ;
        RECT 91.105 152.205 91.275 153.005 ;
        RECT 91.445 152.835 92.615 153.175 ;
        RECT 91.445 152.375 91.775 152.835 ;
        RECT 91.945 152.205 92.115 152.665 ;
        RECT 92.285 152.375 92.615 152.835 ;
        RECT 92.785 152.205 92.955 153.005 ;
        RECT 93.125 152.375 93.455 153.175 ;
        RECT 93.625 152.205 94.315 153.395 ;
        RECT 94.485 152.375 94.825 153.395 ;
        RECT 95.920 154.015 96.175 154.585 ;
        RECT 96.345 154.355 96.675 154.755 ;
        RECT 97.100 154.220 97.630 154.585 ;
        RECT 97.820 154.415 98.095 154.585 ;
        RECT 97.815 154.245 98.095 154.415 ;
        RECT 97.100 154.185 97.275 154.220 ;
        RECT 96.345 154.015 97.275 154.185 ;
        RECT 95.920 153.345 96.090 154.015 ;
        RECT 96.345 153.845 96.515 154.015 ;
        RECT 96.260 153.515 96.515 153.845 ;
        RECT 96.740 153.515 96.935 153.845 ;
        RECT 95.920 152.375 96.255 153.345 ;
        RECT 96.425 152.205 96.595 153.345 ;
        RECT 96.765 152.545 96.935 153.515 ;
        RECT 97.105 152.885 97.275 154.015 ;
        RECT 97.445 153.225 97.615 154.025 ;
        RECT 97.820 153.425 98.095 154.245 ;
        RECT 98.265 153.225 98.455 154.585 ;
        RECT 98.635 154.220 99.145 154.755 ;
        RECT 99.365 153.945 99.610 154.550 ;
        RECT 100.055 154.030 100.345 154.755 ;
        RECT 100.515 154.080 100.775 154.585 ;
        RECT 100.955 154.375 101.285 154.755 ;
        RECT 101.465 154.205 101.635 154.585 ;
        RECT 98.655 153.775 99.885 153.945 ;
        RECT 97.445 153.055 98.455 153.225 ;
        RECT 98.625 153.210 99.375 153.400 ;
        RECT 97.105 152.715 98.230 152.885 ;
        RECT 98.625 152.545 98.795 153.210 ;
        RECT 99.545 152.965 99.885 153.775 ;
        RECT 96.765 152.375 98.795 152.545 ;
        RECT 98.965 152.205 99.135 152.965 ;
        RECT 99.370 152.555 99.885 152.965 ;
        RECT 100.055 152.205 100.345 153.370 ;
        RECT 100.515 153.280 100.685 154.080 ;
        RECT 100.970 154.035 101.635 154.205 ;
        RECT 100.970 153.780 101.140 154.035 ;
        RECT 101.895 153.985 104.485 154.755 ;
        RECT 104.745 154.205 104.915 154.585 ;
        RECT 105.095 154.375 105.425 154.755 ;
        RECT 104.745 154.035 105.410 154.205 ;
        RECT 105.605 154.080 105.865 154.585 ;
        RECT 100.855 153.450 101.140 153.780 ;
        RECT 101.375 153.485 101.705 153.855 ;
        RECT 101.895 153.465 103.105 153.985 ;
        RECT 100.970 153.305 101.140 153.450 ;
        RECT 100.515 152.375 100.785 153.280 ;
        RECT 100.970 153.135 101.635 153.305 ;
        RECT 103.275 153.295 104.485 153.815 ;
        RECT 104.675 153.485 105.005 153.855 ;
        RECT 105.240 153.780 105.410 154.035 ;
        RECT 105.240 153.450 105.525 153.780 ;
        RECT 105.240 153.305 105.410 153.450 ;
        RECT 100.955 152.205 101.285 152.965 ;
        RECT 101.465 152.375 101.635 153.135 ;
        RECT 101.895 152.205 104.485 153.295 ;
        RECT 104.745 153.135 105.410 153.305 ;
        RECT 105.695 153.280 105.865 154.080 ;
        RECT 106.125 154.205 106.295 154.495 ;
        RECT 106.465 154.375 106.795 154.755 ;
        RECT 106.125 154.035 106.790 154.205 ;
        RECT 104.745 152.375 104.915 153.135 ;
        RECT 105.095 152.205 105.425 152.965 ;
        RECT 105.595 152.375 105.865 153.280 ;
        RECT 106.040 153.215 106.390 153.865 ;
        RECT 106.560 153.045 106.790 154.035 ;
        RECT 106.125 152.875 106.790 153.045 ;
        RECT 106.125 152.375 106.295 152.875 ;
        RECT 106.465 152.205 106.795 152.705 ;
        RECT 106.965 152.375 107.150 154.495 ;
        RECT 107.405 154.295 107.655 154.755 ;
        RECT 107.825 154.305 108.160 154.475 ;
        RECT 108.355 154.305 109.030 154.475 ;
        RECT 107.825 154.165 107.995 154.305 ;
        RECT 107.320 153.175 107.600 154.125 ;
        RECT 107.770 154.035 107.995 154.165 ;
        RECT 107.770 152.930 107.940 154.035 ;
        RECT 108.165 153.885 108.690 154.105 ;
        RECT 108.110 153.120 108.350 153.715 ;
        RECT 108.520 153.185 108.690 153.885 ;
        RECT 108.860 153.525 109.030 154.305 ;
        RECT 109.350 154.255 109.720 154.755 ;
        RECT 109.900 154.305 110.305 154.475 ;
        RECT 110.475 154.305 111.260 154.475 ;
        RECT 109.900 154.075 110.070 154.305 ;
        RECT 109.240 153.775 110.070 154.075 ;
        RECT 110.455 153.805 110.920 154.135 ;
        RECT 109.240 153.745 109.440 153.775 ;
        RECT 109.560 153.525 109.730 153.595 ;
        RECT 108.860 153.355 109.730 153.525 ;
        RECT 109.220 153.265 109.730 153.355 ;
        RECT 107.770 152.800 108.075 152.930 ;
        RECT 108.520 152.820 109.050 153.185 ;
        RECT 107.390 152.205 107.655 152.665 ;
        RECT 107.825 152.375 108.075 152.800 ;
        RECT 109.220 152.650 109.390 153.265 ;
        RECT 108.285 152.480 109.390 152.650 ;
        RECT 109.560 152.205 109.730 153.005 ;
        RECT 109.900 152.705 110.070 153.775 ;
        RECT 110.240 152.875 110.430 153.595 ;
        RECT 110.600 152.845 110.920 153.805 ;
        RECT 111.090 153.845 111.260 154.305 ;
        RECT 111.535 154.225 111.745 154.755 ;
        RECT 112.005 154.015 112.335 154.540 ;
        RECT 112.505 154.145 112.675 154.755 ;
        RECT 112.845 154.100 113.175 154.535 ;
        RECT 112.845 154.015 113.225 154.100 ;
        RECT 112.135 153.845 112.335 154.015 ;
        RECT 113.000 153.975 113.225 154.015 ;
        RECT 111.090 153.515 111.965 153.845 ;
        RECT 112.135 153.515 112.885 153.845 ;
        RECT 109.900 152.375 110.150 152.705 ;
        RECT 111.090 152.675 111.260 153.515 ;
        RECT 112.135 153.310 112.325 153.515 ;
        RECT 113.055 153.395 113.225 153.975 ;
        RECT 113.395 153.985 115.065 154.755 ;
        RECT 113.395 153.465 114.145 153.985 ;
        RECT 115.510 153.945 115.755 154.550 ;
        RECT 115.975 154.220 116.485 154.755 ;
        RECT 113.010 153.345 113.225 153.395 ;
        RECT 111.430 152.935 112.325 153.310 ;
        RECT 112.835 153.265 113.225 153.345 ;
        RECT 114.315 153.295 115.065 153.815 ;
        RECT 110.375 152.505 111.260 152.675 ;
        RECT 111.440 152.205 111.755 152.705 ;
        RECT 111.985 152.375 112.325 152.935 ;
        RECT 112.495 152.205 112.665 153.215 ;
        RECT 112.835 152.420 113.165 153.265 ;
        RECT 113.395 152.205 115.065 153.295 ;
        RECT 115.235 153.775 116.465 153.945 ;
        RECT 115.235 152.965 115.575 153.775 ;
        RECT 115.745 153.210 116.495 153.400 ;
        RECT 115.235 152.555 115.750 152.965 ;
        RECT 115.985 152.205 116.155 152.965 ;
        RECT 116.325 152.545 116.495 153.210 ;
        RECT 116.665 153.225 116.855 154.585 ;
        RECT 117.025 154.415 117.300 154.585 ;
        RECT 117.025 154.245 117.305 154.415 ;
        RECT 117.025 153.425 117.300 154.245 ;
        RECT 117.490 154.220 118.020 154.585 ;
        RECT 118.445 154.355 118.775 154.755 ;
        RECT 117.845 154.185 118.020 154.220 ;
        RECT 117.505 153.225 117.675 154.025 ;
        RECT 116.665 153.055 117.675 153.225 ;
        RECT 117.845 154.015 118.775 154.185 ;
        RECT 118.945 154.015 119.200 154.585 ;
        RECT 117.845 152.885 118.015 154.015 ;
        RECT 118.605 153.845 118.775 154.015 ;
        RECT 116.890 152.715 118.015 152.885 ;
        RECT 118.185 153.515 118.380 153.845 ;
        RECT 118.605 153.515 118.860 153.845 ;
        RECT 118.185 152.545 118.355 153.515 ;
        RECT 119.030 153.345 119.200 154.015 ;
        RECT 116.325 152.375 118.355 152.545 ;
        RECT 118.525 152.205 118.695 153.345 ;
        RECT 118.865 152.375 119.200 153.345 ;
        RECT 119.375 154.295 119.935 154.585 ;
        RECT 120.105 154.295 120.355 154.755 ;
        RECT 119.375 152.925 119.625 154.295 ;
        RECT 120.975 154.125 121.305 154.485 ;
        RECT 119.915 153.935 121.305 154.125 ;
        RECT 121.675 154.080 121.935 154.585 ;
        RECT 122.115 154.375 122.445 154.755 ;
        RECT 122.625 154.205 122.795 154.585 ;
        RECT 119.915 153.845 120.085 153.935 ;
        RECT 119.795 153.515 120.085 153.845 ;
        RECT 120.255 153.515 120.595 153.765 ;
        RECT 120.815 153.515 121.490 153.765 ;
        RECT 119.915 153.265 120.085 153.515 ;
        RECT 119.915 153.095 120.855 153.265 ;
        RECT 121.225 153.155 121.490 153.515 ;
        RECT 121.675 153.280 121.845 154.080 ;
        RECT 122.130 154.035 122.795 154.205 ;
        RECT 123.715 154.125 124.045 154.485 ;
        RECT 124.665 154.295 124.915 154.755 ;
        RECT 125.085 154.295 125.645 154.585 ;
        RECT 122.130 153.780 122.300 154.035 ;
        RECT 123.715 153.935 125.105 154.125 ;
        RECT 122.015 153.450 122.300 153.780 ;
        RECT 122.535 153.485 122.865 153.855 ;
        RECT 124.935 153.845 125.105 153.935 ;
        RECT 123.530 153.515 124.205 153.765 ;
        RECT 124.425 153.515 124.765 153.765 ;
        RECT 124.935 153.515 125.225 153.845 ;
        RECT 122.130 153.305 122.300 153.450 ;
        RECT 119.375 152.375 119.835 152.925 ;
        RECT 120.025 152.205 120.355 152.925 ;
        RECT 120.555 152.545 120.855 153.095 ;
        RECT 121.025 152.205 121.305 152.875 ;
        RECT 121.675 152.375 121.945 153.280 ;
        RECT 122.130 153.135 122.795 153.305 ;
        RECT 123.530 153.155 123.795 153.515 ;
        RECT 124.935 153.265 125.105 153.515 ;
        RECT 122.115 152.205 122.445 152.965 ;
        RECT 122.625 152.375 122.795 153.135 ;
        RECT 124.165 153.095 125.105 153.265 ;
        RECT 123.715 152.205 123.995 152.875 ;
        RECT 124.165 152.545 124.465 153.095 ;
        RECT 125.395 152.925 125.645 154.295 ;
        RECT 125.815 154.030 126.105 154.755 ;
        RECT 126.280 154.015 126.535 154.585 ;
        RECT 126.705 154.355 127.035 154.755 ;
        RECT 127.460 154.220 127.990 154.585 ;
        RECT 127.460 154.185 127.635 154.220 ;
        RECT 126.705 154.015 127.635 154.185 ;
        RECT 124.665 152.205 124.995 152.925 ;
        RECT 125.185 152.375 125.645 152.925 ;
        RECT 125.815 152.205 126.105 153.370 ;
        RECT 126.280 153.345 126.450 154.015 ;
        RECT 126.705 153.845 126.875 154.015 ;
        RECT 126.620 153.515 126.875 153.845 ;
        RECT 127.100 153.515 127.295 153.845 ;
        RECT 126.280 152.375 126.615 153.345 ;
        RECT 126.785 152.205 126.955 153.345 ;
        RECT 127.125 152.545 127.295 153.515 ;
        RECT 127.465 152.885 127.635 154.015 ;
        RECT 127.805 153.225 127.975 154.025 ;
        RECT 128.180 153.735 128.455 154.585 ;
        RECT 128.175 153.565 128.455 153.735 ;
        RECT 128.180 153.425 128.455 153.565 ;
        RECT 128.625 153.225 128.815 154.585 ;
        RECT 128.995 154.220 129.505 154.755 ;
        RECT 129.725 153.945 129.970 154.550 ;
        RECT 129.015 153.775 130.245 153.945 ;
        RECT 130.915 153.935 131.145 154.755 ;
        RECT 131.315 153.955 131.645 154.585 ;
        RECT 127.805 153.055 128.815 153.225 ;
        RECT 128.985 153.210 129.735 153.400 ;
        RECT 127.465 152.715 128.590 152.885 ;
        RECT 128.985 152.545 129.155 153.210 ;
        RECT 129.905 152.965 130.245 153.775 ;
        RECT 130.895 153.515 131.225 153.765 ;
        RECT 131.395 153.355 131.645 153.955 ;
        RECT 131.815 153.935 132.025 154.755 ;
        RECT 132.255 153.985 133.925 154.755 ;
        RECT 134.555 154.245 134.860 154.755 ;
        RECT 132.255 153.465 133.005 153.985 ;
        RECT 127.125 152.375 129.155 152.545 ;
        RECT 129.325 152.205 129.495 152.965 ;
        RECT 129.730 152.555 130.245 152.965 ;
        RECT 130.915 152.205 131.145 153.345 ;
        RECT 131.315 152.375 131.645 153.355 ;
        RECT 131.815 152.205 132.025 153.345 ;
        RECT 133.175 153.295 133.925 153.815 ;
        RECT 134.555 153.515 134.870 154.075 ;
        RECT 135.040 153.765 135.290 154.575 ;
        RECT 135.460 154.230 135.720 154.755 ;
        RECT 135.900 153.765 136.150 154.575 ;
        RECT 136.320 154.195 136.580 154.755 ;
        RECT 136.750 154.105 137.010 154.560 ;
        RECT 137.180 154.275 137.440 154.755 ;
        RECT 137.610 154.105 137.870 154.560 ;
        RECT 138.040 154.275 138.300 154.755 ;
        RECT 138.470 154.105 138.730 154.560 ;
        RECT 138.900 154.275 139.145 154.755 ;
        RECT 139.315 154.105 139.590 154.560 ;
        RECT 139.760 154.275 140.005 154.755 ;
        RECT 140.175 154.105 140.435 154.560 ;
        RECT 140.615 154.275 140.865 154.755 ;
        RECT 141.035 154.105 141.295 154.560 ;
        RECT 141.475 154.275 141.725 154.755 ;
        RECT 141.895 154.105 142.155 154.560 ;
        RECT 142.335 154.275 142.595 154.755 ;
        RECT 142.765 154.105 143.025 154.560 ;
        RECT 143.195 154.275 143.495 154.755 ;
        RECT 143.755 154.210 149.100 154.755 ;
        RECT 136.750 153.935 143.495 154.105 ;
        RECT 135.040 153.515 142.160 153.765 ;
        RECT 132.255 152.205 133.925 153.295 ;
        RECT 134.565 152.205 134.860 153.015 ;
        RECT 135.040 152.375 135.285 153.515 ;
        RECT 135.460 152.205 135.720 153.015 ;
        RECT 135.900 152.380 136.150 153.515 ;
        RECT 142.330 153.345 143.495 153.935 ;
        RECT 145.340 153.380 145.680 154.210 ;
        RECT 149.275 153.985 150.945 154.755 ;
        RECT 151.575 154.030 151.865 154.755 ;
        RECT 152.035 154.015 152.420 154.585 ;
        RECT 152.590 154.295 152.915 154.755 ;
        RECT 153.435 154.125 153.715 154.585 ;
        RECT 136.750 153.120 143.495 153.345 ;
        RECT 136.750 153.105 142.155 153.120 ;
        RECT 136.320 152.210 136.580 153.005 ;
        RECT 136.750 152.380 137.010 153.105 ;
        RECT 137.180 152.210 137.440 152.935 ;
        RECT 137.610 152.380 137.870 153.105 ;
        RECT 138.040 152.210 138.300 152.935 ;
        RECT 138.470 152.380 138.730 153.105 ;
        RECT 138.900 152.210 139.160 152.935 ;
        RECT 139.330 152.380 139.590 153.105 ;
        RECT 139.760 152.210 140.005 152.935 ;
        RECT 140.175 152.380 140.435 153.105 ;
        RECT 140.620 152.210 140.865 152.935 ;
        RECT 141.035 152.380 141.295 153.105 ;
        RECT 141.480 152.210 141.725 152.935 ;
        RECT 141.895 152.380 142.155 153.105 ;
        RECT 142.340 152.210 142.595 152.935 ;
        RECT 142.765 152.380 143.055 153.120 ;
        RECT 136.320 152.205 142.595 152.210 ;
        RECT 143.225 152.205 143.495 152.950 ;
        RECT 147.160 152.640 147.510 153.890 ;
        RECT 149.275 153.465 150.025 153.985 ;
        RECT 150.195 153.295 150.945 153.815 ;
        RECT 143.755 152.205 149.100 152.640 ;
        RECT 149.275 152.205 150.945 153.295 ;
        RECT 151.575 152.205 151.865 153.370 ;
        RECT 152.035 153.345 152.315 154.015 ;
        RECT 152.590 153.955 153.715 154.125 ;
        RECT 152.590 153.845 153.040 153.955 ;
        RECT 152.485 153.515 153.040 153.845 ;
        RECT 153.905 153.785 154.305 154.585 ;
        RECT 154.705 154.295 154.975 154.755 ;
        RECT 155.145 154.125 155.430 154.585 ;
        RECT 152.035 152.375 152.420 153.345 ;
        RECT 152.590 153.055 153.040 153.515 ;
        RECT 153.210 153.225 154.305 153.785 ;
        RECT 152.590 152.835 153.715 153.055 ;
        RECT 152.590 152.205 152.915 152.665 ;
        RECT 153.435 152.375 153.715 152.835 ;
        RECT 153.905 152.375 154.305 153.225 ;
        RECT 154.475 153.955 155.430 154.125 ;
        RECT 155.715 154.005 156.925 154.755 ;
        RECT 154.475 153.055 154.685 153.955 ;
        RECT 154.855 153.225 155.545 153.785 ;
        RECT 155.715 153.295 156.235 153.835 ;
        RECT 156.405 153.465 156.925 154.005 ;
        RECT 154.475 152.835 155.430 153.055 ;
        RECT 154.705 152.205 154.975 152.665 ;
        RECT 155.145 152.375 155.430 152.835 ;
        RECT 155.715 152.205 156.925 153.295 ;
        RECT 22.690 152.035 157.010 152.205 ;
        RECT 22.775 150.945 23.985 152.035 ;
        RECT 24.245 151.365 24.415 151.865 ;
        RECT 24.585 151.535 24.915 152.035 ;
        RECT 24.245 151.195 24.910 151.365 ;
        RECT 22.775 150.235 23.295 150.775 ;
        RECT 23.465 150.405 23.985 150.945 ;
        RECT 24.160 150.375 24.510 151.025 ;
        RECT 22.775 149.485 23.985 150.235 ;
        RECT 24.680 150.205 24.910 151.195 ;
        RECT 24.245 150.035 24.910 150.205 ;
        RECT 24.245 149.745 24.415 150.035 ;
        RECT 24.585 149.485 24.915 149.865 ;
        RECT 25.085 149.745 25.270 151.865 ;
        RECT 25.510 151.575 25.775 152.035 ;
        RECT 25.945 151.440 26.195 151.865 ;
        RECT 26.405 151.590 27.510 151.760 ;
        RECT 25.890 151.310 26.195 151.440 ;
        RECT 25.440 150.115 25.720 151.065 ;
        RECT 25.890 150.205 26.060 151.310 ;
        RECT 26.230 150.525 26.470 151.120 ;
        RECT 26.640 151.055 27.170 151.420 ;
        RECT 26.640 150.355 26.810 151.055 ;
        RECT 27.340 150.975 27.510 151.590 ;
        RECT 27.680 151.235 27.850 152.035 ;
        RECT 28.020 151.535 28.270 151.865 ;
        RECT 28.495 151.565 29.380 151.735 ;
        RECT 27.340 150.885 27.850 150.975 ;
        RECT 25.890 150.075 26.115 150.205 ;
        RECT 26.285 150.135 26.810 150.355 ;
        RECT 26.980 150.715 27.850 150.885 ;
        RECT 25.525 149.485 25.775 149.945 ;
        RECT 25.945 149.935 26.115 150.075 ;
        RECT 26.980 149.935 27.150 150.715 ;
        RECT 27.680 150.645 27.850 150.715 ;
        RECT 27.360 150.465 27.560 150.495 ;
        RECT 28.020 150.465 28.190 151.535 ;
        RECT 28.360 150.645 28.550 151.365 ;
        RECT 27.360 150.165 28.190 150.465 ;
        RECT 28.720 150.435 29.040 151.395 ;
        RECT 25.945 149.765 26.280 149.935 ;
        RECT 26.475 149.765 27.150 149.935 ;
        RECT 27.470 149.485 27.840 149.985 ;
        RECT 28.020 149.935 28.190 150.165 ;
        RECT 28.575 150.105 29.040 150.435 ;
        RECT 29.210 150.725 29.380 151.565 ;
        RECT 29.560 151.535 29.875 152.035 ;
        RECT 30.105 151.305 30.445 151.865 ;
        RECT 29.550 150.930 30.445 151.305 ;
        RECT 30.615 151.025 30.785 152.035 ;
        RECT 30.255 150.725 30.445 150.930 ;
        RECT 30.955 150.975 31.285 151.820 ;
        RECT 30.955 150.895 31.345 150.975 ;
        RECT 31.515 150.945 32.725 152.035 ;
        RECT 31.130 150.845 31.345 150.895 ;
        RECT 29.210 150.395 30.085 150.725 ;
        RECT 30.255 150.395 31.005 150.725 ;
        RECT 29.210 149.935 29.380 150.395 ;
        RECT 30.255 150.225 30.455 150.395 ;
        RECT 31.175 150.265 31.345 150.845 ;
        RECT 31.120 150.225 31.345 150.265 ;
        RECT 28.020 149.765 28.425 149.935 ;
        RECT 28.595 149.765 29.380 149.935 ;
        RECT 29.655 149.485 29.865 150.015 ;
        RECT 30.125 149.700 30.455 150.225 ;
        RECT 30.965 150.140 31.345 150.225 ;
        RECT 31.515 150.235 32.035 150.775 ;
        RECT 32.205 150.405 32.725 150.945 ;
        RECT 32.905 150.895 33.235 152.035 ;
        RECT 33.765 151.065 34.095 151.850 ;
        RECT 33.415 150.895 34.095 151.065 ;
        RECT 34.275 150.945 35.485 152.035 ;
        RECT 32.895 150.475 33.245 150.725 ;
        RECT 33.415 150.295 33.585 150.895 ;
        RECT 33.755 150.475 34.105 150.725 ;
        RECT 30.625 149.485 30.795 150.095 ;
        RECT 30.965 149.705 31.295 150.140 ;
        RECT 31.515 149.485 32.725 150.235 ;
        RECT 32.905 149.485 33.175 150.295 ;
        RECT 33.345 149.655 33.675 150.295 ;
        RECT 33.845 149.485 34.085 150.295 ;
        RECT 34.275 150.235 34.795 150.775 ;
        RECT 34.965 150.405 35.485 150.945 ;
        RECT 35.655 150.870 35.945 152.035 ;
        RECT 36.115 150.945 37.325 152.035 ;
        RECT 36.115 150.235 36.635 150.775 ;
        RECT 36.805 150.405 37.325 150.945 ;
        RECT 37.585 151.105 37.755 151.865 ;
        RECT 37.970 151.275 38.300 152.035 ;
        RECT 37.585 150.935 38.300 151.105 ;
        RECT 38.470 150.960 38.725 151.865 ;
        RECT 37.495 150.385 37.850 150.755 ;
        RECT 38.130 150.725 38.300 150.935 ;
        RECT 38.130 150.395 38.385 150.725 ;
        RECT 34.275 149.485 35.485 150.235 ;
        RECT 35.655 149.485 35.945 150.210 ;
        RECT 36.115 149.485 37.325 150.235 ;
        RECT 38.130 150.205 38.300 150.395 ;
        RECT 38.555 150.230 38.725 150.960 ;
        RECT 38.900 150.885 39.160 152.035 ;
        RECT 39.485 150.885 39.815 152.035 ;
        RECT 39.985 151.015 40.155 151.865 ;
        RECT 40.325 151.235 40.655 152.035 ;
        RECT 40.825 151.015 40.995 151.865 ;
        RECT 41.175 151.235 41.415 152.035 ;
        RECT 41.585 151.055 41.915 151.865 ;
        RECT 39.985 150.845 40.995 151.015 ;
        RECT 41.200 150.885 41.915 151.055 ;
        RECT 42.095 150.925 42.355 151.865 ;
        RECT 42.525 151.635 42.855 152.035 ;
        RECT 44.000 151.770 44.255 151.865 ;
        RECT 43.115 151.600 44.255 151.770 ;
        RECT 44.425 151.655 44.755 151.825 ;
        RECT 43.115 151.375 43.285 151.600 ;
        RECT 42.525 151.205 43.285 151.375 ;
        RECT 44.000 151.465 44.255 151.600 ;
        RECT 39.985 150.675 40.480 150.845 ;
        RECT 39.985 150.505 40.485 150.675 ;
        RECT 41.200 150.645 41.370 150.885 ;
        RECT 37.585 150.035 38.300 150.205 ;
        RECT 37.585 149.655 37.755 150.035 ;
        RECT 37.970 149.485 38.300 149.865 ;
        RECT 38.470 149.655 38.725 150.230 ;
        RECT 38.900 149.485 39.160 150.325 ;
        RECT 39.985 150.305 40.480 150.505 ;
        RECT 40.870 150.475 41.370 150.645 ;
        RECT 41.540 150.475 41.920 150.715 ;
        RECT 41.200 150.305 41.370 150.475 ;
        RECT 39.485 149.485 39.815 150.285 ;
        RECT 39.985 150.135 40.995 150.305 ;
        RECT 41.200 150.135 41.835 150.305 ;
        RECT 39.985 149.655 40.155 150.135 ;
        RECT 40.325 149.485 40.655 149.965 ;
        RECT 40.825 149.655 40.995 150.135 ;
        RECT 41.245 149.485 41.485 149.965 ;
        RECT 41.665 149.655 41.835 150.135 ;
        RECT 42.095 150.210 42.270 150.925 ;
        RECT 42.525 150.725 42.695 151.205 ;
        RECT 43.550 151.115 43.720 151.305 ;
        RECT 44.000 151.295 44.410 151.465 ;
        RECT 42.440 150.395 42.695 150.725 ;
        RECT 42.920 150.395 43.250 151.015 ;
        RECT 43.550 150.945 44.070 151.115 ;
        RECT 43.420 150.395 43.710 150.775 ;
        RECT 43.900 150.225 44.070 150.945 ;
        RECT 42.095 149.655 42.355 150.210 ;
        RECT 43.190 150.055 44.070 150.225 ;
        RECT 44.240 150.270 44.410 151.295 ;
        RECT 44.585 151.405 44.755 151.655 ;
        RECT 44.925 151.575 45.175 152.035 ;
        RECT 45.345 151.405 45.525 151.865 ;
        RECT 44.585 151.235 45.525 151.405 ;
        RECT 44.610 150.755 45.090 151.055 ;
        RECT 44.240 150.100 44.590 150.270 ;
        RECT 44.830 150.165 45.090 150.755 ;
        RECT 45.290 150.165 45.550 151.055 ;
        RECT 45.775 150.895 46.160 151.865 ;
        RECT 46.330 151.575 46.655 152.035 ;
        RECT 47.175 151.405 47.455 151.865 ;
        RECT 46.330 151.185 47.455 151.405 ;
        RECT 45.775 150.225 46.055 150.895 ;
        RECT 46.330 150.725 46.780 151.185 ;
        RECT 47.645 151.015 48.045 151.865 ;
        RECT 48.445 151.575 48.715 152.035 ;
        RECT 48.885 151.405 49.170 151.865 ;
        RECT 46.225 150.395 46.780 150.725 ;
        RECT 46.950 150.455 48.045 151.015 ;
        RECT 46.330 150.285 46.780 150.395 ;
        RECT 42.525 149.485 42.955 149.930 ;
        RECT 43.190 149.655 43.360 150.055 ;
        RECT 43.530 149.485 44.250 149.885 ;
        RECT 44.420 149.655 44.590 150.100 ;
        RECT 45.165 149.485 45.565 149.995 ;
        RECT 45.775 149.655 46.160 150.225 ;
        RECT 46.330 150.115 47.455 150.285 ;
        RECT 46.330 149.485 46.655 149.945 ;
        RECT 47.175 149.655 47.455 150.115 ;
        RECT 47.645 149.655 48.045 150.455 ;
        RECT 48.215 151.185 49.170 151.405 ;
        RECT 49.465 151.225 49.760 152.035 ;
        RECT 48.215 150.285 48.425 151.185 ;
        RECT 48.595 150.455 49.285 151.015 ;
        RECT 49.940 150.725 50.185 151.865 ;
        RECT 50.360 151.225 50.620 152.035 ;
        RECT 51.220 152.030 57.495 152.035 ;
        RECT 50.800 150.725 51.050 151.860 ;
        RECT 51.220 151.235 51.480 152.030 ;
        RECT 51.650 151.135 51.910 151.860 ;
        RECT 52.080 151.305 52.340 152.030 ;
        RECT 52.510 151.135 52.770 151.860 ;
        RECT 52.940 151.305 53.200 152.030 ;
        RECT 53.370 151.135 53.630 151.860 ;
        RECT 53.800 151.305 54.060 152.030 ;
        RECT 54.230 151.135 54.490 151.860 ;
        RECT 54.660 151.305 54.905 152.030 ;
        RECT 55.075 151.135 55.335 151.860 ;
        RECT 55.520 151.305 55.765 152.030 ;
        RECT 55.935 151.135 56.195 151.860 ;
        RECT 56.380 151.305 56.625 152.030 ;
        RECT 56.795 151.135 57.055 151.860 ;
        RECT 57.240 151.305 57.495 152.030 ;
        RECT 51.650 151.120 57.055 151.135 ;
        RECT 57.665 151.120 57.955 151.860 ;
        RECT 58.125 151.290 58.395 152.035 ;
        RECT 51.650 150.895 58.395 151.120 ;
        RECT 58.655 150.945 61.245 152.035 ;
        RECT 48.215 150.115 49.170 150.285 ;
        RECT 49.455 150.165 49.770 150.725 ;
        RECT 49.940 150.475 57.060 150.725 ;
        RECT 57.230 150.675 58.395 150.895 ;
        RECT 57.230 150.505 58.425 150.675 ;
        RECT 48.445 149.485 48.715 149.945 ;
        RECT 48.885 149.655 49.170 150.115 ;
        RECT 49.455 149.485 49.760 149.995 ;
        RECT 49.940 149.665 50.190 150.475 ;
        RECT 50.360 149.485 50.620 150.010 ;
        RECT 50.800 149.665 51.050 150.475 ;
        RECT 57.230 150.305 58.395 150.505 ;
        RECT 51.650 150.135 58.395 150.305 ;
        RECT 58.655 150.255 59.865 150.775 ;
        RECT 60.035 150.425 61.245 150.945 ;
        RECT 61.415 150.870 61.705 152.035 ;
        RECT 61.885 150.975 62.215 151.825 ;
        RECT 51.220 149.485 51.480 150.045 ;
        RECT 51.650 149.680 51.910 150.135 ;
        RECT 52.080 149.485 52.340 149.965 ;
        RECT 52.510 149.680 52.770 150.135 ;
        RECT 52.940 149.485 53.200 149.965 ;
        RECT 53.370 149.680 53.630 150.135 ;
        RECT 53.800 149.485 54.045 149.965 ;
        RECT 54.215 149.680 54.490 150.135 ;
        RECT 54.660 149.485 54.905 149.965 ;
        RECT 55.075 149.680 55.335 150.135 ;
        RECT 55.515 149.485 55.765 149.965 ;
        RECT 55.935 149.680 56.195 150.135 ;
        RECT 56.375 149.485 56.625 149.965 ;
        RECT 56.795 149.680 57.055 150.135 ;
        RECT 57.235 149.485 57.495 149.965 ;
        RECT 57.665 149.680 57.925 150.135 ;
        RECT 58.095 149.485 58.395 149.965 ;
        RECT 58.655 149.485 61.245 150.255 ;
        RECT 61.885 150.210 62.075 150.975 ;
        RECT 62.385 150.895 62.635 152.035 ;
        RECT 62.825 151.395 63.075 151.815 ;
        RECT 63.305 151.565 63.635 152.035 ;
        RECT 63.865 151.395 64.115 151.815 ;
        RECT 62.825 151.225 64.115 151.395 ;
        RECT 64.295 151.395 64.625 151.825 ;
        RECT 65.095 151.480 65.700 152.035 ;
        RECT 65.875 151.525 66.355 151.865 ;
        RECT 66.525 151.490 66.780 152.035 ;
        RECT 64.295 151.225 64.750 151.395 ;
        RECT 65.095 151.380 65.710 151.480 ;
        RECT 62.815 150.725 63.030 151.055 ;
        RECT 62.245 150.395 62.555 150.725 ;
        RECT 62.725 150.395 63.030 150.725 ;
        RECT 63.205 150.395 63.490 151.055 ;
        RECT 63.685 150.395 63.950 151.055 ;
        RECT 64.165 150.395 64.410 151.055 ;
        RECT 62.385 150.225 62.555 150.395 ;
        RECT 64.580 150.225 64.750 151.225 ;
        RECT 65.525 151.355 65.710 151.380 ;
        RECT 65.095 150.760 65.355 151.210 ;
        RECT 65.525 151.110 65.855 151.355 ;
        RECT 66.025 151.035 66.780 151.285 ;
        RECT 66.950 151.165 67.225 151.865 ;
        RECT 66.010 151.000 66.780 151.035 ;
        RECT 65.995 150.990 66.780 151.000 ;
        RECT 65.990 150.975 66.885 150.990 ;
        RECT 65.970 150.960 66.885 150.975 ;
        RECT 65.950 150.950 66.885 150.960 ;
        RECT 65.925 150.940 66.885 150.950 ;
        RECT 65.855 150.910 66.885 150.940 ;
        RECT 65.835 150.880 66.885 150.910 ;
        RECT 65.815 150.850 66.885 150.880 ;
        RECT 65.785 150.825 66.885 150.850 ;
        RECT 65.750 150.790 66.885 150.825 ;
        RECT 65.720 150.785 66.885 150.790 ;
        RECT 65.720 150.780 66.110 150.785 ;
        RECT 65.720 150.770 66.085 150.780 ;
        RECT 65.720 150.765 66.070 150.770 ;
        RECT 65.720 150.760 66.055 150.765 ;
        RECT 65.095 150.755 66.055 150.760 ;
        RECT 65.095 150.745 66.045 150.755 ;
        RECT 65.095 150.740 66.035 150.745 ;
        RECT 65.095 150.730 66.025 150.740 ;
        RECT 65.095 150.720 66.020 150.730 ;
        RECT 65.095 150.715 66.015 150.720 ;
        RECT 65.095 150.700 66.005 150.715 ;
        RECT 65.095 150.685 66.000 150.700 ;
        RECT 65.095 150.660 65.990 150.685 ;
        RECT 65.095 150.590 65.985 150.660 ;
        RECT 61.415 149.485 61.705 150.210 ;
        RECT 61.885 149.700 62.215 150.210 ;
        RECT 62.385 150.055 64.750 150.225 ;
        RECT 62.385 149.485 62.715 149.885 ;
        RECT 63.765 149.715 64.095 150.055 ;
        RECT 65.095 150.035 65.645 150.420 ;
        RECT 64.265 149.485 64.595 149.885 ;
        RECT 65.815 149.865 65.985 150.590 ;
        RECT 65.095 149.695 65.985 149.865 ;
        RECT 66.155 150.190 66.485 150.615 ;
        RECT 66.655 150.390 66.885 150.785 ;
        RECT 66.155 149.705 66.375 150.190 ;
        RECT 67.055 150.135 67.225 151.165 ;
        RECT 67.860 151.645 68.195 151.865 ;
        RECT 69.200 151.655 69.555 152.035 ;
        RECT 67.860 151.025 68.115 151.645 ;
        RECT 68.365 151.485 68.595 151.525 ;
        RECT 69.725 151.485 69.975 151.865 ;
        RECT 68.365 151.285 69.975 151.485 ;
        RECT 68.365 151.195 68.550 151.285 ;
        RECT 69.140 151.275 69.975 151.285 ;
        RECT 70.225 151.255 70.475 152.035 ;
        RECT 70.645 151.185 70.905 151.865 ;
        RECT 68.705 151.085 69.035 151.115 ;
        RECT 68.705 151.025 70.505 151.085 ;
        RECT 67.860 150.915 70.565 151.025 ;
        RECT 67.860 150.855 69.035 150.915 ;
        RECT 70.365 150.880 70.565 150.915 ;
        RECT 67.855 150.475 68.345 150.675 ;
        RECT 68.535 150.475 69.010 150.685 ;
        RECT 66.545 149.485 66.795 150.025 ;
        RECT 66.965 149.655 67.225 150.135 ;
        RECT 67.860 149.485 68.315 150.250 ;
        RECT 68.790 150.075 69.010 150.475 ;
        RECT 69.255 150.475 69.585 150.685 ;
        RECT 69.255 150.075 69.465 150.475 ;
        RECT 69.755 150.440 70.165 150.745 ;
        RECT 70.395 150.305 70.565 150.880 ;
        RECT 70.295 150.185 70.565 150.305 ;
        RECT 69.720 150.140 70.565 150.185 ;
        RECT 69.720 150.015 70.475 150.140 ;
        RECT 69.720 149.865 69.890 150.015 ;
        RECT 70.735 149.995 70.905 151.185 ;
        RECT 70.675 149.985 70.905 149.995 ;
        RECT 68.590 149.655 69.890 149.865 ;
        RECT 70.145 149.485 70.475 149.845 ;
        RECT 70.645 149.655 70.905 149.985 ;
        RECT 71.090 149.665 71.370 151.855 ;
        RECT 71.560 150.895 71.845 152.035 ;
        RECT 72.110 151.385 72.280 151.855 ;
        RECT 72.455 151.555 72.785 152.035 ;
        RECT 72.955 151.385 73.135 151.855 ;
        RECT 72.110 151.185 73.135 151.385 ;
        RECT 71.570 150.215 71.830 150.725 ;
        RECT 72.040 150.395 72.300 151.015 ;
        RECT 72.495 150.395 72.920 151.015 ;
        RECT 73.305 150.745 73.635 151.855 ;
        RECT 73.805 151.625 74.155 152.035 ;
        RECT 74.325 151.445 74.565 151.835 ;
        RECT 73.090 150.445 73.635 150.745 ;
        RECT 73.815 151.245 74.565 151.445 ;
        RECT 75.790 151.405 76.075 151.865 ;
        RECT 76.245 151.575 76.515 152.035 ;
        RECT 73.815 150.565 74.155 151.245 ;
        RECT 75.790 151.185 76.745 151.405 ;
        RECT 73.090 150.215 73.310 150.445 ;
        RECT 71.570 150.025 73.310 150.215 ;
        RECT 71.570 149.485 72.300 149.855 ;
        RECT 72.880 149.665 73.310 150.025 ;
        RECT 73.480 149.485 73.725 150.265 ;
        RECT 73.925 149.665 74.155 150.565 ;
        RECT 74.335 149.725 74.565 151.065 ;
        RECT 75.675 150.455 76.365 151.015 ;
        RECT 76.535 150.285 76.745 151.185 ;
        RECT 75.790 150.115 76.745 150.285 ;
        RECT 76.915 151.015 77.315 151.865 ;
        RECT 77.505 151.405 77.785 151.865 ;
        RECT 78.305 151.575 78.630 152.035 ;
        RECT 77.505 151.185 78.630 151.405 ;
        RECT 76.915 150.455 78.010 151.015 ;
        RECT 78.180 150.725 78.630 151.185 ;
        RECT 78.800 150.895 79.185 151.865 ;
        RECT 75.790 149.655 76.075 150.115 ;
        RECT 76.245 149.485 76.515 149.945 ;
        RECT 76.915 149.655 77.315 150.455 ;
        RECT 78.180 150.395 78.735 150.725 ;
        RECT 78.180 150.285 78.630 150.395 ;
        RECT 77.505 150.115 78.630 150.285 ;
        RECT 78.905 150.225 79.185 150.895 ;
        RECT 79.360 151.645 79.695 151.865 ;
        RECT 80.700 151.655 81.055 152.035 ;
        RECT 79.360 151.025 79.615 151.645 ;
        RECT 79.865 151.485 80.095 151.525 ;
        RECT 81.225 151.485 81.475 151.865 ;
        RECT 79.865 151.285 81.475 151.485 ;
        RECT 79.865 151.195 80.050 151.285 ;
        RECT 80.640 151.275 81.475 151.285 ;
        RECT 81.725 151.255 81.975 152.035 ;
        RECT 82.145 151.185 82.405 151.865 ;
        RECT 80.205 151.085 80.535 151.115 ;
        RECT 80.205 151.025 82.005 151.085 ;
        RECT 79.360 150.915 82.065 151.025 ;
        RECT 79.360 150.855 80.535 150.915 ;
        RECT 81.865 150.880 82.065 150.915 ;
        RECT 79.355 150.475 79.845 150.675 ;
        RECT 80.035 150.475 80.510 150.685 ;
        RECT 77.505 149.655 77.785 150.115 ;
        RECT 78.305 149.485 78.630 149.945 ;
        RECT 78.800 149.655 79.185 150.225 ;
        RECT 79.360 149.485 79.815 150.250 ;
        RECT 80.290 150.075 80.510 150.475 ;
        RECT 80.755 150.475 81.085 150.685 ;
        RECT 80.755 150.075 80.965 150.475 ;
        RECT 81.255 150.440 81.665 150.745 ;
        RECT 81.895 150.305 82.065 150.880 ;
        RECT 81.795 150.185 82.065 150.305 ;
        RECT 81.220 150.140 82.065 150.185 ;
        RECT 81.220 150.015 81.975 150.140 ;
        RECT 81.220 149.865 81.390 150.015 ;
        RECT 82.235 149.995 82.405 151.185 ;
        RECT 82.175 149.985 82.405 149.995 ;
        RECT 80.090 149.655 81.390 149.865 ;
        RECT 81.645 149.485 81.975 149.845 ;
        RECT 82.145 149.655 82.405 149.985 ;
        RECT 82.575 150.430 82.855 151.865 ;
        RECT 83.025 151.260 83.735 152.035 ;
        RECT 83.905 151.090 84.235 151.865 ;
        RECT 83.085 150.875 84.235 151.090 ;
        RECT 82.575 149.655 82.915 150.430 ;
        RECT 83.085 150.305 83.370 150.875 ;
        RECT 83.555 150.475 84.025 150.705 ;
        RECT 84.430 150.675 84.645 151.790 ;
        RECT 84.825 151.315 85.155 152.035 ;
        RECT 84.935 150.675 85.165 151.015 ;
        RECT 85.335 150.945 87.005 152.035 ;
        RECT 84.195 150.495 84.645 150.675 ;
        RECT 84.195 150.475 84.525 150.495 ;
        RECT 84.835 150.475 85.165 150.675 ;
        RECT 83.085 150.115 83.795 150.305 ;
        RECT 83.495 149.975 83.795 150.115 ;
        RECT 83.985 150.115 85.165 150.305 ;
        RECT 83.985 150.035 84.315 150.115 ;
        RECT 83.495 149.965 83.810 149.975 ;
        RECT 83.495 149.955 83.820 149.965 ;
        RECT 83.495 149.950 83.830 149.955 ;
        RECT 83.085 149.485 83.255 149.945 ;
        RECT 83.495 149.940 83.835 149.950 ;
        RECT 83.495 149.935 83.840 149.940 ;
        RECT 83.495 149.925 83.845 149.935 ;
        RECT 83.495 149.920 83.850 149.925 ;
        RECT 83.495 149.655 83.855 149.920 ;
        RECT 84.485 149.485 84.655 149.945 ;
        RECT 84.825 149.655 85.165 150.115 ;
        RECT 85.335 150.255 86.085 150.775 ;
        RECT 86.255 150.425 87.005 150.945 ;
        RECT 87.175 150.870 87.465 152.035 ;
        RECT 87.675 151.695 88.815 151.865 ;
        RECT 87.675 151.235 87.975 151.695 ;
        RECT 88.145 151.065 88.475 151.525 ;
        RECT 87.715 150.845 88.475 151.065 ;
        RECT 88.645 151.065 88.815 151.695 ;
        RECT 88.985 151.235 89.315 152.035 ;
        RECT 89.485 151.065 89.760 151.865 ;
        RECT 88.645 150.855 89.760 151.065 ;
        RECT 90.395 151.165 90.670 151.865 ;
        RECT 90.880 151.490 91.095 152.035 ;
        RECT 91.265 151.525 91.740 151.865 ;
        RECT 91.910 151.530 92.525 152.035 ;
        RECT 91.910 151.355 92.105 151.530 ;
        RECT 87.715 150.305 87.930 150.845 ;
        RECT 88.100 150.475 88.870 150.675 ;
        RECT 89.040 150.475 89.760 150.675 ;
        RECT 85.335 149.485 87.005 150.255 ;
        RECT 87.175 149.485 87.465 150.210 ;
        RECT 87.715 150.135 89.315 150.305 ;
        RECT 88.145 150.125 89.315 150.135 ;
        RECT 87.685 149.485 87.975 149.955 ;
        RECT 88.145 149.655 88.475 150.125 ;
        RECT 88.645 149.485 88.815 149.955 ;
        RECT 88.985 149.655 89.315 150.125 ;
        RECT 89.485 149.485 89.760 150.305 ;
        RECT 90.395 150.135 90.565 151.165 ;
        RECT 90.840 150.995 91.555 151.290 ;
        RECT 91.775 151.165 92.105 151.355 ;
        RECT 92.275 150.995 92.525 151.360 ;
        RECT 90.735 150.825 92.525 150.995 ;
        RECT 90.735 150.395 90.965 150.825 ;
        RECT 90.395 149.655 90.655 150.135 ;
        RECT 91.135 150.125 91.545 150.645 ;
        RECT 90.825 149.485 91.155 149.945 ;
        RECT 91.345 149.705 91.545 150.125 ;
        RECT 91.715 149.970 91.970 150.825 ;
        RECT 92.765 150.645 92.935 151.865 ;
        RECT 93.185 151.525 93.445 152.035 ;
        RECT 92.140 150.395 92.935 150.645 ;
        RECT 93.105 150.475 93.445 151.355 ;
        RECT 93.615 150.895 93.945 152.035 ;
        RECT 94.115 151.405 94.470 151.865 ;
        RECT 94.640 151.575 95.215 152.035 ;
        RECT 95.385 151.405 95.715 151.865 ;
        RECT 94.115 151.235 95.715 151.405 ;
        RECT 95.915 151.235 96.170 152.035 ;
        RECT 97.035 151.365 97.315 152.035 ;
        RECT 94.115 150.895 94.390 151.235 ;
        RECT 94.570 151.015 94.760 151.055 ;
        RECT 94.570 150.845 94.765 151.015 ;
        RECT 94.570 150.675 94.760 150.845 ;
        RECT 93.615 150.475 94.760 150.675 ;
        RECT 92.685 150.305 92.935 150.395 ;
        RECT 94.940 150.335 95.220 151.235 ;
        RECT 96.340 151.065 96.640 151.260 ;
        RECT 97.485 151.145 97.785 151.695 ;
        RECT 97.985 151.315 98.315 152.035 ;
        RECT 98.505 151.315 98.965 151.865 ;
        RECT 95.390 150.895 96.640 151.065 ;
        RECT 95.390 150.475 95.720 150.895 ;
        RECT 95.950 150.395 96.295 150.725 ;
        RECT 94.940 150.305 95.225 150.335 ;
        RECT 91.715 149.705 92.505 149.970 ;
        RECT 92.685 149.885 93.015 150.305 ;
        RECT 93.185 149.485 93.445 150.305 ;
        RECT 93.615 150.095 94.725 150.305 ;
        RECT 93.615 149.655 93.965 150.095 ;
        RECT 94.135 149.485 94.305 149.925 ;
        RECT 94.475 149.865 94.725 150.095 ;
        RECT 94.895 150.035 95.225 150.305 ;
        RECT 95.395 149.865 95.670 150.305 ;
        RECT 96.470 150.240 96.640 150.895 ;
        RECT 96.850 150.725 97.115 151.085 ;
        RECT 97.485 150.975 98.425 151.145 ;
        RECT 98.255 150.725 98.425 150.975 ;
        RECT 96.850 150.475 97.525 150.725 ;
        RECT 97.745 150.475 98.085 150.725 ;
        RECT 98.255 150.395 98.545 150.725 ;
        RECT 98.255 150.305 98.425 150.395 ;
        RECT 94.475 149.655 95.670 149.865 ;
        RECT 95.905 149.485 96.235 150.225 ;
        RECT 96.405 149.910 96.640 150.240 ;
        RECT 97.035 150.115 98.425 150.305 ;
        RECT 97.035 149.755 97.365 150.115 ;
        RECT 98.715 149.945 98.965 151.315 ;
        RECT 99.225 151.365 99.395 151.865 ;
        RECT 99.565 151.535 99.895 152.035 ;
        RECT 99.225 151.195 99.890 151.365 ;
        RECT 99.140 150.375 99.490 151.025 ;
        RECT 99.660 150.205 99.890 151.195 ;
        RECT 97.985 149.485 98.235 149.945 ;
        RECT 98.405 149.655 98.965 149.945 ;
        RECT 99.225 150.035 99.890 150.205 ;
        RECT 99.225 149.745 99.395 150.035 ;
        RECT 99.565 149.485 99.895 149.865 ;
        RECT 100.065 149.745 100.250 151.865 ;
        RECT 100.490 151.575 100.755 152.035 ;
        RECT 100.925 151.440 101.175 151.865 ;
        RECT 101.385 151.590 102.490 151.760 ;
        RECT 100.870 151.310 101.175 151.440 ;
        RECT 100.420 150.115 100.700 151.065 ;
        RECT 100.870 150.205 101.040 151.310 ;
        RECT 101.210 150.525 101.450 151.120 ;
        RECT 101.620 151.055 102.150 151.420 ;
        RECT 101.620 150.355 101.790 151.055 ;
        RECT 102.320 150.975 102.490 151.590 ;
        RECT 102.660 151.235 102.830 152.035 ;
        RECT 103.000 151.535 103.250 151.865 ;
        RECT 103.475 151.565 104.360 151.735 ;
        RECT 102.320 150.885 102.830 150.975 ;
        RECT 100.870 150.075 101.095 150.205 ;
        RECT 101.265 150.135 101.790 150.355 ;
        RECT 101.960 150.715 102.830 150.885 ;
        RECT 100.505 149.485 100.755 149.945 ;
        RECT 100.925 149.935 101.095 150.075 ;
        RECT 101.960 149.935 102.130 150.715 ;
        RECT 102.660 150.645 102.830 150.715 ;
        RECT 102.340 150.465 102.540 150.495 ;
        RECT 103.000 150.465 103.170 151.535 ;
        RECT 103.340 150.645 103.530 151.365 ;
        RECT 102.340 150.165 103.170 150.465 ;
        RECT 103.700 150.435 104.020 151.395 ;
        RECT 100.925 149.765 101.260 149.935 ;
        RECT 101.455 149.765 102.130 149.935 ;
        RECT 102.450 149.485 102.820 149.985 ;
        RECT 103.000 149.935 103.170 150.165 ;
        RECT 103.555 150.105 104.020 150.435 ;
        RECT 104.190 150.725 104.360 151.565 ;
        RECT 104.540 151.535 104.855 152.035 ;
        RECT 105.085 151.305 105.425 151.865 ;
        RECT 104.530 150.930 105.425 151.305 ;
        RECT 105.595 151.025 105.765 152.035 ;
        RECT 105.235 150.725 105.425 150.930 ;
        RECT 105.935 150.975 106.265 151.820 ;
        RECT 105.935 150.895 106.325 150.975 ;
        RECT 106.110 150.845 106.325 150.895 ;
        RECT 104.190 150.395 105.065 150.725 ;
        RECT 105.235 150.395 105.985 150.725 ;
        RECT 104.190 149.935 104.360 150.395 ;
        RECT 105.235 150.225 105.435 150.395 ;
        RECT 106.155 150.265 106.325 150.845 ;
        RECT 106.100 150.225 106.325 150.265 ;
        RECT 103.000 149.765 103.405 149.935 ;
        RECT 103.575 149.765 104.360 149.935 ;
        RECT 104.635 149.485 104.845 150.015 ;
        RECT 105.105 149.700 105.435 150.225 ;
        RECT 105.945 150.140 106.325 150.225 ;
        RECT 106.500 150.895 106.835 151.865 ;
        RECT 107.005 150.895 107.175 152.035 ;
        RECT 107.345 151.695 109.375 151.865 ;
        RECT 106.500 150.225 106.670 150.895 ;
        RECT 107.345 150.725 107.515 151.695 ;
        RECT 106.840 150.395 107.095 150.725 ;
        RECT 107.320 150.395 107.515 150.725 ;
        RECT 107.685 151.355 108.810 151.525 ;
        RECT 106.925 150.225 107.095 150.395 ;
        RECT 107.685 150.225 107.855 151.355 ;
        RECT 105.605 149.485 105.775 150.095 ;
        RECT 105.945 149.705 106.275 150.140 ;
        RECT 106.500 149.655 106.755 150.225 ;
        RECT 106.925 150.055 107.855 150.225 ;
        RECT 108.025 151.015 109.035 151.185 ;
        RECT 108.025 150.215 108.195 151.015 ;
        RECT 108.400 150.335 108.675 150.815 ;
        RECT 108.395 150.165 108.675 150.335 ;
        RECT 107.680 150.020 107.855 150.055 ;
        RECT 106.925 149.485 107.255 149.885 ;
        RECT 107.680 149.655 108.210 150.020 ;
        RECT 108.400 149.655 108.675 150.165 ;
        RECT 108.845 149.655 109.035 151.015 ;
        RECT 109.205 151.030 109.375 151.695 ;
        RECT 109.545 151.275 109.715 152.035 ;
        RECT 109.950 151.275 110.465 151.685 ;
        RECT 109.205 150.840 109.955 151.030 ;
        RECT 110.125 150.465 110.465 151.275 ;
        RECT 109.235 150.295 110.465 150.465 ;
        RECT 110.635 151.315 111.095 151.865 ;
        RECT 111.285 151.315 111.615 152.035 ;
        RECT 109.215 149.485 109.725 150.020 ;
        RECT 109.945 149.690 110.190 150.295 ;
        RECT 110.635 149.945 110.885 151.315 ;
        RECT 111.815 151.145 112.115 151.695 ;
        RECT 112.285 151.365 112.565 152.035 ;
        RECT 111.175 150.975 112.115 151.145 ;
        RECT 111.175 150.725 111.345 150.975 ;
        RECT 112.485 150.725 112.750 151.085 ;
        RECT 112.935 150.870 113.225 152.035 ;
        RECT 113.865 151.225 114.160 152.035 ;
        RECT 114.340 150.725 114.585 151.865 ;
        RECT 114.760 151.225 115.020 152.035 ;
        RECT 115.620 152.030 121.895 152.035 ;
        RECT 115.200 150.725 115.450 151.860 ;
        RECT 115.620 151.235 115.880 152.030 ;
        RECT 116.050 151.135 116.310 151.860 ;
        RECT 116.480 151.305 116.740 152.030 ;
        RECT 116.910 151.135 117.170 151.860 ;
        RECT 117.340 151.305 117.600 152.030 ;
        RECT 117.770 151.135 118.030 151.860 ;
        RECT 118.200 151.305 118.460 152.030 ;
        RECT 118.630 151.135 118.890 151.860 ;
        RECT 119.060 151.305 119.305 152.030 ;
        RECT 119.475 151.135 119.735 151.860 ;
        RECT 119.920 151.305 120.165 152.030 ;
        RECT 120.335 151.135 120.595 151.860 ;
        RECT 120.780 151.305 121.025 152.030 ;
        RECT 121.195 151.135 121.455 151.860 ;
        RECT 121.640 151.305 121.895 152.030 ;
        RECT 116.050 151.120 121.455 151.135 ;
        RECT 122.065 151.120 122.355 151.860 ;
        RECT 122.525 151.290 122.795 152.035 ;
        RECT 116.050 150.895 122.795 151.120 ;
        RECT 111.055 150.395 111.345 150.725 ;
        RECT 111.515 150.475 111.855 150.725 ;
        RECT 112.075 150.475 112.750 150.725 ;
        RECT 111.175 150.305 111.345 150.395 ;
        RECT 111.175 150.115 112.565 150.305 ;
        RECT 110.635 149.655 111.195 149.945 ;
        RECT 111.365 149.485 111.615 149.945 ;
        RECT 112.235 149.755 112.565 150.115 ;
        RECT 112.935 149.485 113.225 150.210 ;
        RECT 113.855 150.165 114.170 150.725 ;
        RECT 114.340 150.475 121.460 150.725 ;
        RECT 113.855 149.485 114.160 149.995 ;
        RECT 114.340 149.665 114.590 150.475 ;
        RECT 114.760 149.485 115.020 150.010 ;
        RECT 115.200 149.665 115.450 150.475 ;
        RECT 121.630 150.305 122.795 150.895 ;
        RECT 116.050 150.135 122.795 150.305 ;
        RECT 123.060 150.895 123.395 151.865 ;
        RECT 123.565 150.895 123.735 152.035 ;
        RECT 123.905 151.695 125.935 151.865 ;
        RECT 123.060 150.225 123.230 150.895 ;
        RECT 123.905 150.725 124.075 151.695 ;
        RECT 123.400 150.395 123.655 150.725 ;
        RECT 123.880 150.395 124.075 150.725 ;
        RECT 124.245 151.355 125.370 151.525 ;
        RECT 123.485 150.225 123.655 150.395 ;
        RECT 124.245 150.225 124.415 151.355 ;
        RECT 115.620 149.485 115.880 150.045 ;
        RECT 116.050 149.680 116.310 150.135 ;
        RECT 116.480 149.485 116.740 149.965 ;
        RECT 116.910 149.680 117.170 150.135 ;
        RECT 117.340 149.485 117.600 149.965 ;
        RECT 117.770 149.680 118.030 150.135 ;
        RECT 118.200 149.485 118.445 149.965 ;
        RECT 118.615 149.680 118.890 150.135 ;
        RECT 119.060 149.485 119.305 149.965 ;
        RECT 119.475 149.680 119.735 150.135 ;
        RECT 119.915 149.485 120.165 149.965 ;
        RECT 120.335 149.680 120.595 150.135 ;
        RECT 120.775 149.485 121.025 149.965 ;
        RECT 121.195 149.680 121.455 150.135 ;
        RECT 121.635 149.485 121.895 149.965 ;
        RECT 122.065 149.680 122.325 150.135 ;
        RECT 122.495 149.485 122.795 149.965 ;
        RECT 123.060 149.655 123.315 150.225 ;
        RECT 123.485 150.055 124.415 150.225 ;
        RECT 124.585 151.015 125.595 151.185 ;
        RECT 124.585 150.215 124.755 151.015 ;
        RECT 124.240 150.020 124.415 150.055 ;
        RECT 123.485 149.485 123.815 149.885 ;
        RECT 124.240 149.655 124.770 150.020 ;
        RECT 124.960 149.995 125.235 150.815 ;
        RECT 124.955 149.825 125.235 149.995 ;
        RECT 124.960 149.655 125.235 149.825 ;
        RECT 125.405 149.655 125.595 151.015 ;
        RECT 125.765 151.030 125.935 151.695 ;
        RECT 126.105 151.275 126.275 152.035 ;
        RECT 126.510 151.275 127.025 151.685 ;
        RECT 125.765 150.840 126.515 151.030 ;
        RECT 126.685 150.465 127.025 151.275 ;
        RECT 127.195 150.945 129.785 152.035 ;
        RECT 125.795 150.295 127.025 150.465 ;
        RECT 125.775 149.485 126.285 150.020 ;
        RECT 126.505 149.690 126.750 150.295 ;
        RECT 127.195 150.255 128.405 150.775 ;
        RECT 128.575 150.425 129.785 150.945 ;
        RECT 130.415 150.430 130.695 151.865 ;
        RECT 130.865 151.260 131.575 152.035 ;
        RECT 131.745 151.090 132.075 151.865 ;
        RECT 130.925 150.875 132.075 151.090 ;
        RECT 127.195 149.485 129.785 150.255 ;
        RECT 130.415 149.655 130.755 150.430 ;
        RECT 130.925 150.305 131.210 150.875 ;
        RECT 131.395 150.475 131.865 150.705 ;
        RECT 132.270 150.675 132.485 151.790 ;
        RECT 132.665 151.315 132.995 152.035 ;
        RECT 132.775 150.675 133.005 151.015 ;
        RECT 133.695 150.895 133.905 152.035 ;
        RECT 132.035 150.495 132.485 150.675 ;
        RECT 132.035 150.475 132.365 150.495 ;
        RECT 132.675 150.475 133.005 150.675 ;
        RECT 134.075 150.885 134.405 151.865 ;
        RECT 134.575 150.895 134.805 152.035 ;
        RECT 135.075 150.895 135.285 152.035 ;
        RECT 135.455 150.885 135.785 151.865 ;
        RECT 135.955 150.895 136.185 152.035 ;
        RECT 136.395 151.480 137.000 152.035 ;
        RECT 137.175 151.525 137.655 151.865 ;
        RECT 137.825 151.490 138.080 152.035 ;
        RECT 136.395 151.380 137.010 151.480 ;
        RECT 136.825 151.355 137.010 151.380 ;
        RECT 130.925 150.115 131.635 150.305 ;
        RECT 131.335 149.975 131.635 150.115 ;
        RECT 131.825 150.115 133.005 150.305 ;
        RECT 131.825 150.035 132.155 150.115 ;
        RECT 131.335 149.965 131.650 149.975 ;
        RECT 131.335 149.955 131.660 149.965 ;
        RECT 131.335 149.950 131.670 149.955 ;
        RECT 130.925 149.485 131.095 149.945 ;
        RECT 131.335 149.940 131.675 149.950 ;
        RECT 131.335 149.935 131.680 149.940 ;
        RECT 131.335 149.925 131.685 149.935 ;
        RECT 131.335 149.920 131.690 149.925 ;
        RECT 131.335 149.655 131.695 149.920 ;
        RECT 132.325 149.485 132.495 149.945 ;
        RECT 132.665 149.655 133.005 150.115 ;
        RECT 133.695 149.485 133.905 150.305 ;
        RECT 134.075 150.285 134.325 150.885 ;
        RECT 134.495 150.475 134.825 150.725 ;
        RECT 134.075 149.655 134.405 150.285 ;
        RECT 134.575 149.485 134.805 150.305 ;
        RECT 135.075 149.485 135.285 150.305 ;
        RECT 135.455 150.285 135.705 150.885 ;
        RECT 136.395 150.760 136.655 151.210 ;
        RECT 136.825 151.110 137.155 151.355 ;
        RECT 137.325 151.035 138.080 151.285 ;
        RECT 138.250 151.165 138.525 151.865 ;
        RECT 137.310 151.000 138.080 151.035 ;
        RECT 137.295 150.990 138.080 151.000 ;
        RECT 137.290 150.975 138.185 150.990 ;
        RECT 137.270 150.960 138.185 150.975 ;
        RECT 137.250 150.950 138.185 150.960 ;
        RECT 137.225 150.940 138.185 150.950 ;
        RECT 137.155 150.910 138.185 150.940 ;
        RECT 137.135 150.880 138.185 150.910 ;
        RECT 137.115 150.850 138.185 150.880 ;
        RECT 137.085 150.825 138.185 150.850 ;
        RECT 137.050 150.790 138.185 150.825 ;
        RECT 137.020 150.785 138.185 150.790 ;
        RECT 137.020 150.780 137.410 150.785 ;
        RECT 137.020 150.770 137.385 150.780 ;
        RECT 137.020 150.765 137.370 150.770 ;
        RECT 137.020 150.760 137.355 150.765 ;
        RECT 136.395 150.755 137.355 150.760 ;
        RECT 136.395 150.745 137.345 150.755 ;
        RECT 136.395 150.740 137.335 150.745 ;
        RECT 136.395 150.730 137.325 150.740 ;
        RECT 135.875 150.475 136.205 150.725 ;
        RECT 136.395 150.720 137.320 150.730 ;
        RECT 136.395 150.715 137.315 150.720 ;
        RECT 136.395 150.700 137.305 150.715 ;
        RECT 136.395 150.685 137.300 150.700 ;
        RECT 136.395 150.660 137.290 150.685 ;
        RECT 136.395 150.590 137.285 150.660 ;
        RECT 135.455 149.655 135.785 150.285 ;
        RECT 135.955 149.485 136.185 150.305 ;
        RECT 136.395 150.035 136.945 150.420 ;
        RECT 137.115 149.865 137.285 150.590 ;
        RECT 136.395 149.695 137.285 149.865 ;
        RECT 137.455 150.190 137.785 150.615 ;
        RECT 137.955 150.390 138.185 150.785 ;
        RECT 137.455 150.165 137.705 150.190 ;
        RECT 137.455 149.705 137.675 150.165 ;
        RECT 138.355 150.135 138.525 151.165 ;
        RECT 138.695 150.870 138.985 152.035 ;
        RECT 137.845 149.485 138.095 150.025 ;
        RECT 138.265 149.655 138.525 150.135 ;
        RECT 138.695 149.485 138.985 150.210 ;
        RECT 139.165 149.665 139.425 151.855 ;
        RECT 139.595 151.305 139.935 152.035 ;
        RECT 140.115 151.125 140.385 151.855 ;
        RECT 139.615 150.905 140.385 151.125 ;
        RECT 140.565 151.145 140.795 151.855 ;
        RECT 140.965 151.325 141.295 152.035 ;
        RECT 141.465 151.145 141.725 151.855 ;
        RECT 142.375 151.525 142.675 152.035 ;
        RECT 142.845 151.355 143.175 151.865 ;
        RECT 143.345 151.525 143.975 152.035 ;
        RECT 144.555 151.525 144.935 151.695 ;
        RECT 145.105 151.525 145.405 152.035 ;
        RECT 144.765 151.355 144.935 151.525 ;
        RECT 140.565 150.905 141.725 151.145 ;
        RECT 142.375 151.185 144.595 151.355 ;
        RECT 139.615 150.235 139.905 150.905 ;
        RECT 140.085 150.415 140.550 150.725 ;
        RECT 140.730 150.415 141.255 150.725 ;
        RECT 139.615 150.035 140.845 150.235 ;
        RECT 139.685 149.485 140.355 149.855 ;
        RECT 140.535 149.665 140.845 150.035 ;
        RECT 141.025 149.775 141.255 150.415 ;
        RECT 141.435 150.395 141.735 150.725 ;
        RECT 142.375 150.225 142.545 151.185 ;
        RECT 142.715 150.845 144.255 151.015 ;
        RECT 142.715 150.395 142.960 150.845 ;
        RECT 143.220 150.475 143.915 150.675 ;
        RECT 144.085 150.645 144.255 150.845 ;
        RECT 144.425 150.985 144.595 151.185 ;
        RECT 144.765 151.155 145.425 151.355 ;
        RECT 144.425 150.815 145.085 150.985 ;
        RECT 144.085 150.475 144.685 150.645 ;
        RECT 144.915 150.395 145.085 150.815 ;
        RECT 141.435 149.485 141.725 150.215 ;
        RECT 142.375 149.680 142.840 150.225 ;
        RECT 143.345 149.485 143.515 150.305 ;
        RECT 143.685 150.225 144.595 150.305 ;
        RECT 145.255 150.225 145.425 151.155 ;
        RECT 145.595 150.895 145.875 152.035 ;
        RECT 146.045 150.885 146.375 151.865 ;
        RECT 146.545 150.895 146.805 152.035 ;
        RECT 147.035 150.975 147.365 151.820 ;
        RECT 147.535 151.025 147.705 152.035 ;
        RECT 147.875 151.305 148.215 151.865 ;
        RECT 148.445 151.535 148.760 152.035 ;
        RECT 148.940 151.565 149.825 151.735 ;
        RECT 146.975 150.895 147.365 150.975 ;
        RECT 147.875 150.930 148.770 151.305 ;
        RECT 145.605 150.455 145.940 150.725 ;
        RECT 146.110 150.285 146.280 150.885 ;
        RECT 146.975 150.845 147.190 150.895 ;
        RECT 146.450 150.475 146.785 150.725 ;
        RECT 143.685 150.135 144.935 150.225 ;
        RECT 143.685 149.655 144.015 150.135 ;
        RECT 144.425 150.055 144.935 150.135 ;
        RECT 144.185 149.485 144.535 149.875 ;
        RECT 144.705 149.655 144.935 150.055 ;
        RECT 145.105 149.745 145.425 150.225 ;
        RECT 145.595 149.485 145.905 150.285 ;
        RECT 146.110 149.655 146.805 150.285 ;
        RECT 146.975 150.265 147.145 150.845 ;
        RECT 147.875 150.725 148.065 150.930 ;
        RECT 148.940 150.725 149.110 151.565 ;
        RECT 150.050 151.535 150.300 151.865 ;
        RECT 147.315 150.395 148.065 150.725 ;
        RECT 148.235 150.395 149.110 150.725 ;
        RECT 146.975 150.225 147.200 150.265 ;
        RECT 147.865 150.225 148.065 150.395 ;
        RECT 146.975 150.140 147.355 150.225 ;
        RECT 147.025 149.705 147.355 150.140 ;
        RECT 147.525 149.485 147.695 150.095 ;
        RECT 147.865 149.700 148.195 150.225 ;
        RECT 148.455 149.485 148.665 150.015 ;
        RECT 148.940 149.935 149.110 150.395 ;
        RECT 149.280 150.435 149.600 151.395 ;
        RECT 149.770 150.645 149.960 151.365 ;
        RECT 150.130 150.465 150.300 151.535 ;
        RECT 150.470 151.235 150.640 152.035 ;
        RECT 150.810 151.590 151.915 151.760 ;
        RECT 150.810 150.975 150.980 151.590 ;
        RECT 152.125 151.440 152.375 151.865 ;
        RECT 152.545 151.575 152.810 152.035 ;
        RECT 151.150 151.055 151.680 151.420 ;
        RECT 152.125 151.310 152.430 151.440 ;
        RECT 150.470 150.885 150.980 150.975 ;
        RECT 150.470 150.715 151.340 150.885 ;
        RECT 150.470 150.645 150.640 150.715 ;
        RECT 150.760 150.465 150.960 150.495 ;
        RECT 149.280 150.105 149.745 150.435 ;
        RECT 150.130 150.165 150.960 150.465 ;
        RECT 150.130 149.935 150.300 150.165 ;
        RECT 148.940 149.765 149.725 149.935 ;
        RECT 149.895 149.765 150.300 149.935 ;
        RECT 150.480 149.485 150.850 149.985 ;
        RECT 151.170 149.935 151.340 150.715 ;
        RECT 151.510 150.355 151.680 151.055 ;
        RECT 151.850 150.525 152.090 151.120 ;
        RECT 151.510 150.135 152.035 150.355 ;
        RECT 152.260 150.205 152.430 151.310 ;
        RECT 152.205 150.075 152.430 150.205 ;
        RECT 152.600 150.115 152.880 151.065 ;
        RECT 152.205 149.935 152.375 150.075 ;
        RECT 151.170 149.765 151.845 149.935 ;
        RECT 152.040 149.765 152.375 149.935 ;
        RECT 152.545 149.485 152.795 149.945 ;
        RECT 153.050 149.745 153.235 151.865 ;
        RECT 153.405 151.535 153.735 152.035 ;
        RECT 153.905 151.365 154.075 151.865 ;
        RECT 153.410 151.195 154.075 151.365 ;
        RECT 153.410 150.205 153.640 151.195 ;
        RECT 153.810 150.375 154.160 151.025 ;
        RECT 154.335 150.945 155.545 152.035 ;
        RECT 154.335 150.235 154.855 150.775 ;
        RECT 155.025 150.405 155.545 150.945 ;
        RECT 155.715 150.945 156.925 152.035 ;
        RECT 155.715 150.405 156.235 150.945 ;
        RECT 156.405 150.235 156.925 150.775 ;
        RECT 153.410 150.035 154.075 150.205 ;
        RECT 153.405 149.485 153.735 149.865 ;
        RECT 153.905 149.745 154.075 150.035 ;
        RECT 154.335 149.485 155.545 150.235 ;
        RECT 155.715 149.485 156.925 150.235 ;
        RECT 22.690 149.315 157.010 149.485 ;
        RECT 22.775 148.565 23.985 149.315 ;
        RECT 25.080 148.810 25.415 149.315 ;
        RECT 25.585 148.745 25.825 149.120 ;
        RECT 26.105 148.985 26.275 149.130 ;
        RECT 26.105 148.790 26.480 148.985 ;
        RECT 26.840 148.820 27.235 149.315 ;
        RECT 22.775 148.025 23.295 148.565 ;
        RECT 23.465 147.855 23.985 148.395 ;
        RECT 22.775 146.765 23.985 147.855 ;
        RECT 25.135 147.785 25.435 148.635 ;
        RECT 25.605 148.595 25.825 148.745 ;
        RECT 25.605 148.265 26.140 148.595 ;
        RECT 26.310 148.455 26.480 148.790 ;
        RECT 27.405 148.625 27.645 149.145 ;
        RECT 25.605 147.615 25.840 148.265 ;
        RECT 26.310 148.095 27.295 148.455 ;
        RECT 25.165 147.385 25.840 147.615 ;
        RECT 26.010 148.075 27.295 148.095 ;
        RECT 26.010 147.925 26.870 148.075 ;
        RECT 25.165 146.955 25.335 147.385 ;
        RECT 25.505 146.765 25.835 147.215 ;
        RECT 26.010 146.980 26.295 147.925 ;
        RECT 27.470 147.820 27.645 148.625 ;
        RECT 27.835 148.545 29.505 149.315 ;
        RECT 29.675 148.855 30.235 149.145 ;
        RECT 30.405 148.855 30.655 149.315 ;
        RECT 27.835 148.025 28.585 148.545 ;
        RECT 28.755 147.855 29.505 148.375 ;
        RECT 26.470 147.445 27.165 147.755 ;
        RECT 26.475 146.765 27.160 147.235 ;
        RECT 27.340 147.035 27.645 147.820 ;
        RECT 27.835 146.765 29.505 147.855 ;
        RECT 29.675 147.485 29.925 148.855 ;
        RECT 31.275 148.685 31.605 149.045 ;
        RECT 30.215 148.495 31.605 148.685 ;
        RECT 32.065 148.765 32.235 149.055 ;
        RECT 32.405 148.935 32.735 149.315 ;
        RECT 32.065 148.595 32.730 148.765 ;
        RECT 30.215 148.405 30.385 148.495 ;
        RECT 30.095 148.075 30.385 148.405 ;
        RECT 30.555 148.075 30.895 148.325 ;
        RECT 31.115 148.075 31.790 148.325 ;
        RECT 30.215 147.825 30.385 148.075 ;
        RECT 30.215 147.655 31.155 147.825 ;
        RECT 31.525 147.715 31.790 148.075 ;
        RECT 31.980 147.775 32.330 148.425 ;
        RECT 29.675 146.935 30.135 147.485 ;
        RECT 30.325 146.765 30.655 147.485 ;
        RECT 30.855 147.105 31.155 147.655 ;
        RECT 32.500 147.605 32.730 148.595 ;
        RECT 32.065 147.435 32.730 147.605 ;
        RECT 31.325 146.765 31.605 147.435 ;
        RECT 32.065 146.935 32.235 147.435 ;
        RECT 32.405 146.765 32.735 147.265 ;
        RECT 32.905 146.935 33.090 149.055 ;
        RECT 33.345 148.855 33.595 149.315 ;
        RECT 33.765 148.865 34.100 149.035 ;
        RECT 34.295 148.865 34.970 149.035 ;
        RECT 33.765 148.725 33.935 148.865 ;
        RECT 33.260 147.735 33.540 148.685 ;
        RECT 33.710 148.595 33.935 148.725 ;
        RECT 33.710 147.490 33.880 148.595 ;
        RECT 34.105 148.445 34.630 148.665 ;
        RECT 34.050 147.680 34.290 148.275 ;
        RECT 34.460 147.745 34.630 148.445 ;
        RECT 34.800 148.085 34.970 148.865 ;
        RECT 35.290 148.815 35.660 149.315 ;
        RECT 35.840 148.865 36.245 149.035 ;
        RECT 36.415 148.865 37.200 149.035 ;
        RECT 35.840 148.635 36.010 148.865 ;
        RECT 35.180 148.335 36.010 148.635 ;
        RECT 36.395 148.365 36.860 148.695 ;
        RECT 35.180 148.305 35.380 148.335 ;
        RECT 35.500 148.085 35.670 148.155 ;
        RECT 34.800 147.915 35.670 148.085 ;
        RECT 35.160 147.825 35.670 147.915 ;
        RECT 33.710 147.360 34.015 147.490 ;
        RECT 34.460 147.380 34.990 147.745 ;
        RECT 33.330 146.765 33.595 147.225 ;
        RECT 33.765 146.935 34.015 147.360 ;
        RECT 35.160 147.210 35.330 147.825 ;
        RECT 34.225 147.040 35.330 147.210 ;
        RECT 35.500 146.765 35.670 147.565 ;
        RECT 35.840 147.265 36.010 148.335 ;
        RECT 36.180 147.435 36.370 148.155 ;
        RECT 36.540 147.405 36.860 148.365 ;
        RECT 37.030 148.405 37.200 148.865 ;
        RECT 37.475 148.785 37.685 149.315 ;
        RECT 37.945 148.575 38.275 149.100 ;
        RECT 38.445 148.705 38.615 149.315 ;
        RECT 38.785 148.660 39.115 149.095 ;
        RECT 39.885 148.765 40.055 149.055 ;
        RECT 40.225 148.935 40.555 149.315 ;
        RECT 38.785 148.575 39.165 148.660 ;
        RECT 39.885 148.595 40.550 148.765 ;
        RECT 38.075 148.405 38.275 148.575 ;
        RECT 38.940 148.535 39.165 148.575 ;
        RECT 37.030 148.075 37.905 148.405 ;
        RECT 38.075 148.075 38.825 148.405 ;
        RECT 35.840 146.935 36.090 147.265 ;
        RECT 37.030 147.235 37.200 148.075 ;
        RECT 38.075 147.870 38.265 148.075 ;
        RECT 38.995 147.955 39.165 148.535 ;
        RECT 38.950 147.905 39.165 147.955 ;
        RECT 37.370 147.495 38.265 147.870 ;
        RECT 38.775 147.825 39.165 147.905 ;
        RECT 36.315 147.065 37.200 147.235 ;
        RECT 37.380 146.765 37.695 147.265 ;
        RECT 37.925 146.935 38.265 147.495 ;
        RECT 38.435 146.765 38.605 147.775 ;
        RECT 38.775 146.980 39.105 147.825 ;
        RECT 39.800 147.775 40.150 148.425 ;
        RECT 40.320 147.605 40.550 148.595 ;
        RECT 39.885 147.435 40.550 147.605 ;
        RECT 39.885 146.935 40.055 147.435 ;
        RECT 40.225 146.765 40.555 147.265 ;
        RECT 40.725 146.935 40.910 149.055 ;
        RECT 41.165 148.855 41.415 149.315 ;
        RECT 41.585 148.865 41.920 149.035 ;
        RECT 42.115 148.865 42.790 149.035 ;
        RECT 41.585 148.725 41.755 148.865 ;
        RECT 41.080 147.735 41.360 148.685 ;
        RECT 41.530 148.595 41.755 148.725 ;
        RECT 41.530 147.490 41.700 148.595 ;
        RECT 41.925 148.445 42.450 148.665 ;
        RECT 41.870 147.680 42.110 148.275 ;
        RECT 42.280 147.745 42.450 148.445 ;
        RECT 42.620 148.085 42.790 148.865 ;
        RECT 43.110 148.815 43.480 149.315 ;
        RECT 43.660 148.865 44.065 149.035 ;
        RECT 44.235 148.865 45.020 149.035 ;
        RECT 43.660 148.635 43.830 148.865 ;
        RECT 43.000 148.335 43.830 148.635 ;
        RECT 44.215 148.365 44.680 148.695 ;
        RECT 43.000 148.305 43.200 148.335 ;
        RECT 43.320 148.085 43.490 148.155 ;
        RECT 42.620 147.915 43.490 148.085 ;
        RECT 42.980 147.825 43.490 147.915 ;
        RECT 41.530 147.360 41.835 147.490 ;
        RECT 42.280 147.380 42.810 147.745 ;
        RECT 41.150 146.765 41.415 147.225 ;
        RECT 41.585 146.935 41.835 147.360 ;
        RECT 42.980 147.210 43.150 147.825 ;
        RECT 42.045 147.040 43.150 147.210 ;
        RECT 43.320 146.765 43.490 147.565 ;
        RECT 43.660 147.265 43.830 148.335 ;
        RECT 44.000 147.435 44.190 148.155 ;
        RECT 44.360 147.405 44.680 148.365 ;
        RECT 44.850 148.405 45.020 148.865 ;
        RECT 45.295 148.785 45.505 149.315 ;
        RECT 45.765 148.575 46.095 149.100 ;
        RECT 46.265 148.705 46.435 149.315 ;
        RECT 46.605 148.660 46.935 149.095 ;
        RECT 46.605 148.575 46.985 148.660 ;
        RECT 45.895 148.405 46.095 148.575 ;
        RECT 46.760 148.535 46.985 148.575 ;
        RECT 44.850 148.075 45.725 148.405 ;
        RECT 45.895 148.075 46.645 148.405 ;
        RECT 43.660 146.935 43.910 147.265 ;
        RECT 44.850 147.235 45.020 148.075 ;
        RECT 45.895 147.870 46.085 148.075 ;
        RECT 46.815 147.955 46.985 148.535 ;
        RECT 47.155 148.515 47.850 149.145 ;
        RECT 48.055 148.515 48.365 149.315 ;
        RECT 48.535 148.590 48.825 149.315 ;
        RECT 48.995 148.545 50.665 149.315 ;
        RECT 50.925 148.765 51.095 149.055 ;
        RECT 51.265 148.935 51.595 149.315 ;
        RECT 50.925 148.595 51.590 148.765 ;
        RECT 47.175 148.075 47.510 148.325 ;
        RECT 46.770 147.905 46.985 147.955 ;
        RECT 47.680 147.915 47.850 148.515 ;
        RECT 48.020 148.075 48.355 148.345 ;
        RECT 48.995 148.025 49.745 148.545 ;
        RECT 45.190 147.495 46.085 147.870 ;
        RECT 46.595 147.825 46.985 147.905 ;
        RECT 44.135 147.065 45.020 147.235 ;
        RECT 45.200 146.765 45.515 147.265 ;
        RECT 45.745 146.935 46.085 147.495 ;
        RECT 46.255 146.765 46.425 147.775 ;
        RECT 46.595 146.980 46.925 147.825 ;
        RECT 47.155 146.765 47.415 147.905 ;
        RECT 47.585 146.935 47.915 147.915 ;
        RECT 48.085 146.765 48.365 147.905 ;
        RECT 48.535 146.765 48.825 147.930 ;
        RECT 49.915 147.855 50.665 148.375 ;
        RECT 48.995 146.765 50.665 147.855 ;
        RECT 50.840 147.775 51.190 148.425 ;
        RECT 51.360 147.605 51.590 148.595 ;
        RECT 50.925 147.435 51.590 147.605 ;
        RECT 50.925 146.935 51.095 147.435 ;
        RECT 51.265 146.765 51.595 147.265 ;
        RECT 51.765 146.935 51.950 149.055 ;
        RECT 52.205 148.855 52.455 149.315 ;
        RECT 52.625 148.865 52.960 149.035 ;
        RECT 53.155 148.865 53.830 149.035 ;
        RECT 52.625 148.725 52.795 148.865 ;
        RECT 52.120 147.735 52.400 148.685 ;
        RECT 52.570 148.595 52.795 148.725 ;
        RECT 52.570 147.490 52.740 148.595 ;
        RECT 52.965 148.445 53.490 148.665 ;
        RECT 52.910 147.680 53.150 148.275 ;
        RECT 53.320 147.745 53.490 148.445 ;
        RECT 53.660 148.085 53.830 148.865 ;
        RECT 54.150 148.815 54.520 149.315 ;
        RECT 54.700 148.865 55.105 149.035 ;
        RECT 55.275 148.865 56.060 149.035 ;
        RECT 54.700 148.635 54.870 148.865 ;
        RECT 54.040 148.335 54.870 148.635 ;
        RECT 55.255 148.365 55.720 148.695 ;
        RECT 54.040 148.305 54.240 148.335 ;
        RECT 54.360 148.085 54.530 148.155 ;
        RECT 53.660 147.915 54.530 148.085 ;
        RECT 54.020 147.825 54.530 147.915 ;
        RECT 52.570 147.360 52.875 147.490 ;
        RECT 53.320 147.380 53.850 147.745 ;
        RECT 52.190 146.765 52.455 147.225 ;
        RECT 52.625 146.935 52.875 147.360 ;
        RECT 54.020 147.210 54.190 147.825 ;
        RECT 53.085 147.040 54.190 147.210 ;
        RECT 54.360 146.765 54.530 147.565 ;
        RECT 54.700 147.265 54.870 148.335 ;
        RECT 55.040 147.435 55.230 148.155 ;
        RECT 55.400 147.405 55.720 148.365 ;
        RECT 55.890 148.405 56.060 148.865 ;
        RECT 56.335 148.785 56.545 149.315 ;
        RECT 56.805 148.575 57.135 149.100 ;
        RECT 57.305 148.705 57.475 149.315 ;
        RECT 57.645 148.660 57.975 149.095 ;
        RECT 57.645 148.575 58.025 148.660 ;
        RECT 56.935 148.405 57.135 148.575 ;
        RECT 57.800 148.535 58.025 148.575 ;
        RECT 55.890 148.075 56.765 148.405 ;
        RECT 56.935 148.075 57.685 148.405 ;
        RECT 54.700 146.935 54.950 147.265 ;
        RECT 55.890 147.235 56.060 148.075 ;
        RECT 56.935 147.870 57.125 148.075 ;
        RECT 57.855 147.955 58.025 148.535 ;
        RECT 57.810 147.905 58.025 147.955 ;
        RECT 56.230 147.495 57.125 147.870 ;
        RECT 57.635 147.825 58.025 147.905 ;
        RECT 59.115 148.595 59.455 149.105 ;
        RECT 55.175 147.065 56.060 147.235 ;
        RECT 56.240 146.765 56.555 147.265 ;
        RECT 56.785 146.935 57.125 147.495 ;
        RECT 57.295 146.765 57.465 147.775 ;
        RECT 57.635 146.980 57.965 147.825 ;
        RECT 59.115 147.195 59.375 148.595 ;
        RECT 59.625 148.515 59.895 149.315 ;
        RECT 59.550 148.075 59.880 148.325 ;
        RECT 60.075 148.075 60.355 149.045 ;
        RECT 60.535 148.075 60.835 149.045 ;
        RECT 61.015 148.075 61.365 149.040 ;
        RECT 61.585 148.815 62.080 149.145 ;
        RECT 62.340 148.825 62.595 149.315 ;
        RECT 59.565 147.905 59.880 148.075 ;
        RECT 61.585 147.905 61.755 148.815 ;
        RECT 62.765 148.805 63.995 149.145 ;
        RECT 59.565 147.735 61.755 147.905 ;
        RECT 59.115 146.935 59.455 147.195 ;
        RECT 59.625 146.765 59.955 147.565 ;
        RECT 60.420 146.935 60.670 147.735 ;
        RECT 60.855 146.765 61.185 147.485 ;
        RECT 61.405 146.935 61.655 147.735 ;
        RECT 61.925 147.325 62.165 148.635 ;
        RECT 62.360 148.075 62.580 148.655 ;
        RECT 62.765 147.905 62.945 148.805 ;
        RECT 63.115 148.075 63.490 148.635 ;
        RECT 63.665 148.575 63.995 148.805 ;
        RECT 64.225 148.660 64.555 149.095 ;
        RECT 64.725 148.705 64.895 149.315 ;
        RECT 64.175 148.575 64.555 148.660 ;
        RECT 65.065 148.575 65.395 149.100 ;
        RECT 65.655 148.785 65.865 149.315 ;
        RECT 66.140 148.865 66.925 149.035 ;
        RECT 67.095 148.865 67.500 149.035 ;
        RECT 64.175 148.535 64.400 148.575 ;
        RECT 63.695 148.075 64.005 148.405 ;
        RECT 64.175 147.955 64.345 148.535 ;
        RECT 65.065 148.405 65.265 148.575 ;
        RECT 66.140 148.405 66.310 148.865 ;
        RECT 64.515 148.075 65.265 148.405 ;
        RECT 65.435 148.075 66.310 148.405 ;
        RECT 64.175 147.905 64.390 147.955 ;
        RECT 61.825 146.765 62.160 147.145 ;
        RECT 62.340 146.765 62.595 147.905 ;
        RECT 62.765 147.735 63.995 147.905 ;
        RECT 64.175 147.825 64.565 147.905 ;
        RECT 62.765 146.935 63.095 147.735 ;
        RECT 63.265 146.765 63.495 147.565 ;
        RECT 63.665 146.935 63.995 147.735 ;
        RECT 64.235 146.980 64.565 147.825 ;
        RECT 65.075 147.870 65.265 148.075 ;
        RECT 64.735 146.765 64.905 147.775 ;
        RECT 65.075 147.495 65.970 147.870 ;
        RECT 65.075 146.935 65.415 147.495 ;
        RECT 65.645 146.765 65.960 147.265 ;
        RECT 66.140 147.235 66.310 148.075 ;
        RECT 66.480 148.365 66.945 148.695 ;
        RECT 67.330 148.635 67.500 148.865 ;
        RECT 67.680 148.815 68.050 149.315 ;
        RECT 68.370 148.865 69.045 149.035 ;
        RECT 69.240 148.865 69.575 149.035 ;
        RECT 66.480 147.405 66.800 148.365 ;
        RECT 67.330 148.335 68.160 148.635 ;
        RECT 66.970 147.435 67.160 148.155 ;
        RECT 67.330 147.265 67.500 148.335 ;
        RECT 67.960 148.305 68.160 148.335 ;
        RECT 67.670 148.085 67.840 148.155 ;
        RECT 68.370 148.085 68.540 148.865 ;
        RECT 69.405 148.725 69.575 148.865 ;
        RECT 69.745 148.855 69.995 149.315 ;
        RECT 67.670 147.915 68.540 148.085 ;
        RECT 68.710 148.445 69.235 148.665 ;
        RECT 69.405 148.595 69.630 148.725 ;
        RECT 67.670 147.825 68.180 147.915 ;
        RECT 66.140 147.065 67.025 147.235 ;
        RECT 67.250 146.935 67.500 147.265 ;
        RECT 67.670 146.765 67.840 147.565 ;
        RECT 68.010 147.210 68.180 147.825 ;
        RECT 68.710 147.745 68.880 148.445 ;
        RECT 68.350 147.380 68.880 147.745 ;
        RECT 69.050 147.680 69.290 148.275 ;
        RECT 69.460 147.490 69.630 148.595 ;
        RECT 69.800 147.735 70.080 148.685 ;
        RECT 69.325 147.360 69.630 147.490 ;
        RECT 68.010 147.040 69.115 147.210 ;
        RECT 69.325 146.935 69.575 147.360 ;
        RECT 69.745 146.765 70.010 147.225 ;
        RECT 70.250 146.935 70.435 149.055 ;
        RECT 70.605 148.935 70.935 149.315 ;
        RECT 71.105 148.765 71.275 149.055 ;
        RECT 70.610 148.595 71.275 148.765 ;
        RECT 71.535 148.640 71.795 149.145 ;
        RECT 71.975 148.935 72.305 149.315 ;
        RECT 72.485 148.765 72.655 149.145 ;
        RECT 70.610 147.605 70.840 148.595 ;
        RECT 71.010 147.775 71.360 148.425 ;
        RECT 71.535 147.840 71.705 148.640 ;
        RECT 71.990 148.595 72.655 148.765 ;
        RECT 71.990 148.340 72.160 148.595 ;
        RECT 72.915 148.565 74.125 149.315 ;
        RECT 74.295 148.590 74.585 149.315 ;
        RECT 75.265 148.660 75.595 149.095 ;
        RECT 75.765 148.705 75.935 149.315 ;
        RECT 75.215 148.575 75.595 148.660 ;
        RECT 76.105 148.575 76.435 149.100 ;
        RECT 76.695 148.785 76.905 149.315 ;
        RECT 77.180 148.865 77.965 149.035 ;
        RECT 78.135 148.865 78.540 149.035 ;
        RECT 71.875 148.010 72.160 148.340 ;
        RECT 72.395 148.045 72.725 148.415 ;
        RECT 72.915 148.025 73.435 148.565 ;
        RECT 75.215 148.535 75.440 148.575 ;
        RECT 71.990 147.865 72.160 148.010 ;
        RECT 70.610 147.435 71.275 147.605 ;
        RECT 70.605 146.765 70.935 147.265 ;
        RECT 71.105 146.935 71.275 147.435 ;
        RECT 71.535 146.935 71.805 147.840 ;
        RECT 71.990 147.695 72.655 147.865 ;
        RECT 73.605 147.855 74.125 148.395 ;
        RECT 75.215 147.955 75.385 148.535 ;
        RECT 76.105 148.405 76.305 148.575 ;
        RECT 77.180 148.405 77.350 148.865 ;
        RECT 75.555 148.075 76.305 148.405 ;
        RECT 76.475 148.075 77.350 148.405 ;
        RECT 71.975 146.765 72.305 147.525 ;
        RECT 72.485 146.935 72.655 147.695 ;
        RECT 72.915 146.765 74.125 147.855 ;
        RECT 74.295 146.765 74.585 147.930 ;
        RECT 75.215 147.905 75.430 147.955 ;
        RECT 75.215 147.825 75.605 147.905 ;
        RECT 75.275 146.980 75.605 147.825 ;
        RECT 76.115 147.870 76.305 148.075 ;
        RECT 75.775 146.765 75.945 147.775 ;
        RECT 76.115 147.495 77.010 147.870 ;
        RECT 76.115 146.935 76.455 147.495 ;
        RECT 76.685 146.765 77.000 147.265 ;
        RECT 77.180 147.235 77.350 148.075 ;
        RECT 77.520 148.365 77.985 148.695 ;
        RECT 78.370 148.635 78.540 148.865 ;
        RECT 78.720 148.815 79.090 149.315 ;
        RECT 79.410 148.865 80.085 149.035 ;
        RECT 80.280 148.865 80.615 149.035 ;
        RECT 77.520 147.405 77.840 148.365 ;
        RECT 78.370 148.335 79.200 148.635 ;
        RECT 78.010 147.435 78.200 148.155 ;
        RECT 78.370 147.265 78.540 148.335 ;
        RECT 79.000 148.305 79.200 148.335 ;
        RECT 78.710 148.085 78.880 148.155 ;
        RECT 79.410 148.085 79.580 148.865 ;
        RECT 80.445 148.725 80.615 148.865 ;
        RECT 80.785 148.855 81.035 149.315 ;
        RECT 78.710 147.915 79.580 148.085 ;
        RECT 79.750 148.445 80.275 148.665 ;
        RECT 80.445 148.595 80.670 148.725 ;
        RECT 78.710 147.825 79.220 147.915 ;
        RECT 77.180 147.065 78.065 147.235 ;
        RECT 78.290 146.935 78.540 147.265 ;
        RECT 78.710 146.765 78.880 147.565 ;
        RECT 79.050 147.210 79.220 147.825 ;
        RECT 79.750 147.745 79.920 148.445 ;
        RECT 79.390 147.380 79.920 147.745 ;
        RECT 80.090 147.680 80.330 148.275 ;
        RECT 80.500 147.490 80.670 148.595 ;
        RECT 80.840 147.735 81.120 148.685 ;
        RECT 80.365 147.360 80.670 147.490 ;
        RECT 79.050 147.040 80.155 147.210 ;
        RECT 80.365 146.935 80.615 147.360 ;
        RECT 80.785 146.765 81.050 147.225 ;
        RECT 81.290 146.935 81.475 149.055 ;
        RECT 81.645 148.935 81.975 149.315 ;
        RECT 82.145 148.765 82.315 149.055 ;
        RECT 81.650 148.595 82.315 148.765 ;
        RECT 81.650 147.605 81.880 148.595 ;
        RECT 82.615 148.495 82.845 149.315 ;
        RECT 83.015 148.515 83.345 149.145 ;
        RECT 82.050 147.775 82.400 148.425 ;
        RECT 82.595 148.075 82.925 148.325 ;
        RECT 83.095 147.915 83.345 148.515 ;
        RECT 83.515 148.495 83.725 149.315 ;
        RECT 83.955 148.545 87.465 149.315 ;
        RECT 88.755 148.685 89.085 149.045 ;
        RECT 89.705 148.855 89.955 149.315 ;
        RECT 90.125 148.855 90.685 149.145 ;
        RECT 83.955 148.025 85.605 148.545 ;
        RECT 88.755 148.495 90.145 148.685 ;
        RECT 89.975 148.405 90.145 148.495 ;
        RECT 81.650 147.435 82.315 147.605 ;
        RECT 81.645 146.765 81.975 147.265 ;
        RECT 82.145 146.935 82.315 147.435 ;
        RECT 82.615 146.765 82.845 147.905 ;
        RECT 83.015 146.935 83.345 147.915 ;
        RECT 83.515 146.765 83.725 147.905 ;
        RECT 85.775 147.855 87.465 148.375 ;
        RECT 83.955 146.765 87.465 147.855 ;
        RECT 88.570 148.075 89.245 148.325 ;
        RECT 89.465 148.075 89.805 148.325 ;
        RECT 89.975 148.075 90.265 148.405 ;
        RECT 88.570 147.715 88.835 148.075 ;
        RECT 89.975 147.825 90.145 148.075 ;
        RECT 89.205 147.655 90.145 147.825 ;
        RECT 88.755 146.765 89.035 147.435 ;
        RECT 89.205 147.105 89.505 147.655 ;
        RECT 90.435 147.485 90.685 148.855 ;
        RECT 89.705 146.765 90.035 147.485 ;
        RECT 90.225 146.935 90.685 147.485 ;
        RECT 90.860 148.575 91.115 149.145 ;
        RECT 91.285 148.915 91.615 149.315 ;
        RECT 92.040 148.780 92.570 149.145 ;
        RECT 92.040 148.745 92.215 148.780 ;
        RECT 91.285 148.575 92.215 148.745 ;
        RECT 92.760 148.635 93.035 149.145 ;
        RECT 90.860 147.905 91.030 148.575 ;
        RECT 91.285 148.405 91.455 148.575 ;
        RECT 91.200 148.075 91.455 148.405 ;
        RECT 91.680 148.075 91.875 148.405 ;
        RECT 90.860 146.935 91.195 147.905 ;
        RECT 91.365 146.765 91.535 147.905 ;
        RECT 91.705 147.105 91.875 148.075 ;
        RECT 92.045 147.445 92.215 148.575 ;
        RECT 92.385 147.785 92.555 148.585 ;
        RECT 92.755 148.465 93.035 148.635 ;
        RECT 92.760 147.985 93.035 148.465 ;
        RECT 93.205 147.785 93.395 149.145 ;
        RECT 93.575 148.780 94.085 149.315 ;
        RECT 94.305 148.505 94.550 149.110 ;
        RECT 94.995 148.545 98.505 149.315 ;
        RECT 98.675 148.565 99.885 149.315 ;
        RECT 100.055 148.590 100.345 149.315 ;
        RECT 100.520 148.575 100.775 149.145 ;
        RECT 100.945 148.915 101.275 149.315 ;
        RECT 101.700 148.780 102.230 149.145 ;
        RECT 101.700 148.745 101.875 148.780 ;
        RECT 100.945 148.575 101.875 148.745 ;
        RECT 93.595 148.335 94.825 148.505 ;
        RECT 92.385 147.615 93.395 147.785 ;
        RECT 93.565 147.770 94.315 147.960 ;
        RECT 92.045 147.275 93.170 147.445 ;
        RECT 93.565 147.105 93.735 147.770 ;
        RECT 94.485 147.525 94.825 148.335 ;
        RECT 94.995 148.025 96.645 148.545 ;
        RECT 96.815 147.855 98.505 148.375 ;
        RECT 98.675 148.025 99.195 148.565 ;
        RECT 99.365 147.855 99.885 148.395 ;
        RECT 91.705 146.935 93.735 147.105 ;
        RECT 93.905 146.765 94.075 147.525 ;
        RECT 94.310 147.115 94.825 147.525 ;
        RECT 94.995 146.765 98.505 147.855 ;
        RECT 98.675 146.765 99.885 147.855 ;
        RECT 100.055 146.765 100.345 147.930 ;
        RECT 100.520 147.905 100.690 148.575 ;
        RECT 100.945 148.405 101.115 148.575 ;
        RECT 100.860 148.075 101.115 148.405 ;
        RECT 101.340 148.075 101.535 148.405 ;
        RECT 100.520 146.935 100.855 147.905 ;
        RECT 101.025 146.765 101.195 147.905 ;
        RECT 101.365 147.105 101.535 148.075 ;
        RECT 101.705 147.445 101.875 148.575 ;
        RECT 102.045 147.785 102.215 148.585 ;
        RECT 102.420 148.295 102.695 149.145 ;
        RECT 102.415 148.125 102.695 148.295 ;
        RECT 102.420 147.985 102.695 148.125 ;
        RECT 102.865 147.785 103.055 149.145 ;
        RECT 103.235 148.780 103.745 149.315 ;
        RECT 103.965 148.505 104.210 149.110 ;
        RECT 105.205 148.765 105.375 149.145 ;
        RECT 105.555 148.935 105.885 149.315 ;
        RECT 105.205 148.595 105.870 148.765 ;
        RECT 106.065 148.640 106.325 149.145 ;
        RECT 103.255 148.335 104.485 148.505 ;
        RECT 102.045 147.615 103.055 147.785 ;
        RECT 103.225 147.770 103.975 147.960 ;
        RECT 101.705 147.275 102.830 147.445 ;
        RECT 103.225 147.105 103.395 147.770 ;
        RECT 104.145 147.525 104.485 148.335 ;
        RECT 105.135 148.045 105.465 148.415 ;
        RECT 105.700 148.340 105.870 148.595 ;
        RECT 105.700 148.010 105.985 148.340 ;
        RECT 105.700 147.865 105.870 148.010 ;
        RECT 101.365 146.935 103.395 147.105 ;
        RECT 103.565 146.765 103.735 147.525 ;
        RECT 103.970 147.115 104.485 147.525 ;
        RECT 105.205 147.695 105.870 147.865 ;
        RECT 106.155 147.840 106.325 148.640 ;
        RECT 106.585 148.765 106.755 149.055 ;
        RECT 106.925 148.935 107.255 149.315 ;
        RECT 106.585 148.595 107.250 148.765 ;
        RECT 105.205 146.935 105.375 147.695 ;
        RECT 105.555 146.765 105.885 147.525 ;
        RECT 106.055 146.935 106.325 147.840 ;
        RECT 106.500 147.775 106.850 148.425 ;
        RECT 107.020 147.605 107.250 148.595 ;
        RECT 106.585 147.435 107.250 147.605 ;
        RECT 106.585 146.935 106.755 147.435 ;
        RECT 106.925 146.765 107.255 147.265 ;
        RECT 107.425 146.935 107.610 149.055 ;
        RECT 107.865 148.855 108.115 149.315 ;
        RECT 108.285 148.865 108.620 149.035 ;
        RECT 108.815 148.865 109.490 149.035 ;
        RECT 108.285 148.725 108.455 148.865 ;
        RECT 107.780 147.735 108.060 148.685 ;
        RECT 108.230 148.595 108.455 148.725 ;
        RECT 108.230 147.490 108.400 148.595 ;
        RECT 108.625 148.445 109.150 148.665 ;
        RECT 108.570 147.680 108.810 148.275 ;
        RECT 108.980 147.745 109.150 148.445 ;
        RECT 109.320 148.085 109.490 148.865 ;
        RECT 109.810 148.815 110.180 149.315 ;
        RECT 110.360 148.865 110.765 149.035 ;
        RECT 110.935 148.865 111.720 149.035 ;
        RECT 110.360 148.635 110.530 148.865 ;
        RECT 109.700 148.335 110.530 148.635 ;
        RECT 110.915 148.365 111.380 148.695 ;
        RECT 109.700 148.305 109.900 148.335 ;
        RECT 110.020 148.085 110.190 148.155 ;
        RECT 109.320 147.915 110.190 148.085 ;
        RECT 109.680 147.825 110.190 147.915 ;
        RECT 108.230 147.360 108.535 147.490 ;
        RECT 108.980 147.380 109.510 147.745 ;
        RECT 107.850 146.765 108.115 147.225 ;
        RECT 108.285 146.935 108.535 147.360 ;
        RECT 109.680 147.210 109.850 147.825 ;
        RECT 108.745 147.040 109.850 147.210 ;
        RECT 110.020 146.765 110.190 147.565 ;
        RECT 110.360 147.265 110.530 148.335 ;
        RECT 110.700 147.435 110.890 148.155 ;
        RECT 111.060 147.405 111.380 148.365 ;
        RECT 111.550 148.405 111.720 148.865 ;
        RECT 111.995 148.785 112.205 149.315 ;
        RECT 112.465 148.575 112.795 149.100 ;
        RECT 112.965 148.705 113.135 149.315 ;
        RECT 113.305 148.660 113.635 149.095 ;
        RECT 114.865 148.765 115.035 149.055 ;
        RECT 115.205 148.935 115.535 149.315 ;
        RECT 113.305 148.575 113.685 148.660 ;
        RECT 114.865 148.595 115.530 148.765 ;
        RECT 112.595 148.405 112.795 148.575 ;
        RECT 113.460 148.535 113.685 148.575 ;
        RECT 111.550 148.075 112.425 148.405 ;
        RECT 112.595 148.075 113.345 148.405 ;
        RECT 110.360 146.935 110.610 147.265 ;
        RECT 111.550 147.235 111.720 148.075 ;
        RECT 112.595 147.870 112.785 148.075 ;
        RECT 113.515 147.955 113.685 148.535 ;
        RECT 113.470 147.905 113.685 147.955 ;
        RECT 111.890 147.495 112.785 147.870 ;
        RECT 113.295 147.825 113.685 147.905 ;
        RECT 110.835 147.065 111.720 147.235 ;
        RECT 111.900 146.765 112.215 147.265 ;
        RECT 112.445 146.935 112.785 147.495 ;
        RECT 112.955 146.765 113.125 147.775 ;
        RECT 113.295 146.980 113.625 147.825 ;
        RECT 114.780 147.775 115.130 148.425 ;
        RECT 115.300 147.605 115.530 148.595 ;
        RECT 114.865 147.435 115.530 147.605 ;
        RECT 114.865 146.935 115.035 147.435 ;
        RECT 115.205 146.765 115.535 147.265 ;
        RECT 115.705 146.935 115.890 149.055 ;
        RECT 116.145 148.855 116.395 149.315 ;
        RECT 116.565 148.865 116.900 149.035 ;
        RECT 117.095 148.865 117.770 149.035 ;
        RECT 116.565 148.725 116.735 148.865 ;
        RECT 116.060 147.735 116.340 148.685 ;
        RECT 116.510 148.595 116.735 148.725 ;
        RECT 116.510 147.490 116.680 148.595 ;
        RECT 116.905 148.445 117.430 148.665 ;
        RECT 116.850 147.680 117.090 148.275 ;
        RECT 117.260 147.745 117.430 148.445 ;
        RECT 117.600 148.085 117.770 148.865 ;
        RECT 118.090 148.815 118.460 149.315 ;
        RECT 118.640 148.865 119.045 149.035 ;
        RECT 119.215 148.865 120.000 149.035 ;
        RECT 118.640 148.635 118.810 148.865 ;
        RECT 117.980 148.335 118.810 148.635 ;
        RECT 119.195 148.365 119.660 148.695 ;
        RECT 117.980 148.305 118.180 148.335 ;
        RECT 118.300 148.085 118.470 148.155 ;
        RECT 117.600 147.915 118.470 148.085 ;
        RECT 117.960 147.825 118.470 147.915 ;
        RECT 116.510 147.360 116.815 147.490 ;
        RECT 117.260 147.380 117.790 147.745 ;
        RECT 116.130 146.765 116.395 147.225 ;
        RECT 116.565 146.935 116.815 147.360 ;
        RECT 117.960 147.210 118.130 147.825 ;
        RECT 117.025 147.040 118.130 147.210 ;
        RECT 118.300 146.765 118.470 147.565 ;
        RECT 118.640 147.265 118.810 148.335 ;
        RECT 118.980 147.435 119.170 148.155 ;
        RECT 119.340 147.405 119.660 148.365 ;
        RECT 119.830 148.405 120.000 148.865 ;
        RECT 120.275 148.785 120.485 149.315 ;
        RECT 120.745 148.575 121.075 149.100 ;
        RECT 121.245 148.705 121.415 149.315 ;
        RECT 121.585 148.660 121.915 149.095 ;
        RECT 121.585 148.575 121.965 148.660 ;
        RECT 120.875 148.405 121.075 148.575 ;
        RECT 121.740 148.535 121.965 148.575 ;
        RECT 119.830 148.075 120.705 148.405 ;
        RECT 120.875 148.075 121.625 148.405 ;
        RECT 118.640 146.935 118.890 147.265 ;
        RECT 119.830 147.235 120.000 148.075 ;
        RECT 120.875 147.870 121.065 148.075 ;
        RECT 121.795 147.955 121.965 148.535 ;
        RECT 121.750 147.905 121.965 147.955 ;
        RECT 120.170 147.495 121.065 147.870 ;
        RECT 121.575 147.825 121.965 147.905 ;
        RECT 122.135 148.640 122.395 149.145 ;
        RECT 122.575 148.935 122.905 149.315 ;
        RECT 123.085 148.765 123.255 149.145 ;
        RECT 122.135 147.840 122.305 148.640 ;
        RECT 122.590 148.595 123.255 148.765 ;
        RECT 123.515 148.855 124.075 149.145 ;
        RECT 124.245 148.855 124.495 149.315 ;
        RECT 122.590 148.340 122.760 148.595 ;
        RECT 122.475 148.010 122.760 148.340 ;
        RECT 122.995 148.045 123.325 148.415 ;
        RECT 122.590 147.865 122.760 148.010 ;
        RECT 119.115 147.065 120.000 147.235 ;
        RECT 120.180 146.765 120.495 147.265 ;
        RECT 120.725 146.935 121.065 147.495 ;
        RECT 121.235 146.765 121.405 147.775 ;
        RECT 121.575 146.980 121.905 147.825 ;
        RECT 122.135 146.935 122.405 147.840 ;
        RECT 122.590 147.695 123.255 147.865 ;
        RECT 122.575 146.765 122.905 147.525 ;
        RECT 123.085 146.935 123.255 147.695 ;
        RECT 123.515 147.485 123.765 148.855 ;
        RECT 125.115 148.685 125.445 149.045 ;
        RECT 124.055 148.495 125.445 148.685 ;
        RECT 125.815 148.590 126.105 149.315 ;
        RECT 126.275 148.545 128.865 149.315 ;
        RECT 124.055 148.405 124.225 148.495 ;
        RECT 123.935 148.075 124.225 148.405 ;
        RECT 124.395 148.075 124.735 148.325 ;
        RECT 124.955 148.075 125.630 148.325 ;
        RECT 124.055 147.825 124.225 148.075 ;
        RECT 124.055 147.655 124.995 147.825 ;
        RECT 125.365 147.715 125.630 148.075 ;
        RECT 126.275 148.025 127.485 148.545 ;
        RECT 129.700 148.535 130.200 149.145 ;
        RECT 123.515 146.935 123.975 147.485 ;
        RECT 124.165 146.765 124.495 147.485 ;
        RECT 124.695 147.105 124.995 147.655 ;
        RECT 125.165 146.765 125.445 147.435 ;
        RECT 125.815 146.765 126.105 147.930 ;
        RECT 127.655 147.855 128.865 148.375 ;
        RECT 129.495 148.075 129.845 148.325 ;
        RECT 130.030 147.905 130.200 148.535 ;
        RECT 130.830 148.665 131.160 149.145 ;
        RECT 131.330 148.855 131.555 149.315 ;
        RECT 131.725 148.665 132.055 149.145 ;
        RECT 130.830 148.495 132.055 148.665 ;
        RECT 132.245 148.515 132.495 149.315 ;
        RECT 132.665 148.515 133.005 149.145 ;
        RECT 130.370 148.125 130.700 148.325 ;
        RECT 130.870 148.125 131.200 148.325 ;
        RECT 131.370 148.125 131.790 148.325 ;
        RECT 131.965 148.155 132.660 148.325 ;
        RECT 131.965 147.905 132.135 148.155 ;
        RECT 132.830 147.905 133.005 148.515 ;
        RECT 133.175 148.565 134.385 149.315 ;
        RECT 134.645 148.765 134.815 149.055 ;
        RECT 134.985 148.935 135.315 149.315 ;
        RECT 134.645 148.595 135.310 148.765 ;
        RECT 133.175 148.025 133.695 148.565 ;
        RECT 126.275 146.765 128.865 147.855 ;
        RECT 129.700 147.735 132.135 147.905 ;
        RECT 129.700 146.935 130.030 147.735 ;
        RECT 130.200 146.765 130.530 147.565 ;
        RECT 130.830 146.935 131.160 147.735 ;
        RECT 131.805 146.765 132.055 147.565 ;
        RECT 132.325 146.765 132.495 147.905 ;
        RECT 132.665 146.935 133.005 147.905 ;
        RECT 133.865 147.855 134.385 148.395 ;
        RECT 133.175 146.765 134.385 147.855 ;
        RECT 134.560 147.775 134.910 148.425 ;
        RECT 135.080 147.605 135.310 148.595 ;
        RECT 134.645 147.435 135.310 147.605 ;
        RECT 134.645 146.935 134.815 147.435 ;
        RECT 134.985 146.765 135.315 147.265 ;
        RECT 135.485 146.935 135.670 149.055 ;
        RECT 135.925 148.855 136.175 149.315 ;
        RECT 136.345 148.865 136.680 149.035 ;
        RECT 136.875 148.865 137.550 149.035 ;
        RECT 136.345 148.725 136.515 148.865 ;
        RECT 135.840 147.735 136.120 148.685 ;
        RECT 136.290 148.595 136.515 148.725 ;
        RECT 136.290 147.490 136.460 148.595 ;
        RECT 136.685 148.445 137.210 148.665 ;
        RECT 136.630 147.680 136.870 148.275 ;
        RECT 137.040 147.745 137.210 148.445 ;
        RECT 137.380 148.085 137.550 148.865 ;
        RECT 137.870 148.815 138.240 149.315 ;
        RECT 138.420 148.865 138.825 149.035 ;
        RECT 138.995 148.865 139.780 149.035 ;
        RECT 138.420 148.635 138.590 148.865 ;
        RECT 137.760 148.335 138.590 148.635 ;
        RECT 138.975 148.365 139.440 148.695 ;
        RECT 137.760 148.305 137.960 148.335 ;
        RECT 138.080 148.085 138.250 148.155 ;
        RECT 137.380 147.915 138.250 148.085 ;
        RECT 137.740 147.825 138.250 147.915 ;
        RECT 136.290 147.360 136.595 147.490 ;
        RECT 137.040 147.380 137.570 147.745 ;
        RECT 135.910 146.765 136.175 147.225 ;
        RECT 136.345 146.935 136.595 147.360 ;
        RECT 137.740 147.210 137.910 147.825 ;
        RECT 136.805 147.040 137.910 147.210 ;
        RECT 138.080 146.765 138.250 147.565 ;
        RECT 138.420 147.265 138.590 148.335 ;
        RECT 138.760 147.435 138.950 148.155 ;
        RECT 139.120 147.405 139.440 148.365 ;
        RECT 139.610 148.405 139.780 148.865 ;
        RECT 140.055 148.785 140.265 149.315 ;
        RECT 140.525 148.575 140.855 149.100 ;
        RECT 141.025 148.705 141.195 149.315 ;
        RECT 141.365 148.660 141.695 149.095 ;
        RECT 142.000 148.815 142.495 149.145 ;
        RECT 141.365 148.575 141.745 148.660 ;
        RECT 140.655 148.405 140.855 148.575 ;
        RECT 141.520 148.535 141.745 148.575 ;
        RECT 139.610 148.075 140.485 148.405 ;
        RECT 140.655 148.075 141.405 148.405 ;
        RECT 138.420 146.935 138.670 147.265 ;
        RECT 139.610 147.235 139.780 148.075 ;
        RECT 140.655 147.870 140.845 148.075 ;
        RECT 141.575 147.955 141.745 148.535 ;
        RECT 141.530 147.905 141.745 147.955 ;
        RECT 139.950 147.495 140.845 147.870 ;
        RECT 141.355 147.825 141.745 147.905 ;
        RECT 138.895 147.065 139.780 147.235 ;
        RECT 139.960 146.765 140.275 147.265 ;
        RECT 140.505 146.935 140.845 147.495 ;
        RECT 141.015 146.765 141.185 147.775 ;
        RECT 141.355 146.980 141.685 147.825 ;
        RECT 141.915 147.325 142.155 148.635 ;
        RECT 142.325 147.905 142.495 148.815 ;
        RECT 142.715 148.075 143.065 149.040 ;
        RECT 143.245 148.075 143.545 149.045 ;
        RECT 143.725 148.075 144.005 149.045 ;
        RECT 144.185 148.515 144.455 149.315 ;
        RECT 144.625 148.595 144.965 149.105 ;
        RECT 144.200 148.075 144.530 148.325 ;
        RECT 144.200 147.905 144.515 148.075 ;
        RECT 142.325 147.735 144.515 147.905 ;
        RECT 141.920 146.765 142.255 147.145 ;
        RECT 142.425 146.935 142.675 147.735 ;
        RECT 142.895 146.765 143.225 147.485 ;
        RECT 143.410 146.935 143.660 147.735 ;
        RECT 144.125 146.765 144.455 147.565 ;
        RECT 144.705 147.195 144.965 148.595 ;
        RECT 145.135 148.495 145.395 149.315 ;
        RECT 145.565 148.495 145.895 148.915 ;
        RECT 146.075 148.830 146.865 149.095 ;
        RECT 145.645 148.405 145.895 148.495 ;
        RECT 145.135 147.445 145.475 148.325 ;
        RECT 145.645 148.155 146.440 148.405 ;
        RECT 144.625 146.935 144.965 147.195 ;
        RECT 145.135 146.765 145.395 147.275 ;
        RECT 145.645 146.935 145.815 148.155 ;
        RECT 146.610 147.975 146.865 148.830 ;
        RECT 147.035 148.675 147.235 149.095 ;
        RECT 147.425 148.855 147.755 149.315 ;
        RECT 147.035 148.155 147.445 148.675 ;
        RECT 147.925 148.665 148.185 149.145 ;
        RECT 147.615 147.975 147.845 148.405 ;
        RECT 146.055 147.805 147.845 147.975 ;
        RECT 146.055 147.440 146.305 147.805 ;
        RECT 146.475 147.445 146.805 147.635 ;
        RECT 147.025 147.510 147.740 147.805 ;
        RECT 148.015 147.635 148.185 148.665 ;
        RECT 148.445 148.765 148.615 149.145 ;
        RECT 148.795 148.935 149.125 149.315 ;
        RECT 148.445 148.595 149.110 148.765 ;
        RECT 149.305 148.640 149.565 149.145 ;
        RECT 148.375 148.045 148.705 148.415 ;
        RECT 148.940 148.340 149.110 148.595 ;
        RECT 148.940 148.010 149.225 148.340 ;
        RECT 148.940 147.865 149.110 148.010 ;
        RECT 146.475 147.270 146.670 147.445 ;
        RECT 146.055 146.765 146.670 147.270 ;
        RECT 146.840 146.935 147.315 147.275 ;
        RECT 147.485 146.765 147.700 147.310 ;
        RECT 147.910 146.935 148.185 147.635 ;
        RECT 148.445 147.695 149.110 147.865 ;
        RECT 149.395 147.840 149.565 148.640 ;
        RECT 149.735 148.545 151.405 149.315 ;
        RECT 151.575 148.590 151.865 149.315 ;
        RECT 152.035 148.545 155.545 149.315 ;
        RECT 155.715 148.565 156.925 149.315 ;
        RECT 149.735 148.025 150.485 148.545 ;
        RECT 150.655 147.855 151.405 148.375 ;
        RECT 152.035 148.025 153.685 148.545 ;
        RECT 148.445 146.935 148.615 147.695 ;
        RECT 148.795 146.765 149.125 147.525 ;
        RECT 149.295 146.935 149.565 147.840 ;
        RECT 149.735 146.765 151.405 147.855 ;
        RECT 151.575 146.765 151.865 147.930 ;
        RECT 153.855 147.855 155.545 148.375 ;
        RECT 152.035 146.765 155.545 147.855 ;
        RECT 155.715 147.855 156.235 148.395 ;
        RECT 156.405 148.025 156.925 148.565 ;
        RECT 155.715 146.765 156.925 147.855 ;
        RECT 22.690 146.595 157.010 146.765 ;
        RECT 22.775 145.505 23.985 146.595 ;
        RECT 24.155 145.505 26.745 146.595 ;
        RECT 26.925 146.005 27.185 146.395 ;
        RECT 27.355 146.185 27.685 146.595 ;
        RECT 26.925 145.805 27.685 146.005 ;
        RECT 22.775 144.795 23.295 145.335 ;
        RECT 23.465 144.965 23.985 145.505 ;
        RECT 24.155 144.815 25.365 145.335 ;
        RECT 25.535 144.985 26.745 145.505 ;
        RECT 26.935 144.935 27.165 145.625 ;
        RECT 27.345 145.125 27.685 145.805 ;
        RECT 27.875 145.305 28.205 146.415 ;
        RECT 28.375 145.685 28.565 146.415 ;
        RECT 28.735 145.865 29.065 146.595 ;
        RECT 29.245 145.685 29.415 146.415 ;
        RECT 28.375 145.485 29.415 145.685 ;
        RECT 29.675 145.505 33.185 146.595 ;
        RECT 33.360 145.795 33.615 146.595 ;
        RECT 33.815 145.745 34.145 146.425 ;
        RECT 22.775 144.045 23.985 144.795 ;
        RECT 24.155 144.045 26.745 144.815 ;
        RECT 27.345 144.675 27.575 145.125 ;
        RECT 27.875 145.005 28.410 145.305 ;
        RECT 27.195 144.225 27.575 144.675 ;
        RECT 27.755 144.045 27.985 144.825 ;
        RECT 28.165 144.755 28.410 145.005 ;
        RECT 28.590 144.955 28.985 145.305 ;
        RECT 29.180 144.955 29.470 145.305 ;
        RECT 28.165 144.225 28.595 144.755 ;
        RECT 28.775 144.335 28.985 144.955 ;
        RECT 29.675 144.815 31.325 145.335 ;
        RECT 31.495 144.985 33.185 145.505 ;
        RECT 33.360 145.255 33.605 145.615 ;
        RECT 33.795 145.465 34.145 145.745 ;
        RECT 33.795 145.085 33.965 145.465 ;
        RECT 34.325 145.285 34.520 146.335 ;
        RECT 34.700 145.455 35.020 146.595 ;
        RECT 35.655 145.430 35.945 146.595 ;
        RECT 37.035 145.455 37.420 146.425 ;
        RECT 37.590 146.135 37.915 146.595 ;
        RECT 38.435 145.965 38.715 146.425 ;
        RECT 37.590 145.745 38.715 145.965 ;
        RECT 33.445 144.915 33.965 145.085 ;
        RECT 34.135 144.955 34.520 145.285 ;
        RECT 34.700 145.235 34.960 145.285 ;
        RECT 34.700 145.065 34.965 145.235 ;
        RECT 34.700 144.955 34.960 145.065 ;
        RECT 29.155 144.045 29.485 144.775 ;
        RECT 29.675 144.045 33.185 144.815 ;
        RECT 33.445 144.350 33.615 144.915 ;
        RECT 37.035 144.785 37.315 145.455 ;
        RECT 37.590 145.285 38.040 145.745 ;
        RECT 38.905 145.575 39.305 146.425 ;
        RECT 39.705 146.135 39.975 146.595 ;
        RECT 40.145 145.965 40.430 146.425 ;
        RECT 37.485 144.955 38.040 145.285 ;
        RECT 38.210 145.015 39.305 145.575 ;
        RECT 37.590 144.845 38.040 144.955 ;
        RECT 33.805 144.575 35.020 144.745 ;
        RECT 33.805 144.270 34.035 144.575 ;
        RECT 34.205 144.045 34.535 144.405 ;
        RECT 34.730 144.225 35.020 144.575 ;
        RECT 35.655 144.045 35.945 144.770 ;
        RECT 37.035 144.215 37.420 144.785 ;
        RECT 37.590 144.675 38.715 144.845 ;
        RECT 37.590 144.045 37.915 144.505 ;
        RECT 38.435 144.215 38.715 144.675 ;
        RECT 38.905 144.215 39.305 145.015 ;
        RECT 39.475 145.745 40.430 145.965 ;
        RECT 39.475 144.845 39.685 145.745 ;
        RECT 39.855 145.015 40.545 145.575 ;
        RECT 40.715 145.505 44.225 146.595 ;
        RECT 44.435 145.965 44.765 146.425 ;
        RECT 44.935 146.135 45.195 146.595 ;
        RECT 45.470 146.175 47.405 146.425 ;
        RECT 47.575 146.235 47.905 146.595 ;
        RECT 48.435 146.235 48.765 146.595 ;
        RECT 44.435 145.745 45.300 145.965 ;
        RECT 45.470 145.755 45.665 146.175 ;
        RECT 46.245 146.165 47.405 146.175 ;
        RECT 47.205 146.065 47.405 146.165 ;
        RECT 48.935 146.065 49.125 146.425 ;
        RECT 49.295 146.235 49.625 146.595 ;
        RECT 49.795 146.065 49.975 146.425 ;
        RECT 50.155 146.235 50.485 146.595 ;
        RECT 50.655 146.065 50.915 146.425 ;
        RECT 45.870 145.915 47.035 145.995 ;
        RECT 45.835 145.745 47.035 145.915 ;
        RECT 47.205 145.835 50.915 146.065 ;
        RECT 39.475 144.675 40.430 144.845 ;
        RECT 39.705 144.045 39.975 144.505 ;
        RECT 40.145 144.215 40.430 144.675 ;
        RECT 40.715 144.815 42.365 145.335 ;
        RECT 42.535 144.985 44.225 145.505 ;
        RECT 44.455 145.035 44.960 145.575 ;
        RECT 44.790 144.955 44.960 145.035 ;
        RECT 45.130 145.305 45.300 145.745 ;
        RECT 45.870 145.665 47.035 145.745 ;
        RECT 45.870 145.545 47.170 145.665 ;
        RECT 45.130 144.995 46.710 145.305 ;
        RECT 40.715 144.045 44.225 144.815 ;
        RECT 45.130 144.755 45.415 144.995 ;
        RECT 46.880 144.855 47.170 145.545 ;
        RECT 47.340 145.440 50.760 145.665 ;
        RECT 52.215 145.455 52.495 146.595 ;
        RECT 52.665 145.445 52.995 146.425 ;
        RECT 53.165 145.455 53.425 146.595 ;
        RECT 53.595 145.505 55.265 146.595 ;
        RECT 47.340 145.025 47.685 145.440 ;
        RECT 47.855 145.025 49.280 145.270 ;
        RECT 49.515 145.035 50.760 145.440 ;
        RECT 52.225 145.015 52.560 145.285 ;
        RECT 46.880 144.825 49.195 144.855 ;
        RECT 44.400 144.575 45.415 144.755 ;
        RECT 45.585 144.655 49.195 144.825 ;
        RECT 45.585 144.575 46.635 144.655 ;
        RECT 47.565 144.635 49.195 144.655 ;
        RECT 49.365 144.695 50.485 144.865 ;
        RECT 52.730 144.845 52.900 145.445 ;
        RECT 53.070 145.035 53.405 145.285 ;
        RECT 44.400 144.215 44.755 144.575 ;
        RECT 45.030 144.045 45.415 144.405 ;
        RECT 45.585 144.330 45.775 144.575 ;
        RECT 45.945 144.045 46.275 144.405 ;
        RECT 46.445 144.215 46.635 144.575 ;
        RECT 46.805 144.045 47.395 144.485 ;
        RECT 49.365 144.465 49.625 144.695 ;
        RECT 47.575 144.215 49.625 144.465 ;
        RECT 49.795 144.045 49.985 144.525 ;
        RECT 50.155 144.215 50.485 144.695 ;
        RECT 50.655 144.045 50.915 144.845 ;
        RECT 52.215 144.045 52.525 144.845 ;
        RECT 52.730 144.215 53.425 144.845 ;
        RECT 53.595 144.815 54.345 145.335 ;
        RECT 54.515 144.985 55.265 145.505 ;
        RECT 55.435 145.725 55.710 146.425 ;
        RECT 55.920 146.050 56.135 146.595 ;
        RECT 56.305 146.085 56.780 146.425 ;
        RECT 56.950 146.090 57.565 146.595 ;
        RECT 56.950 145.915 57.145 146.090 ;
        RECT 53.595 144.045 55.265 144.815 ;
        RECT 55.435 144.695 55.605 145.725 ;
        RECT 55.880 145.555 56.595 145.850 ;
        RECT 56.815 145.725 57.145 145.915 ;
        RECT 57.315 145.555 57.565 145.920 ;
        RECT 55.775 145.385 57.565 145.555 ;
        RECT 55.775 144.955 56.005 145.385 ;
        RECT 55.435 144.215 55.695 144.695 ;
        RECT 56.175 144.685 56.585 145.205 ;
        RECT 55.865 144.045 56.195 144.505 ;
        RECT 56.385 144.265 56.585 144.685 ;
        RECT 56.755 144.530 57.010 145.385 ;
        RECT 57.805 145.205 57.975 146.425 ;
        RECT 58.225 146.085 58.485 146.595 ;
        RECT 57.180 144.955 57.975 145.205 ;
        RECT 58.145 145.035 58.485 145.915 ;
        RECT 58.655 145.505 61.245 146.595 ;
        RECT 57.725 144.865 57.975 144.955 ;
        RECT 56.755 144.265 57.545 144.530 ;
        RECT 57.725 144.445 58.055 144.865 ;
        RECT 58.225 144.045 58.485 144.865 ;
        RECT 58.655 144.815 59.865 145.335 ;
        RECT 60.035 144.985 61.245 145.505 ;
        RECT 61.415 145.430 61.705 146.595 ;
        RECT 61.875 145.505 63.545 146.595 ;
        RECT 61.875 144.815 62.625 145.335 ;
        RECT 62.795 144.985 63.545 145.505 ;
        RECT 58.655 144.045 61.245 144.815 ;
        RECT 61.415 144.045 61.705 144.770 ;
        RECT 61.875 144.045 63.545 144.815 ;
        RECT 63.730 144.225 64.010 146.415 ;
        RECT 64.200 145.455 64.485 146.595 ;
        RECT 64.750 145.945 64.920 146.415 ;
        RECT 65.095 146.115 65.425 146.595 ;
        RECT 65.595 145.945 65.775 146.415 ;
        RECT 64.750 145.745 65.775 145.945 ;
        RECT 64.210 144.775 64.470 145.285 ;
        RECT 64.680 144.955 64.940 145.575 ;
        RECT 65.135 144.955 65.560 145.575 ;
        RECT 65.945 145.305 66.275 146.415 ;
        RECT 66.445 146.185 66.795 146.595 ;
        RECT 66.965 146.005 67.205 146.395 ;
        RECT 65.730 145.005 66.275 145.305 ;
        RECT 66.455 145.805 67.205 146.005 ;
        RECT 66.455 145.125 66.795 145.805 ;
        RECT 65.730 144.775 65.950 145.005 ;
        RECT 64.210 144.585 65.950 144.775 ;
        RECT 64.210 144.045 64.940 144.415 ;
        RECT 65.520 144.225 65.950 144.585 ;
        RECT 66.120 144.045 66.365 144.825 ;
        RECT 66.565 144.225 66.795 145.125 ;
        RECT 66.975 144.285 67.205 145.625 ;
        RECT 67.395 145.455 67.780 146.425 ;
        RECT 67.950 146.135 68.275 146.595 ;
        RECT 68.795 145.965 69.075 146.425 ;
        RECT 67.950 145.745 69.075 145.965 ;
        RECT 67.395 144.785 67.675 145.455 ;
        RECT 67.950 145.285 68.400 145.745 ;
        RECT 69.265 145.575 69.665 146.425 ;
        RECT 70.065 146.135 70.335 146.595 ;
        RECT 70.505 145.965 70.790 146.425 ;
        RECT 67.845 144.955 68.400 145.285 ;
        RECT 68.570 145.015 69.665 145.575 ;
        RECT 67.950 144.845 68.400 144.955 ;
        RECT 67.395 144.215 67.780 144.785 ;
        RECT 67.950 144.675 69.075 144.845 ;
        RECT 67.950 144.045 68.275 144.505 ;
        RECT 68.795 144.215 69.075 144.675 ;
        RECT 69.265 144.215 69.665 145.015 ;
        RECT 69.835 145.745 70.790 145.965 ;
        RECT 69.835 144.845 70.045 145.745 ;
        RECT 70.215 145.015 70.905 145.575 ;
        RECT 71.995 145.455 72.380 146.425 ;
        RECT 72.550 146.135 72.875 146.595 ;
        RECT 73.395 145.965 73.675 146.425 ;
        RECT 72.550 145.745 73.675 145.965 ;
        RECT 69.835 144.675 70.790 144.845 ;
        RECT 70.065 144.045 70.335 144.505 ;
        RECT 70.505 144.215 70.790 144.675 ;
        RECT 71.995 144.785 72.275 145.455 ;
        RECT 72.550 145.285 73.000 145.745 ;
        RECT 73.865 145.575 74.265 146.425 ;
        RECT 74.665 146.135 74.935 146.595 ;
        RECT 75.105 145.965 75.390 146.425 ;
        RECT 72.445 144.955 73.000 145.285 ;
        RECT 73.170 145.015 74.265 145.575 ;
        RECT 72.550 144.845 73.000 144.955 ;
        RECT 71.995 144.215 72.380 144.785 ;
        RECT 72.550 144.675 73.675 144.845 ;
        RECT 72.550 144.045 72.875 144.505 ;
        RECT 73.395 144.215 73.675 144.675 ;
        RECT 73.865 144.215 74.265 145.015 ;
        RECT 74.435 145.745 75.390 145.965 ;
        RECT 75.685 145.785 75.980 146.595 ;
        RECT 74.435 144.845 74.645 145.745 ;
        RECT 74.815 145.015 75.505 145.575 ;
        RECT 76.160 145.285 76.405 146.425 ;
        RECT 76.580 145.785 76.840 146.595 ;
        RECT 77.440 146.590 83.715 146.595 ;
        RECT 77.020 145.285 77.270 146.420 ;
        RECT 77.440 145.795 77.700 146.590 ;
        RECT 77.870 145.695 78.130 146.420 ;
        RECT 78.300 145.865 78.560 146.590 ;
        RECT 78.730 145.695 78.990 146.420 ;
        RECT 79.160 145.865 79.420 146.590 ;
        RECT 79.590 145.695 79.850 146.420 ;
        RECT 80.020 145.865 80.280 146.590 ;
        RECT 80.450 145.695 80.710 146.420 ;
        RECT 80.880 145.865 81.125 146.590 ;
        RECT 81.295 145.695 81.555 146.420 ;
        RECT 81.740 145.865 81.985 146.590 ;
        RECT 82.155 145.695 82.415 146.420 ;
        RECT 82.600 145.865 82.845 146.590 ;
        RECT 83.015 145.695 83.275 146.420 ;
        RECT 83.460 145.865 83.715 146.590 ;
        RECT 77.870 145.680 83.275 145.695 ;
        RECT 83.885 145.680 84.175 146.420 ;
        RECT 84.345 145.850 84.615 146.595 ;
        RECT 77.870 145.455 84.615 145.680 ;
        RECT 84.875 145.505 86.545 146.595 ;
        RECT 74.435 144.675 75.390 144.845 ;
        RECT 75.675 144.725 75.990 145.285 ;
        RECT 76.160 145.035 83.280 145.285 ;
        RECT 74.665 144.045 74.935 144.505 ;
        RECT 75.105 144.215 75.390 144.675 ;
        RECT 75.675 144.045 75.980 144.555 ;
        RECT 76.160 144.225 76.410 145.035 ;
        RECT 76.580 144.045 76.840 144.570 ;
        RECT 77.020 144.225 77.270 145.035 ;
        RECT 83.450 144.865 84.615 145.455 ;
        RECT 77.870 144.695 84.615 144.865 ;
        RECT 84.875 144.815 85.625 145.335 ;
        RECT 85.795 144.985 86.545 145.505 ;
        RECT 87.175 145.430 87.465 146.595 ;
        RECT 88.645 145.925 88.815 146.425 ;
        RECT 88.985 146.095 89.315 146.595 ;
        RECT 88.645 145.755 89.310 145.925 ;
        RECT 88.560 144.935 88.910 145.585 ;
        RECT 77.440 144.045 77.700 144.605 ;
        RECT 77.870 144.240 78.130 144.695 ;
        RECT 78.300 144.045 78.560 144.525 ;
        RECT 78.730 144.240 78.990 144.695 ;
        RECT 79.160 144.045 79.420 144.525 ;
        RECT 79.590 144.240 79.850 144.695 ;
        RECT 80.020 144.045 80.265 144.525 ;
        RECT 80.435 144.240 80.710 144.695 ;
        RECT 80.880 144.045 81.125 144.525 ;
        RECT 81.295 144.240 81.555 144.695 ;
        RECT 81.735 144.045 81.985 144.525 ;
        RECT 82.155 144.240 82.415 144.695 ;
        RECT 82.595 144.045 82.845 144.525 ;
        RECT 83.015 144.240 83.275 144.695 ;
        RECT 83.455 144.045 83.715 144.525 ;
        RECT 83.885 144.240 84.145 144.695 ;
        RECT 84.315 144.045 84.615 144.525 ;
        RECT 84.875 144.045 86.545 144.815 ;
        RECT 87.175 144.045 87.465 144.770 ;
        RECT 89.080 144.765 89.310 145.755 ;
        RECT 88.645 144.595 89.310 144.765 ;
        RECT 88.645 144.305 88.815 144.595 ;
        RECT 88.985 144.045 89.315 144.425 ;
        RECT 89.485 144.305 89.670 146.425 ;
        RECT 89.910 146.135 90.175 146.595 ;
        RECT 90.345 146.000 90.595 146.425 ;
        RECT 90.805 146.150 91.910 146.320 ;
        RECT 90.290 145.870 90.595 146.000 ;
        RECT 89.840 144.675 90.120 145.625 ;
        RECT 90.290 144.765 90.460 145.870 ;
        RECT 90.630 145.085 90.870 145.680 ;
        RECT 91.040 145.615 91.570 145.980 ;
        RECT 91.040 144.915 91.210 145.615 ;
        RECT 91.740 145.535 91.910 146.150 ;
        RECT 92.080 145.795 92.250 146.595 ;
        RECT 92.420 146.095 92.670 146.425 ;
        RECT 92.895 146.125 93.780 146.295 ;
        RECT 91.740 145.445 92.250 145.535 ;
        RECT 90.290 144.635 90.515 144.765 ;
        RECT 90.685 144.695 91.210 144.915 ;
        RECT 91.380 145.275 92.250 145.445 ;
        RECT 89.925 144.045 90.175 144.505 ;
        RECT 90.345 144.495 90.515 144.635 ;
        RECT 91.380 144.495 91.550 145.275 ;
        RECT 92.080 145.205 92.250 145.275 ;
        RECT 91.760 145.025 91.960 145.055 ;
        RECT 92.420 145.025 92.590 146.095 ;
        RECT 92.760 145.205 92.950 145.925 ;
        RECT 91.760 144.725 92.590 145.025 ;
        RECT 93.120 144.995 93.440 145.955 ;
        RECT 90.345 144.325 90.680 144.495 ;
        RECT 90.875 144.325 91.550 144.495 ;
        RECT 91.870 144.045 92.240 144.545 ;
        RECT 92.420 144.495 92.590 144.725 ;
        RECT 92.975 144.665 93.440 144.995 ;
        RECT 93.610 145.285 93.780 146.125 ;
        RECT 93.960 146.095 94.275 146.595 ;
        RECT 94.505 145.865 94.845 146.425 ;
        RECT 93.950 145.490 94.845 145.865 ;
        RECT 95.015 145.585 95.185 146.595 ;
        RECT 94.655 145.285 94.845 145.490 ;
        RECT 95.355 145.535 95.685 146.380 ;
        RECT 96.100 145.625 96.490 145.800 ;
        RECT 96.975 145.795 97.305 146.595 ;
        RECT 97.475 145.805 98.010 146.425 ;
        RECT 95.355 145.455 95.745 145.535 ;
        RECT 96.100 145.455 97.525 145.625 ;
        RECT 95.530 145.405 95.745 145.455 ;
        RECT 93.610 144.955 94.485 145.285 ;
        RECT 94.655 144.955 95.405 145.285 ;
        RECT 93.610 144.495 93.780 144.955 ;
        RECT 94.655 144.785 94.855 144.955 ;
        RECT 95.575 144.825 95.745 145.405 ;
        RECT 95.520 144.785 95.745 144.825 ;
        RECT 92.420 144.325 92.825 144.495 ;
        RECT 92.995 144.325 93.780 144.495 ;
        RECT 94.055 144.045 94.265 144.575 ;
        RECT 94.525 144.260 94.855 144.785 ;
        RECT 95.365 144.700 95.745 144.785 ;
        RECT 95.975 144.725 96.330 145.285 ;
        RECT 95.025 144.045 95.195 144.655 ;
        RECT 95.365 144.265 95.695 144.700 ;
        RECT 96.500 144.555 96.670 145.455 ;
        RECT 96.840 144.725 97.105 145.285 ;
        RECT 97.355 144.955 97.525 145.455 ;
        RECT 97.695 144.785 98.010 145.805 ;
        RECT 98.305 145.665 98.475 146.425 ;
        RECT 98.690 145.835 99.020 146.595 ;
        RECT 98.305 145.495 99.020 145.665 ;
        RECT 99.190 145.520 99.445 146.425 ;
        RECT 98.215 144.945 98.570 145.315 ;
        RECT 98.850 145.285 99.020 145.495 ;
        RECT 98.850 144.955 99.105 145.285 ;
        RECT 96.080 144.045 96.320 144.555 ;
        RECT 96.500 144.225 96.780 144.555 ;
        RECT 97.010 144.045 97.225 144.555 ;
        RECT 97.395 144.215 98.010 144.785 ;
        RECT 98.850 144.765 99.020 144.955 ;
        RECT 99.275 144.790 99.445 145.520 ;
        RECT 99.620 145.445 99.880 146.595 ;
        RECT 100.055 145.505 103.565 146.595 ;
        RECT 98.305 144.595 99.020 144.765 ;
        RECT 98.305 144.215 98.475 144.595 ;
        RECT 98.690 144.045 99.020 144.425 ;
        RECT 99.190 144.215 99.445 144.790 ;
        RECT 99.620 144.045 99.880 144.885 ;
        RECT 100.055 144.815 101.705 145.335 ;
        RECT 101.875 144.985 103.565 145.505 ;
        RECT 103.740 145.625 104.015 146.425 ;
        RECT 104.185 145.795 104.515 146.595 ;
        RECT 104.685 145.625 104.855 146.425 ;
        RECT 105.025 145.795 105.275 146.595 ;
        RECT 105.445 146.255 107.540 146.425 ;
        RECT 105.445 145.625 105.775 146.255 ;
        RECT 103.740 145.415 105.775 145.625 ;
        RECT 105.945 145.705 106.115 146.085 ;
        RECT 106.285 145.895 106.615 146.255 ;
        RECT 106.785 145.705 106.955 146.085 ;
        RECT 107.125 145.875 107.540 146.255 ;
        RECT 105.945 145.405 107.705 145.705 ;
        RECT 103.790 145.035 105.450 145.235 ;
        RECT 105.770 145.035 107.135 145.235 ;
        RECT 107.305 144.865 107.705 145.405 ;
        RECT 100.055 144.045 103.565 144.815 ;
        RECT 103.740 144.045 104.015 144.865 ;
        RECT 104.185 144.685 107.705 144.865 ;
        RECT 108.800 145.455 109.135 146.425 ;
        RECT 109.305 145.455 109.475 146.595 ;
        RECT 109.645 146.255 111.675 146.425 ;
        RECT 108.800 144.785 108.970 145.455 ;
        RECT 109.645 145.285 109.815 146.255 ;
        RECT 109.140 144.955 109.395 145.285 ;
        RECT 109.620 144.955 109.815 145.285 ;
        RECT 109.985 145.915 111.110 146.085 ;
        RECT 109.225 144.785 109.395 144.955 ;
        RECT 109.985 144.785 110.155 145.915 ;
        RECT 104.185 144.215 104.515 144.685 ;
        RECT 104.685 144.045 104.855 144.515 ;
        RECT 105.025 144.215 105.355 144.685 ;
        RECT 105.525 144.045 105.695 144.515 ;
        RECT 105.865 144.215 106.195 144.685 ;
        RECT 106.365 144.045 106.535 144.515 ;
        RECT 106.705 144.215 107.035 144.685 ;
        RECT 107.205 144.045 107.490 144.515 ;
        RECT 108.800 144.215 109.055 144.785 ;
        RECT 109.225 144.615 110.155 144.785 ;
        RECT 110.325 145.575 111.335 145.745 ;
        RECT 110.325 144.775 110.495 145.575 ;
        RECT 109.980 144.580 110.155 144.615 ;
        RECT 109.225 144.045 109.555 144.445 ;
        RECT 109.980 144.215 110.510 144.580 ;
        RECT 110.700 144.555 110.975 145.375 ;
        RECT 110.695 144.385 110.975 144.555 ;
        RECT 110.700 144.215 110.975 144.385 ;
        RECT 111.145 144.215 111.335 145.575 ;
        RECT 111.505 145.590 111.675 146.255 ;
        RECT 111.845 145.835 112.015 146.595 ;
        RECT 112.250 145.835 112.765 146.245 ;
        RECT 111.505 145.400 112.255 145.590 ;
        RECT 112.425 145.025 112.765 145.835 ;
        RECT 112.935 145.430 113.225 146.595 ;
        RECT 113.395 145.505 115.065 146.595 ;
        RECT 111.535 144.855 112.765 145.025 ;
        RECT 111.515 144.045 112.025 144.580 ;
        RECT 112.245 144.250 112.490 144.855 ;
        RECT 113.395 144.815 114.145 145.335 ;
        RECT 114.315 144.985 115.065 145.505 ;
        RECT 115.235 145.835 115.750 146.245 ;
        RECT 115.985 145.835 116.155 146.595 ;
        RECT 116.325 146.255 118.355 146.425 ;
        RECT 115.235 145.025 115.575 145.835 ;
        RECT 116.325 145.590 116.495 146.255 ;
        RECT 116.890 145.915 118.015 146.085 ;
        RECT 115.745 145.400 116.495 145.590 ;
        RECT 116.665 145.575 117.675 145.745 ;
        RECT 115.235 144.855 116.465 145.025 ;
        RECT 112.935 144.045 113.225 144.770 ;
        RECT 113.395 144.045 115.065 144.815 ;
        RECT 115.510 144.250 115.755 144.855 ;
        RECT 115.975 144.045 116.485 144.580 ;
        RECT 116.665 144.215 116.855 145.575 ;
        RECT 117.025 144.895 117.300 145.375 ;
        RECT 117.025 144.725 117.305 144.895 ;
        RECT 117.505 144.775 117.675 145.575 ;
        RECT 117.845 144.785 118.015 145.915 ;
        RECT 118.185 145.285 118.355 146.255 ;
        RECT 118.525 145.455 118.695 146.595 ;
        RECT 118.865 145.455 119.200 146.425 ;
        RECT 119.375 145.505 121.045 146.595 ;
        RECT 121.765 145.925 121.935 146.425 ;
        RECT 122.105 146.095 122.435 146.595 ;
        RECT 121.765 145.755 122.430 145.925 ;
        RECT 118.185 144.955 118.380 145.285 ;
        RECT 118.605 144.955 118.860 145.285 ;
        RECT 118.605 144.785 118.775 144.955 ;
        RECT 119.030 144.785 119.200 145.455 ;
        RECT 117.025 144.215 117.300 144.725 ;
        RECT 117.845 144.615 118.775 144.785 ;
        RECT 117.845 144.580 118.020 144.615 ;
        RECT 117.490 144.215 118.020 144.580 ;
        RECT 118.445 144.045 118.775 144.445 ;
        RECT 118.945 144.215 119.200 144.785 ;
        RECT 119.375 144.815 120.125 145.335 ;
        RECT 120.295 144.985 121.045 145.505 ;
        RECT 121.680 144.935 122.030 145.585 ;
        RECT 119.375 144.045 121.045 144.815 ;
        RECT 122.200 144.765 122.430 145.755 ;
        RECT 121.765 144.595 122.430 144.765 ;
        RECT 121.765 144.305 121.935 144.595 ;
        RECT 122.105 144.045 122.435 144.425 ;
        RECT 122.605 144.305 122.790 146.425 ;
        RECT 123.030 146.135 123.295 146.595 ;
        RECT 123.465 146.000 123.715 146.425 ;
        RECT 123.925 146.150 125.030 146.320 ;
        RECT 123.410 145.870 123.715 146.000 ;
        RECT 122.960 144.675 123.240 145.625 ;
        RECT 123.410 144.765 123.580 145.870 ;
        RECT 123.750 145.085 123.990 145.680 ;
        RECT 124.160 145.615 124.690 145.980 ;
        RECT 124.160 144.915 124.330 145.615 ;
        RECT 124.860 145.535 125.030 146.150 ;
        RECT 125.200 145.795 125.370 146.595 ;
        RECT 125.540 146.095 125.790 146.425 ;
        RECT 126.015 146.125 126.900 146.295 ;
        RECT 124.860 145.445 125.370 145.535 ;
        RECT 123.410 144.635 123.635 144.765 ;
        RECT 123.805 144.695 124.330 144.915 ;
        RECT 124.500 145.275 125.370 145.445 ;
        RECT 123.045 144.045 123.295 144.505 ;
        RECT 123.465 144.495 123.635 144.635 ;
        RECT 124.500 144.495 124.670 145.275 ;
        RECT 125.200 145.205 125.370 145.275 ;
        RECT 124.880 145.025 125.080 145.055 ;
        RECT 125.540 145.025 125.710 146.095 ;
        RECT 125.880 145.205 126.070 145.925 ;
        RECT 124.880 144.725 125.710 145.025 ;
        RECT 126.240 144.995 126.560 145.955 ;
        RECT 123.465 144.325 123.800 144.495 ;
        RECT 123.995 144.325 124.670 144.495 ;
        RECT 124.990 144.045 125.360 144.545 ;
        RECT 125.540 144.495 125.710 144.725 ;
        RECT 126.095 144.665 126.560 144.995 ;
        RECT 126.730 145.285 126.900 146.125 ;
        RECT 127.080 146.095 127.395 146.595 ;
        RECT 127.625 145.865 127.965 146.425 ;
        RECT 127.070 145.490 127.965 145.865 ;
        RECT 128.135 145.585 128.305 146.595 ;
        RECT 127.775 145.285 127.965 145.490 ;
        RECT 128.475 145.535 128.805 146.380 ;
        RECT 129.960 146.205 130.295 146.425 ;
        RECT 131.300 146.215 131.655 146.595 ;
        RECT 129.960 145.585 130.215 146.205 ;
        RECT 130.465 146.045 130.695 146.085 ;
        RECT 131.825 146.045 132.075 146.425 ;
        RECT 130.465 145.845 132.075 146.045 ;
        RECT 130.465 145.755 130.650 145.845 ;
        RECT 131.240 145.835 132.075 145.845 ;
        RECT 132.325 145.815 132.575 146.595 ;
        RECT 132.745 145.745 133.005 146.425 ;
        RECT 130.805 145.645 131.135 145.675 ;
        RECT 130.805 145.585 132.605 145.645 ;
        RECT 128.475 145.455 128.865 145.535 ;
        RECT 128.650 145.405 128.865 145.455 ;
        RECT 129.960 145.475 132.665 145.585 ;
        RECT 129.960 145.415 131.135 145.475 ;
        RECT 132.465 145.440 132.665 145.475 ;
        RECT 126.730 144.955 127.605 145.285 ;
        RECT 127.775 144.955 128.525 145.285 ;
        RECT 126.730 144.495 126.900 144.955 ;
        RECT 127.775 144.785 127.975 144.955 ;
        RECT 128.695 144.825 128.865 145.405 ;
        RECT 129.955 145.035 130.445 145.235 ;
        RECT 130.635 145.035 131.110 145.245 ;
        RECT 128.640 144.785 128.865 144.825 ;
        RECT 125.540 144.325 125.945 144.495 ;
        RECT 126.115 144.325 126.900 144.495 ;
        RECT 127.175 144.045 127.385 144.575 ;
        RECT 127.645 144.260 127.975 144.785 ;
        RECT 128.485 144.700 128.865 144.785 ;
        RECT 128.145 144.045 128.315 144.655 ;
        RECT 128.485 144.265 128.815 144.700 ;
        RECT 129.960 144.045 130.415 144.810 ;
        RECT 130.890 144.635 131.110 145.035 ;
        RECT 131.355 145.035 131.685 145.245 ;
        RECT 131.355 144.635 131.565 145.035 ;
        RECT 131.855 145.000 132.265 145.305 ;
        RECT 132.495 144.865 132.665 145.440 ;
        RECT 132.395 144.745 132.665 144.865 ;
        RECT 131.820 144.700 132.665 144.745 ;
        RECT 131.820 144.575 132.575 144.700 ;
        RECT 131.820 144.425 131.990 144.575 ;
        RECT 132.835 144.545 133.005 145.745 ;
        RECT 130.690 144.215 131.990 144.425 ;
        RECT 132.245 144.045 132.575 144.405 ;
        RECT 132.745 144.215 133.005 144.545 ;
        RECT 133.175 144.325 133.455 146.425 ;
        RECT 133.645 145.835 134.430 146.595 ;
        RECT 134.825 145.765 135.210 146.425 ;
        RECT 134.825 145.665 135.235 145.765 ;
        RECT 133.625 145.455 135.235 145.665 ;
        RECT 135.535 145.575 135.735 146.365 ;
        RECT 133.625 144.855 133.900 145.455 ;
        RECT 135.405 145.405 135.735 145.575 ;
        RECT 135.905 145.415 136.225 146.595 ;
        RECT 136.395 146.085 137.585 146.375 ;
        RECT 136.415 145.745 137.585 145.915 ;
        RECT 137.755 145.795 138.035 146.595 ;
        RECT 136.415 145.455 136.740 145.745 ;
        RECT 137.415 145.625 137.585 145.745 ;
        RECT 135.405 145.285 135.585 145.405 ;
        RECT 136.910 145.285 137.105 145.575 ;
        RECT 137.415 145.455 138.075 145.625 ;
        RECT 138.245 145.455 138.520 146.425 ;
        RECT 137.905 145.285 138.075 145.455 ;
        RECT 134.070 145.035 134.425 145.285 ;
        RECT 134.620 145.235 135.085 145.285 ;
        RECT 134.615 145.065 135.085 145.235 ;
        RECT 134.620 145.035 135.085 145.065 ;
        RECT 135.255 145.035 135.585 145.285 ;
        RECT 135.760 145.035 136.225 145.235 ;
        RECT 136.395 144.955 136.740 145.285 ;
        RECT 136.910 144.955 137.735 145.285 ;
        RECT 137.905 144.955 138.180 145.285 ;
        RECT 133.625 144.675 134.875 144.855 ;
        RECT 134.510 144.605 134.875 144.675 ;
        RECT 135.045 144.655 136.225 144.825 ;
        RECT 137.905 144.785 138.075 144.955 ;
        RECT 133.685 144.045 133.855 144.505 ;
        RECT 135.045 144.435 135.375 144.655 ;
        RECT 134.125 144.255 135.375 144.435 ;
        RECT 135.545 144.045 135.715 144.485 ;
        RECT 135.885 144.240 136.225 144.655 ;
        RECT 136.410 144.615 138.075 144.785 ;
        RECT 138.350 144.720 138.520 145.455 ;
        RECT 138.695 145.430 138.985 146.595 ;
        RECT 139.215 145.455 139.425 146.595 ;
        RECT 139.595 145.445 139.925 146.425 ;
        RECT 140.095 145.455 140.325 146.595 ;
        RECT 140.535 145.455 140.815 146.595 ;
        RECT 140.985 145.445 141.315 146.425 ;
        RECT 141.485 145.455 141.745 146.595 ;
        RECT 141.975 145.455 142.185 146.595 ;
        RECT 142.355 145.445 142.685 146.425 ;
        RECT 142.855 145.455 143.085 146.595 ;
        RECT 143.295 145.505 146.805 146.595 ;
        RECT 146.975 145.505 148.185 146.595 ;
        RECT 148.445 145.925 148.615 146.425 ;
        RECT 148.785 146.095 149.115 146.595 ;
        RECT 148.445 145.755 149.110 145.925 ;
        RECT 136.410 144.265 136.665 144.615 ;
        RECT 136.835 144.045 137.165 144.445 ;
        RECT 137.335 144.265 137.505 144.615 ;
        RECT 137.675 144.045 138.055 144.445 ;
        RECT 138.245 144.375 138.520 144.720 ;
        RECT 138.695 144.045 138.985 144.770 ;
        RECT 139.215 144.045 139.425 144.865 ;
        RECT 139.595 144.845 139.845 145.445 ;
        RECT 140.015 145.035 140.345 145.285 ;
        RECT 140.545 145.015 140.880 145.285 ;
        RECT 139.595 144.215 139.925 144.845 ;
        RECT 140.095 144.045 140.325 144.865 ;
        RECT 141.050 144.845 141.220 145.445 ;
        RECT 141.390 145.035 141.725 145.285 ;
        RECT 140.535 144.045 140.845 144.845 ;
        RECT 141.050 144.215 141.745 144.845 ;
        RECT 141.975 144.045 142.185 144.865 ;
        RECT 142.355 144.845 142.605 145.445 ;
        RECT 142.775 145.035 143.105 145.285 ;
        RECT 142.355 144.215 142.685 144.845 ;
        RECT 142.855 144.045 143.085 144.865 ;
        RECT 143.295 144.815 144.945 145.335 ;
        RECT 145.115 144.985 146.805 145.505 ;
        RECT 143.295 144.045 146.805 144.815 ;
        RECT 146.975 144.795 147.495 145.335 ;
        RECT 147.665 144.965 148.185 145.505 ;
        RECT 148.360 144.935 148.710 145.585 ;
        RECT 146.975 144.045 148.185 144.795 ;
        RECT 148.880 144.765 149.110 145.755 ;
        RECT 148.445 144.595 149.110 144.765 ;
        RECT 148.445 144.305 148.615 144.595 ;
        RECT 148.785 144.045 149.115 144.425 ;
        RECT 149.285 144.305 149.470 146.425 ;
        RECT 149.710 146.135 149.975 146.595 ;
        RECT 150.145 146.000 150.395 146.425 ;
        RECT 150.605 146.150 151.710 146.320 ;
        RECT 150.090 145.870 150.395 146.000 ;
        RECT 149.640 144.675 149.920 145.625 ;
        RECT 150.090 144.765 150.260 145.870 ;
        RECT 150.430 145.085 150.670 145.680 ;
        RECT 150.840 145.615 151.370 145.980 ;
        RECT 150.840 144.915 151.010 145.615 ;
        RECT 151.540 145.535 151.710 146.150 ;
        RECT 151.880 145.795 152.050 146.595 ;
        RECT 152.220 146.095 152.470 146.425 ;
        RECT 152.695 146.125 153.580 146.295 ;
        RECT 151.540 145.445 152.050 145.535 ;
        RECT 150.090 144.635 150.315 144.765 ;
        RECT 150.485 144.695 151.010 144.915 ;
        RECT 151.180 145.275 152.050 145.445 ;
        RECT 149.725 144.045 149.975 144.505 ;
        RECT 150.145 144.495 150.315 144.635 ;
        RECT 151.180 144.495 151.350 145.275 ;
        RECT 151.880 145.205 152.050 145.275 ;
        RECT 151.560 145.025 151.760 145.055 ;
        RECT 152.220 145.025 152.390 146.095 ;
        RECT 152.560 145.205 152.750 145.925 ;
        RECT 151.560 144.725 152.390 145.025 ;
        RECT 152.920 144.995 153.240 145.955 ;
        RECT 150.145 144.325 150.480 144.495 ;
        RECT 150.675 144.325 151.350 144.495 ;
        RECT 151.670 144.045 152.040 144.545 ;
        RECT 152.220 144.495 152.390 144.725 ;
        RECT 152.775 144.665 153.240 144.995 ;
        RECT 153.410 145.285 153.580 146.125 ;
        RECT 153.760 146.095 154.075 146.595 ;
        RECT 154.305 145.865 154.645 146.425 ;
        RECT 153.750 145.490 154.645 145.865 ;
        RECT 154.815 145.585 154.985 146.595 ;
        RECT 154.455 145.285 154.645 145.490 ;
        RECT 155.155 145.535 155.485 146.380 ;
        RECT 155.155 145.455 155.545 145.535 ;
        RECT 155.330 145.405 155.545 145.455 ;
        RECT 153.410 144.955 154.285 145.285 ;
        RECT 154.455 144.955 155.205 145.285 ;
        RECT 153.410 144.495 153.580 144.955 ;
        RECT 154.455 144.785 154.655 144.955 ;
        RECT 155.375 144.825 155.545 145.405 ;
        RECT 155.715 145.505 156.925 146.595 ;
        RECT 155.715 144.965 156.235 145.505 ;
        RECT 155.320 144.785 155.545 144.825 ;
        RECT 156.405 144.795 156.925 145.335 ;
        RECT 152.220 144.325 152.625 144.495 ;
        RECT 152.795 144.325 153.580 144.495 ;
        RECT 153.855 144.045 154.065 144.575 ;
        RECT 154.325 144.260 154.655 144.785 ;
        RECT 155.165 144.700 155.545 144.785 ;
        RECT 154.825 144.045 154.995 144.655 ;
        RECT 155.165 144.265 155.495 144.700 ;
        RECT 155.715 144.045 156.925 144.795 ;
        RECT 22.690 143.875 157.010 144.045 ;
        RECT 22.775 143.125 23.985 143.875 ;
        RECT 24.245 143.325 24.415 143.615 ;
        RECT 24.585 143.495 24.915 143.875 ;
        RECT 24.245 143.155 24.910 143.325 ;
        RECT 22.775 142.585 23.295 143.125 ;
        RECT 23.465 142.415 23.985 142.955 ;
        RECT 22.775 141.325 23.985 142.415 ;
        RECT 24.160 142.335 24.510 142.985 ;
        RECT 24.680 142.165 24.910 143.155 ;
        RECT 24.245 141.995 24.910 142.165 ;
        RECT 24.245 141.495 24.415 141.995 ;
        RECT 24.585 141.325 24.915 141.825 ;
        RECT 25.085 141.495 25.270 143.615 ;
        RECT 25.525 143.415 25.775 143.875 ;
        RECT 25.945 143.425 26.280 143.595 ;
        RECT 26.475 143.425 27.150 143.595 ;
        RECT 25.945 143.285 26.115 143.425 ;
        RECT 25.440 142.295 25.720 143.245 ;
        RECT 25.890 143.155 26.115 143.285 ;
        RECT 25.890 142.050 26.060 143.155 ;
        RECT 26.285 143.005 26.810 143.225 ;
        RECT 26.230 142.240 26.470 142.835 ;
        RECT 26.640 142.305 26.810 143.005 ;
        RECT 26.980 142.645 27.150 143.425 ;
        RECT 27.470 143.375 27.840 143.875 ;
        RECT 28.020 143.425 28.425 143.595 ;
        RECT 28.595 143.425 29.380 143.595 ;
        RECT 28.020 143.195 28.190 143.425 ;
        RECT 27.360 142.895 28.190 143.195 ;
        RECT 28.575 142.925 29.040 143.255 ;
        RECT 27.360 142.865 27.560 142.895 ;
        RECT 27.680 142.645 27.850 142.715 ;
        RECT 26.980 142.475 27.850 142.645 ;
        RECT 27.340 142.385 27.850 142.475 ;
        RECT 25.890 141.920 26.195 142.050 ;
        RECT 26.640 141.940 27.170 142.305 ;
        RECT 25.510 141.325 25.775 141.785 ;
        RECT 25.945 141.495 26.195 141.920 ;
        RECT 27.340 141.770 27.510 142.385 ;
        RECT 26.405 141.600 27.510 141.770 ;
        RECT 27.680 141.325 27.850 142.125 ;
        RECT 28.020 141.825 28.190 142.895 ;
        RECT 28.360 141.995 28.550 142.715 ;
        RECT 28.720 141.965 29.040 142.925 ;
        RECT 29.210 142.965 29.380 143.425 ;
        RECT 29.655 143.345 29.865 143.875 ;
        RECT 30.125 143.135 30.455 143.660 ;
        RECT 30.625 143.265 30.795 143.875 ;
        RECT 30.965 143.220 31.295 143.655 ;
        RECT 30.965 143.135 31.345 143.220 ;
        RECT 30.255 142.965 30.455 143.135 ;
        RECT 31.120 143.095 31.345 143.135 ;
        RECT 29.210 142.635 30.085 142.965 ;
        RECT 30.255 142.635 31.005 142.965 ;
        RECT 28.020 141.495 28.270 141.825 ;
        RECT 29.210 141.795 29.380 142.635 ;
        RECT 30.255 142.430 30.445 142.635 ;
        RECT 31.175 142.515 31.345 143.095 ;
        RECT 31.130 142.465 31.345 142.515 ;
        RECT 29.550 142.055 30.445 142.430 ;
        RECT 30.955 142.385 31.345 142.465 ;
        RECT 31.515 143.135 31.900 143.705 ;
        RECT 32.070 143.415 32.395 143.875 ;
        RECT 32.915 143.245 33.195 143.705 ;
        RECT 31.515 142.465 31.795 143.135 ;
        RECT 32.070 143.075 33.195 143.245 ;
        RECT 32.070 142.965 32.520 143.075 ;
        RECT 31.965 142.635 32.520 142.965 ;
        RECT 33.385 142.905 33.785 143.705 ;
        RECT 34.185 143.415 34.455 143.875 ;
        RECT 34.625 143.245 34.910 143.705 ;
        RECT 36.445 143.475 36.775 143.875 ;
        RECT 36.945 143.305 37.275 143.645 ;
        RECT 38.325 143.475 38.655 143.875 ;
        RECT 28.495 141.625 29.380 141.795 ;
        RECT 29.560 141.325 29.875 141.825 ;
        RECT 30.105 141.495 30.445 142.055 ;
        RECT 30.615 141.325 30.785 142.335 ;
        RECT 30.955 141.540 31.285 142.385 ;
        RECT 31.515 141.495 31.900 142.465 ;
        RECT 32.070 142.175 32.520 142.635 ;
        RECT 32.690 142.345 33.785 142.905 ;
        RECT 32.070 141.955 33.195 142.175 ;
        RECT 32.070 141.325 32.395 141.785 ;
        RECT 32.915 141.495 33.195 141.955 ;
        RECT 33.385 141.495 33.785 142.345 ;
        RECT 33.955 143.075 34.910 143.245 ;
        RECT 36.290 143.135 38.655 143.305 ;
        RECT 38.825 143.150 39.155 143.660 ;
        RECT 39.345 143.375 39.675 143.875 ;
        RECT 39.875 143.305 40.045 143.655 ;
        RECT 40.245 143.475 40.575 143.875 ;
        RECT 40.745 143.305 40.915 143.655 ;
        RECT 41.085 143.475 41.465 143.875 ;
        RECT 33.955 142.175 34.165 143.075 ;
        RECT 34.335 142.345 35.025 142.905 ;
        RECT 33.955 141.955 34.910 142.175 ;
        RECT 36.290 142.135 36.460 143.135 ;
        RECT 38.485 142.965 38.655 143.135 ;
        RECT 36.630 142.305 36.875 142.965 ;
        RECT 37.090 142.305 37.355 142.965 ;
        RECT 37.550 142.305 37.835 142.965 ;
        RECT 38.010 142.635 38.315 142.965 ;
        RECT 38.485 142.635 38.795 142.965 ;
        RECT 38.010 142.305 38.225 142.635 ;
        RECT 36.290 141.965 36.745 142.135 ;
        RECT 34.185 141.325 34.455 141.785 ;
        RECT 34.625 141.495 34.910 141.955 ;
        RECT 36.415 141.535 36.745 141.965 ;
        RECT 36.925 141.965 38.215 142.135 ;
        RECT 36.925 141.545 37.175 141.965 ;
        RECT 37.405 141.325 37.735 141.795 ;
        RECT 37.965 141.545 38.215 141.965 ;
        RECT 38.405 141.325 38.655 142.465 ;
        RECT 38.965 142.385 39.155 143.150 ;
        RECT 39.340 142.635 39.690 143.205 ;
        RECT 39.875 143.135 41.485 143.305 ;
        RECT 41.655 143.200 41.925 143.545 ;
        RECT 41.315 142.965 41.485 143.135 ;
        RECT 39.860 142.515 40.570 142.965 ;
        RECT 40.740 142.635 41.145 142.965 ;
        RECT 41.315 142.635 41.585 142.965 ;
        RECT 38.825 141.535 39.155 142.385 ;
        RECT 39.340 142.175 39.660 142.465 ;
        RECT 39.855 142.345 40.570 142.515 ;
        RECT 41.315 142.465 41.485 142.635 ;
        RECT 41.755 142.465 41.925 143.200 ;
        RECT 40.760 142.295 41.485 142.465 ;
        RECT 40.760 142.175 40.930 142.295 ;
        RECT 39.340 142.005 40.930 142.175 ;
        RECT 39.340 141.545 40.995 141.835 ;
        RECT 41.165 141.325 41.445 142.125 ;
        RECT 41.655 141.495 41.925 142.465 ;
        RECT 42.095 143.200 42.355 143.705 ;
        RECT 42.535 143.495 42.865 143.875 ;
        RECT 43.045 143.325 43.215 143.705 ;
        RECT 42.095 142.400 42.265 143.200 ;
        RECT 42.550 143.155 43.215 143.325 ;
        RECT 42.550 142.900 42.720 143.155 ;
        RECT 43.475 143.125 44.685 143.875 ;
        RECT 45.055 143.245 45.385 143.605 ;
        RECT 46.005 143.415 46.255 143.875 ;
        RECT 46.425 143.415 46.985 143.705 ;
        RECT 42.435 142.570 42.720 142.900 ;
        RECT 42.955 142.605 43.285 142.975 ;
        RECT 43.475 142.585 43.995 143.125 ;
        RECT 45.055 143.055 46.445 143.245 ;
        RECT 46.275 142.965 46.445 143.055 ;
        RECT 42.550 142.425 42.720 142.570 ;
        RECT 42.095 141.495 42.365 142.400 ;
        RECT 42.550 142.255 43.215 142.425 ;
        RECT 44.165 142.415 44.685 142.955 ;
        RECT 42.535 141.325 42.865 142.085 ;
        RECT 43.045 141.495 43.215 142.255 ;
        RECT 43.475 141.325 44.685 142.415 ;
        RECT 44.870 142.635 45.545 142.885 ;
        RECT 45.765 142.635 46.105 142.885 ;
        RECT 46.275 142.635 46.565 142.965 ;
        RECT 44.870 142.275 45.135 142.635 ;
        RECT 46.275 142.385 46.445 142.635 ;
        RECT 45.505 142.215 46.445 142.385 ;
        RECT 45.055 141.325 45.335 141.995 ;
        RECT 45.505 141.665 45.805 142.215 ;
        RECT 46.735 142.045 46.985 143.415 ;
        RECT 46.005 141.325 46.335 142.045 ;
        RECT 46.525 141.495 46.985 142.045 ;
        RECT 47.155 143.200 47.415 143.705 ;
        RECT 47.595 143.495 47.925 143.875 ;
        RECT 48.105 143.325 48.275 143.705 ;
        RECT 47.155 142.400 47.325 143.200 ;
        RECT 47.610 143.155 48.275 143.325 ;
        RECT 47.610 142.900 47.780 143.155 ;
        RECT 48.535 143.150 48.825 143.875 ;
        RECT 48.995 143.105 51.585 143.875 ;
        RECT 51.845 143.325 52.015 143.615 ;
        RECT 52.185 143.495 52.515 143.875 ;
        RECT 51.845 143.155 52.510 143.325 ;
        RECT 47.495 142.570 47.780 142.900 ;
        RECT 48.015 142.605 48.345 142.975 ;
        RECT 48.995 142.585 50.205 143.105 ;
        RECT 47.610 142.425 47.780 142.570 ;
        RECT 47.155 141.495 47.425 142.400 ;
        RECT 47.610 142.255 48.275 142.425 ;
        RECT 47.595 141.325 47.925 142.085 ;
        RECT 48.105 141.495 48.275 142.255 ;
        RECT 48.535 141.325 48.825 142.490 ;
        RECT 50.375 142.415 51.585 142.935 ;
        RECT 48.995 141.325 51.585 142.415 ;
        RECT 51.760 142.335 52.110 142.985 ;
        RECT 52.280 142.165 52.510 143.155 ;
        RECT 51.845 141.995 52.510 142.165 ;
        RECT 51.845 141.495 52.015 141.995 ;
        RECT 52.185 141.325 52.515 141.825 ;
        RECT 52.685 141.495 52.870 143.615 ;
        RECT 53.125 143.415 53.375 143.875 ;
        RECT 53.545 143.425 53.880 143.595 ;
        RECT 54.075 143.425 54.750 143.595 ;
        RECT 53.545 143.285 53.715 143.425 ;
        RECT 53.040 142.295 53.320 143.245 ;
        RECT 53.490 143.155 53.715 143.285 ;
        RECT 53.490 142.050 53.660 143.155 ;
        RECT 53.885 143.005 54.410 143.225 ;
        RECT 53.830 142.240 54.070 142.835 ;
        RECT 54.240 142.305 54.410 143.005 ;
        RECT 54.580 142.645 54.750 143.425 ;
        RECT 55.070 143.375 55.440 143.875 ;
        RECT 55.620 143.425 56.025 143.595 ;
        RECT 56.195 143.425 56.980 143.595 ;
        RECT 55.620 143.195 55.790 143.425 ;
        RECT 54.960 142.895 55.790 143.195 ;
        RECT 56.175 142.925 56.640 143.255 ;
        RECT 54.960 142.865 55.160 142.895 ;
        RECT 55.280 142.645 55.450 142.715 ;
        RECT 54.580 142.475 55.450 142.645 ;
        RECT 54.940 142.385 55.450 142.475 ;
        RECT 53.490 141.920 53.795 142.050 ;
        RECT 54.240 141.940 54.770 142.305 ;
        RECT 53.110 141.325 53.375 141.785 ;
        RECT 53.545 141.495 53.795 141.920 ;
        RECT 54.940 141.770 55.110 142.385 ;
        RECT 54.005 141.600 55.110 141.770 ;
        RECT 55.280 141.325 55.450 142.125 ;
        RECT 55.620 141.825 55.790 142.895 ;
        RECT 55.960 141.995 56.150 142.715 ;
        RECT 56.320 141.965 56.640 142.925 ;
        RECT 56.810 142.965 56.980 143.425 ;
        RECT 57.255 143.345 57.465 143.875 ;
        RECT 57.725 143.135 58.055 143.660 ;
        RECT 58.225 143.265 58.395 143.875 ;
        RECT 58.565 143.220 58.895 143.655 ;
        RECT 58.565 143.135 58.945 143.220 ;
        RECT 57.855 142.965 58.055 143.135 ;
        RECT 58.720 143.095 58.945 143.135 ;
        RECT 56.810 142.635 57.685 142.965 ;
        RECT 57.855 142.635 58.605 142.965 ;
        RECT 55.620 141.495 55.870 141.825 ;
        RECT 56.810 141.795 56.980 142.635 ;
        RECT 57.855 142.430 58.045 142.635 ;
        RECT 58.775 142.515 58.945 143.095 ;
        RECT 59.115 143.125 60.325 143.875 ;
        RECT 59.115 142.585 59.635 143.125 ;
        RECT 60.555 143.055 60.765 143.875 ;
        RECT 60.935 143.075 61.265 143.705 ;
        RECT 58.730 142.465 58.945 142.515 ;
        RECT 57.150 142.055 58.045 142.430 ;
        RECT 58.555 142.385 58.945 142.465 ;
        RECT 59.805 142.415 60.325 142.955 ;
        RECT 60.935 142.475 61.185 143.075 ;
        RECT 61.435 143.055 61.665 143.875 ;
        RECT 61.895 143.145 62.185 143.875 ;
        RECT 61.355 142.635 61.685 142.885 ;
        RECT 61.885 142.635 62.185 142.965 ;
        RECT 62.365 142.945 62.595 143.585 ;
        RECT 62.775 143.325 63.085 143.695 ;
        RECT 63.265 143.505 63.935 143.875 ;
        RECT 62.775 143.125 64.005 143.325 ;
        RECT 62.365 142.635 62.890 142.945 ;
        RECT 63.070 142.635 63.535 142.945 ;
        RECT 56.095 141.625 56.980 141.795 ;
        RECT 57.160 141.325 57.475 141.825 ;
        RECT 57.705 141.495 58.045 142.055 ;
        RECT 58.215 141.325 58.385 142.335 ;
        RECT 58.555 141.540 58.885 142.385 ;
        RECT 59.115 141.325 60.325 142.415 ;
        RECT 60.555 141.325 60.765 142.465 ;
        RECT 60.935 141.495 61.265 142.475 ;
        RECT 61.435 141.325 61.665 142.465 ;
        RECT 63.715 142.455 64.005 143.125 ;
        RECT 61.895 142.215 63.055 142.455 ;
        RECT 61.895 141.505 62.155 142.215 ;
        RECT 62.325 141.325 62.655 142.035 ;
        RECT 62.825 141.505 63.055 142.215 ;
        RECT 63.235 142.235 64.005 142.455 ;
        RECT 63.235 141.505 63.505 142.235 ;
        RECT 63.685 141.325 64.025 142.055 ;
        RECT 64.195 141.505 64.455 143.695 ;
        RECT 64.635 141.495 64.915 143.595 ;
        RECT 65.145 143.415 65.315 143.875 ;
        RECT 65.585 143.485 66.835 143.665 ;
        RECT 65.970 143.245 66.335 143.315 ;
        RECT 65.085 143.065 66.335 143.245 ;
        RECT 66.505 143.265 66.835 143.485 ;
        RECT 67.005 143.435 67.175 143.875 ;
        RECT 67.345 143.265 67.685 143.680 ;
        RECT 66.505 143.095 67.685 143.265 ;
        RECT 68.475 143.315 68.805 143.705 ;
        RECT 68.975 143.485 70.160 143.655 ;
        RECT 70.420 143.405 70.590 143.875 ;
        RECT 68.475 143.135 68.985 143.315 ;
        RECT 65.085 142.465 65.360 143.065 ;
        RECT 65.530 142.635 65.885 142.885 ;
        RECT 66.080 142.855 66.545 142.885 ;
        RECT 66.075 142.685 66.545 142.855 ;
        RECT 66.080 142.635 66.545 142.685 ;
        RECT 66.715 142.635 67.045 142.885 ;
        RECT 67.220 142.685 67.685 142.885 ;
        RECT 68.315 142.675 68.645 142.965 ;
        RECT 66.865 142.515 67.045 142.635 ;
        RECT 65.085 142.255 66.695 142.465 ;
        RECT 66.865 142.345 67.195 142.515 ;
        RECT 68.815 142.505 68.985 143.135 ;
        RECT 69.390 143.225 69.775 143.315 ;
        RECT 70.760 143.225 71.090 143.690 ;
        RECT 69.390 143.055 71.090 143.225 ;
        RECT 71.260 143.055 71.430 143.875 ;
        RECT 71.600 143.055 72.285 143.695 ;
        RECT 69.155 142.675 69.485 142.885 ;
        RECT 69.665 142.635 70.045 142.885 ;
        RECT 66.285 142.155 66.695 142.255 ;
        RECT 65.105 141.325 65.890 142.085 ;
        RECT 66.285 141.495 66.670 142.155 ;
        RECT 66.995 141.555 67.195 142.345 ;
        RECT 67.365 141.325 67.685 142.505 ;
        RECT 68.470 142.335 69.555 142.505 ;
        RECT 68.470 141.495 68.770 142.335 ;
        RECT 68.965 141.325 69.215 142.165 ;
        RECT 69.385 142.085 69.555 142.335 ;
        RECT 69.725 142.255 70.045 142.635 ;
        RECT 70.235 142.675 70.720 142.885 ;
        RECT 70.910 142.675 71.360 142.885 ;
        RECT 71.530 142.675 71.865 142.885 ;
        RECT 70.235 142.515 70.610 142.675 ;
        RECT 70.215 142.345 70.610 142.515 ;
        RECT 71.530 142.505 71.700 142.675 ;
        RECT 70.235 142.255 70.610 142.345 ;
        RECT 70.780 142.335 71.700 142.505 ;
        RECT 70.780 142.085 70.950 142.335 ;
        RECT 69.385 141.915 70.950 142.085 ;
        RECT 69.805 141.495 70.610 141.915 ;
        RECT 71.120 141.325 71.450 142.165 ;
        RECT 72.035 142.085 72.285 143.055 ;
        RECT 72.455 143.105 74.125 143.875 ;
        RECT 74.295 143.150 74.585 143.875 ;
        RECT 75.790 143.245 76.075 143.705 ;
        RECT 76.245 143.415 76.515 143.875 ;
        RECT 72.455 142.585 73.205 143.105 ;
        RECT 75.790 143.075 76.745 143.245 ;
        RECT 73.375 142.415 74.125 142.935 ;
        RECT 71.620 141.495 72.285 142.085 ;
        RECT 72.455 141.325 74.125 142.415 ;
        RECT 74.295 141.325 74.585 142.490 ;
        RECT 75.675 142.345 76.365 142.905 ;
        RECT 76.535 142.175 76.745 143.075 ;
        RECT 75.790 141.955 76.745 142.175 ;
        RECT 76.915 142.905 77.315 143.705 ;
        RECT 77.505 143.245 77.785 143.705 ;
        RECT 78.305 143.415 78.630 143.875 ;
        RECT 77.505 143.075 78.630 143.245 ;
        RECT 78.800 143.135 79.185 143.705 ;
        RECT 79.405 143.220 79.735 143.655 ;
        RECT 79.905 143.265 80.075 143.875 ;
        RECT 78.180 142.965 78.630 143.075 ;
        RECT 76.915 142.345 78.010 142.905 ;
        RECT 78.180 142.635 78.735 142.965 ;
        RECT 75.790 141.495 76.075 141.955 ;
        RECT 76.245 141.325 76.515 141.785 ;
        RECT 76.915 141.495 77.315 142.345 ;
        RECT 78.180 142.175 78.630 142.635 ;
        RECT 78.905 142.465 79.185 143.135 ;
        RECT 77.505 141.955 78.630 142.175 ;
        RECT 77.505 141.495 77.785 141.955 ;
        RECT 78.305 141.325 78.630 141.785 ;
        RECT 78.800 141.495 79.185 142.465 ;
        RECT 79.355 143.135 79.735 143.220 ;
        RECT 80.245 143.135 80.575 143.660 ;
        RECT 80.835 143.345 81.045 143.875 ;
        RECT 81.320 143.425 82.105 143.595 ;
        RECT 82.275 143.425 82.680 143.595 ;
        RECT 79.355 143.095 79.580 143.135 ;
        RECT 79.355 142.515 79.525 143.095 ;
        RECT 80.245 142.965 80.445 143.135 ;
        RECT 81.320 142.965 81.490 143.425 ;
        RECT 79.695 142.635 80.445 142.965 ;
        RECT 80.615 142.635 81.490 142.965 ;
        RECT 79.355 142.465 79.570 142.515 ;
        RECT 79.355 142.385 79.745 142.465 ;
        RECT 79.415 141.540 79.745 142.385 ;
        RECT 80.255 142.430 80.445 142.635 ;
        RECT 79.915 141.325 80.085 142.335 ;
        RECT 80.255 142.055 81.150 142.430 ;
        RECT 80.255 141.495 80.595 142.055 ;
        RECT 80.825 141.325 81.140 141.825 ;
        RECT 81.320 141.795 81.490 142.635 ;
        RECT 81.660 142.925 82.125 143.255 ;
        RECT 82.510 143.195 82.680 143.425 ;
        RECT 82.860 143.375 83.230 143.875 ;
        RECT 83.550 143.425 84.225 143.595 ;
        RECT 84.420 143.425 84.755 143.595 ;
        RECT 81.660 141.965 81.980 142.925 ;
        RECT 82.510 142.895 83.340 143.195 ;
        RECT 82.150 141.995 82.340 142.715 ;
        RECT 82.510 141.825 82.680 142.895 ;
        RECT 83.140 142.865 83.340 142.895 ;
        RECT 82.850 142.645 83.020 142.715 ;
        RECT 83.550 142.645 83.720 143.425 ;
        RECT 84.585 143.285 84.755 143.425 ;
        RECT 84.925 143.415 85.175 143.875 ;
        RECT 82.850 142.475 83.720 142.645 ;
        RECT 83.890 143.005 84.415 143.225 ;
        RECT 84.585 143.155 84.810 143.285 ;
        RECT 82.850 142.385 83.360 142.475 ;
        RECT 81.320 141.625 82.205 141.795 ;
        RECT 82.430 141.495 82.680 141.825 ;
        RECT 82.850 141.325 83.020 142.125 ;
        RECT 83.190 141.770 83.360 142.385 ;
        RECT 83.890 142.305 84.060 143.005 ;
        RECT 83.530 141.940 84.060 142.305 ;
        RECT 84.230 142.240 84.470 142.835 ;
        RECT 84.640 142.050 84.810 143.155 ;
        RECT 84.980 142.295 85.260 143.245 ;
        RECT 84.505 141.920 84.810 142.050 ;
        RECT 83.190 141.600 84.295 141.770 ;
        RECT 84.505 141.495 84.755 141.920 ;
        RECT 84.925 141.325 85.190 141.785 ;
        RECT 85.430 141.495 85.615 143.615 ;
        RECT 85.785 143.495 86.115 143.875 ;
        RECT 86.285 143.325 86.455 143.615 ;
        RECT 85.790 143.155 86.455 143.325 ;
        RECT 85.790 142.165 86.020 143.155 ;
        RECT 86.720 143.110 87.175 143.875 ;
        RECT 87.450 143.495 88.750 143.705 ;
        RECT 89.005 143.515 89.335 143.875 ;
        RECT 88.580 143.345 88.750 143.495 ;
        RECT 89.505 143.375 89.765 143.705 ;
        RECT 89.960 143.475 90.290 143.875 ;
        RECT 86.190 142.335 86.540 142.985 ;
        RECT 87.650 142.885 87.870 143.285 ;
        RECT 86.715 142.685 87.205 142.885 ;
        RECT 87.395 142.675 87.870 142.885 ;
        RECT 88.115 142.885 88.325 143.285 ;
        RECT 88.580 143.220 89.335 143.345 ;
        RECT 88.580 143.175 89.425 143.220 ;
        RECT 89.155 143.055 89.425 143.175 ;
        RECT 88.115 142.675 88.445 142.885 ;
        RECT 88.615 142.615 89.025 142.920 ;
        RECT 86.720 142.445 87.895 142.505 ;
        RECT 89.255 142.480 89.425 143.055 ;
        RECT 89.225 142.445 89.425 142.480 ;
        RECT 86.720 142.335 89.425 142.445 ;
        RECT 85.790 141.995 86.455 142.165 ;
        RECT 85.785 141.325 86.115 141.825 ;
        RECT 86.285 141.495 86.455 141.995 ;
        RECT 86.720 141.715 86.975 142.335 ;
        RECT 87.565 142.275 89.365 142.335 ;
        RECT 87.565 142.245 87.895 142.275 ;
        RECT 89.595 142.175 89.765 143.375 ;
        RECT 90.460 143.305 90.630 143.575 ;
        RECT 90.800 143.365 91.115 143.875 ;
        RECT 91.345 143.365 91.635 143.705 ;
        RECT 91.805 143.365 92.045 143.875 ;
        RECT 87.225 142.075 87.410 142.165 ;
        RECT 88.000 142.075 88.835 142.085 ;
        RECT 87.225 141.875 88.835 142.075 ;
        RECT 87.225 141.835 87.455 141.875 ;
        RECT 86.720 141.495 87.055 141.715 ;
        RECT 88.060 141.325 88.415 141.705 ;
        RECT 88.585 141.495 88.835 141.875 ;
        RECT 89.085 141.325 89.335 142.105 ;
        RECT 89.505 141.495 89.765 142.175 ;
        RECT 89.935 143.135 90.630 143.305 ;
        RECT 89.935 142.125 90.365 143.135 ;
        RECT 90.535 142.465 90.705 142.965 ;
        RECT 90.875 142.635 91.285 143.195 ;
        RECT 91.455 142.465 91.635 143.365 ;
        RECT 91.805 142.855 92.000 143.195 ;
        RECT 92.235 143.075 92.930 143.705 ;
        RECT 93.135 143.075 93.445 143.875 ;
        RECT 94.075 143.200 94.345 143.545 ;
        RECT 94.535 143.475 94.915 143.875 ;
        RECT 95.085 143.305 95.255 143.655 ;
        RECT 95.425 143.395 96.160 143.875 ;
        RECT 91.805 142.685 92.005 142.855 ;
        RECT 91.805 142.635 92.000 142.685 ;
        RECT 92.255 142.635 92.590 142.885 ;
        RECT 92.760 142.475 92.930 143.075 ;
        RECT 93.100 142.635 93.435 142.905 ;
        RECT 90.535 142.295 91.995 142.465 ;
        RECT 89.935 141.955 90.710 142.125 ;
        RECT 90.040 141.325 90.210 141.785 ;
        RECT 90.380 141.495 90.710 141.955 ;
        RECT 90.880 141.325 91.050 142.125 ;
        RECT 91.635 142.120 91.995 142.295 ;
        RECT 92.235 141.325 92.495 142.465 ;
        RECT 92.665 141.495 92.995 142.475 ;
        RECT 94.075 142.465 94.245 143.200 ;
        RECT 94.515 143.135 95.255 143.305 ;
        RECT 96.330 143.225 96.640 143.695 ;
        RECT 94.515 142.965 94.685 143.135 ;
        RECT 95.905 143.055 96.640 143.225 ;
        RECT 96.835 143.055 97.095 143.875 ;
        RECT 97.265 143.055 97.595 143.475 ;
        RECT 97.775 143.390 98.565 143.655 ;
        RECT 95.905 142.965 96.155 143.055 ;
        RECT 94.455 142.635 94.685 142.965 ;
        RECT 95.415 142.635 96.155 142.965 ;
        RECT 97.345 142.965 97.595 143.055 ;
        RECT 96.325 142.635 96.660 142.885 ;
        RECT 94.515 142.465 94.685 142.635 ;
        RECT 93.165 141.325 93.445 142.465 ;
        RECT 94.075 141.495 94.345 142.465 ;
        RECT 94.515 142.295 95.760 142.465 ;
        RECT 94.555 141.325 94.835 142.125 ;
        RECT 95.340 142.045 95.760 142.295 ;
        RECT 95.985 142.075 96.155 142.635 ;
        RECT 95.015 141.545 96.210 141.875 ;
        RECT 96.405 141.325 96.660 142.465 ;
        RECT 96.835 142.005 97.175 142.885 ;
        RECT 97.345 142.715 98.140 142.965 ;
        RECT 96.835 141.325 97.095 141.835 ;
        RECT 97.345 141.495 97.515 142.715 ;
        RECT 98.310 142.535 98.565 143.390 ;
        RECT 98.735 143.235 98.935 143.655 ;
        RECT 99.125 143.415 99.455 143.875 ;
        RECT 98.735 142.715 99.145 143.235 ;
        RECT 99.625 143.225 99.885 143.705 ;
        RECT 99.315 142.535 99.545 142.965 ;
        RECT 97.755 142.365 99.545 142.535 ;
        RECT 97.755 142.000 98.005 142.365 ;
        RECT 98.175 142.005 98.505 142.195 ;
        RECT 98.725 142.070 99.440 142.365 ;
        RECT 99.715 142.195 99.885 143.225 ;
        RECT 100.055 143.150 100.345 143.875 ;
        RECT 100.515 143.125 101.725 143.875 ;
        RECT 100.515 142.585 101.035 143.125 ;
        RECT 102.000 143.115 102.255 143.875 ;
        RECT 102.465 143.235 102.635 143.515 ;
        RECT 102.465 143.065 102.815 143.235 ;
        RECT 102.985 143.065 103.155 143.875 ;
        RECT 103.325 143.235 103.655 143.705 ;
        RECT 103.825 143.405 103.995 143.875 ;
        RECT 104.165 143.235 104.495 143.705 ;
        RECT 103.325 143.065 104.495 143.235 ;
        RECT 104.665 143.065 104.945 143.875 ;
        RECT 105.115 143.375 105.415 143.705 ;
        RECT 105.585 143.395 105.860 143.875 ;
        RECT 98.175 141.830 98.370 142.005 ;
        RECT 97.755 141.325 98.370 141.830 ;
        RECT 98.540 141.495 99.015 141.835 ;
        RECT 99.185 141.325 99.400 141.870 ;
        RECT 99.610 141.495 99.885 142.195 ;
        RECT 100.055 141.325 100.345 142.490 ;
        RECT 101.205 142.415 101.725 142.955 ;
        RECT 100.515 141.325 101.725 142.415 ;
        RECT 101.905 142.685 102.430 142.895 ;
        RECT 102.600 142.885 102.815 143.065 ;
        RECT 102.600 142.715 103.155 142.885 ;
        RECT 101.905 141.995 102.120 142.685 ;
        RECT 102.600 142.515 102.770 142.715 ;
        RECT 102.465 142.345 102.770 142.515 ;
        RECT 102.005 141.325 102.255 141.815 ;
        RECT 102.465 141.500 102.635 142.345 ;
        RECT 102.940 142.070 103.195 142.515 ;
        RECT 102.905 141.665 103.195 142.070 ;
        RECT 103.365 141.835 103.615 143.065 ;
        RECT 103.795 143.025 103.965 143.065 ;
        RECT 104.110 142.685 104.550 142.895 ;
        RECT 103.785 142.305 104.945 142.515 ;
        RECT 103.785 141.665 104.035 142.305 ;
        RECT 102.905 141.495 104.035 141.665 ;
        RECT 104.205 141.325 104.455 142.135 ;
        RECT 104.625 141.495 104.945 142.305 ;
        RECT 105.115 142.465 105.285 143.375 ;
        RECT 106.040 143.225 106.335 143.615 ;
        RECT 106.505 143.395 106.760 143.875 ;
        RECT 106.935 143.225 107.195 143.615 ;
        RECT 107.365 143.395 107.645 143.875 ;
        RECT 105.455 142.635 105.805 143.205 ;
        RECT 106.040 143.055 107.690 143.225 ;
        RECT 105.975 142.715 107.115 142.885 ;
        RECT 105.975 142.465 106.145 142.715 ;
        RECT 107.285 142.545 107.690 143.055 ;
        RECT 105.115 142.295 106.145 142.465 ;
        RECT 106.935 142.375 107.690 142.545 ;
        RECT 107.875 143.200 108.135 143.705 ;
        RECT 108.315 143.495 108.645 143.875 ;
        RECT 108.825 143.325 108.995 143.705 ;
        RECT 107.875 142.400 108.045 143.200 ;
        RECT 108.330 143.155 108.995 143.325 ;
        RECT 108.330 142.900 108.500 143.155 ;
        RECT 109.255 143.105 110.925 143.875 ;
        RECT 111.555 143.415 112.115 143.705 ;
        RECT 112.285 143.415 112.535 143.875 ;
        RECT 108.215 142.570 108.500 142.900 ;
        RECT 108.735 142.605 109.065 142.975 ;
        RECT 109.255 142.585 110.005 143.105 ;
        RECT 108.330 142.425 108.500 142.570 ;
        RECT 105.115 141.495 105.425 142.295 ;
        RECT 106.935 142.125 107.195 142.375 ;
        RECT 105.595 141.325 105.905 142.125 ;
        RECT 106.075 141.955 107.195 142.125 ;
        RECT 106.075 141.495 106.335 141.955 ;
        RECT 106.505 141.325 106.760 141.785 ;
        RECT 106.935 141.495 107.195 141.955 ;
        RECT 107.365 141.325 107.650 142.195 ;
        RECT 107.875 141.495 108.145 142.400 ;
        RECT 108.330 142.255 108.995 142.425 ;
        RECT 110.175 142.415 110.925 142.935 ;
        RECT 108.315 141.325 108.645 142.085 ;
        RECT 108.825 141.495 108.995 142.255 ;
        RECT 109.255 141.325 110.925 142.415 ;
        RECT 111.555 142.045 111.805 143.415 ;
        RECT 113.155 143.245 113.485 143.605 ;
        RECT 112.095 143.055 113.485 143.245 ;
        RECT 113.855 143.125 115.065 143.875 ;
        RECT 115.325 143.325 115.495 143.705 ;
        RECT 115.675 143.495 116.005 143.875 ;
        RECT 115.325 143.155 115.990 143.325 ;
        RECT 116.185 143.200 116.445 143.705 ;
        RECT 112.095 142.965 112.265 143.055 ;
        RECT 111.975 142.635 112.265 142.965 ;
        RECT 112.435 142.635 112.775 142.885 ;
        RECT 112.995 142.635 113.670 142.885 ;
        RECT 112.095 142.385 112.265 142.635 ;
        RECT 112.095 142.215 113.035 142.385 ;
        RECT 113.405 142.275 113.670 142.635 ;
        RECT 113.855 142.585 114.375 143.125 ;
        RECT 114.545 142.415 115.065 142.955 ;
        RECT 115.255 142.605 115.585 142.975 ;
        RECT 115.820 142.900 115.990 143.155 ;
        RECT 115.820 142.570 116.105 142.900 ;
        RECT 115.820 142.425 115.990 142.570 ;
        RECT 111.555 141.495 112.015 142.045 ;
        RECT 112.205 141.325 112.535 142.045 ;
        RECT 112.735 141.665 113.035 142.215 ;
        RECT 113.205 141.325 113.485 141.995 ;
        RECT 113.855 141.325 115.065 142.415 ;
        RECT 115.325 142.255 115.990 142.425 ;
        RECT 116.275 142.400 116.445 143.200 ;
        RECT 116.615 143.125 117.825 143.875 ;
        RECT 117.995 143.415 118.555 143.705 ;
        RECT 118.725 143.415 118.975 143.875 ;
        RECT 116.615 142.585 117.135 143.125 ;
        RECT 117.305 142.415 117.825 142.955 ;
        RECT 115.325 141.495 115.495 142.255 ;
        RECT 115.675 141.325 116.005 142.085 ;
        RECT 116.175 141.495 116.445 142.400 ;
        RECT 116.615 141.325 117.825 142.415 ;
        RECT 117.995 142.045 118.245 143.415 ;
        RECT 119.595 143.245 119.925 143.605 ;
        RECT 120.295 143.330 125.640 143.875 ;
        RECT 118.535 143.055 119.925 143.245 ;
        RECT 118.535 142.965 118.705 143.055 ;
        RECT 118.415 142.635 118.705 142.965 ;
        RECT 118.875 142.635 119.215 142.885 ;
        RECT 119.435 142.635 120.110 142.885 ;
        RECT 118.535 142.385 118.705 142.635 ;
        RECT 118.535 142.215 119.475 142.385 ;
        RECT 119.845 142.275 120.110 142.635 ;
        RECT 121.880 142.500 122.220 143.330 ;
        RECT 125.815 143.150 126.105 143.875 ;
        RECT 126.475 143.245 126.805 143.605 ;
        RECT 127.425 143.415 127.675 143.875 ;
        RECT 127.845 143.415 128.405 143.705 ;
        RECT 126.475 143.055 127.865 143.245 ;
        RECT 117.995 141.495 118.455 142.045 ;
        RECT 118.645 141.325 118.975 142.045 ;
        RECT 119.175 141.665 119.475 142.215 ;
        RECT 119.645 141.325 119.925 141.995 ;
        RECT 123.700 141.760 124.050 143.010 ;
        RECT 127.695 142.965 127.865 143.055 ;
        RECT 126.290 142.635 126.965 142.885 ;
        RECT 127.185 142.635 127.525 142.885 ;
        RECT 127.695 142.635 127.985 142.965 ;
        RECT 120.295 141.325 125.640 141.760 ;
        RECT 125.815 141.325 126.105 142.490 ;
        RECT 126.290 142.275 126.555 142.635 ;
        RECT 127.695 142.385 127.865 142.635 ;
        RECT 126.925 142.215 127.865 142.385 ;
        RECT 126.475 141.325 126.755 141.995 ;
        RECT 126.925 141.665 127.225 142.215 ;
        RECT 128.155 142.045 128.405 143.415 ;
        RECT 128.575 143.105 130.245 143.875 ;
        RECT 128.575 142.585 129.325 143.105 ;
        RECT 129.495 142.415 130.245 142.935 ;
        RECT 127.425 141.325 127.755 142.045 ;
        RECT 127.945 141.495 128.405 142.045 ;
        RECT 128.575 141.325 130.245 142.415 ;
        RECT 130.875 141.495 131.155 143.595 ;
        RECT 131.385 143.415 131.555 143.875 ;
        RECT 131.825 143.485 133.075 143.665 ;
        RECT 132.210 143.245 132.575 143.315 ;
        RECT 131.325 143.065 132.575 143.245 ;
        RECT 132.745 143.265 133.075 143.485 ;
        RECT 133.245 143.435 133.415 143.875 ;
        RECT 133.585 143.265 133.925 143.680 ;
        RECT 132.745 143.095 133.925 143.265 ;
        RECT 131.325 142.465 131.600 143.065 ;
        RECT 135.075 143.055 135.285 143.875 ;
        RECT 135.455 143.075 135.785 143.705 ;
        RECT 131.770 142.635 132.125 142.885 ;
        RECT 132.320 142.855 132.785 142.885 ;
        RECT 132.315 142.685 132.785 142.855 ;
        RECT 132.320 142.635 132.785 142.685 ;
        RECT 132.955 142.635 133.285 142.885 ;
        RECT 133.460 142.685 133.925 142.885 ;
        RECT 133.105 142.515 133.285 142.635 ;
        RECT 131.325 142.255 132.935 142.465 ;
        RECT 133.105 142.345 133.435 142.515 ;
        RECT 132.525 142.155 132.935 142.255 ;
        RECT 131.345 141.325 132.130 142.085 ;
        RECT 132.525 141.495 132.910 142.155 ;
        RECT 133.235 141.555 133.435 142.345 ;
        RECT 133.605 141.325 133.925 142.505 ;
        RECT 135.455 142.475 135.705 143.075 ;
        RECT 135.955 143.055 136.185 143.875 ;
        RECT 136.395 143.105 138.985 143.875 ;
        RECT 135.875 142.635 136.205 142.885 ;
        RECT 136.395 142.585 137.605 143.105 ;
        RECT 139.615 143.075 140.310 143.705 ;
        RECT 140.515 143.075 140.825 143.875 ;
        RECT 140.995 143.495 141.885 143.665 ;
        RECT 135.075 141.325 135.285 142.465 ;
        RECT 135.455 141.495 135.785 142.475 ;
        RECT 135.955 141.325 136.185 142.465 ;
        RECT 137.775 142.415 138.985 142.935 ;
        RECT 139.635 142.635 139.970 142.885 ;
        RECT 140.140 142.475 140.310 143.075 ;
        RECT 140.995 142.940 141.545 143.325 ;
        RECT 140.480 142.635 140.815 142.905 ;
        RECT 141.715 142.770 141.885 143.495 ;
        RECT 140.995 142.700 141.885 142.770 ;
        RECT 142.055 143.170 142.275 143.655 ;
        RECT 142.445 143.335 142.695 143.875 ;
        RECT 142.865 143.225 143.125 143.705 ;
        RECT 143.920 143.365 144.160 143.875 ;
        RECT 144.340 143.365 144.620 143.695 ;
        RECT 144.850 143.365 145.065 143.875 ;
        RECT 142.055 142.745 142.385 143.170 ;
        RECT 140.995 142.675 141.890 142.700 ;
        RECT 140.995 142.660 141.900 142.675 ;
        RECT 140.995 142.645 141.905 142.660 ;
        RECT 140.995 142.640 141.915 142.645 ;
        RECT 140.995 142.630 141.920 142.640 ;
        RECT 140.995 142.620 141.925 142.630 ;
        RECT 140.995 142.615 141.935 142.620 ;
        RECT 140.995 142.605 141.945 142.615 ;
        RECT 140.995 142.600 141.955 142.605 ;
        RECT 136.395 141.325 138.985 142.415 ;
        RECT 139.615 141.325 139.875 142.465 ;
        RECT 140.045 141.495 140.375 142.475 ;
        RECT 140.545 141.325 140.825 142.465 ;
        RECT 140.995 142.150 141.255 142.600 ;
        RECT 141.620 142.595 141.955 142.600 ;
        RECT 141.620 142.590 141.970 142.595 ;
        RECT 141.620 142.580 141.985 142.590 ;
        RECT 141.620 142.575 142.010 142.580 ;
        RECT 142.555 142.575 142.785 142.970 ;
        RECT 141.620 142.570 142.785 142.575 ;
        RECT 141.650 142.535 142.785 142.570 ;
        RECT 141.685 142.510 142.785 142.535 ;
        RECT 141.715 142.480 142.785 142.510 ;
        RECT 141.735 142.450 142.785 142.480 ;
        RECT 141.755 142.420 142.785 142.450 ;
        RECT 141.825 142.410 142.785 142.420 ;
        RECT 141.850 142.400 142.785 142.410 ;
        RECT 141.870 142.385 142.785 142.400 ;
        RECT 141.890 142.370 142.785 142.385 ;
        RECT 141.895 142.360 142.680 142.370 ;
        RECT 141.910 142.325 142.680 142.360 ;
        RECT 141.425 142.005 141.755 142.250 ;
        RECT 141.925 142.075 142.680 142.325 ;
        RECT 142.955 142.195 143.125 143.225 ;
        RECT 143.815 142.635 144.170 143.195 ;
        RECT 144.340 142.465 144.510 143.365 ;
        RECT 144.680 142.635 144.945 143.195 ;
        RECT 145.235 143.135 145.850 143.705 ;
        RECT 146.055 143.495 146.945 143.665 ;
        RECT 145.195 142.465 145.365 142.965 ;
        RECT 141.425 141.980 141.610 142.005 ;
        RECT 140.995 141.880 141.610 141.980 ;
        RECT 140.995 141.325 141.600 141.880 ;
        RECT 141.775 141.495 142.255 141.835 ;
        RECT 142.425 141.325 142.680 141.870 ;
        RECT 142.850 141.495 143.125 142.195 ;
        RECT 143.940 142.295 145.365 142.465 ;
        RECT 143.940 142.120 144.330 142.295 ;
        RECT 144.815 141.325 145.145 142.125 ;
        RECT 145.535 142.115 145.850 143.135 ;
        RECT 146.055 142.940 146.605 143.325 ;
        RECT 146.775 142.770 146.945 143.495 ;
        RECT 146.055 142.700 146.945 142.770 ;
        RECT 147.115 143.170 147.335 143.655 ;
        RECT 147.505 143.335 147.755 143.875 ;
        RECT 147.925 143.225 148.185 143.705 ;
        RECT 147.115 142.745 147.445 143.170 ;
        RECT 146.055 142.675 146.950 142.700 ;
        RECT 146.055 142.660 146.960 142.675 ;
        RECT 146.055 142.645 146.965 142.660 ;
        RECT 146.055 142.640 146.975 142.645 ;
        RECT 146.055 142.630 146.980 142.640 ;
        RECT 146.055 142.620 146.985 142.630 ;
        RECT 146.055 142.615 146.995 142.620 ;
        RECT 146.055 142.605 147.005 142.615 ;
        RECT 146.055 142.600 147.015 142.605 ;
        RECT 146.055 142.150 146.315 142.600 ;
        RECT 146.680 142.595 147.015 142.600 ;
        RECT 146.680 142.590 147.030 142.595 ;
        RECT 146.680 142.580 147.045 142.590 ;
        RECT 146.680 142.575 147.070 142.580 ;
        RECT 147.615 142.575 147.845 142.970 ;
        RECT 146.680 142.570 147.845 142.575 ;
        RECT 146.710 142.535 147.845 142.570 ;
        RECT 146.745 142.510 147.845 142.535 ;
        RECT 146.775 142.480 147.845 142.510 ;
        RECT 146.795 142.450 147.845 142.480 ;
        RECT 146.815 142.420 147.845 142.450 ;
        RECT 146.885 142.410 147.845 142.420 ;
        RECT 146.910 142.400 147.845 142.410 ;
        RECT 146.930 142.385 147.845 142.400 ;
        RECT 146.950 142.370 147.845 142.385 ;
        RECT 146.955 142.360 147.740 142.370 ;
        RECT 146.970 142.325 147.740 142.360 ;
        RECT 145.315 141.495 145.850 142.115 ;
        RECT 146.485 142.005 146.815 142.250 ;
        RECT 146.985 142.075 147.740 142.325 ;
        RECT 148.015 142.195 148.185 143.225 ;
        RECT 148.445 143.325 148.615 143.705 ;
        RECT 148.795 143.495 149.125 143.875 ;
        RECT 148.445 143.155 149.110 143.325 ;
        RECT 149.305 143.200 149.565 143.705 ;
        RECT 148.375 142.605 148.705 142.975 ;
        RECT 148.940 142.900 149.110 143.155 ;
        RECT 148.940 142.570 149.225 142.900 ;
        RECT 148.940 142.425 149.110 142.570 ;
        RECT 146.485 141.980 146.670 142.005 ;
        RECT 146.055 141.880 146.670 141.980 ;
        RECT 146.055 141.325 146.660 141.880 ;
        RECT 146.835 141.495 147.315 141.835 ;
        RECT 147.485 141.325 147.740 141.870 ;
        RECT 147.910 141.495 148.185 142.195 ;
        RECT 148.445 142.255 149.110 142.425 ;
        RECT 149.395 142.400 149.565 143.200 ;
        RECT 149.735 143.105 151.405 143.875 ;
        RECT 151.575 143.150 151.865 143.875 ;
        RECT 152.035 143.105 155.545 143.875 ;
        RECT 155.715 143.125 156.925 143.875 ;
        RECT 149.735 142.585 150.485 143.105 ;
        RECT 150.655 142.415 151.405 142.935 ;
        RECT 152.035 142.585 153.685 143.105 ;
        RECT 148.445 141.495 148.615 142.255 ;
        RECT 148.795 141.325 149.125 142.085 ;
        RECT 149.295 141.495 149.565 142.400 ;
        RECT 149.735 141.325 151.405 142.415 ;
        RECT 151.575 141.325 151.865 142.490 ;
        RECT 153.855 142.415 155.545 142.935 ;
        RECT 152.035 141.325 155.545 142.415 ;
        RECT 155.715 142.415 156.235 142.955 ;
        RECT 156.405 142.585 156.925 143.125 ;
        RECT 155.715 141.325 156.925 142.415 ;
        RECT 22.690 141.155 157.010 141.325 ;
        RECT 22.775 140.065 23.985 141.155 ;
        RECT 24.155 140.065 26.745 141.155 ;
        RECT 22.775 139.355 23.295 139.895 ;
        RECT 23.465 139.525 23.985 140.065 ;
        RECT 24.155 139.375 25.365 139.895 ;
        RECT 25.535 139.545 26.745 140.065 ;
        RECT 26.915 139.550 27.195 140.985 ;
        RECT 27.365 140.380 28.075 141.155 ;
        RECT 28.245 140.210 28.575 140.985 ;
        RECT 27.425 139.995 28.575 140.210 ;
        RECT 22.775 138.605 23.985 139.355 ;
        RECT 24.155 138.605 26.745 139.375 ;
        RECT 26.915 138.775 27.255 139.550 ;
        RECT 27.425 139.425 27.710 139.995 ;
        RECT 27.895 139.595 28.365 139.825 ;
        RECT 28.770 139.795 28.985 140.910 ;
        RECT 29.165 140.435 29.495 141.155 ;
        RECT 29.275 139.795 29.505 140.135 ;
        RECT 29.675 140.065 32.265 141.155 ;
        RECT 28.535 139.615 28.985 139.795 ;
        RECT 28.535 139.595 28.865 139.615 ;
        RECT 29.175 139.595 29.505 139.795 ;
        RECT 27.425 139.235 28.135 139.425 ;
        RECT 27.835 139.095 28.135 139.235 ;
        RECT 28.325 139.235 29.505 139.425 ;
        RECT 28.325 139.155 28.655 139.235 ;
        RECT 27.835 139.085 28.150 139.095 ;
        RECT 27.835 139.075 28.160 139.085 ;
        RECT 27.835 139.070 28.170 139.075 ;
        RECT 27.425 138.605 27.595 139.065 ;
        RECT 27.835 139.060 28.175 139.070 ;
        RECT 27.835 139.055 28.180 139.060 ;
        RECT 27.835 139.045 28.185 139.055 ;
        RECT 27.835 139.040 28.190 139.045 ;
        RECT 27.835 138.775 28.195 139.040 ;
        RECT 28.825 138.605 28.995 139.065 ;
        RECT 29.165 138.775 29.505 139.235 ;
        RECT 29.675 139.375 30.885 139.895 ;
        RECT 31.055 139.545 32.265 140.065 ;
        RECT 32.895 140.285 33.170 140.985 ;
        RECT 33.340 140.610 33.595 141.155 ;
        RECT 33.765 140.645 34.245 140.985 ;
        RECT 34.420 140.600 35.025 141.155 ;
        RECT 34.410 140.500 35.025 140.600 ;
        RECT 34.410 140.475 34.595 140.500 ;
        RECT 29.675 138.605 32.265 139.375 ;
        RECT 32.895 139.255 33.065 140.285 ;
        RECT 33.340 140.155 34.095 140.405 ;
        RECT 34.265 140.230 34.595 140.475 ;
        RECT 33.340 140.120 34.110 140.155 ;
        RECT 33.340 140.110 34.125 140.120 ;
        RECT 33.235 140.095 34.130 140.110 ;
        RECT 33.235 140.080 34.150 140.095 ;
        RECT 33.235 140.070 34.170 140.080 ;
        RECT 33.235 140.060 34.195 140.070 ;
        RECT 33.235 140.030 34.265 140.060 ;
        RECT 33.235 140.000 34.285 140.030 ;
        RECT 33.235 139.970 34.305 140.000 ;
        RECT 33.235 139.945 34.335 139.970 ;
        RECT 33.235 139.910 34.370 139.945 ;
        RECT 33.235 139.905 34.400 139.910 ;
        RECT 33.235 139.510 33.465 139.905 ;
        RECT 34.010 139.900 34.400 139.905 ;
        RECT 34.035 139.890 34.400 139.900 ;
        RECT 34.050 139.885 34.400 139.890 ;
        RECT 34.065 139.880 34.400 139.885 ;
        RECT 34.765 139.880 35.025 140.330 ;
        RECT 35.655 139.990 35.945 141.155 ;
        RECT 36.115 140.015 36.500 140.985 ;
        RECT 36.670 140.695 36.995 141.155 ;
        RECT 37.515 140.525 37.795 140.985 ;
        RECT 36.670 140.305 37.795 140.525 ;
        RECT 34.065 139.875 35.025 139.880 ;
        RECT 34.075 139.865 35.025 139.875 ;
        RECT 34.085 139.860 35.025 139.865 ;
        RECT 34.095 139.850 35.025 139.860 ;
        RECT 34.100 139.840 35.025 139.850 ;
        RECT 34.105 139.835 35.025 139.840 ;
        RECT 34.115 139.820 35.025 139.835 ;
        RECT 34.120 139.805 35.025 139.820 ;
        RECT 34.130 139.780 35.025 139.805 ;
        RECT 33.635 139.310 33.965 139.735 ;
        RECT 32.895 138.775 33.155 139.255 ;
        RECT 33.325 138.605 33.575 139.145 ;
        RECT 33.745 138.825 33.965 139.310 ;
        RECT 34.135 139.710 35.025 139.780 ;
        RECT 34.135 138.985 34.305 139.710 ;
        RECT 34.475 139.155 35.025 139.540 ;
        RECT 36.115 139.345 36.395 140.015 ;
        RECT 36.670 139.845 37.120 140.305 ;
        RECT 37.985 140.135 38.385 140.985 ;
        RECT 38.785 140.695 39.055 141.155 ;
        RECT 39.225 140.525 39.510 140.985 ;
        RECT 39.795 140.645 40.055 141.155 ;
        RECT 36.565 139.515 37.120 139.845 ;
        RECT 37.290 139.575 38.385 140.135 ;
        RECT 36.670 139.405 37.120 139.515 ;
        RECT 34.135 138.815 35.025 138.985 ;
        RECT 35.655 138.605 35.945 139.330 ;
        RECT 36.115 138.775 36.500 139.345 ;
        RECT 36.670 139.235 37.795 139.405 ;
        RECT 36.670 138.605 36.995 139.065 ;
        RECT 37.515 138.775 37.795 139.235 ;
        RECT 37.985 138.775 38.385 139.575 ;
        RECT 38.555 140.305 39.510 140.525 ;
        RECT 38.555 139.405 38.765 140.305 ;
        RECT 38.935 139.575 39.625 140.135 ;
        RECT 39.795 139.595 40.135 140.475 ;
        RECT 40.305 139.765 40.475 140.985 ;
        RECT 40.715 140.650 41.330 141.155 ;
        RECT 40.715 140.115 40.965 140.480 ;
        RECT 41.135 140.475 41.330 140.650 ;
        RECT 41.500 140.645 41.975 140.985 ;
        RECT 42.145 140.610 42.360 141.155 ;
        RECT 41.135 140.285 41.465 140.475 ;
        RECT 41.685 140.115 42.400 140.410 ;
        RECT 42.570 140.285 42.845 140.985 ;
        RECT 43.105 140.485 43.275 140.985 ;
        RECT 43.445 140.655 43.775 141.155 ;
        RECT 43.105 140.315 43.770 140.485 ;
        RECT 40.715 139.945 42.505 140.115 ;
        RECT 40.305 139.515 41.100 139.765 ;
        RECT 40.305 139.425 40.555 139.515 ;
        RECT 38.555 139.235 39.510 139.405 ;
        RECT 38.785 138.605 39.055 139.065 ;
        RECT 39.225 138.775 39.510 139.235 ;
        RECT 39.795 138.605 40.055 139.425 ;
        RECT 40.225 139.005 40.555 139.425 ;
        RECT 41.270 139.090 41.525 139.945 ;
        RECT 40.735 138.825 41.525 139.090 ;
        RECT 41.695 139.245 42.105 139.765 ;
        RECT 42.275 139.515 42.505 139.945 ;
        RECT 42.675 139.255 42.845 140.285 ;
        RECT 43.020 139.495 43.370 140.145 ;
        RECT 43.540 139.325 43.770 140.315 ;
        RECT 41.695 138.825 41.895 139.245 ;
        RECT 42.085 138.605 42.415 139.065 ;
        RECT 42.585 138.775 42.845 139.255 ;
        RECT 43.105 139.155 43.770 139.325 ;
        RECT 43.105 138.865 43.275 139.155 ;
        RECT 43.445 138.605 43.775 138.985 ;
        RECT 43.945 138.865 44.130 140.985 ;
        RECT 44.370 140.695 44.635 141.155 ;
        RECT 44.805 140.560 45.055 140.985 ;
        RECT 45.265 140.710 46.370 140.880 ;
        RECT 44.750 140.430 45.055 140.560 ;
        RECT 44.300 139.235 44.580 140.185 ;
        RECT 44.750 139.325 44.920 140.430 ;
        RECT 45.090 139.645 45.330 140.240 ;
        RECT 45.500 140.175 46.030 140.540 ;
        RECT 45.500 139.475 45.670 140.175 ;
        RECT 46.200 140.095 46.370 140.710 ;
        RECT 46.540 140.355 46.710 141.155 ;
        RECT 46.880 140.655 47.130 140.985 ;
        RECT 47.355 140.685 48.240 140.855 ;
        RECT 46.200 140.005 46.710 140.095 ;
        RECT 44.750 139.195 44.975 139.325 ;
        RECT 45.145 139.255 45.670 139.475 ;
        RECT 45.840 139.835 46.710 140.005 ;
        RECT 44.385 138.605 44.635 139.065 ;
        RECT 44.805 139.055 44.975 139.195 ;
        RECT 45.840 139.055 46.010 139.835 ;
        RECT 46.540 139.765 46.710 139.835 ;
        RECT 46.220 139.585 46.420 139.615 ;
        RECT 46.880 139.585 47.050 140.655 ;
        RECT 47.220 139.765 47.410 140.485 ;
        RECT 46.220 139.285 47.050 139.585 ;
        RECT 47.580 139.555 47.900 140.515 ;
        RECT 44.805 138.885 45.140 139.055 ;
        RECT 45.335 138.885 46.010 139.055 ;
        RECT 46.330 138.605 46.700 139.105 ;
        RECT 46.880 139.055 47.050 139.285 ;
        RECT 47.435 139.225 47.900 139.555 ;
        RECT 48.070 139.845 48.240 140.685 ;
        RECT 48.420 140.655 48.735 141.155 ;
        RECT 48.965 140.425 49.305 140.985 ;
        RECT 48.410 140.050 49.305 140.425 ;
        RECT 49.475 140.145 49.645 141.155 ;
        RECT 49.115 139.845 49.305 140.050 ;
        RECT 49.815 140.095 50.145 140.940 ;
        RECT 49.815 140.015 50.205 140.095 ;
        RECT 50.380 140.015 50.635 141.155 ;
        RECT 50.830 140.605 52.025 140.935 ;
        RECT 49.990 139.965 50.205 140.015 ;
        RECT 48.070 139.515 48.945 139.845 ;
        RECT 49.115 139.515 49.865 139.845 ;
        RECT 48.070 139.055 48.240 139.515 ;
        RECT 49.115 139.345 49.315 139.515 ;
        RECT 50.035 139.385 50.205 139.965 ;
        RECT 50.885 139.845 51.055 140.405 ;
        RECT 51.280 140.185 51.700 140.435 ;
        RECT 52.205 140.355 52.485 141.155 ;
        RECT 51.280 140.015 52.525 140.185 ;
        RECT 52.695 140.015 52.965 140.985 ;
        RECT 52.355 139.845 52.525 140.015 ;
        RECT 52.735 139.965 52.965 140.015 ;
        RECT 50.380 139.595 50.715 139.845 ;
        RECT 50.885 139.515 51.625 139.845 ;
        RECT 52.355 139.515 52.585 139.845 ;
        RECT 50.885 139.425 51.135 139.515 ;
        RECT 49.980 139.345 50.205 139.385 ;
        RECT 46.880 138.885 47.285 139.055 ;
        RECT 47.455 138.885 48.240 139.055 ;
        RECT 48.515 138.605 48.725 139.135 ;
        RECT 48.985 138.820 49.315 139.345 ;
        RECT 49.825 139.260 50.205 139.345 ;
        RECT 49.485 138.605 49.655 139.215 ;
        RECT 49.825 138.825 50.155 139.260 ;
        RECT 50.400 139.255 51.135 139.425 ;
        RECT 52.355 139.345 52.525 139.515 ;
        RECT 50.400 138.785 50.710 139.255 ;
        RECT 51.785 139.175 52.525 139.345 ;
        RECT 52.795 139.280 52.965 139.965 ;
        RECT 50.880 138.605 51.615 139.085 ;
        RECT 51.785 138.825 51.955 139.175 ;
        RECT 52.125 138.605 52.505 139.005 ;
        RECT 52.695 138.935 52.965 139.280 ;
        RECT 54.055 140.080 54.325 140.985 ;
        RECT 54.495 140.395 54.825 141.155 ;
        RECT 55.005 140.225 55.175 140.985 ;
        RECT 54.055 139.280 54.225 140.080 ;
        RECT 54.510 140.055 55.175 140.225 ;
        RECT 55.435 140.065 58.025 141.155 ;
        RECT 58.665 140.565 58.925 140.955 ;
        RECT 59.095 140.745 59.425 141.155 ;
        RECT 58.665 140.365 59.425 140.565 ;
        RECT 54.510 139.910 54.680 140.055 ;
        RECT 54.395 139.580 54.680 139.910 ;
        RECT 54.510 139.325 54.680 139.580 ;
        RECT 54.915 139.505 55.245 139.875 ;
        RECT 55.435 139.375 56.645 139.895 ;
        RECT 56.815 139.545 58.025 140.065 ;
        RECT 58.675 139.495 58.905 140.185 ;
        RECT 59.085 139.685 59.425 140.365 ;
        RECT 59.615 139.865 59.945 140.975 ;
        RECT 60.115 140.245 60.305 140.975 ;
        RECT 60.475 140.425 60.805 141.155 ;
        RECT 60.985 140.245 61.155 140.975 ;
        RECT 60.115 140.045 61.155 140.245 ;
        RECT 61.415 139.990 61.705 141.155 ;
        RECT 61.965 140.485 62.135 140.985 ;
        RECT 62.305 140.655 62.635 141.155 ;
        RECT 61.965 140.315 62.630 140.485 ;
        RECT 54.055 138.775 54.315 139.280 ;
        RECT 54.510 139.155 55.175 139.325 ;
        RECT 54.495 138.605 54.825 138.985 ;
        RECT 55.005 138.775 55.175 139.155 ;
        RECT 55.435 138.605 58.025 139.375 ;
        RECT 59.085 139.235 59.315 139.685 ;
        RECT 59.615 139.565 60.150 139.865 ;
        RECT 58.935 138.785 59.315 139.235 ;
        RECT 59.495 138.605 59.725 139.385 ;
        RECT 59.905 139.315 60.150 139.565 ;
        RECT 60.330 139.515 60.725 139.865 ;
        RECT 60.920 139.515 61.210 139.865 ;
        RECT 59.905 138.785 60.335 139.315 ;
        RECT 60.515 138.895 60.725 139.515 ;
        RECT 61.880 139.495 62.230 140.145 ;
        RECT 60.895 138.605 61.225 139.335 ;
        RECT 61.415 138.605 61.705 139.330 ;
        RECT 62.400 139.325 62.630 140.315 ;
        RECT 61.965 139.155 62.630 139.325 ;
        RECT 61.965 138.865 62.135 139.155 ;
        RECT 62.305 138.605 62.635 138.985 ;
        RECT 62.805 138.865 62.990 140.985 ;
        RECT 63.230 140.695 63.495 141.155 ;
        RECT 63.665 140.560 63.915 140.985 ;
        RECT 64.125 140.710 65.230 140.880 ;
        RECT 63.610 140.430 63.915 140.560 ;
        RECT 63.160 139.235 63.440 140.185 ;
        RECT 63.610 139.325 63.780 140.430 ;
        RECT 63.950 139.645 64.190 140.240 ;
        RECT 64.360 140.175 64.890 140.540 ;
        RECT 64.360 139.475 64.530 140.175 ;
        RECT 65.060 140.095 65.230 140.710 ;
        RECT 65.400 140.355 65.570 141.155 ;
        RECT 65.740 140.655 65.990 140.985 ;
        RECT 66.215 140.685 67.100 140.855 ;
        RECT 65.060 140.005 65.570 140.095 ;
        RECT 63.610 139.195 63.835 139.325 ;
        RECT 64.005 139.255 64.530 139.475 ;
        RECT 64.700 139.835 65.570 140.005 ;
        RECT 63.245 138.605 63.495 139.065 ;
        RECT 63.665 139.055 63.835 139.195 ;
        RECT 64.700 139.055 64.870 139.835 ;
        RECT 65.400 139.765 65.570 139.835 ;
        RECT 65.080 139.585 65.280 139.615 ;
        RECT 65.740 139.585 65.910 140.655 ;
        RECT 66.080 139.765 66.270 140.485 ;
        RECT 65.080 139.285 65.910 139.585 ;
        RECT 66.440 139.555 66.760 140.515 ;
        RECT 63.665 138.885 64.000 139.055 ;
        RECT 64.195 138.885 64.870 139.055 ;
        RECT 65.190 138.605 65.560 139.105 ;
        RECT 65.740 139.055 65.910 139.285 ;
        RECT 66.295 139.225 66.760 139.555 ;
        RECT 66.930 139.845 67.100 140.685 ;
        RECT 67.280 140.655 67.595 141.155 ;
        RECT 67.825 140.425 68.165 140.985 ;
        RECT 67.270 140.050 68.165 140.425 ;
        RECT 68.335 140.145 68.505 141.155 ;
        RECT 67.975 139.845 68.165 140.050 ;
        RECT 68.675 140.095 69.005 140.940 ;
        RECT 69.235 140.395 69.900 140.985 ;
        RECT 68.675 140.015 69.065 140.095 ;
        RECT 68.850 139.965 69.065 140.015 ;
        RECT 66.930 139.515 67.805 139.845 ;
        RECT 67.975 139.515 68.725 139.845 ;
        RECT 66.930 139.055 67.100 139.515 ;
        RECT 67.975 139.345 68.175 139.515 ;
        RECT 68.895 139.385 69.065 139.965 ;
        RECT 68.840 139.345 69.065 139.385 ;
        RECT 65.740 138.885 66.145 139.055 ;
        RECT 66.315 138.885 67.100 139.055 ;
        RECT 67.375 138.605 67.585 139.135 ;
        RECT 67.845 138.820 68.175 139.345 ;
        RECT 68.685 139.260 69.065 139.345 ;
        RECT 69.235 139.425 69.485 140.395 ;
        RECT 70.070 140.315 70.400 141.155 ;
        RECT 70.910 140.565 71.715 140.985 ;
        RECT 70.570 140.395 72.135 140.565 ;
        RECT 70.570 140.145 70.740 140.395 ;
        RECT 69.820 139.975 70.740 140.145 ;
        RECT 70.910 140.135 71.285 140.225 ;
        RECT 69.820 139.805 69.990 139.975 ;
        RECT 70.910 139.965 71.305 140.135 ;
        RECT 70.910 139.805 71.285 139.965 ;
        RECT 69.655 139.595 69.990 139.805 ;
        RECT 70.160 139.595 70.610 139.805 ;
        RECT 70.800 139.595 71.285 139.805 ;
        RECT 71.475 139.845 71.795 140.225 ;
        RECT 71.965 140.145 72.135 140.395 ;
        RECT 72.305 140.315 72.555 141.155 ;
        RECT 72.750 140.145 73.050 140.985 ;
        RECT 71.965 139.975 73.050 140.145 ;
        RECT 73.435 140.015 73.645 141.155 ;
        RECT 73.815 140.005 74.145 140.985 ;
        RECT 74.315 140.015 74.545 141.155 ;
        RECT 74.815 140.015 75.025 141.155 ;
        RECT 75.195 140.005 75.525 140.985 ;
        RECT 75.695 140.015 75.925 141.155 ;
        RECT 76.250 140.525 76.535 140.985 ;
        RECT 76.705 140.695 76.975 141.155 ;
        RECT 76.250 140.305 77.205 140.525 ;
        RECT 71.475 139.595 71.855 139.845 ;
        RECT 72.035 139.595 72.365 139.805 ;
        RECT 68.345 138.605 68.515 139.215 ;
        RECT 68.685 138.825 69.015 139.260 ;
        RECT 69.235 138.785 69.920 139.425 ;
        RECT 70.090 138.605 70.260 139.425 ;
        RECT 70.430 139.255 72.130 139.425 ;
        RECT 70.430 138.790 70.760 139.255 ;
        RECT 71.745 139.165 72.130 139.255 ;
        RECT 72.535 139.345 72.705 139.975 ;
        RECT 72.875 139.515 73.205 139.805 ;
        RECT 72.535 139.165 73.045 139.345 ;
        RECT 70.930 138.605 71.100 139.075 ;
        RECT 71.360 138.825 72.545 138.995 ;
        RECT 72.715 138.775 73.045 139.165 ;
        RECT 73.435 138.605 73.645 139.425 ;
        RECT 73.815 139.405 74.065 140.005 ;
        RECT 74.235 139.595 74.565 139.845 ;
        RECT 73.815 138.775 74.145 139.405 ;
        RECT 74.315 138.605 74.545 139.425 ;
        RECT 74.815 138.605 75.025 139.425 ;
        RECT 75.195 139.405 75.445 140.005 ;
        RECT 75.615 139.595 75.945 139.845 ;
        RECT 76.135 139.575 76.825 140.135 ;
        RECT 75.195 138.775 75.525 139.405 ;
        RECT 75.695 138.605 75.925 139.425 ;
        RECT 76.995 139.405 77.205 140.305 ;
        RECT 76.250 139.235 77.205 139.405 ;
        RECT 77.375 140.135 77.775 140.985 ;
        RECT 77.965 140.525 78.245 140.985 ;
        RECT 78.765 140.695 79.090 141.155 ;
        RECT 77.965 140.305 79.090 140.525 ;
        RECT 77.375 139.575 78.470 140.135 ;
        RECT 78.640 139.845 79.090 140.305 ;
        RECT 79.260 140.015 79.645 140.985 ;
        RECT 79.875 140.095 80.205 140.940 ;
        RECT 80.375 140.145 80.545 141.155 ;
        RECT 80.715 140.425 81.055 140.985 ;
        RECT 81.285 140.655 81.600 141.155 ;
        RECT 81.780 140.685 82.665 140.855 ;
        RECT 76.250 138.775 76.535 139.235 ;
        RECT 76.705 138.605 76.975 139.065 ;
        RECT 77.375 138.775 77.775 139.575 ;
        RECT 78.640 139.515 79.195 139.845 ;
        RECT 78.640 139.405 79.090 139.515 ;
        RECT 77.965 139.235 79.090 139.405 ;
        RECT 79.365 139.345 79.645 140.015 ;
        RECT 77.965 138.775 78.245 139.235 ;
        RECT 78.765 138.605 79.090 139.065 ;
        RECT 79.260 138.775 79.645 139.345 ;
        RECT 79.815 140.015 80.205 140.095 ;
        RECT 80.715 140.050 81.610 140.425 ;
        RECT 79.815 139.965 80.030 140.015 ;
        RECT 79.815 139.385 79.985 139.965 ;
        RECT 80.715 139.845 80.905 140.050 ;
        RECT 81.780 139.845 81.950 140.685 ;
        RECT 82.890 140.655 83.140 140.985 ;
        RECT 80.155 139.515 80.905 139.845 ;
        RECT 81.075 139.515 81.950 139.845 ;
        RECT 79.815 139.345 80.040 139.385 ;
        RECT 80.705 139.345 80.905 139.515 ;
        RECT 79.815 139.260 80.195 139.345 ;
        RECT 79.865 138.825 80.195 139.260 ;
        RECT 80.365 138.605 80.535 139.215 ;
        RECT 80.705 138.820 81.035 139.345 ;
        RECT 81.295 138.605 81.505 139.135 ;
        RECT 81.780 139.055 81.950 139.515 ;
        RECT 82.120 139.555 82.440 140.515 ;
        RECT 82.610 139.765 82.800 140.485 ;
        RECT 82.970 139.585 83.140 140.655 ;
        RECT 83.310 140.355 83.480 141.155 ;
        RECT 83.650 140.710 84.755 140.880 ;
        RECT 83.650 140.095 83.820 140.710 ;
        RECT 84.965 140.560 85.215 140.985 ;
        RECT 85.385 140.695 85.650 141.155 ;
        RECT 83.990 140.175 84.520 140.540 ;
        RECT 84.965 140.430 85.270 140.560 ;
        RECT 83.310 140.005 83.820 140.095 ;
        RECT 83.310 139.835 84.180 140.005 ;
        RECT 83.310 139.765 83.480 139.835 ;
        RECT 83.600 139.585 83.800 139.615 ;
        RECT 82.120 139.225 82.585 139.555 ;
        RECT 82.970 139.285 83.800 139.585 ;
        RECT 82.970 139.055 83.140 139.285 ;
        RECT 81.780 138.885 82.565 139.055 ;
        RECT 82.735 138.885 83.140 139.055 ;
        RECT 83.320 138.605 83.690 139.105 ;
        RECT 84.010 139.055 84.180 139.835 ;
        RECT 84.350 139.475 84.520 140.175 ;
        RECT 84.690 139.645 84.930 140.240 ;
        RECT 84.350 139.255 84.875 139.475 ;
        RECT 85.100 139.325 85.270 140.430 ;
        RECT 85.045 139.195 85.270 139.325 ;
        RECT 85.440 139.235 85.720 140.185 ;
        RECT 85.045 139.055 85.215 139.195 ;
        RECT 84.010 138.885 84.685 139.055 ;
        RECT 84.880 138.885 85.215 139.055 ;
        RECT 85.385 138.605 85.635 139.065 ;
        RECT 85.890 138.865 86.075 140.985 ;
        RECT 86.245 140.655 86.575 141.155 ;
        RECT 86.745 140.485 86.915 140.985 ;
        RECT 86.250 140.315 86.915 140.485 ;
        RECT 86.250 139.325 86.480 140.315 ;
        RECT 86.650 139.495 87.000 140.145 ;
        RECT 87.175 139.990 87.465 141.155 ;
        RECT 87.740 140.695 87.910 141.155 ;
        RECT 88.080 140.525 88.410 140.985 ;
        RECT 87.635 140.355 88.410 140.525 ;
        RECT 88.580 140.355 88.750 141.155 ;
        RECT 87.635 139.345 88.065 140.355 ;
        RECT 89.335 140.185 89.695 140.360 ;
        RECT 88.235 140.015 89.695 140.185 ;
        RECT 89.935 140.080 90.205 140.985 ;
        RECT 90.375 140.395 90.705 141.155 ;
        RECT 90.885 140.225 91.055 140.985 ;
        RECT 91.865 140.410 92.135 141.155 ;
        RECT 92.765 141.150 99.040 141.155 ;
        RECT 92.305 140.240 92.595 140.980 ;
        RECT 92.765 140.425 93.020 141.150 ;
        RECT 93.205 140.255 93.465 140.980 ;
        RECT 93.635 140.425 93.880 141.150 ;
        RECT 94.065 140.255 94.325 140.980 ;
        RECT 94.495 140.425 94.740 141.150 ;
        RECT 94.925 140.255 95.185 140.980 ;
        RECT 95.355 140.425 95.600 141.150 ;
        RECT 95.770 140.255 96.030 140.980 ;
        RECT 96.200 140.425 96.460 141.150 ;
        RECT 96.630 140.255 96.890 140.980 ;
        RECT 97.060 140.425 97.320 141.150 ;
        RECT 97.490 140.255 97.750 140.980 ;
        RECT 97.920 140.425 98.180 141.150 ;
        RECT 98.350 140.255 98.610 140.980 ;
        RECT 98.780 140.355 99.040 141.150 ;
        RECT 93.205 140.240 98.610 140.255 ;
        RECT 88.235 139.515 88.405 140.015 ;
        RECT 86.250 139.155 86.915 139.325 ;
        RECT 86.245 138.605 86.575 138.985 ;
        RECT 86.745 138.865 86.915 139.155 ;
        RECT 87.175 138.605 87.465 139.330 ;
        RECT 87.635 139.175 88.330 139.345 ;
        RECT 88.575 139.285 88.985 139.845 ;
        RECT 87.660 138.605 87.990 139.005 ;
        RECT 88.160 138.905 88.330 139.175 ;
        RECT 89.155 139.115 89.335 140.015 ;
        RECT 89.505 139.455 89.700 139.845 ;
        RECT 89.505 139.285 89.705 139.455 ;
        RECT 89.935 139.280 90.105 140.080 ;
        RECT 90.390 140.055 91.055 140.225 ;
        RECT 90.390 139.910 90.560 140.055 ;
        RECT 90.275 139.580 90.560 139.910 ;
        RECT 91.865 140.015 98.610 140.240 ;
        RECT 90.390 139.325 90.560 139.580 ;
        RECT 90.795 139.505 91.125 139.875 ;
        RECT 91.865 139.425 93.030 140.015 ;
        RECT 99.210 139.845 99.460 140.980 ;
        RECT 99.640 140.345 99.900 141.155 ;
        RECT 100.075 139.845 100.320 140.985 ;
        RECT 100.500 140.345 100.795 141.155 ;
        RECT 101.015 140.815 102.155 140.985 ;
        RECT 101.015 140.355 101.315 140.815 ;
        RECT 101.485 140.185 101.815 140.645 ;
        RECT 101.055 139.965 101.815 140.185 ;
        RECT 101.985 140.185 102.155 140.815 ;
        RECT 102.325 140.355 102.655 141.155 ;
        RECT 102.825 140.185 103.100 140.985 ;
        RECT 101.985 139.975 103.100 140.185 ;
        RECT 103.280 140.185 103.555 140.985 ;
        RECT 103.725 140.355 104.055 141.155 ;
        RECT 104.225 140.815 105.365 140.985 ;
        RECT 104.225 140.185 104.395 140.815 ;
        RECT 103.280 139.975 104.395 140.185 ;
        RECT 104.565 140.185 104.895 140.645 ;
        RECT 105.065 140.355 105.365 140.815 ;
        RECT 105.665 140.225 105.835 140.985 ;
        RECT 106.050 140.395 106.380 141.155 ;
        RECT 104.565 139.965 105.325 140.185 ;
        RECT 105.665 140.055 106.380 140.225 ;
        RECT 106.550 140.080 106.805 140.985 ;
        RECT 93.200 139.595 100.320 139.845 ;
        RECT 88.500 138.605 88.815 139.115 ;
        RECT 89.045 138.775 89.335 139.115 ;
        RECT 89.505 138.605 89.745 139.115 ;
        RECT 89.935 138.775 90.195 139.280 ;
        RECT 90.390 139.155 91.055 139.325 ;
        RECT 91.865 139.255 98.610 139.425 ;
        RECT 90.375 138.605 90.705 138.985 ;
        RECT 90.885 138.775 91.055 139.155 ;
        RECT 91.865 138.605 92.165 139.085 ;
        RECT 92.335 138.800 92.595 139.255 ;
        RECT 92.765 138.605 93.025 139.085 ;
        RECT 93.205 138.800 93.465 139.255 ;
        RECT 93.635 138.605 93.885 139.085 ;
        RECT 94.065 138.800 94.325 139.255 ;
        RECT 94.495 138.605 94.745 139.085 ;
        RECT 94.925 138.800 95.185 139.255 ;
        RECT 95.355 138.605 95.600 139.085 ;
        RECT 95.770 138.800 96.045 139.255 ;
        RECT 96.215 138.605 96.460 139.085 ;
        RECT 96.630 138.800 96.890 139.255 ;
        RECT 97.060 138.605 97.320 139.085 ;
        RECT 97.490 138.800 97.750 139.255 ;
        RECT 97.920 138.605 98.180 139.085 ;
        RECT 98.350 138.800 98.610 139.255 ;
        RECT 98.780 138.605 99.040 139.165 ;
        RECT 99.210 138.785 99.460 139.595 ;
        RECT 99.640 138.605 99.900 139.130 ;
        RECT 100.070 138.785 100.320 139.595 ;
        RECT 100.490 139.285 100.805 139.845 ;
        RECT 101.055 139.425 101.270 139.965 ;
        RECT 101.440 139.595 102.210 139.795 ;
        RECT 102.380 139.595 103.100 139.795 ;
        RECT 103.280 139.595 104.000 139.795 ;
        RECT 104.170 139.595 104.940 139.795 ;
        RECT 105.110 139.425 105.325 139.965 ;
        RECT 105.575 139.505 105.930 139.875 ;
        RECT 106.210 139.845 106.380 140.055 ;
        RECT 106.210 139.515 106.465 139.845 ;
        RECT 101.055 139.255 102.655 139.425 ;
        RECT 101.485 139.245 102.655 139.255 ;
        RECT 100.500 138.605 100.805 139.115 ;
        RECT 101.025 138.605 101.315 139.075 ;
        RECT 101.485 138.775 101.815 139.245 ;
        RECT 101.985 138.605 102.155 139.075 ;
        RECT 102.325 138.775 102.655 139.245 ;
        RECT 102.825 138.605 103.100 139.425 ;
        RECT 103.280 138.605 103.555 139.425 ;
        RECT 103.725 139.255 105.325 139.425 ;
        RECT 106.210 139.325 106.380 139.515 ;
        RECT 106.635 139.350 106.805 140.080 ;
        RECT 106.980 140.005 107.240 141.155 ;
        RECT 107.420 140.015 107.755 140.985 ;
        RECT 107.925 140.015 108.095 141.155 ;
        RECT 108.265 140.815 110.295 140.985 ;
        RECT 103.725 139.245 104.895 139.255 ;
        RECT 103.725 138.775 104.055 139.245 ;
        RECT 104.225 138.605 104.395 139.075 ;
        RECT 104.565 138.775 104.895 139.245 ;
        RECT 105.665 139.155 106.380 139.325 ;
        RECT 105.065 138.605 105.355 139.075 ;
        RECT 105.665 138.775 105.835 139.155 ;
        RECT 106.050 138.605 106.380 138.985 ;
        RECT 106.550 138.775 106.805 139.350 ;
        RECT 106.980 138.605 107.240 139.445 ;
        RECT 107.420 139.345 107.590 140.015 ;
        RECT 108.265 139.845 108.435 140.815 ;
        RECT 107.760 139.515 108.015 139.845 ;
        RECT 108.240 139.515 108.435 139.845 ;
        RECT 108.605 140.475 109.730 140.645 ;
        RECT 107.845 139.345 108.015 139.515 ;
        RECT 108.605 139.345 108.775 140.475 ;
        RECT 107.420 138.775 107.675 139.345 ;
        RECT 107.845 139.175 108.775 139.345 ;
        RECT 108.945 140.135 109.955 140.305 ;
        RECT 108.945 139.335 109.115 140.135 ;
        RECT 108.600 139.140 108.775 139.175 ;
        RECT 107.845 138.605 108.175 139.005 ;
        RECT 108.600 138.775 109.130 139.140 ;
        RECT 109.320 139.115 109.595 139.935 ;
        RECT 109.315 138.945 109.595 139.115 ;
        RECT 109.320 138.775 109.595 138.945 ;
        RECT 109.765 138.775 109.955 140.135 ;
        RECT 110.125 140.150 110.295 140.815 ;
        RECT 110.465 140.395 110.635 141.155 ;
        RECT 110.870 140.395 111.385 140.805 ;
        RECT 110.125 139.960 110.875 140.150 ;
        RECT 111.045 139.585 111.385 140.395 ;
        RECT 111.555 140.065 112.765 141.155 ;
        RECT 110.155 139.415 111.385 139.585 ;
        RECT 110.135 138.605 110.645 139.140 ;
        RECT 110.865 138.810 111.110 139.415 ;
        RECT 111.555 139.355 112.075 139.895 ;
        RECT 112.245 139.525 112.765 140.065 ;
        RECT 112.935 139.990 113.225 141.155 ;
        RECT 114.405 140.485 114.575 140.985 ;
        RECT 114.745 140.655 115.075 141.155 ;
        RECT 114.405 140.315 115.070 140.485 ;
        RECT 114.320 139.495 114.670 140.145 ;
        RECT 111.555 138.605 112.765 139.355 ;
        RECT 112.935 138.605 113.225 139.330 ;
        RECT 114.840 139.325 115.070 140.315 ;
        RECT 114.405 139.155 115.070 139.325 ;
        RECT 114.405 138.865 114.575 139.155 ;
        RECT 114.745 138.605 115.075 138.985 ;
        RECT 115.245 138.865 115.430 140.985 ;
        RECT 115.670 140.695 115.935 141.155 ;
        RECT 116.105 140.560 116.355 140.985 ;
        RECT 116.565 140.710 117.670 140.880 ;
        RECT 116.050 140.430 116.355 140.560 ;
        RECT 115.600 139.235 115.880 140.185 ;
        RECT 116.050 139.325 116.220 140.430 ;
        RECT 116.390 139.645 116.630 140.240 ;
        RECT 116.800 140.175 117.330 140.540 ;
        RECT 116.800 139.475 116.970 140.175 ;
        RECT 117.500 140.095 117.670 140.710 ;
        RECT 117.840 140.355 118.010 141.155 ;
        RECT 118.180 140.655 118.430 140.985 ;
        RECT 118.655 140.685 119.540 140.855 ;
        RECT 117.500 140.005 118.010 140.095 ;
        RECT 116.050 139.195 116.275 139.325 ;
        RECT 116.445 139.255 116.970 139.475 ;
        RECT 117.140 139.835 118.010 140.005 ;
        RECT 115.685 138.605 115.935 139.065 ;
        RECT 116.105 139.055 116.275 139.195 ;
        RECT 117.140 139.055 117.310 139.835 ;
        RECT 117.840 139.765 118.010 139.835 ;
        RECT 117.520 139.585 117.720 139.615 ;
        RECT 118.180 139.585 118.350 140.655 ;
        RECT 118.520 139.765 118.710 140.485 ;
        RECT 117.520 139.285 118.350 139.585 ;
        RECT 118.880 139.555 119.200 140.515 ;
        RECT 116.105 138.885 116.440 139.055 ;
        RECT 116.635 138.885 117.310 139.055 ;
        RECT 117.630 138.605 118.000 139.105 ;
        RECT 118.180 139.055 118.350 139.285 ;
        RECT 118.735 139.225 119.200 139.555 ;
        RECT 119.370 139.845 119.540 140.685 ;
        RECT 119.720 140.655 120.035 141.155 ;
        RECT 120.265 140.425 120.605 140.985 ;
        RECT 119.710 140.050 120.605 140.425 ;
        RECT 120.775 140.145 120.945 141.155 ;
        RECT 120.415 139.845 120.605 140.050 ;
        RECT 121.115 140.095 121.445 140.940 ;
        RECT 122.225 140.485 122.395 140.985 ;
        RECT 122.565 140.655 122.895 141.155 ;
        RECT 122.225 140.315 122.890 140.485 ;
        RECT 121.115 140.015 121.505 140.095 ;
        RECT 121.290 139.965 121.505 140.015 ;
        RECT 119.370 139.515 120.245 139.845 ;
        RECT 120.415 139.515 121.165 139.845 ;
        RECT 119.370 139.055 119.540 139.515 ;
        RECT 120.415 139.345 120.615 139.515 ;
        RECT 121.335 139.385 121.505 139.965 ;
        RECT 122.140 139.495 122.490 140.145 ;
        RECT 121.280 139.345 121.505 139.385 ;
        RECT 118.180 138.885 118.585 139.055 ;
        RECT 118.755 138.885 119.540 139.055 ;
        RECT 119.815 138.605 120.025 139.135 ;
        RECT 120.285 138.820 120.615 139.345 ;
        RECT 121.125 139.260 121.505 139.345 ;
        RECT 122.660 139.325 122.890 140.315 ;
        RECT 120.785 138.605 120.955 139.215 ;
        RECT 121.125 138.825 121.455 139.260 ;
        RECT 122.225 139.155 122.890 139.325 ;
        RECT 122.225 138.865 122.395 139.155 ;
        RECT 122.565 138.605 122.895 138.985 ;
        RECT 123.065 138.865 123.250 140.985 ;
        RECT 123.490 140.695 123.755 141.155 ;
        RECT 123.925 140.560 124.175 140.985 ;
        RECT 124.385 140.710 125.490 140.880 ;
        RECT 123.870 140.430 124.175 140.560 ;
        RECT 123.420 139.235 123.700 140.185 ;
        RECT 123.870 139.325 124.040 140.430 ;
        RECT 124.210 139.645 124.450 140.240 ;
        RECT 124.620 140.175 125.150 140.540 ;
        RECT 124.620 139.475 124.790 140.175 ;
        RECT 125.320 140.095 125.490 140.710 ;
        RECT 125.660 140.355 125.830 141.155 ;
        RECT 126.000 140.655 126.250 140.985 ;
        RECT 126.475 140.685 127.360 140.855 ;
        RECT 125.320 140.005 125.830 140.095 ;
        RECT 123.870 139.195 124.095 139.325 ;
        RECT 124.265 139.255 124.790 139.475 ;
        RECT 124.960 139.835 125.830 140.005 ;
        RECT 123.505 138.605 123.755 139.065 ;
        RECT 123.925 139.055 124.095 139.195 ;
        RECT 124.960 139.055 125.130 139.835 ;
        RECT 125.660 139.765 125.830 139.835 ;
        RECT 125.340 139.585 125.540 139.615 ;
        RECT 126.000 139.585 126.170 140.655 ;
        RECT 126.340 139.765 126.530 140.485 ;
        RECT 125.340 139.285 126.170 139.585 ;
        RECT 126.700 139.555 127.020 140.515 ;
        RECT 123.925 138.885 124.260 139.055 ;
        RECT 124.455 138.885 125.130 139.055 ;
        RECT 125.450 138.605 125.820 139.105 ;
        RECT 126.000 139.055 126.170 139.285 ;
        RECT 126.555 139.225 127.020 139.555 ;
        RECT 127.190 139.845 127.360 140.685 ;
        RECT 127.540 140.655 127.855 141.155 ;
        RECT 128.085 140.425 128.425 140.985 ;
        RECT 127.530 140.050 128.425 140.425 ;
        RECT 128.595 140.145 128.765 141.155 ;
        RECT 128.235 139.845 128.425 140.050 ;
        RECT 128.935 140.095 129.265 140.940 ;
        RECT 128.935 140.015 129.325 140.095 ;
        RECT 129.495 140.065 131.165 141.155 ;
        RECT 129.110 139.965 129.325 140.015 ;
        RECT 127.190 139.515 128.065 139.845 ;
        RECT 128.235 139.515 128.985 139.845 ;
        RECT 127.190 139.055 127.360 139.515 ;
        RECT 128.235 139.345 128.435 139.515 ;
        RECT 129.155 139.385 129.325 139.965 ;
        RECT 129.100 139.345 129.325 139.385 ;
        RECT 126.000 138.885 126.405 139.055 ;
        RECT 126.575 138.885 127.360 139.055 ;
        RECT 127.635 138.605 127.845 139.135 ;
        RECT 128.105 138.820 128.435 139.345 ;
        RECT 128.945 139.260 129.325 139.345 ;
        RECT 129.495 139.375 130.245 139.895 ;
        RECT 130.415 139.545 131.165 140.065 ;
        RECT 131.815 140.315 132.070 140.985 ;
        RECT 132.240 140.395 132.570 141.155 ;
        RECT 132.740 140.555 132.990 140.985 ;
        RECT 133.160 140.735 133.515 141.155 ;
        RECT 133.705 140.815 134.875 140.985 ;
        RECT 133.705 140.775 134.035 140.815 ;
        RECT 134.145 140.555 134.375 140.645 ;
        RECT 132.740 140.315 134.375 140.555 ;
        RECT 134.545 140.315 134.875 140.815 ;
        RECT 128.605 138.605 128.775 139.215 ;
        RECT 128.945 138.825 129.275 139.260 ;
        RECT 129.495 138.605 131.165 139.375 ;
        RECT 131.815 139.185 131.985 140.315 ;
        RECT 135.045 140.145 135.215 140.985 ;
        RECT 132.155 139.975 135.215 140.145 ;
        RECT 135.475 140.435 135.935 140.985 ;
        RECT 136.125 140.435 136.455 141.155 ;
        RECT 132.155 139.425 132.325 139.975 ;
        RECT 132.545 139.625 132.920 139.795 ;
        RECT 132.555 139.595 132.920 139.625 ;
        RECT 133.090 139.595 133.420 139.795 ;
        RECT 132.155 139.255 132.955 139.425 ;
        RECT 131.815 139.115 132.000 139.185 ;
        RECT 131.815 139.105 132.025 139.115 ;
        RECT 131.815 138.775 132.070 139.105 ;
        RECT 132.285 138.605 132.615 139.085 ;
        RECT 132.785 139.025 132.955 139.255 ;
        RECT 133.135 139.195 133.420 139.595 ;
        RECT 133.690 139.595 134.165 139.795 ;
        RECT 134.335 139.595 134.780 139.795 ;
        RECT 134.950 139.595 135.300 139.805 ;
        RECT 133.690 139.195 133.970 139.595 ;
        RECT 134.150 139.255 135.215 139.425 ;
        RECT 134.150 139.025 134.320 139.255 ;
        RECT 132.785 138.775 134.320 139.025 ;
        RECT 134.545 138.605 134.875 139.085 ;
        RECT 135.045 138.775 135.215 139.255 ;
        RECT 135.475 139.065 135.725 140.435 ;
        RECT 136.655 140.265 136.955 140.815 ;
        RECT 137.125 140.485 137.405 141.155 ;
        RECT 136.015 140.095 136.955 140.265 ;
        RECT 136.015 139.845 136.185 140.095 ;
        RECT 137.325 139.845 137.590 140.205 ;
        RECT 138.695 139.990 138.985 141.155 ;
        RECT 139.215 140.015 139.425 141.155 ;
        RECT 139.595 140.005 139.925 140.985 ;
        RECT 140.095 140.015 140.325 141.155 ;
        RECT 140.535 140.725 140.875 140.985 ;
        RECT 135.895 139.515 136.185 139.845 ;
        RECT 136.355 139.595 136.695 139.845 ;
        RECT 136.915 139.595 137.590 139.845 ;
        RECT 136.015 139.425 136.185 139.515 ;
        RECT 136.015 139.235 137.405 139.425 ;
        RECT 135.475 138.775 136.035 139.065 ;
        RECT 136.205 138.605 136.455 139.065 ;
        RECT 137.075 138.875 137.405 139.235 ;
        RECT 138.695 138.605 138.985 139.330 ;
        RECT 139.215 138.605 139.425 139.425 ;
        RECT 139.595 139.405 139.845 140.005 ;
        RECT 140.015 139.595 140.345 139.845 ;
        RECT 139.595 138.775 139.925 139.405 ;
        RECT 140.095 138.605 140.325 139.425 ;
        RECT 140.535 139.325 140.795 140.725 ;
        RECT 141.045 140.355 141.375 141.155 ;
        RECT 141.840 140.185 142.090 140.985 ;
        RECT 142.275 140.435 142.605 141.155 ;
        RECT 142.825 140.185 143.075 140.985 ;
        RECT 143.245 140.775 143.580 141.155 ;
        RECT 140.985 140.015 143.175 140.185 ;
        RECT 140.985 139.845 141.300 140.015 ;
        RECT 140.970 139.595 141.300 139.845 ;
        RECT 140.535 138.815 140.875 139.325 ;
        RECT 141.045 138.605 141.315 139.405 ;
        RECT 141.495 138.875 141.775 139.845 ;
        RECT 141.955 138.875 142.255 139.845 ;
        RECT 142.435 138.880 142.785 139.845 ;
        RECT 143.005 139.105 143.175 140.015 ;
        RECT 143.345 139.285 143.585 140.595 ;
        RECT 143.940 140.185 144.330 140.360 ;
        RECT 144.815 140.355 145.145 141.155 ;
        RECT 145.315 140.365 145.850 140.985 ;
        RECT 143.940 140.015 145.365 140.185 ;
        RECT 143.815 139.285 144.170 139.845 ;
        RECT 144.340 139.115 144.510 140.015 ;
        RECT 144.680 139.285 144.945 139.845 ;
        RECT 145.195 139.515 145.365 140.015 ;
        RECT 145.535 139.345 145.850 140.365 ;
        RECT 146.055 140.015 146.315 141.155 ;
        RECT 146.485 140.005 146.815 140.985 ;
        RECT 146.985 140.015 147.265 141.155 ;
        RECT 147.525 140.485 147.695 140.985 ;
        RECT 147.865 140.655 148.195 141.155 ;
        RECT 147.525 140.315 148.190 140.485 ;
        RECT 146.075 139.595 146.410 139.845 ;
        RECT 146.580 139.405 146.750 140.005 ;
        RECT 146.920 139.575 147.255 139.845 ;
        RECT 147.440 139.495 147.790 140.145 ;
        RECT 143.005 138.775 143.500 139.105 ;
        RECT 143.920 138.605 144.160 139.115 ;
        RECT 144.340 138.785 144.620 139.115 ;
        RECT 144.850 138.605 145.065 139.115 ;
        RECT 145.235 138.775 145.850 139.345 ;
        RECT 146.055 138.775 146.750 139.405 ;
        RECT 146.955 138.605 147.265 139.405 ;
        RECT 147.960 139.325 148.190 140.315 ;
        RECT 147.525 139.155 148.190 139.325 ;
        RECT 147.525 138.865 147.695 139.155 ;
        RECT 147.865 138.605 148.195 138.985 ;
        RECT 148.365 138.865 148.550 140.985 ;
        RECT 148.790 140.695 149.055 141.155 ;
        RECT 149.225 140.560 149.475 140.985 ;
        RECT 149.685 140.710 150.790 140.880 ;
        RECT 149.170 140.430 149.475 140.560 ;
        RECT 148.720 139.235 149.000 140.185 ;
        RECT 149.170 139.325 149.340 140.430 ;
        RECT 149.510 139.645 149.750 140.240 ;
        RECT 149.920 140.175 150.450 140.540 ;
        RECT 149.920 139.475 150.090 140.175 ;
        RECT 150.620 140.095 150.790 140.710 ;
        RECT 150.960 140.355 151.130 141.155 ;
        RECT 151.300 140.655 151.550 140.985 ;
        RECT 151.775 140.685 152.660 140.855 ;
        RECT 150.620 140.005 151.130 140.095 ;
        RECT 149.170 139.195 149.395 139.325 ;
        RECT 149.565 139.255 150.090 139.475 ;
        RECT 150.260 139.835 151.130 140.005 ;
        RECT 148.805 138.605 149.055 139.065 ;
        RECT 149.225 139.055 149.395 139.195 ;
        RECT 150.260 139.055 150.430 139.835 ;
        RECT 150.960 139.765 151.130 139.835 ;
        RECT 150.640 139.585 150.840 139.615 ;
        RECT 151.300 139.585 151.470 140.655 ;
        RECT 151.640 139.765 151.830 140.485 ;
        RECT 150.640 139.285 151.470 139.585 ;
        RECT 152.000 139.555 152.320 140.515 ;
        RECT 149.225 138.885 149.560 139.055 ;
        RECT 149.755 138.885 150.430 139.055 ;
        RECT 150.750 138.605 151.120 139.105 ;
        RECT 151.300 139.055 151.470 139.285 ;
        RECT 151.855 139.225 152.320 139.555 ;
        RECT 152.490 139.845 152.660 140.685 ;
        RECT 152.840 140.655 153.155 141.155 ;
        RECT 153.385 140.425 153.725 140.985 ;
        RECT 152.830 140.050 153.725 140.425 ;
        RECT 153.895 140.145 154.065 141.155 ;
        RECT 153.535 139.845 153.725 140.050 ;
        RECT 154.235 140.095 154.565 140.940 ;
        RECT 154.235 140.015 154.625 140.095 ;
        RECT 154.410 139.965 154.625 140.015 ;
        RECT 152.490 139.515 153.365 139.845 ;
        RECT 153.535 139.515 154.285 139.845 ;
        RECT 152.490 139.055 152.660 139.515 ;
        RECT 153.535 139.345 153.735 139.515 ;
        RECT 154.455 139.385 154.625 139.965 ;
        RECT 155.715 140.065 156.925 141.155 ;
        RECT 155.715 139.525 156.235 140.065 ;
        RECT 154.400 139.345 154.625 139.385 ;
        RECT 156.405 139.355 156.925 139.895 ;
        RECT 151.300 138.885 151.705 139.055 ;
        RECT 151.875 138.885 152.660 139.055 ;
        RECT 152.935 138.605 153.145 139.135 ;
        RECT 153.405 138.820 153.735 139.345 ;
        RECT 154.245 139.260 154.625 139.345 ;
        RECT 153.905 138.605 154.075 139.215 ;
        RECT 154.245 138.825 154.575 139.260 ;
        RECT 155.715 138.605 156.925 139.355 ;
        RECT 22.690 138.435 157.010 138.605 ;
        RECT 22.775 137.685 23.985 138.435 ;
        RECT 25.165 137.885 25.335 138.175 ;
        RECT 25.505 138.055 25.835 138.435 ;
        RECT 25.165 137.715 25.830 137.885 ;
        RECT 22.775 137.145 23.295 137.685 ;
        RECT 23.465 136.975 23.985 137.515 ;
        RECT 22.775 135.885 23.985 136.975 ;
        RECT 25.080 136.895 25.430 137.545 ;
        RECT 25.600 136.725 25.830 137.715 ;
        RECT 25.165 136.555 25.830 136.725 ;
        RECT 25.165 136.055 25.335 136.555 ;
        RECT 25.505 135.885 25.835 136.385 ;
        RECT 26.005 136.055 26.190 138.175 ;
        RECT 26.445 137.975 26.695 138.435 ;
        RECT 26.865 137.985 27.200 138.155 ;
        RECT 27.395 137.985 28.070 138.155 ;
        RECT 26.865 137.845 27.035 137.985 ;
        RECT 26.360 136.855 26.640 137.805 ;
        RECT 26.810 137.715 27.035 137.845 ;
        RECT 26.810 136.610 26.980 137.715 ;
        RECT 27.205 137.565 27.730 137.785 ;
        RECT 27.150 136.800 27.390 137.395 ;
        RECT 27.560 136.865 27.730 137.565 ;
        RECT 27.900 137.205 28.070 137.985 ;
        RECT 28.390 137.935 28.760 138.435 ;
        RECT 28.940 137.985 29.345 138.155 ;
        RECT 29.515 137.985 30.300 138.155 ;
        RECT 28.940 137.755 29.110 137.985 ;
        RECT 28.280 137.455 29.110 137.755 ;
        RECT 29.495 137.485 29.960 137.815 ;
        RECT 28.280 137.425 28.480 137.455 ;
        RECT 28.600 137.205 28.770 137.275 ;
        RECT 27.900 137.035 28.770 137.205 ;
        RECT 28.260 136.945 28.770 137.035 ;
        RECT 26.810 136.480 27.115 136.610 ;
        RECT 27.560 136.500 28.090 136.865 ;
        RECT 26.430 135.885 26.695 136.345 ;
        RECT 26.865 136.055 27.115 136.480 ;
        RECT 28.260 136.330 28.430 136.945 ;
        RECT 27.325 136.160 28.430 136.330 ;
        RECT 28.600 135.885 28.770 136.685 ;
        RECT 28.940 136.385 29.110 137.455 ;
        RECT 29.280 136.555 29.470 137.275 ;
        RECT 29.640 136.525 29.960 137.485 ;
        RECT 30.130 137.525 30.300 137.985 ;
        RECT 30.575 137.905 30.785 138.435 ;
        RECT 31.045 137.695 31.375 138.220 ;
        RECT 31.545 137.825 31.715 138.435 ;
        RECT 31.885 137.780 32.215 138.215 ;
        RECT 31.885 137.695 32.265 137.780 ;
        RECT 31.175 137.525 31.375 137.695 ;
        RECT 32.040 137.655 32.265 137.695 ;
        RECT 30.130 137.195 31.005 137.525 ;
        RECT 31.175 137.195 31.925 137.525 ;
        RECT 28.940 136.055 29.190 136.385 ;
        RECT 30.130 136.355 30.300 137.195 ;
        RECT 31.175 136.990 31.365 137.195 ;
        RECT 32.095 137.075 32.265 137.655 ;
        RECT 32.050 137.025 32.265 137.075 ;
        RECT 30.470 136.615 31.365 136.990 ;
        RECT 31.875 136.945 32.265 137.025 ;
        RECT 32.435 137.490 32.775 138.265 ;
        RECT 32.945 137.975 33.115 138.435 ;
        RECT 33.355 138.000 33.715 138.265 ;
        RECT 33.355 137.995 33.710 138.000 ;
        RECT 33.355 137.985 33.705 137.995 ;
        RECT 33.355 137.980 33.700 137.985 ;
        RECT 33.355 137.970 33.695 137.980 ;
        RECT 34.345 137.975 34.515 138.435 ;
        RECT 33.355 137.965 33.690 137.970 ;
        RECT 33.355 137.955 33.680 137.965 ;
        RECT 33.355 137.945 33.670 137.955 ;
        RECT 33.355 137.805 33.655 137.945 ;
        RECT 32.945 137.615 33.655 137.805 ;
        RECT 33.845 137.805 34.175 137.885 ;
        RECT 34.685 137.805 35.025 138.265 ;
        RECT 33.845 137.615 35.025 137.805 ;
        RECT 36.165 137.780 36.495 138.215 ;
        RECT 36.665 137.825 36.835 138.435 ;
        RECT 36.115 137.695 36.495 137.780 ;
        RECT 37.005 137.695 37.335 138.220 ;
        RECT 37.595 137.905 37.805 138.435 ;
        RECT 38.080 137.985 38.865 138.155 ;
        RECT 39.035 137.985 39.440 138.155 ;
        RECT 36.115 137.655 36.340 137.695 ;
        RECT 29.415 136.185 30.300 136.355 ;
        RECT 30.480 135.885 30.795 136.385 ;
        RECT 31.025 136.055 31.365 136.615 ;
        RECT 31.535 135.885 31.705 136.895 ;
        RECT 31.875 136.100 32.205 136.945 ;
        RECT 32.435 136.055 32.715 137.490 ;
        RECT 32.945 137.045 33.230 137.615 ;
        RECT 33.415 137.215 33.885 137.445 ;
        RECT 34.055 137.425 34.385 137.445 ;
        RECT 34.055 137.245 34.505 137.425 ;
        RECT 34.695 137.245 35.025 137.445 ;
        RECT 32.945 136.830 34.095 137.045 ;
        RECT 32.885 135.885 33.595 136.660 ;
        RECT 33.765 136.055 34.095 136.830 ;
        RECT 34.290 136.130 34.505 137.245 ;
        RECT 34.795 136.905 35.025 137.245 ;
        RECT 36.115 137.075 36.285 137.655 ;
        RECT 37.005 137.525 37.205 137.695 ;
        RECT 38.080 137.525 38.250 137.985 ;
        RECT 36.455 137.195 37.205 137.525 ;
        RECT 37.375 137.195 38.250 137.525 ;
        RECT 36.115 137.025 36.330 137.075 ;
        RECT 36.115 136.945 36.505 137.025 ;
        RECT 34.685 135.885 35.015 136.605 ;
        RECT 36.175 136.100 36.505 136.945 ;
        RECT 37.015 136.990 37.205 137.195 ;
        RECT 36.675 135.885 36.845 136.895 ;
        RECT 37.015 136.615 37.910 136.990 ;
        RECT 37.015 136.055 37.355 136.615 ;
        RECT 37.585 135.885 37.900 136.385 ;
        RECT 38.080 136.355 38.250 137.195 ;
        RECT 38.420 137.485 38.885 137.815 ;
        RECT 39.270 137.755 39.440 137.985 ;
        RECT 39.620 137.935 39.990 138.435 ;
        RECT 40.310 137.985 40.985 138.155 ;
        RECT 41.180 137.985 41.515 138.155 ;
        RECT 38.420 136.525 38.740 137.485 ;
        RECT 39.270 137.455 40.100 137.755 ;
        RECT 38.910 136.555 39.100 137.275 ;
        RECT 39.270 136.385 39.440 137.455 ;
        RECT 39.900 137.425 40.100 137.455 ;
        RECT 39.610 137.205 39.780 137.275 ;
        RECT 40.310 137.205 40.480 137.985 ;
        RECT 41.345 137.845 41.515 137.985 ;
        RECT 41.685 137.975 41.935 138.435 ;
        RECT 39.610 137.035 40.480 137.205 ;
        RECT 40.650 137.565 41.175 137.785 ;
        RECT 41.345 137.715 41.570 137.845 ;
        RECT 39.610 136.945 40.120 137.035 ;
        RECT 38.080 136.185 38.965 136.355 ;
        RECT 39.190 136.055 39.440 136.385 ;
        RECT 39.610 135.885 39.780 136.685 ;
        RECT 39.950 136.330 40.120 136.945 ;
        RECT 40.650 136.865 40.820 137.565 ;
        RECT 40.290 136.500 40.820 136.865 ;
        RECT 40.990 136.800 41.230 137.395 ;
        RECT 41.400 136.610 41.570 137.715 ;
        RECT 41.740 136.855 42.020 137.805 ;
        RECT 41.265 136.480 41.570 136.610 ;
        RECT 39.950 136.160 41.055 136.330 ;
        RECT 41.265 136.055 41.515 136.480 ;
        RECT 41.685 135.885 41.950 136.345 ;
        RECT 42.190 136.055 42.375 138.175 ;
        RECT 42.545 138.055 42.875 138.435 ;
        RECT 43.045 137.885 43.215 138.175 ;
        RECT 42.550 137.715 43.215 137.885 ;
        RECT 42.550 136.725 42.780 137.715 ;
        RECT 43.475 137.665 46.985 138.435 ;
        RECT 47.155 137.685 48.365 138.435 ;
        RECT 48.535 137.710 48.825 138.435 ;
        RECT 42.950 136.895 43.300 137.545 ;
        RECT 43.475 137.145 45.125 137.665 ;
        RECT 45.295 136.975 46.985 137.495 ;
        RECT 47.155 137.145 47.675 137.685 ;
        RECT 48.995 137.665 52.505 138.435 ;
        RECT 53.135 137.760 53.395 138.265 ;
        RECT 53.575 138.055 53.905 138.435 ;
        RECT 54.085 137.885 54.255 138.265 ;
        RECT 47.845 136.975 48.365 137.515 ;
        RECT 48.995 137.145 50.645 137.665 ;
        RECT 42.550 136.555 43.215 136.725 ;
        RECT 42.545 135.885 42.875 136.385 ;
        RECT 43.045 136.055 43.215 136.555 ;
        RECT 43.475 135.885 46.985 136.975 ;
        RECT 47.155 135.885 48.365 136.975 ;
        RECT 48.535 135.885 48.825 137.050 ;
        RECT 50.815 136.975 52.505 137.495 ;
        RECT 48.995 135.885 52.505 136.975 ;
        RECT 53.135 136.960 53.305 137.760 ;
        RECT 53.590 137.715 54.255 137.885 ;
        RECT 53.590 137.460 53.760 137.715 ;
        RECT 54.515 137.625 54.795 138.435 ;
        RECT 54.965 137.795 55.295 138.265 ;
        RECT 55.465 137.965 55.635 138.435 ;
        RECT 55.805 137.795 56.135 138.265 ;
        RECT 54.965 137.625 56.135 137.795 ;
        RECT 56.305 137.625 56.475 138.435 ;
        RECT 56.825 137.795 56.995 138.075 ;
        RECT 56.645 137.625 56.995 137.795 ;
        RECT 57.205 137.675 57.460 138.435 ;
        RECT 58.195 137.635 58.505 138.435 ;
        RECT 58.710 137.635 59.405 138.265 ;
        RECT 59.740 137.925 59.980 138.435 ;
        RECT 60.160 137.925 60.440 138.255 ;
        RECT 60.670 137.925 60.885 138.435 ;
        RECT 53.475 137.130 53.760 137.460 ;
        RECT 53.995 137.165 54.325 137.535 ;
        RECT 54.910 137.245 55.350 137.455 ;
        RECT 53.590 136.985 53.760 137.130 ;
        RECT 53.135 136.055 53.405 136.960 ;
        RECT 53.590 136.815 54.255 136.985 ;
        RECT 53.575 135.885 53.905 136.645 ;
        RECT 54.085 136.055 54.255 136.815 ;
        RECT 54.515 136.865 55.675 137.075 ;
        RECT 54.515 136.055 54.835 136.865 ;
        RECT 55.005 135.885 55.255 136.695 ;
        RECT 55.425 136.225 55.675 136.865 ;
        RECT 55.845 136.395 56.095 137.625 ;
        RECT 56.645 137.445 56.860 137.625 ;
        RECT 56.305 137.275 56.860 137.445 ;
        RECT 56.690 137.075 56.860 137.275 ;
        RECT 57.030 137.245 57.555 137.455 ;
        RECT 57.340 137.075 57.555 137.245 ;
        RECT 58.205 137.195 58.540 137.465 ;
        RECT 56.265 136.630 56.520 137.075 ;
        RECT 56.690 136.905 56.995 137.075 ;
        RECT 57.335 136.905 57.555 137.075 ;
        RECT 58.710 137.035 58.880 137.635 ;
        RECT 59.050 137.195 59.385 137.445 ;
        RECT 59.635 137.195 59.990 137.755 ;
        RECT 56.265 136.225 56.555 136.630 ;
        RECT 55.425 136.055 56.555 136.225 ;
        RECT 56.825 136.060 56.995 136.905 ;
        RECT 57.340 136.555 57.555 136.905 ;
        RECT 57.205 135.885 57.455 136.375 ;
        RECT 58.195 135.885 58.475 137.025 ;
        RECT 58.645 136.055 58.975 137.035 ;
        RECT 60.160 137.025 60.330 137.925 ;
        RECT 60.500 137.195 60.765 137.755 ;
        RECT 61.055 137.695 61.670 138.265 ;
        RECT 61.015 137.025 61.185 137.525 ;
        RECT 59.145 135.885 59.405 137.025 ;
        RECT 59.760 136.855 61.185 137.025 ;
        RECT 59.760 136.680 60.150 136.855 ;
        RECT 60.635 135.885 60.965 136.685 ;
        RECT 61.355 136.675 61.670 137.695 ;
        RECT 61.990 137.805 62.275 138.265 ;
        RECT 62.445 137.975 62.715 138.435 ;
        RECT 61.990 137.635 62.945 137.805 ;
        RECT 61.875 136.905 62.565 137.465 ;
        RECT 62.735 136.735 62.945 137.635 ;
        RECT 61.135 136.055 61.670 136.675 ;
        RECT 61.990 136.515 62.945 136.735 ;
        RECT 63.115 137.465 63.515 138.265 ;
        RECT 63.705 137.805 63.985 138.265 ;
        RECT 64.505 137.975 64.830 138.435 ;
        RECT 63.705 137.635 64.830 137.805 ;
        RECT 65.000 137.695 65.385 138.265 ;
        RECT 65.555 138.055 66.445 138.225 ;
        RECT 64.380 137.525 64.830 137.635 ;
        RECT 63.115 136.905 64.210 137.465 ;
        RECT 64.380 137.195 64.935 137.525 ;
        RECT 61.990 136.055 62.275 136.515 ;
        RECT 62.445 135.885 62.715 136.345 ;
        RECT 63.115 136.055 63.515 136.905 ;
        RECT 64.380 136.735 64.830 137.195 ;
        RECT 65.105 137.025 65.385 137.695 ;
        RECT 65.555 137.500 66.105 137.885 ;
        RECT 66.275 137.330 66.445 138.055 ;
        RECT 63.705 136.515 64.830 136.735 ;
        RECT 63.705 136.055 63.985 136.515 ;
        RECT 64.505 135.885 64.830 136.345 ;
        RECT 65.000 136.055 65.385 137.025 ;
        RECT 65.555 137.260 66.445 137.330 ;
        RECT 66.615 137.730 66.835 138.215 ;
        RECT 67.005 137.895 67.255 138.435 ;
        RECT 67.425 137.785 67.685 138.265 ;
        RECT 66.615 137.305 66.945 137.730 ;
        RECT 65.555 137.235 66.450 137.260 ;
        RECT 65.555 137.220 66.460 137.235 ;
        RECT 65.555 137.205 66.465 137.220 ;
        RECT 65.555 137.200 66.475 137.205 ;
        RECT 65.555 137.190 66.480 137.200 ;
        RECT 65.555 137.180 66.485 137.190 ;
        RECT 65.555 137.175 66.495 137.180 ;
        RECT 65.555 137.165 66.505 137.175 ;
        RECT 65.555 137.160 66.515 137.165 ;
        RECT 65.555 136.710 65.815 137.160 ;
        RECT 66.180 137.155 66.515 137.160 ;
        RECT 66.180 137.150 66.530 137.155 ;
        RECT 66.180 137.140 66.545 137.150 ;
        RECT 66.180 137.135 66.570 137.140 ;
        RECT 67.115 137.135 67.345 137.530 ;
        RECT 66.180 137.130 67.345 137.135 ;
        RECT 66.210 137.095 67.345 137.130 ;
        RECT 66.245 137.070 67.345 137.095 ;
        RECT 66.275 137.040 67.345 137.070 ;
        RECT 66.295 137.010 67.345 137.040 ;
        RECT 66.315 136.980 67.345 137.010 ;
        RECT 66.385 136.970 67.345 136.980 ;
        RECT 66.410 136.960 67.345 136.970 ;
        RECT 66.430 136.945 67.345 136.960 ;
        RECT 66.450 136.930 67.345 136.945 ;
        RECT 66.455 136.920 67.240 136.930 ;
        RECT 66.470 136.885 67.240 136.920 ;
        RECT 65.985 136.565 66.315 136.810 ;
        RECT 66.485 136.635 67.240 136.885 ;
        RECT 67.515 136.755 67.685 137.785 ;
        RECT 67.855 137.665 69.525 138.435 ;
        RECT 69.700 137.670 70.155 138.435 ;
        RECT 70.430 138.055 71.730 138.265 ;
        RECT 71.985 138.075 72.315 138.435 ;
        RECT 71.560 137.905 71.730 138.055 ;
        RECT 72.485 137.935 72.745 138.265 ;
        RECT 72.515 137.925 72.745 137.935 ;
        RECT 67.855 137.145 68.605 137.665 ;
        RECT 68.775 136.975 69.525 137.495 ;
        RECT 70.630 137.445 70.850 137.845 ;
        RECT 69.695 137.245 70.185 137.445 ;
        RECT 70.375 137.235 70.850 137.445 ;
        RECT 71.095 137.445 71.305 137.845 ;
        RECT 71.560 137.780 72.315 137.905 ;
        RECT 71.560 137.735 72.405 137.780 ;
        RECT 72.135 137.615 72.405 137.735 ;
        RECT 71.095 137.235 71.425 137.445 ;
        RECT 71.595 137.175 72.005 137.480 ;
        RECT 65.985 136.540 66.170 136.565 ;
        RECT 65.555 136.440 66.170 136.540 ;
        RECT 65.555 135.885 66.160 136.440 ;
        RECT 66.335 136.055 66.815 136.395 ;
        RECT 66.985 135.885 67.240 136.430 ;
        RECT 67.410 136.055 67.685 136.755 ;
        RECT 67.855 135.885 69.525 136.975 ;
        RECT 69.700 137.005 70.875 137.065 ;
        RECT 72.235 137.040 72.405 137.615 ;
        RECT 72.205 137.005 72.405 137.040 ;
        RECT 69.700 136.895 72.405 137.005 ;
        RECT 69.700 136.275 69.955 136.895 ;
        RECT 70.545 136.835 72.345 136.895 ;
        RECT 70.545 136.805 70.875 136.835 ;
        RECT 72.575 136.735 72.745 137.925 ;
        RECT 72.915 137.685 74.125 138.435 ;
        RECT 74.295 137.710 74.585 138.435 ;
        RECT 74.805 137.780 75.135 138.215 ;
        RECT 75.305 137.825 75.475 138.435 ;
        RECT 74.755 137.695 75.135 137.780 ;
        RECT 75.645 137.695 75.975 138.220 ;
        RECT 76.235 137.905 76.445 138.435 ;
        RECT 76.720 137.985 77.505 138.155 ;
        RECT 77.675 137.985 78.080 138.155 ;
        RECT 72.915 137.145 73.435 137.685 ;
        RECT 74.755 137.655 74.980 137.695 ;
        RECT 73.605 136.975 74.125 137.515 ;
        RECT 74.755 137.075 74.925 137.655 ;
        RECT 75.645 137.525 75.845 137.695 ;
        RECT 76.720 137.525 76.890 137.985 ;
        RECT 75.095 137.195 75.845 137.525 ;
        RECT 76.015 137.195 76.890 137.525 ;
        RECT 70.205 136.635 70.390 136.725 ;
        RECT 70.980 136.635 71.815 136.645 ;
        RECT 70.205 136.435 71.815 136.635 ;
        RECT 70.205 136.395 70.435 136.435 ;
        RECT 69.700 136.055 70.035 136.275 ;
        RECT 71.040 135.885 71.395 136.265 ;
        RECT 71.565 136.055 71.815 136.435 ;
        RECT 72.065 135.885 72.315 136.665 ;
        RECT 72.485 136.055 72.745 136.735 ;
        RECT 72.915 135.885 74.125 136.975 ;
        RECT 74.295 135.885 74.585 137.050 ;
        RECT 74.755 137.025 74.970 137.075 ;
        RECT 74.755 136.945 75.145 137.025 ;
        RECT 74.815 136.100 75.145 136.945 ;
        RECT 75.655 136.990 75.845 137.195 ;
        RECT 75.315 135.885 75.485 136.895 ;
        RECT 75.655 136.615 76.550 136.990 ;
        RECT 75.655 136.055 75.995 136.615 ;
        RECT 76.225 135.885 76.540 136.385 ;
        RECT 76.720 136.355 76.890 137.195 ;
        RECT 77.060 137.485 77.525 137.815 ;
        RECT 77.910 137.755 78.080 137.985 ;
        RECT 78.260 137.935 78.630 138.435 ;
        RECT 78.950 137.985 79.625 138.155 ;
        RECT 79.820 137.985 80.155 138.155 ;
        RECT 77.060 136.525 77.380 137.485 ;
        RECT 77.910 137.455 78.740 137.755 ;
        RECT 77.550 136.555 77.740 137.275 ;
        RECT 77.910 136.385 78.080 137.455 ;
        RECT 78.540 137.425 78.740 137.455 ;
        RECT 78.250 137.205 78.420 137.275 ;
        RECT 78.950 137.205 79.120 137.985 ;
        RECT 79.985 137.845 80.155 137.985 ;
        RECT 80.325 137.975 80.575 138.435 ;
        RECT 78.250 137.035 79.120 137.205 ;
        RECT 79.290 137.565 79.815 137.785 ;
        RECT 79.985 137.715 80.210 137.845 ;
        RECT 78.250 136.945 78.760 137.035 ;
        RECT 76.720 136.185 77.605 136.355 ;
        RECT 77.830 136.055 78.080 136.385 ;
        RECT 78.250 135.885 78.420 136.685 ;
        RECT 78.590 136.330 78.760 136.945 ;
        RECT 79.290 136.865 79.460 137.565 ;
        RECT 78.930 136.500 79.460 136.865 ;
        RECT 79.630 136.800 79.870 137.395 ;
        RECT 80.040 136.610 80.210 137.715 ;
        RECT 80.380 136.855 80.660 137.805 ;
        RECT 79.905 136.480 80.210 136.610 ;
        RECT 78.590 136.160 79.695 136.330 ;
        RECT 79.905 136.055 80.155 136.480 ;
        RECT 80.325 135.885 80.590 136.345 ;
        RECT 80.830 136.055 81.015 138.175 ;
        RECT 81.185 138.055 81.515 138.435 ;
        RECT 81.685 137.885 81.855 138.175 ;
        RECT 81.190 137.715 81.855 137.885 ;
        RECT 81.190 136.725 81.420 137.715 ;
        RECT 82.115 137.665 84.705 138.435 ;
        RECT 85.425 137.885 85.595 138.265 ;
        RECT 85.810 138.055 86.140 138.435 ;
        RECT 85.425 137.715 86.140 137.885 ;
        RECT 81.590 136.895 81.940 137.545 ;
        RECT 82.115 137.145 83.325 137.665 ;
        RECT 83.495 136.975 84.705 137.495 ;
        RECT 85.335 137.165 85.690 137.535 ;
        RECT 85.970 137.525 86.140 137.715 ;
        RECT 86.310 137.690 86.565 138.265 ;
        RECT 85.970 137.195 86.225 137.525 ;
        RECT 85.970 136.985 86.140 137.195 ;
        RECT 81.190 136.555 81.855 136.725 ;
        RECT 81.185 135.885 81.515 136.385 ;
        RECT 81.685 136.055 81.855 136.555 ;
        RECT 82.115 135.885 84.705 136.975 ;
        RECT 85.425 136.815 86.140 136.985 ;
        RECT 86.395 136.960 86.565 137.690 ;
        RECT 86.740 137.595 87.000 138.435 ;
        RECT 87.175 137.665 88.845 138.435 ;
        RECT 89.105 137.885 89.275 138.175 ;
        RECT 89.445 138.055 89.775 138.435 ;
        RECT 89.105 137.715 89.770 137.885 ;
        RECT 87.175 137.145 87.925 137.665 ;
        RECT 85.425 136.055 85.595 136.815 ;
        RECT 85.810 135.885 86.140 136.645 ;
        RECT 86.310 136.055 86.565 136.960 ;
        RECT 86.740 135.885 87.000 137.035 ;
        RECT 88.095 136.975 88.845 137.495 ;
        RECT 87.175 135.885 88.845 136.975 ;
        RECT 89.020 136.895 89.370 137.545 ;
        RECT 89.540 136.725 89.770 137.715 ;
        RECT 89.105 136.555 89.770 136.725 ;
        RECT 89.105 136.055 89.275 136.555 ;
        RECT 89.445 135.885 89.775 136.385 ;
        RECT 89.945 136.055 90.130 138.175 ;
        RECT 90.385 137.975 90.635 138.435 ;
        RECT 90.805 137.985 91.140 138.155 ;
        RECT 91.335 137.985 92.010 138.155 ;
        RECT 90.805 137.845 90.975 137.985 ;
        RECT 90.300 136.855 90.580 137.805 ;
        RECT 90.750 137.715 90.975 137.845 ;
        RECT 90.750 136.610 90.920 137.715 ;
        RECT 91.145 137.565 91.670 137.785 ;
        RECT 91.090 136.800 91.330 137.395 ;
        RECT 91.500 136.865 91.670 137.565 ;
        RECT 91.840 137.205 92.010 137.985 ;
        RECT 92.330 137.935 92.700 138.435 ;
        RECT 92.880 137.985 93.285 138.155 ;
        RECT 93.455 137.985 94.240 138.155 ;
        RECT 92.880 137.755 93.050 137.985 ;
        RECT 92.220 137.455 93.050 137.755 ;
        RECT 93.435 137.485 93.900 137.815 ;
        RECT 92.220 137.425 92.420 137.455 ;
        RECT 92.540 137.205 92.710 137.275 ;
        RECT 91.840 137.035 92.710 137.205 ;
        RECT 92.200 136.945 92.710 137.035 ;
        RECT 90.750 136.480 91.055 136.610 ;
        RECT 91.500 136.500 92.030 136.865 ;
        RECT 90.370 135.885 90.635 136.345 ;
        RECT 90.805 136.055 91.055 136.480 ;
        RECT 92.200 136.330 92.370 136.945 ;
        RECT 91.265 136.160 92.370 136.330 ;
        RECT 92.540 135.885 92.710 136.685 ;
        RECT 92.880 136.385 93.050 137.455 ;
        RECT 93.220 136.555 93.410 137.275 ;
        RECT 93.580 136.525 93.900 137.485 ;
        RECT 94.070 137.525 94.240 137.985 ;
        RECT 94.515 137.905 94.725 138.435 ;
        RECT 94.985 137.695 95.315 138.220 ;
        RECT 95.485 137.825 95.655 138.435 ;
        RECT 95.825 137.780 96.155 138.215 ;
        RECT 96.375 137.975 96.935 138.265 ;
        RECT 97.105 137.975 97.355 138.435 ;
        RECT 95.825 137.695 96.205 137.780 ;
        RECT 95.115 137.525 95.315 137.695 ;
        RECT 95.980 137.655 96.205 137.695 ;
        RECT 94.070 137.195 94.945 137.525 ;
        RECT 95.115 137.195 95.865 137.525 ;
        RECT 92.880 136.055 93.130 136.385 ;
        RECT 94.070 136.355 94.240 137.195 ;
        RECT 95.115 136.990 95.305 137.195 ;
        RECT 96.035 137.075 96.205 137.655 ;
        RECT 95.990 137.025 96.205 137.075 ;
        RECT 94.410 136.615 95.305 136.990 ;
        RECT 95.815 136.945 96.205 137.025 ;
        RECT 93.355 136.185 94.240 136.355 ;
        RECT 94.420 135.885 94.735 136.385 ;
        RECT 94.965 136.055 95.305 136.615 ;
        RECT 95.475 135.885 95.645 136.895 ;
        RECT 95.815 136.100 96.145 136.945 ;
        RECT 96.375 136.605 96.625 137.975 ;
        RECT 97.975 137.805 98.305 138.165 ;
        RECT 96.915 137.615 98.305 137.805 ;
        RECT 98.675 137.685 99.885 138.435 ;
        RECT 100.055 137.710 100.345 138.435 ;
        RECT 100.605 137.885 100.775 138.265 ;
        RECT 100.990 138.055 101.320 138.435 ;
        RECT 100.605 137.715 101.320 137.885 ;
        RECT 96.915 137.525 97.085 137.615 ;
        RECT 96.795 137.195 97.085 137.525 ;
        RECT 97.255 137.195 97.595 137.445 ;
        RECT 97.815 137.195 98.490 137.445 ;
        RECT 96.915 136.945 97.085 137.195 ;
        RECT 96.915 136.775 97.855 136.945 ;
        RECT 98.225 136.835 98.490 137.195 ;
        RECT 98.675 137.145 99.195 137.685 ;
        RECT 99.365 136.975 99.885 137.515 ;
        RECT 100.515 137.165 100.870 137.535 ;
        RECT 101.150 137.525 101.320 137.715 ;
        RECT 101.490 137.690 101.745 138.265 ;
        RECT 101.150 137.195 101.405 137.525 ;
        RECT 96.375 136.055 96.835 136.605 ;
        RECT 97.025 135.885 97.355 136.605 ;
        RECT 97.555 136.225 97.855 136.775 ;
        RECT 98.025 135.885 98.305 136.555 ;
        RECT 98.675 135.885 99.885 136.975 ;
        RECT 100.055 135.885 100.345 137.050 ;
        RECT 101.150 136.985 101.320 137.195 ;
        RECT 100.605 136.815 101.320 136.985 ;
        RECT 101.575 136.960 101.745 137.690 ;
        RECT 101.920 137.595 102.180 138.435 ;
        RECT 102.360 137.595 102.620 138.435 ;
        RECT 102.795 137.690 103.050 138.265 ;
        RECT 103.220 138.055 103.550 138.435 ;
        RECT 103.765 137.885 103.935 138.265 ;
        RECT 103.220 137.715 103.935 137.885 ;
        RECT 105.205 137.885 105.375 138.175 ;
        RECT 105.545 138.055 105.875 138.435 ;
        RECT 105.205 137.715 105.870 137.885 ;
        RECT 100.605 136.055 100.775 136.815 ;
        RECT 100.990 135.885 101.320 136.645 ;
        RECT 101.490 136.055 101.745 136.960 ;
        RECT 101.920 135.885 102.180 137.035 ;
        RECT 102.360 135.885 102.620 137.035 ;
        RECT 102.795 136.960 102.965 137.690 ;
        RECT 103.220 137.525 103.390 137.715 ;
        RECT 103.135 137.195 103.390 137.525 ;
        RECT 103.220 136.985 103.390 137.195 ;
        RECT 103.670 137.165 104.025 137.535 ;
        RECT 102.795 136.055 103.050 136.960 ;
        RECT 103.220 136.815 103.935 136.985 ;
        RECT 105.120 136.895 105.470 137.545 ;
        RECT 103.220 135.885 103.550 136.645 ;
        RECT 103.765 136.055 103.935 136.815 ;
        RECT 105.640 136.725 105.870 137.715 ;
        RECT 105.205 136.555 105.870 136.725 ;
        RECT 105.205 136.055 105.375 136.555 ;
        RECT 105.545 135.885 105.875 136.385 ;
        RECT 106.045 136.055 106.230 138.175 ;
        RECT 106.485 137.975 106.735 138.435 ;
        RECT 106.905 137.985 107.240 138.155 ;
        RECT 107.435 137.985 108.110 138.155 ;
        RECT 106.905 137.845 107.075 137.985 ;
        RECT 106.400 136.855 106.680 137.805 ;
        RECT 106.850 137.715 107.075 137.845 ;
        RECT 106.850 136.610 107.020 137.715 ;
        RECT 107.245 137.565 107.770 137.785 ;
        RECT 107.190 136.800 107.430 137.395 ;
        RECT 107.600 136.865 107.770 137.565 ;
        RECT 107.940 137.205 108.110 137.985 ;
        RECT 108.430 137.935 108.800 138.435 ;
        RECT 108.980 137.985 109.385 138.155 ;
        RECT 109.555 137.985 110.340 138.155 ;
        RECT 108.980 137.755 109.150 137.985 ;
        RECT 108.320 137.455 109.150 137.755 ;
        RECT 109.535 137.485 110.000 137.815 ;
        RECT 108.320 137.425 108.520 137.455 ;
        RECT 108.640 137.205 108.810 137.275 ;
        RECT 107.940 137.035 108.810 137.205 ;
        RECT 108.300 136.945 108.810 137.035 ;
        RECT 106.850 136.480 107.155 136.610 ;
        RECT 107.600 136.500 108.130 136.865 ;
        RECT 106.470 135.885 106.735 136.345 ;
        RECT 106.905 136.055 107.155 136.480 ;
        RECT 108.300 136.330 108.470 136.945 ;
        RECT 107.365 136.160 108.470 136.330 ;
        RECT 108.640 135.885 108.810 136.685 ;
        RECT 108.980 136.385 109.150 137.455 ;
        RECT 109.320 136.555 109.510 137.275 ;
        RECT 109.680 136.525 110.000 137.485 ;
        RECT 110.170 137.525 110.340 137.985 ;
        RECT 110.615 137.905 110.825 138.435 ;
        RECT 111.085 137.695 111.415 138.220 ;
        RECT 111.585 137.825 111.755 138.435 ;
        RECT 111.925 137.780 112.255 138.215 ;
        RECT 112.475 137.975 113.035 138.265 ;
        RECT 113.205 137.975 113.455 138.435 ;
        RECT 111.925 137.695 112.305 137.780 ;
        RECT 111.215 137.525 111.415 137.695 ;
        RECT 112.080 137.655 112.305 137.695 ;
        RECT 110.170 137.195 111.045 137.525 ;
        RECT 111.215 137.195 111.965 137.525 ;
        RECT 108.980 136.055 109.230 136.385 ;
        RECT 110.170 136.355 110.340 137.195 ;
        RECT 111.215 136.990 111.405 137.195 ;
        RECT 112.135 137.075 112.305 137.655 ;
        RECT 112.090 137.025 112.305 137.075 ;
        RECT 110.510 136.615 111.405 136.990 ;
        RECT 111.915 136.945 112.305 137.025 ;
        RECT 109.455 136.185 110.340 136.355 ;
        RECT 110.520 135.885 110.835 136.385 ;
        RECT 111.065 136.055 111.405 136.615 ;
        RECT 111.575 135.885 111.745 136.895 ;
        RECT 111.915 136.100 112.245 136.945 ;
        RECT 112.475 136.605 112.725 137.975 ;
        RECT 114.075 137.805 114.405 138.165 ;
        RECT 113.015 137.615 114.405 137.805 ;
        RECT 115.240 137.695 115.495 138.265 ;
        RECT 115.665 138.035 115.995 138.435 ;
        RECT 116.420 137.900 116.950 138.265 ;
        RECT 117.140 138.095 117.415 138.265 ;
        RECT 117.135 137.925 117.415 138.095 ;
        RECT 116.420 137.865 116.595 137.900 ;
        RECT 115.665 137.695 116.595 137.865 ;
        RECT 113.015 137.525 113.185 137.615 ;
        RECT 112.895 137.195 113.185 137.525 ;
        RECT 113.355 137.195 113.695 137.445 ;
        RECT 113.915 137.195 114.590 137.445 ;
        RECT 113.015 136.945 113.185 137.195 ;
        RECT 113.015 136.775 113.955 136.945 ;
        RECT 114.325 136.835 114.590 137.195 ;
        RECT 115.240 137.025 115.410 137.695 ;
        RECT 115.665 137.525 115.835 137.695 ;
        RECT 115.580 137.195 115.835 137.525 ;
        RECT 116.060 137.195 116.255 137.525 ;
        RECT 112.475 136.055 112.935 136.605 ;
        RECT 113.125 135.885 113.455 136.605 ;
        RECT 113.655 136.225 113.955 136.775 ;
        RECT 114.125 135.885 114.405 136.555 ;
        RECT 115.240 136.055 115.575 137.025 ;
        RECT 115.745 135.885 115.915 137.025 ;
        RECT 116.085 136.225 116.255 137.195 ;
        RECT 116.425 136.565 116.595 137.695 ;
        RECT 116.765 136.905 116.935 137.705 ;
        RECT 117.140 137.105 117.415 137.925 ;
        RECT 117.585 136.905 117.775 138.265 ;
        RECT 117.955 137.900 118.465 138.435 ;
        RECT 118.685 137.625 118.930 138.230 ;
        RECT 119.375 137.665 121.965 138.435 ;
        RECT 122.595 137.760 122.855 138.265 ;
        RECT 123.035 138.055 123.365 138.435 ;
        RECT 123.545 137.885 123.715 138.265 ;
        RECT 117.975 137.455 119.205 137.625 ;
        RECT 116.765 136.735 117.775 136.905 ;
        RECT 117.945 136.890 118.695 137.080 ;
        RECT 116.425 136.395 117.550 136.565 ;
        RECT 117.945 136.225 118.115 136.890 ;
        RECT 118.865 136.645 119.205 137.455 ;
        RECT 119.375 137.145 120.585 137.665 ;
        RECT 120.755 136.975 121.965 137.495 ;
        RECT 116.085 136.055 118.115 136.225 ;
        RECT 118.285 135.885 118.455 136.645 ;
        RECT 118.690 136.235 119.205 136.645 ;
        RECT 119.375 135.885 121.965 136.975 ;
        RECT 122.595 136.960 122.765 137.760 ;
        RECT 123.050 137.715 123.715 137.885 ;
        RECT 123.050 137.460 123.220 137.715 ;
        RECT 123.975 137.665 125.645 138.435 ;
        RECT 125.815 137.710 126.105 138.435 ;
        RECT 126.280 137.695 126.535 138.265 ;
        RECT 126.705 138.035 127.035 138.435 ;
        RECT 127.460 137.900 127.990 138.265 ;
        RECT 128.180 138.095 128.455 138.265 ;
        RECT 128.175 137.925 128.455 138.095 ;
        RECT 127.460 137.865 127.635 137.900 ;
        RECT 126.705 137.695 127.635 137.865 ;
        RECT 122.935 137.130 123.220 137.460 ;
        RECT 123.455 137.165 123.785 137.535 ;
        RECT 123.975 137.145 124.725 137.665 ;
        RECT 123.050 136.985 123.220 137.130 ;
        RECT 122.595 136.055 122.865 136.960 ;
        RECT 123.050 136.815 123.715 136.985 ;
        RECT 124.895 136.975 125.645 137.495 ;
        RECT 123.035 135.885 123.365 136.645 ;
        RECT 123.545 136.055 123.715 136.815 ;
        RECT 123.975 135.885 125.645 136.975 ;
        RECT 125.815 135.885 126.105 137.050 ;
        RECT 126.280 137.025 126.450 137.695 ;
        RECT 126.705 137.525 126.875 137.695 ;
        RECT 126.620 137.195 126.875 137.525 ;
        RECT 127.100 137.195 127.295 137.525 ;
        RECT 126.280 136.055 126.615 137.025 ;
        RECT 126.785 135.885 126.955 137.025 ;
        RECT 127.125 136.225 127.295 137.195 ;
        RECT 127.465 136.565 127.635 137.695 ;
        RECT 127.805 136.905 127.975 137.705 ;
        RECT 128.180 137.105 128.455 137.925 ;
        RECT 128.625 136.905 128.815 138.265 ;
        RECT 128.995 137.900 129.505 138.435 ;
        RECT 129.725 137.625 129.970 138.230 ;
        RECT 131.335 137.760 131.610 138.105 ;
        RECT 131.800 138.035 132.180 138.435 ;
        RECT 132.350 137.865 132.520 138.215 ;
        RECT 132.690 138.035 133.020 138.435 ;
        RECT 133.195 137.865 133.365 138.215 ;
        RECT 133.565 137.935 133.895 138.435 ;
        RECT 129.015 137.455 130.245 137.625 ;
        RECT 127.805 136.735 128.815 136.905 ;
        RECT 128.985 136.890 129.735 137.080 ;
        RECT 127.465 136.395 128.590 136.565 ;
        RECT 128.985 136.225 129.155 136.890 ;
        RECT 129.905 136.645 130.245 137.455 ;
        RECT 127.125 136.055 129.155 136.225 ;
        RECT 129.325 135.885 129.495 136.645 ;
        RECT 129.730 136.235 130.245 136.645 ;
        RECT 131.335 137.025 131.505 137.760 ;
        RECT 131.780 137.695 133.365 137.865 ;
        RECT 131.780 137.525 131.950 137.695 ;
        RECT 134.090 137.525 134.335 138.215 ;
        RECT 134.505 137.935 134.845 138.435 ;
        RECT 135.030 137.865 135.285 138.215 ;
        RECT 135.455 138.035 135.785 138.435 ;
        RECT 135.955 137.865 136.125 138.215 ;
        RECT 136.295 138.035 136.675 138.435 ;
        RECT 131.675 137.195 131.950 137.525 ;
        RECT 132.120 137.195 132.500 137.525 ;
        RECT 131.780 137.025 131.950 137.195 ;
        RECT 131.335 136.055 131.610 137.025 ;
        RECT 131.780 136.855 132.440 137.025 ;
        RECT 132.670 136.905 133.410 137.525 ;
        RECT 133.680 137.195 134.335 137.525 ;
        RECT 134.505 137.195 134.845 137.765 ;
        RECT 135.030 137.695 136.695 137.865 ;
        RECT 136.865 137.760 137.140 138.105 ;
        RECT 136.525 137.525 136.695 137.695 ;
        RECT 135.015 137.195 135.360 137.525 ;
        RECT 135.530 137.195 136.355 137.525 ;
        RECT 136.525 137.195 136.800 137.525 ;
        RECT 132.270 136.735 132.440 136.855 ;
        RECT 133.580 136.735 133.900 137.025 ;
        RECT 131.820 135.885 132.100 136.685 ;
        RECT 132.270 136.565 133.900 136.735 ;
        RECT 134.095 136.600 134.335 137.195 ;
        RECT 132.270 136.225 134.325 136.395 ;
        RECT 132.270 136.105 134.320 136.225 ;
        RECT 134.505 135.885 134.845 136.960 ;
        RECT 135.035 136.735 135.360 137.025 ;
        RECT 135.530 136.905 135.725 137.195 ;
        RECT 136.525 137.025 136.695 137.195 ;
        RECT 136.970 137.025 137.140 137.760 ;
        RECT 137.315 137.665 139.905 138.435 ;
        RECT 137.315 137.145 138.525 137.665 ;
        RECT 140.075 137.635 140.385 138.435 ;
        RECT 140.590 137.635 141.285 138.265 ;
        RECT 136.035 136.855 136.695 137.025 ;
        RECT 136.035 136.735 136.205 136.855 ;
        RECT 135.035 136.565 136.205 136.735 ;
        RECT 135.015 136.105 136.205 136.395 ;
        RECT 136.375 135.885 136.655 136.685 ;
        RECT 136.865 136.055 137.140 137.025 ;
        RECT 138.695 136.975 139.905 137.495 ;
        RECT 140.085 137.195 140.420 137.465 ;
        RECT 140.590 137.035 140.760 137.635 ;
        RECT 141.455 137.615 141.715 138.435 ;
        RECT 141.885 137.615 142.215 138.035 ;
        RECT 142.395 137.950 143.185 138.215 ;
        RECT 141.965 137.525 142.215 137.615 ;
        RECT 140.930 137.195 141.265 137.445 ;
        RECT 137.315 135.885 139.905 136.975 ;
        RECT 140.075 135.885 140.355 137.025 ;
        RECT 140.525 136.055 140.855 137.035 ;
        RECT 141.025 135.885 141.285 137.025 ;
        RECT 141.455 136.565 141.795 137.445 ;
        RECT 141.965 137.275 142.760 137.525 ;
        RECT 141.455 135.885 141.715 136.395 ;
        RECT 141.965 136.055 142.135 137.275 ;
        RECT 142.930 137.095 143.185 137.950 ;
        RECT 143.355 137.795 143.555 138.215 ;
        RECT 143.745 137.975 144.075 138.435 ;
        RECT 143.355 137.275 143.765 137.795 ;
        RECT 144.245 137.785 144.505 138.265 ;
        RECT 143.935 137.095 144.165 137.525 ;
        RECT 142.375 136.925 144.165 137.095 ;
        RECT 142.375 136.560 142.625 136.925 ;
        RECT 142.795 136.565 143.125 136.755 ;
        RECT 143.345 136.630 144.060 136.925 ;
        RECT 144.335 136.755 144.505 137.785 ;
        RECT 144.735 137.615 144.945 138.435 ;
        RECT 145.115 137.635 145.445 138.265 ;
        RECT 145.115 137.035 145.365 137.635 ;
        RECT 145.615 137.615 145.845 138.435 ;
        RECT 146.605 137.885 146.775 138.265 ;
        RECT 146.955 138.055 147.285 138.435 ;
        RECT 146.605 137.715 147.270 137.885 ;
        RECT 147.465 137.760 147.725 138.265 ;
        RECT 145.535 137.195 145.865 137.445 ;
        RECT 146.535 137.165 146.865 137.535 ;
        RECT 147.100 137.460 147.270 137.715 ;
        RECT 147.100 137.130 147.385 137.460 ;
        RECT 142.795 136.390 142.990 136.565 ;
        RECT 142.375 135.885 142.990 136.390 ;
        RECT 143.160 136.055 143.635 136.395 ;
        RECT 143.805 135.885 144.020 136.430 ;
        RECT 144.230 136.055 144.505 136.755 ;
        RECT 144.735 135.885 144.945 137.025 ;
        RECT 145.115 136.055 145.445 137.035 ;
        RECT 145.615 135.885 145.845 137.025 ;
        RECT 147.100 136.985 147.270 137.130 ;
        RECT 146.605 136.815 147.270 136.985 ;
        RECT 147.555 136.960 147.725 137.760 ;
        RECT 147.985 137.885 148.155 138.265 ;
        RECT 148.335 138.055 148.665 138.435 ;
        RECT 147.985 137.715 148.650 137.885 ;
        RECT 148.845 137.760 149.105 138.265 ;
        RECT 147.915 137.165 148.245 137.535 ;
        RECT 148.480 137.460 148.650 137.715 ;
        RECT 148.480 137.130 148.765 137.460 ;
        RECT 148.480 136.985 148.650 137.130 ;
        RECT 146.605 136.055 146.775 136.815 ;
        RECT 146.955 135.885 147.285 136.645 ;
        RECT 147.455 136.055 147.725 136.960 ;
        RECT 147.985 136.815 148.650 136.985 ;
        RECT 148.935 136.960 149.105 137.760 ;
        RECT 149.275 137.665 150.945 138.435 ;
        RECT 151.575 137.710 151.865 138.435 ;
        RECT 152.035 137.665 155.545 138.435 ;
        RECT 155.715 137.685 156.925 138.435 ;
        RECT 149.275 137.145 150.025 137.665 ;
        RECT 150.195 136.975 150.945 137.495 ;
        RECT 152.035 137.145 153.685 137.665 ;
        RECT 147.985 136.055 148.155 136.815 ;
        RECT 148.335 135.885 148.665 136.645 ;
        RECT 148.835 136.055 149.105 136.960 ;
        RECT 149.275 135.885 150.945 136.975 ;
        RECT 151.575 135.885 151.865 137.050 ;
        RECT 153.855 136.975 155.545 137.495 ;
        RECT 152.035 135.885 155.545 136.975 ;
        RECT 155.715 136.975 156.235 137.515 ;
        RECT 156.405 137.145 156.925 137.685 ;
        RECT 155.715 135.885 156.925 136.975 ;
        RECT 22.690 135.715 157.010 135.885 ;
        RECT 22.775 134.625 23.985 135.715 ;
        RECT 24.155 134.625 27.665 135.715 ;
        RECT 22.775 133.915 23.295 134.455 ;
        RECT 23.465 134.085 23.985 134.625 ;
        RECT 24.155 133.935 25.805 134.455 ;
        RECT 25.975 134.105 27.665 134.625 ;
        RECT 28.755 134.575 29.095 135.545 ;
        RECT 29.265 134.575 29.435 135.715 ;
        RECT 29.705 134.915 29.955 135.715 ;
        RECT 30.600 134.745 30.930 135.545 ;
        RECT 31.230 134.915 31.560 135.715 ;
        RECT 31.730 134.745 32.060 135.545 ;
        RECT 32.445 135.125 32.705 135.515 ;
        RECT 32.875 135.305 33.205 135.715 ;
        RECT 32.445 134.925 33.205 135.125 ;
        RECT 29.625 134.575 32.060 134.745 ;
        RECT 28.755 133.965 28.930 134.575 ;
        RECT 29.625 134.325 29.795 134.575 ;
        RECT 29.100 134.155 29.795 134.325 ;
        RECT 29.970 134.155 30.390 134.355 ;
        RECT 30.560 134.155 30.890 134.355 ;
        RECT 31.060 134.155 31.390 134.355 ;
        RECT 22.775 133.165 23.985 133.915 ;
        RECT 24.155 133.165 27.665 133.935 ;
        RECT 28.755 133.335 29.095 133.965 ;
        RECT 29.265 133.165 29.515 133.965 ;
        RECT 29.705 133.815 30.930 133.985 ;
        RECT 29.705 133.335 30.035 133.815 ;
        RECT 30.205 133.165 30.430 133.625 ;
        RECT 30.600 133.335 30.930 133.815 ;
        RECT 31.560 133.945 31.730 134.575 ;
        RECT 31.915 134.155 32.265 134.405 ;
        RECT 32.455 134.055 32.685 134.745 ;
        RECT 32.865 134.245 33.205 134.925 ;
        RECT 33.395 134.425 33.725 135.535 ;
        RECT 33.895 134.805 34.085 135.535 ;
        RECT 34.255 134.985 34.585 135.715 ;
        RECT 34.765 134.805 34.935 135.535 ;
        RECT 33.895 134.605 34.935 134.805 ;
        RECT 35.655 134.550 35.945 135.715 ;
        RECT 36.150 134.925 36.685 135.545 ;
        RECT 31.560 133.335 32.060 133.945 ;
        RECT 32.865 133.795 33.095 134.245 ;
        RECT 33.395 134.125 33.930 134.425 ;
        RECT 32.715 133.345 33.095 133.795 ;
        RECT 33.275 133.165 33.505 133.945 ;
        RECT 33.685 133.875 33.930 134.125 ;
        RECT 34.110 134.075 34.505 134.425 ;
        RECT 34.700 134.075 34.990 134.425 ;
        RECT 33.685 133.345 34.115 133.875 ;
        RECT 34.295 133.455 34.505 134.075 ;
        RECT 36.150 133.905 36.465 134.925 ;
        RECT 36.855 134.915 37.185 135.715 ;
        RECT 37.670 134.745 38.060 134.920 ;
        RECT 36.635 134.575 38.060 134.745 ;
        RECT 38.415 134.625 41.925 135.715 ;
        RECT 42.645 135.045 42.815 135.545 ;
        RECT 42.985 135.215 43.315 135.715 ;
        RECT 42.645 134.875 43.310 135.045 ;
        RECT 36.635 134.075 36.805 134.575 ;
        RECT 34.675 133.165 35.005 133.895 ;
        RECT 35.655 133.165 35.945 133.890 ;
        RECT 36.150 133.335 36.765 133.905 ;
        RECT 37.055 133.845 37.320 134.405 ;
        RECT 37.490 133.675 37.660 134.575 ;
        RECT 37.830 133.845 38.185 134.405 ;
        RECT 38.415 133.935 40.065 134.455 ;
        RECT 40.235 134.105 41.925 134.625 ;
        RECT 42.560 134.055 42.910 134.705 ;
        RECT 36.935 133.165 37.150 133.675 ;
        RECT 37.380 133.345 37.660 133.675 ;
        RECT 37.840 133.165 38.080 133.675 ;
        RECT 38.415 133.165 41.925 133.935 ;
        RECT 43.080 133.885 43.310 134.875 ;
        RECT 42.645 133.715 43.310 133.885 ;
        RECT 42.645 133.425 42.815 133.715 ;
        RECT 42.985 133.165 43.315 133.545 ;
        RECT 43.485 133.425 43.670 135.545 ;
        RECT 43.910 135.255 44.175 135.715 ;
        RECT 44.345 135.120 44.595 135.545 ;
        RECT 44.805 135.270 45.910 135.440 ;
        RECT 44.290 134.990 44.595 135.120 ;
        RECT 43.840 133.795 44.120 134.745 ;
        RECT 44.290 133.885 44.460 134.990 ;
        RECT 44.630 134.205 44.870 134.800 ;
        RECT 45.040 134.735 45.570 135.100 ;
        RECT 45.040 134.035 45.210 134.735 ;
        RECT 45.740 134.655 45.910 135.270 ;
        RECT 46.080 134.915 46.250 135.715 ;
        RECT 46.420 135.215 46.670 135.545 ;
        RECT 46.895 135.245 47.780 135.415 ;
        RECT 45.740 134.565 46.250 134.655 ;
        RECT 44.290 133.755 44.515 133.885 ;
        RECT 44.685 133.815 45.210 134.035 ;
        RECT 45.380 134.395 46.250 134.565 ;
        RECT 43.925 133.165 44.175 133.625 ;
        RECT 44.345 133.615 44.515 133.755 ;
        RECT 45.380 133.615 45.550 134.395 ;
        RECT 46.080 134.325 46.250 134.395 ;
        RECT 45.760 134.145 45.960 134.175 ;
        RECT 46.420 134.145 46.590 135.215 ;
        RECT 46.760 134.325 46.950 135.045 ;
        RECT 45.760 133.845 46.590 134.145 ;
        RECT 47.120 134.115 47.440 135.075 ;
        RECT 44.345 133.445 44.680 133.615 ;
        RECT 44.875 133.445 45.550 133.615 ;
        RECT 45.870 133.165 46.240 133.665 ;
        RECT 46.420 133.615 46.590 133.845 ;
        RECT 46.975 133.785 47.440 134.115 ;
        RECT 47.610 134.405 47.780 135.245 ;
        RECT 47.960 135.215 48.275 135.715 ;
        RECT 48.505 134.985 48.845 135.545 ;
        RECT 47.950 134.610 48.845 134.985 ;
        RECT 49.015 134.705 49.185 135.715 ;
        RECT 48.655 134.405 48.845 134.610 ;
        RECT 49.355 134.655 49.685 135.500 ;
        RECT 50.005 135.045 50.175 135.545 ;
        RECT 50.345 135.215 50.675 135.715 ;
        RECT 50.005 134.875 50.670 135.045 ;
        RECT 49.355 134.575 49.745 134.655 ;
        RECT 49.530 134.525 49.745 134.575 ;
        RECT 47.610 134.075 48.485 134.405 ;
        RECT 48.655 134.075 49.405 134.405 ;
        RECT 47.610 133.615 47.780 134.075 ;
        RECT 48.655 133.905 48.855 134.075 ;
        RECT 49.575 133.945 49.745 134.525 ;
        RECT 49.920 134.055 50.270 134.705 ;
        RECT 49.520 133.905 49.745 133.945 ;
        RECT 46.420 133.445 46.825 133.615 ;
        RECT 46.995 133.445 47.780 133.615 ;
        RECT 48.055 133.165 48.265 133.695 ;
        RECT 48.525 133.380 48.855 133.905 ;
        RECT 49.365 133.820 49.745 133.905 ;
        RECT 50.440 133.885 50.670 134.875 ;
        RECT 49.025 133.165 49.195 133.775 ;
        RECT 49.365 133.385 49.695 133.820 ;
        RECT 50.005 133.715 50.670 133.885 ;
        RECT 50.005 133.425 50.175 133.715 ;
        RECT 50.345 133.165 50.675 133.545 ;
        RECT 50.845 133.425 51.030 135.545 ;
        RECT 51.270 135.255 51.535 135.715 ;
        RECT 51.705 135.120 51.955 135.545 ;
        RECT 52.165 135.270 53.270 135.440 ;
        RECT 51.650 134.990 51.955 135.120 ;
        RECT 51.200 133.795 51.480 134.745 ;
        RECT 51.650 133.885 51.820 134.990 ;
        RECT 51.990 134.205 52.230 134.800 ;
        RECT 52.400 134.735 52.930 135.100 ;
        RECT 52.400 134.035 52.570 134.735 ;
        RECT 53.100 134.655 53.270 135.270 ;
        RECT 53.440 134.915 53.610 135.715 ;
        RECT 53.780 135.215 54.030 135.545 ;
        RECT 54.255 135.245 55.140 135.415 ;
        RECT 53.100 134.565 53.610 134.655 ;
        RECT 51.650 133.755 51.875 133.885 ;
        RECT 52.045 133.815 52.570 134.035 ;
        RECT 52.740 134.395 53.610 134.565 ;
        RECT 51.285 133.165 51.535 133.625 ;
        RECT 51.705 133.615 51.875 133.755 ;
        RECT 52.740 133.615 52.910 134.395 ;
        RECT 53.440 134.325 53.610 134.395 ;
        RECT 53.120 134.145 53.320 134.175 ;
        RECT 53.780 134.145 53.950 135.215 ;
        RECT 54.120 134.325 54.310 135.045 ;
        RECT 53.120 133.845 53.950 134.145 ;
        RECT 54.480 134.115 54.800 135.075 ;
        RECT 51.705 133.445 52.040 133.615 ;
        RECT 52.235 133.445 52.910 133.615 ;
        RECT 53.230 133.165 53.600 133.665 ;
        RECT 53.780 133.615 53.950 133.845 ;
        RECT 54.335 133.785 54.800 134.115 ;
        RECT 54.970 134.405 55.140 135.245 ;
        RECT 55.320 135.215 55.635 135.715 ;
        RECT 55.865 134.985 56.205 135.545 ;
        RECT 55.310 134.610 56.205 134.985 ;
        RECT 56.375 134.705 56.545 135.715 ;
        RECT 56.015 134.405 56.205 134.610 ;
        RECT 56.715 134.655 57.045 135.500 ;
        RECT 56.715 134.575 57.105 134.655 ;
        RECT 56.890 134.525 57.105 134.575 ;
        RECT 54.970 134.075 55.845 134.405 ;
        RECT 56.015 134.075 56.765 134.405 ;
        RECT 54.970 133.615 55.140 134.075 ;
        RECT 56.015 133.905 56.215 134.075 ;
        RECT 56.935 133.945 57.105 134.525 ;
        RECT 56.880 133.905 57.105 133.945 ;
        RECT 53.780 133.445 54.185 133.615 ;
        RECT 54.355 133.445 55.140 133.615 ;
        RECT 55.415 133.165 55.625 133.695 ;
        RECT 55.885 133.380 56.215 133.905 ;
        RECT 56.725 133.820 57.105 133.905 ;
        RECT 57.275 134.575 57.660 135.545 ;
        RECT 57.830 135.255 58.155 135.715 ;
        RECT 58.675 135.085 58.955 135.545 ;
        RECT 57.830 134.865 58.955 135.085 ;
        RECT 57.275 133.905 57.555 134.575 ;
        RECT 57.830 134.405 58.280 134.865 ;
        RECT 59.145 134.695 59.545 135.545 ;
        RECT 59.945 135.255 60.215 135.715 ;
        RECT 60.385 135.085 60.670 135.545 ;
        RECT 57.725 134.075 58.280 134.405 ;
        RECT 58.450 134.135 59.545 134.695 ;
        RECT 57.830 133.965 58.280 134.075 ;
        RECT 56.385 133.165 56.555 133.775 ;
        RECT 56.725 133.385 57.055 133.820 ;
        RECT 57.275 133.335 57.660 133.905 ;
        RECT 57.830 133.795 58.955 133.965 ;
        RECT 57.830 133.165 58.155 133.625 ;
        RECT 58.675 133.335 58.955 133.795 ;
        RECT 59.145 133.335 59.545 134.135 ;
        RECT 59.715 134.865 60.670 135.085 ;
        RECT 59.715 133.965 59.925 134.865 ;
        RECT 60.095 134.135 60.785 134.695 ;
        RECT 61.415 134.550 61.705 135.715 ;
        RECT 61.965 134.970 62.235 135.715 ;
        RECT 62.865 135.710 69.140 135.715 ;
        RECT 62.405 134.800 62.695 135.540 ;
        RECT 62.865 134.985 63.120 135.710 ;
        RECT 63.305 134.815 63.565 135.540 ;
        RECT 63.735 134.985 63.980 135.710 ;
        RECT 64.165 134.815 64.425 135.540 ;
        RECT 64.595 134.985 64.840 135.710 ;
        RECT 65.025 134.815 65.285 135.540 ;
        RECT 65.455 134.985 65.700 135.710 ;
        RECT 65.870 134.815 66.130 135.540 ;
        RECT 66.300 134.985 66.560 135.710 ;
        RECT 66.730 134.815 66.990 135.540 ;
        RECT 67.160 134.985 67.420 135.710 ;
        RECT 67.590 134.815 67.850 135.540 ;
        RECT 68.020 134.985 68.280 135.710 ;
        RECT 68.450 134.815 68.710 135.540 ;
        RECT 68.880 134.915 69.140 135.710 ;
        RECT 63.305 134.800 68.710 134.815 ;
        RECT 61.965 134.575 68.710 134.800 ;
        RECT 61.965 133.985 63.130 134.575 ;
        RECT 69.310 134.405 69.560 135.540 ;
        RECT 69.740 134.905 70.000 135.715 ;
        RECT 70.175 134.405 70.420 135.545 ;
        RECT 70.600 134.905 70.895 135.715 ;
        RECT 71.075 134.625 72.285 135.715 ;
        RECT 63.300 134.155 70.420 134.405 ;
        RECT 59.715 133.795 60.670 133.965 ;
        RECT 59.945 133.165 60.215 133.625 ;
        RECT 60.385 133.335 60.670 133.795 ;
        RECT 61.415 133.165 61.705 133.890 ;
        RECT 61.965 133.815 68.710 133.985 ;
        RECT 61.965 133.165 62.265 133.645 ;
        RECT 62.435 133.360 62.695 133.815 ;
        RECT 62.865 133.165 63.125 133.645 ;
        RECT 63.305 133.360 63.565 133.815 ;
        RECT 63.735 133.165 63.985 133.645 ;
        RECT 64.165 133.360 64.425 133.815 ;
        RECT 64.595 133.165 64.845 133.645 ;
        RECT 65.025 133.360 65.285 133.815 ;
        RECT 65.455 133.165 65.700 133.645 ;
        RECT 65.870 133.360 66.145 133.815 ;
        RECT 66.315 133.165 66.560 133.645 ;
        RECT 66.730 133.360 66.990 133.815 ;
        RECT 67.160 133.165 67.420 133.645 ;
        RECT 67.590 133.360 67.850 133.815 ;
        RECT 68.020 133.165 68.280 133.645 ;
        RECT 68.450 133.360 68.710 133.815 ;
        RECT 68.880 133.165 69.140 133.725 ;
        RECT 69.310 133.345 69.560 134.155 ;
        RECT 69.740 133.165 70.000 133.690 ;
        RECT 70.170 133.345 70.420 134.155 ;
        RECT 70.590 133.845 70.905 134.405 ;
        RECT 71.075 133.915 71.595 134.455 ;
        RECT 71.765 134.085 72.285 134.625 ;
        RECT 72.605 134.565 72.935 135.715 ;
        RECT 73.105 134.695 73.275 135.545 ;
        RECT 73.445 134.915 73.775 135.715 ;
        RECT 73.945 134.695 74.115 135.545 ;
        RECT 74.295 134.915 74.535 135.715 ;
        RECT 74.705 134.735 75.035 135.545 ;
        RECT 73.105 134.525 74.115 134.695 ;
        RECT 74.320 134.565 75.035 134.735 ;
        RECT 75.215 134.865 75.475 135.545 ;
        RECT 75.645 134.935 75.895 135.715 ;
        RECT 76.145 135.165 76.395 135.545 ;
        RECT 76.565 135.335 76.920 135.715 ;
        RECT 77.925 135.325 78.260 135.545 ;
        RECT 77.525 135.165 77.755 135.205 ;
        RECT 76.145 134.965 77.755 135.165 ;
        RECT 76.145 134.955 76.980 134.965 ;
        RECT 77.570 134.875 77.755 134.965 ;
        RECT 73.105 134.015 73.600 134.525 ;
        RECT 74.320 134.325 74.490 134.565 ;
        RECT 73.990 134.155 74.490 134.325 ;
        RECT 74.660 134.155 75.040 134.395 ;
        RECT 73.105 133.985 73.605 134.015 ;
        RECT 74.320 133.985 74.490 134.155 ;
        RECT 70.600 133.165 70.905 133.675 ;
        RECT 71.075 133.165 72.285 133.915 ;
        RECT 72.605 133.165 72.935 133.965 ;
        RECT 73.105 133.815 74.115 133.985 ;
        RECT 74.320 133.815 74.955 133.985 ;
        RECT 73.105 133.335 73.275 133.815 ;
        RECT 73.445 133.165 73.775 133.645 ;
        RECT 73.945 133.335 74.115 133.815 ;
        RECT 74.365 133.165 74.605 133.645 ;
        RECT 74.785 133.335 74.955 133.815 ;
        RECT 75.215 133.665 75.385 134.865 ;
        RECT 77.085 134.765 77.415 134.795 ;
        RECT 75.615 134.705 77.415 134.765 ;
        RECT 78.005 134.705 78.260 135.325 ;
        RECT 75.555 134.595 78.260 134.705 ;
        RECT 78.435 134.625 79.645 135.715 ;
        RECT 75.555 134.560 75.755 134.595 ;
        RECT 75.555 133.985 75.725 134.560 ;
        RECT 77.085 134.535 78.260 134.595 ;
        RECT 75.955 134.120 76.365 134.425 ;
        RECT 76.535 134.155 76.865 134.365 ;
        RECT 75.555 133.865 75.825 133.985 ;
        RECT 75.555 133.820 76.400 133.865 ;
        RECT 75.645 133.695 76.400 133.820 ;
        RECT 76.655 133.755 76.865 134.155 ;
        RECT 77.110 134.155 77.585 134.365 ;
        RECT 77.775 134.155 78.265 134.355 ;
        RECT 77.110 133.755 77.330 134.155 ;
        RECT 75.215 133.335 75.475 133.665 ;
        RECT 76.230 133.545 76.400 133.695 ;
        RECT 75.645 133.165 75.975 133.525 ;
        RECT 76.230 133.335 77.530 133.545 ;
        RECT 77.805 133.165 78.260 133.930 ;
        RECT 78.435 133.915 78.955 134.455 ;
        RECT 79.125 134.085 79.645 134.625 ;
        RECT 79.815 134.745 80.125 135.545 ;
        RECT 80.295 134.915 80.605 135.715 ;
        RECT 80.775 135.085 81.035 135.545 ;
        RECT 81.205 135.255 81.460 135.715 ;
        RECT 81.635 135.085 81.895 135.545 ;
        RECT 80.775 134.915 81.895 135.085 ;
        RECT 79.815 134.575 80.845 134.745 ;
        RECT 78.435 133.165 79.645 133.915 ;
        RECT 79.815 133.665 79.985 134.575 ;
        RECT 80.155 133.835 80.505 134.405 ;
        RECT 80.675 134.325 80.845 134.575 ;
        RECT 81.635 134.665 81.895 134.915 ;
        RECT 82.065 134.845 82.350 135.715 ;
        RECT 81.635 134.495 82.390 134.665 ;
        RECT 82.575 134.625 86.085 135.715 ;
        RECT 80.675 134.155 81.815 134.325 ;
        RECT 81.985 133.985 82.390 134.495 ;
        RECT 80.740 133.815 82.390 133.985 ;
        RECT 82.575 133.935 84.225 134.455 ;
        RECT 84.395 134.105 86.085 134.625 ;
        RECT 87.175 134.550 87.465 135.715 ;
        RECT 87.635 134.625 91.145 135.715 ;
        RECT 87.635 133.935 89.285 134.455 ;
        RECT 89.455 134.105 91.145 134.625 ;
        RECT 91.315 134.640 91.585 135.545 ;
        RECT 91.755 134.955 92.085 135.715 ;
        RECT 92.265 134.785 92.435 135.545 ;
        RECT 79.815 133.335 80.115 133.665 ;
        RECT 80.285 133.165 80.560 133.645 ;
        RECT 80.740 133.425 81.035 133.815 ;
        RECT 81.205 133.165 81.460 133.645 ;
        RECT 81.635 133.425 81.895 133.815 ;
        RECT 82.065 133.165 82.345 133.645 ;
        RECT 82.575 133.165 86.085 133.935 ;
        RECT 87.175 133.165 87.465 133.890 ;
        RECT 87.635 133.165 91.145 133.935 ;
        RECT 91.315 133.840 91.485 134.640 ;
        RECT 91.770 134.615 92.435 134.785 ;
        RECT 91.770 134.470 91.940 134.615 ;
        RECT 91.655 134.140 91.940 134.470 ;
        RECT 93.160 134.575 93.495 135.545 ;
        RECT 93.665 134.575 93.835 135.715 ;
        RECT 94.005 135.375 96.035 135.545 ;
        RECT 91.770 133.885 91.940 134.140 ;
        RECT 92.175 134.065 92.505 134.435 ;
        RECT 93.160 133.905 93.330 134.575 ;
        RECT 94.005 134.405 94.175 135.375 ;
        RECT 93.500 134.075 93.755 134.405 ;
        RECT 93.980 134.075 94.175 134.405 ;
        RECT 94.345 135.035 95.470 135.205 ;
        RECT 93.585 133.905 93.755 134.075 ;
        RECT 94.345 133.905 94.515 135.035 ;
        RECT 91.315 133.335 91.575 133.840 ;
        RECT 91.770 133.715 92.435 133.885 ;
        RECT 91.755 133.165 92.085 133.545 ;
        RECT 92.265 133.335 92.435 133.715 ;
        RECT 93.160 133.335 93.415 133.905 ;
        RECT 93.585 133.735 94.515 133.905 ;
        RECT 94.685 134.695 95.695 134.865 ;
        RECT 94.685 133.895 94.855 134.695 ;
        RECT 95.060 134.355 95.335 134.495 ;
        RECT 95.055 134.185 95.335 134.355 ;
        RECT 94.340 133.700 94.515 133.735 ;
        RECT 93.585 133.165 93.915 133.565 ;
        RECT 94.340 133.335 94.870 133.700 ;
        RECT 95.060 133.335 95.335 134.185 ;
        RECT 95.505 133.335 95.695 134.695 ;
        RECT 95.865 134.710 96.035 135.375 ;
        RECT 96.205 134.955 96.375 135.715 ;
        RECT 96.610 134.955 97.125 135.365 ;
        RECT 97.315 135.205 97.615 135.715 ;
        RECT 97.785 135.205 98.165 135.375 ;
        RECT 98.745 135.205 99.375 135.715 ;
        RECT 97.785 135.035 97.955 135.205 ;
        RECT 99.545 135.035 99.875 135.545 ;
        RECT 100.045 135.205 100.345 135.715 ;
        RECT 95.865 134.520 96.615 134.710 ;
        RECT 96.785 134.145 97.125 134.955 ;
        RECT 95.895 133.975 97.125 134.145 ;
        RECT 97.295 134.835 97.955 135.035 ;
        RECT 98.125 134.865 100.345 135.035 ;
        RECT 95.875 133.165 96.385 133.700 ;
        RECT 96.605 133.370 96.850 133.975 ;
        RECT 97.295 133.905 97.465 134.835 ;
        RECT 98.125 134.665 98.295 134.865 ;
        RECT 97.635 134.495 98.295 134.665 ;
        RECT 98.465 134.525 100.005 134.695 ;
        RECT 97.635 134.075 97.805 134.495 ;
        RECT 98.465 134.325 98.635 134.525 ;
        RECT 98.035 134.155 98.635 134.325 ;
        RECT 98.805 134.155 99.500 134.355 ;
        RECT 99.760 134.075 100.005 134.525 ;
        RECT 98.125 133.905 99.035 133.985 ;
        RECT 97.295 133.425 97.615 133.905 ;
        RECT 97.785 133.815 99.035 133.905 ;
        RECT 97.785 133.735 98.295 133.815 ;
        RECT 97.785 133.335 98.015 133.735 ;
        RECT 98.185 133.165 98.535 133.555 ;
        RECT 98.705 133.335 99.035 133.815 ;
        RECT 99.205 133.165 99.375 133.985 ;
        RECT 100.175 133.905 100.345 134.865 ;
        RECT 99.880 133.360 100.345 133.905 ;
        RECT 100.515 134.575 100.900 135.545 ;
        RECT 101.070 135.255 101.395 135.715 ;
        RECT 101.915 135.085 102.195 135.545 ;
        RECT 101.070 134.865 102.195 135.085 ;
        RECT 100.515 133.905 100.795 134.575 ;
        RECT 101.070 134.405 101.520 134.865 ;
        RECT 102.385 134.695 102.785 135.545 ;
        RECT 103.185 135.255 103.455 135.715 ;
        RECT 103.625 135.085 103.910 135.545 ;
        RECT 100.965 134.075 101.520 134.405 ;
        RECT 101.690 134.135 102.785 134.695 ;
        RECT 101.070 133.965 101.520 134.075 ;
        RECT 100.515 133.335 100.900 133.905 ;
        RECT 101.070 133.795 102.195 133.965 ;
        RECT 101.070 133.165 101.395 133.625 ;
        RECT 101.915 133.335 102.195 133.795 ;
        RECT 102.385 133.335 102.785 134.135 ;
        RECT 102.955 134.865 103.910 135.085 ;
        RECT 102.955 133.965 103.165 134.865 ;
        RECT 103.335 134.135 104.025 134.695 ;
        RECT 104.195 134.625 106.785 135.715 ;
        RECT 102.955 133.795 103.910 133.965 ;
        RECT 103.185 133.165 103.455 133.625 ;
        RECT 103.625 133.335 103.910 133.795 ;
        RECT 104.195 133.935 105.405 134.455 ;
        RECT 105.575 134.105 106.785 134.625 ;
        RECT 107.505 134.785 107.675 135.545 ;
        RECT 107.855 134.955 108.185 135.715 ;
        RECT 107.505 134.615 108.170 134.785 ;
        RECT 108.355 134.640 108.625 135.545 ;
        RECT 108.000 134.470 108.170 134.615 ;
        RECT 107.435 134.065 107.765 134.435 ;
        RECT 108.000 134.140 108.285 134.470 ;
        RECT 104.195 133.165 106.785 133.935 ;
        RECT 108.000 133.885 108.170 134.140 ;
        RECT 107.505 133.715 108.170 133.885 ;
        RECT 108.455 133.840 108.625 134.640 ;
        RECT 108.795 134.625 110.465 135.715 ;
        RECT 107.505 133.335 107.675 133.715 ;
        RECT 107.855 133.165 108.185 133.545 ;
        RECT 108.365 133.335 108.625 133.840 ;
        RECT 108.795 133.935 109.545 134.455 ;
        RECT 109.715 134.105 110.465 134.625 ;
        RECT 110.635 134.995 111.095 135.545 ;
        RECT 111.285 134.995 111.615 135.715 ;
        RECT 108.795 133.165 110.465 133.935 ;
        RECT 110.635 133.625 110.885 134.995 ;
        RECT 111.815 134.825 112.115 135.375 ;
        RECT 112.285 135.045 112.565 135.715 ;
        RECT 111.175 134.655 112.115 134.825 ;
        RECT 111.175 134.405 111.345 134.655 ;
        RECT 112.485 134.405 112.750 134.765 ;
        RECT 112.935 134.550 113.225 135.715 ;
        RECT 113.405 134.905 113.700 135.715 ;
        RECT 113.880 134.405 114.125 135.545 ;
        RECT 114.300 134.905 114.560 135.715 ;
        RECT 115.160 135.710 121.435 135.715 ;
        RECT 114.740 134.405 114.990 135.540 ;
        RECT 115.160 134.915 115.420 135.710 ;
        RECT 115.590 134.815 115.850 135.540 ;
        RECT 116.020 134.985 116.280 135.710 ;
        RECT 116.450 134.815 116.710 135.540 ;
        RECT 116.880 134.985 117.140 135.710 ;
        RECT 117.310 134.815 117.570 135.540 ;
        RECT 117.740 134.985 118.000 135.710 ;
        RECT 118.170 134.815 118.430 135.540 ;
        RECT 118.600 134.985 118.845 135.710 ;
        RECT 119.015 134.815 119.275 135.540 ;
        RECT 119.460 134.985 119.705 135.710 ;
        RECT 119.875 134.815 120.135 135.540 ;
        RECT 120.320 134.985 120.565 135.710 ;
        RECT 120.735 134.815 120.995 135.540 ;
        RECT 121.180 134.985 121.435 135.710 ;
        RECT 115.590 134.800 120.995 134.815 ;
        RECT 121.605 134.800 121.895 135.540 ;
        RECT 122.065 134.970 122.335 135.715 ;
        RECT 115.590 134.575 122.335 134.800 ;
        RECT 122.685 134.785 122.855 135.545 ;
        RECT 123.070 134.955 123.400 135.715 ;
        RECT 122.685 134.615 123.400 134.785 ;
        RECT 123.570 134.640 123.825 135.545 ;
        RECT 111.055 134.075 111.345 134.405 ;
        RECT 111.515 134.155 111.855 134.405 ;
        RECT 112.075 134.155 112.750 134.405 ;
        RECT 111.175 133.985 111.345 134.075 ;
        RECT 111.175 133.795 112.565 133.985 ;
        RECT 110.635 133.335 111.195 133.625 ;
        RECT 111.365 133.165 111.615 133.625 ;
        RECT 112.235 133.435 112.565 133.795 ;
        RECT 112.935 133.165 113.225 133.890 ;
        RECT 113.395 133.845 113.710 134.405 ;
        RECT 113.880 134.155 121.000 134.405 ;
        RECT 113.395 133.165 113.700 133.675 ;
        RECT 113.880 133.345 114.130 134.155 ;
        RECT 114.300 133.165 114.560 133.690 ;
        RECT 114.740 133.345 114.990 134.155 ;
        RECT 121.170 133.985 122.335 134.575 ;
        RECT 122.595 134.065 122.950 134.435 ;
        RECT 123.230 134.405 123.400 134.615 ;
        RECT 123.230 134.075 123.485 134.405 ;
        RECT 115.590 133.815 122.335 133.985 ;
        RECT 123.230 133.885 123.400 134.075 ;
        RECT 123.655 133.910 123.825 134.640 ;
        RECT 124.000 134.565 124.260 135.715 ;
        RECT 124.435 134.575 124.695 135.715 ;
        RECT 124.865 134.565 125.195 135.545 ;
        RECT 125.365 134.575 125.645 135.715 ;
        RECT 125.815 135.280 131.160 135.715 ;
        RECT 131.335 135.280 136.680 135.715 ;
        RECT 124.455 134.155 124.790 134.405 ;
        RECT 115.160 133.165 115.420 133.725 ;
        RECT 115.590 133.360 115.850 133.815 ;
        RECT 116.020 133.165 116.280 133.645 ;
        RECT 116.450 133.360 116.710 133.815 ;
        RECT 116.880 133.165 117.140 133.645 ;
        RECT 117.310 133.360 117.570 133.815 ;
        RECT 117.740 133.165 117.985 133.645 ;
        RECT 118.155 133.360 118.430 133.815 ;
        RECT 118.600 133.165 118.845 133.645 ;
        RECT 119.015 133.360 119.275 133.815 ;
        RECT 119.455 133.165 119.705 133.645 ;
        RECT 119.875 133.360 120.135 133.815 ;
        RECT 120.315 133.165 120.565 133.645 ;
        RECT 120.735 133.360 120.995 133.815 ;
        RECT 121.175 133.165 121.435 133.645 ;
        RECT 121.605 133.360 121.865 133.815 ;
        RECT 122.685 133.715 123.400 133.885 ;
        RECT 122.035 133.165 122.335 133.645 ;
        RECT 122.685 133.335 122.855 133.715 ;
        RECT 123.070 133.165 123.400 133.545 ;
        RECT 123.570 133.335 123.825 133.910 ;
        RECT 124.000 133.165 124.260 134.005 ;
        RECT 124.960 133.965 125.130 134.565 ;
        RECT 125.300 134.135 125.635 134.405 ;
        RECT 124.435 133.335 125.130 133.965 ;
        RECT 125.335 133.165 125.645 133.965 ;
        RECT 127.400 133.710 127.740 134.540 ;
        RECT 129.220 134.030 129.570 135.280 ;
        RECT 132.920 133.710 133.260 134.540 ;
        RECT 134.740 134.030 135.090 135.280 ;
        RECT 136.855 134.625 138.525 135.715 ;
        RECT 136.855 133.935 137.605 134.455 ;
        RECT 137.775 134.105 138.525 134.625 ;
        RECT 138.695 134.550 138.985 135.715 ;
        RECT 140.075 134.745 140.345 135.515 ;
        RECT 140.515 134.935 140.845 135.715 ;
        RECT 141.050 135.110 141.235 135.515 ;
        RECT 141.405 135.290 141.740 135.715 ;
        RECT 141.050 134.935 141.715 135.110 ;
        RECT 140.075 134.575 141.205 134.745 ;
        RECT 125.815 133.165 131.160 133.710 ;
        RECT 131.335 133.165 136.680 133.710 ;
        RECT 136.855 133.165 138.525 133.935 ;
        RECT 138.695 133.165 138.985 133.890 ;
        RECT 140.075 133.665 140.245 134.575 ;
        RECT 140.415 133.825 140.775 134.405 ;
        RECT 140.955 134.075 141.205 134.575 ;
        RECT 141.375 133.905 141.715 134.935 ;
        RECT 141.915 134.625 145.425 135.715 ;
        RECT 145.595 134.625 146.805 135.715 ;
        RECT 147.035 134.655 147.365 135.500 ;
        RECT 147.535 134.705 147.705 135.715 ;
        RECT 147.875 134.985 148.215 135.545 ;
        RECT 148.445 135.215 148.760 135.715 ;
        RECT 148.940 135.245 149.825 135.415 ;
        RECT 141.030 133.735 141.715 133.905 ;
        RECT 141.915 133.935 143.565 134.455 ;
        RECT 143.735 134.105 145.425 134.625 ;
        RECT 140.075 133.335 140.335 133.665 ;
        RECT 140.545 133.165 140.820 133.645 ;
        RECT 141.030 133.335 141.235 133.735 ;
        RECT 141.405 133.165 141.740 133.565 ;
        RECT 141.915 133.165 145.425 133.935 ;
        RECT 145.595 133.915 146.115 134.455 ;
        RECT 146.285 134.085 146.805 134.625 ;
        RECT 146.975 134.575 147.365 134.655 ;
        RECT 147.875 134.610 148.770 134.985 ;
        RECT 146.975 134.525 147.190 134.575 ;
        RECT 146.975 133.945 147.145 134.525 ;
        RECT 147.875 134.405 148.065 134.610 ;
        RECT 148.940 134.405 149.110 135.245 ;
        RECT 150.050 135.215 150.300 135.545 ;
        RECT 147.315 134.075 148.065 134.405 ;
        RECT 148.235 134.075 149.110 134.405 ;
        RECT 145.595 133.165 146.805 133.915 ;
        RECT 146.975 133.905 147.200 133.945 ;
        RECT 147.865 133.905 148.065 134.075 ;
        RECT 146.975 133.820 147.355 133.905 ;
        RECT 147.025 133.385 147.355 133.820 ;
        RECT 147.525 133.165 147.695 133.775 ;
        RECT 147.865 133.380 148.195 133.905 ;
        RECT 148.455 133.165 148.665 133.695 ;
        RECT 148.940 133.615 149.110 134.075 ;
        RECT 149.280 134.115 149.600 135.075 ;
        RECT 149.770 134.325 149.960 135.045 ;
        RECT 150.130 134.145 150.300 135.215 ;
        RECT 150.470 134.915 150.640 135.715 ;
        RECT 150.810 135.270 151.915 135.440 ;
        RECT 150.810 134.655 150.980 135.270 ;
        RECT 152.125 135.120 152.375 135.545 ;
        RECT 152.545 135.255 152.810 135.715 ;
        RECT 151.150 134.735 151.680 135.100 ;
        RECT 152.125 134.990 152.430 135.120 ;
        RECT 150.470 134.565 150.980 134.655 ;
        RECT 150.470 134.395 151.340 134.565 ;
        RECT 150.470 134.325 150.640 134.395 ;
        RECT 150.760 134.145 150.960 134.175 ;
        RECT 149.280 133.785 149.745 134.115 ;
        RECT 150.130 133.845 150.960 134.145 ;
        RECT 150.130 133.615 150.300 133.845 ;
        RECT 148.940 133.445 149.725 133.615 ;
        RECT 149.895 133.445 150.300 133.615 ;
        RECT 150.480 133.165 150.850 133.665 ;
        RECT 151.170 133.615 151.340 134.395 ;
        RECT 151.510 134.035 151.680 134.735 ;
        RECT 151.850 134.205 152.090 134.800 ;
        RECT 151.510 133.815 152.035 134.035 ;
        RECT 152.260 133.885 152.430 134.990 ;
        RECT 152.205 133.755 152.430 133.885 ;
        RECT 152.600 133.795 152.880 134.745 ;
        RECT 152.205 133.615 152.375 133.755 ;
        RECT 151.170 133.445 151.845 133.615 ;
        RECT 152.040 133.445 152.375 133.615 ;
        RECT 152.545 133.165 152.795 133.625 ;
        RECT 153.050 133.425 153.235 135.545 ;
        RECT 153.405 135.215 153.735 135.715 ;
        RECT 153.905 135.045 154.075 135.545 ;
        RECT 153.410 134.875 154.075 135.045 ;
        RECT 153.410 133.885 153.640 134.875 ;
        RECT 153.810 134.055 154.160 134.705 ;
        RECT 154.335 134.625 155.545 135.715 ;
        RECT 154.335 133.915 154.855 134.455 ;
        RECT 155.025 134.085 155.545 134.625 ;
        RECT 155.715 134.625 156.925 135.715 ;
        RECT 155.715 134.085 156.235 134.625 ;
        RECT 156.405 133.915 156.925 134.455 ;
        RECT 153.410 133.715 154.075 133.885 ;
        RECT 153.405 133.165 153.735 133.545 ;
        RECT 153.905 133.425 154.075 133.715 ;
        RECT 154.335 133.165 155.545 133.915 ;
        RECT 155.715 133.165 156.925 133.915 ;
        RECT 22.690 132.995 157.010 133.165 ;
        RECT 22.775 132.245 23.985 132.995 ;
        RECT 22.775 131.705 23.295 132.245 ;
        RECT 24.615 132.195 24.955 132.825 ;
        RECT 25.125 132.195 25.375 132.995 ;
        RECT 25.565 132.345 25.895 132.825 ;
        RECT 26.065 132.535 26.290 132.995 ;
        RECT 26.460 132.345 26.790 132.825 ;
        RECT 23.465 131.535 23.985 132.075 ;
        RECT 22.775 130.445 23.985 131.535 ;
        RECT 24.615 131.585 24.790 132.195 ;
        RECT 25.565 132.175 26.790 132.345 ;
        RECT 27.420 132.215 27.920 132.825 ;
        RECT 28.870 132.365 29.155 132.825 ;
        RECT 29.325 132.535 29.595 132.995 ;
        RECT 24.960 131.835 25.655 132.005 ;
        RECT 25.485 131.585 25.655 131.835 ;
        RECT 25.830 131.805 26.250 132.005 ;
        RECT 26.420 131.805 26.750 132.005 ;
        RECT 26.920 131.805 27.250 132.005 ;
        RECT 27.420 131.585 27.590 132.215 ;
        RECT 28.870 132.195 29.825 132.365 ;
        RECT 27.775 131.755 28.125 132.005 ;
        RECT 24.615 130.615 24.955 131.585 ;
        RECT 25.125 130.445 25.295 131.585 ;
        RECT 25.485 131.415 27.920 131.585 ;
        RECT 28.755 131.465 29.445 132.025 ;
        RECT 25.565 130.445 25.815 131.245 ;
        RECT 26.460 130.615 26.790 131.415 ;
        RECT 27.090 130.445 27.420 131.245 ;
        RECT 27.590 130.615 27.920 131.415 ;
        RECT 29.615 131.295 29.825 132.195 ;
        RECT 28.870 131.075 29.825 131.295 ;
        RECT 29.995 132.025 30.395 132.825 ;
        RECT 30.585 132.365 30.865 132.825 ;
        RECT 31.385 132.535 31.710 132.995 ;
        RECT 30.585 132.195 31.710 132.365 ;
        RECT 31.880 132.255 32.265 132.825 ;
        RECT 31.260 132.085 31.710 132.195 ;
        RECT 29.995 131.465 31.090 132.025 ;
        RECT 31.260 131.755 31.815 132.085 ;
        RECT 28.870 130.615 29.155 131.075 ;
        RECT 29.325 130.445 29.595 130.905 ;
        RECT 29.995 130.615 30.395 131.465 ;
        RECT 31.260 131.295 31.710 131.755 ;
        RECT 31.985 131.585 32.265 132.255 ;
        RECT 30.585 131.075 31.710 131.295 ;
        RECT 30.585 130.615 30.865 131.075 ;
        RECT 31.385 130.445 31.710 130.905 ;
        RECT 31.880 130.615 32.265 131.585 ;
        RECT 32.435 132.255 32.820 132.825 ;
        RECT 32.990 132.535 33.315 132.995 ;
        RECT 33.835 132.365 34.115 132.825 ;
        RECT 32.435 131.585 32.715 132.255 ;
        RECT 32.990 132.195 34.115 132.365 ;
        RECT 32.990 132.085 33.440 132.195 ;
        RECT 32.885 131.755 33.440 132.085 ;
        RECT 34.305 132.025 34.705 132.825 ;
        RECT 35.105 132.535 35.375 132.995 ;
        RECT 35.545 132.365 35.830 132.825 ;
        RECT 32.435 130.615 32.820 131.585 ;
        RECT 32.990 131.295 33.440 131.755 ;
        RECT 33.610 131.465 34.705 132.025 ;
        RECT 32.990 131.075 34.115 131.295 ;
        RECT 32.990 130.445 33.315 130.905 ;
        RECT 33.835 130.615 34.115 131.075 ;
        RECT 34.305 130.615 34.705 131.465 ;
        RECT 34.875 132.195 35.830 132.365 ;
        RECT 36.205 132.445 36.375 132.735 ;
        RECT 36.545 132.615 36.875 132.995 ;
        RECT 36.205 132.275 36.870 132.445 ;
        RECT 34.875 131.295 35.085 132.195 ;
        RECT 35.255 131.465 35.945 132.025 ;
        RECT 36.120 131.455 36.470 132.105 ;
        RECT 34.875 131.075 35.830 131.295 ;
        RECT 36.640 131.285 36.870 132.275 ;
        RECT 35.105 130.445 35.375 130.905 ;
        RECT 35.545 130.615 35.830 131.075 ;
        RECT 36.205 131.115 36.870 131.285 ;
        RECT 36.205 130.615 36.375 131.115 ;
        RECT 36.545 130.445 36.875 130.945 ;
        RECT 37.045 130.615 37.230 132.735 ;
        RECT 37.485 132.535 37.735 132.995 ;
        RECT 37.905 132.545 38.240 132.715 ;
        RECT 38.435 132.545 39.110 132.715 ;
        RECT 37.905 132.405 38.075 132.545 ;
        RECT 37.400 131.415 37.680 132.365 ;
        RECT 37.850 132.275 38.075 132.405 ;
        RECT 37.850 131.170 38.020 132.275 ;
        RECT 38.245 132.125 38.770 132.345 ;
        RECT 38.190 131.360 38.430 131.955 ;
        RECT 38.600 131.425 38.770 132.125 ;
        RECT 38.940 131.765 39.110 132.545 ;
        RECT 39.430 132.495 39.800 132.995 ;
        RECT 39.980 132.545 40.385 132.715 ;
        RECT 40.555 132.545 41.340 132.715 ;
        RECT 39.980 132.315 40.150 132.545 ;
        RECT 39.320 132.015 40.150 132.315 ;
        RECT 40.535 132.045 41.000 132.375 ;
        RECT 39.320 131.985 39.520 132.015 ;
        RECT 39.640 131.765 39.810 131.835 ;
        RECT 38.940 131.595 39.810 131.765 ;
        RECT 39.300 131.505 39.810 131.595 ;
        RECT 37.850 131.040 38.155 131.170 ;
        RECT 38.600 131.060 39.130 131.425 ;
        RECT 37.470 130.445 37.735 130.905 ;
        RECT 37.905 130.615 38.155 131.040 ;
        RECT 39.300 130.890 39.470 131.505 ;
        RECT 38.365 130.720 39.470 130.890 ;
        RECT 39.640 130.445 39.810 131.245 ;
        RECT 39.980 130.945 40.150 132.015 ;
        RECT 40.320 131.115 40.510 131.835 ;
        RECT 40.680 131.085 41.000 132.045 ;
        RECT 41.170 132.085 41.340 132.545 ;
        RECT 41.615 132.465 41.825 132.995 ;
        RECT 42.085 132.255 42.415 132.780 ;
        RECT 42.585 132.385 42.755 132.995 ;
        RECT 42.925 132.340 43.255 132.775 ;
        RECT 42.925 132.255 43.305 132.340 ;
        RECT 42.215 132.085 42.415 132.255 ;
        RECT 43.080 132.215 43.305 132.255 ;
        RECT 41.170 131.755 42.045 132.085 ;
        RECT 42.215 131.755 42.965 132.085 ;
        RECT 39.980 130.615 40.230 130.945 ;
        RECT 41.170 130.915 41.340 131.755 ;
        RECT 42.215 131.550 42.405 131.755 ;
        RECT 43.135 131.635 43.305 132.215 ;
        RECT 43.090 131.585 43.305 131.635 ;
        RECT 41.510 131.175 42.405 131.550 ;
        RECT 42.915 131.505 43.305 131.585 ;
        RECT 43.475 132.255 43.860 132.825 ;
        RECT 44.030 132.535 44.355 132.995 ;
        RECT 44.875 132.365 45.155 132.825 ;
        RECT 43.475 131.585 43.755 132.255 ;
        RECT 44.030 132.195 45.155 132.365 ;
        RECT 44.030 132.085 44.480 132.195 ;
        RECT 43.925 131.755 44.480 132.085 ;
        RECT 45.345 132.025 45.745 132.825 ;
        RECT 46.145 132.535 46.415 132.995 ;
        RECT 46.585 132.365 46.870 132.825 ;
        RECT 40.455 130.745 41.340 130.915 ;
        RECT 41.520 130.445 41.835 130.945 ;
        RECT 42.065 130.615 42.405 131.175 ;
        RECT 42.575 130.445 42.745 131.455 ;
        RECT 42.915 130.660 43.245 131.505 ;
        RECT 43.475 130.615 43.860 131.585 ;
        RECT 44.030 131.295 44.480 131.755 ;
        RECT 44.650 131.465 45.745 132.025 ;
        RECT 44.030 131.075 45.155 131.295 ;
        RECT 44.030 130.445 44.355 130.905 ;
        RECT 44.875 130.615 45.155 131.075 ;
        RECT 45.345 130.615 45.745 131.465 ;
        RECT 45.915 132.195 46.870 132.365 ;
        RECT 45.915 131.295 46.125 132.195 ;
        RECT 47.215 132.175 47.425 132.995 ;
        RECT 47.595 132.195 47.925 132.825 ;
        RECT 46.295 131.465 46.985 132.025 ;
        RECT 47.595 131.595 47.845 132.195 ;
        RECT 48.095 132.175 48.325 132.995 ;
        RECT 48.535 132.270 48.825 132.995 ;
        RECT 48.995 132.495 49.295 132.825 ;
        RECT 49.465 132.515 49.740 132.995 ;
        RECT 48.015 131.755 48.345 132.005 ;
        RECT 45.915 131.075 46.870 131.295 ;
        RECT 46.145 130.445 46.415 130.905 ;
        RECT 46.585 130.615 46.870 131.075 ;
        RECT 47.215 130.445 47.425 131.585 ;
        RECT 47.595 130.615 47.925 131.595 ;
        RECT 48.095 130.445 48.325 131.585 ;
        RECT 48.535 130.445 48.825 131.610 ;
        RECT 48.995 131.585 49.165 132.495 ;
        RECT 49.920 132.345 50.215 132.735 ;
        RECT 50.385 132.515 50.640 132.995 ;
        RECT 50.815 132.345 51.075 132.735 ;
        RECT 51.245 132.515 51.525 132.995 ;
        RECT 51.955 132.365 52.285 132.725 ;
        RECT 52.905 132.535 53.155 132.995 ;
        RECT 53.325 132.535 53.885 132.825 ;
        RECT 49.335 131.755 49.685 132.325 ;
        RECT 49.920 132.175 51.570 132.345 ;
        RECT 51.955 132.175 53.345 132.365 ;
        RECT 49.855 131.835 50.995 132.005 ;
        RECT 49.855 131.585 50.025 131.835 ;
        RECT 51.165 131.665 51.570 132.175 ;
        RECT 53.175 132.085 53.345 132.175 ;
        RECT 48.995 131.415 50.025 131.585 ;
        RECT 50.815 131.495 51.570 131.665 ;
        RECT 51.770 131.755 52.445 132.005 ;
        RECT 52.665 131.755 53.005 132.005 ;
        RECT 53.175 131.755 53.465 132.085 ;
        RECT 48.995 130.615 49.305 131.415 ;
        RECT 50.815 131.245 51.075 131.495 ;
        RECT 51.770 131.395 52.035 131.755 ;
        RECT 53.175 131.505 53.345 131.755 ;
        RECT 52.405 131.335 53.345 131.505 ;
        RECT 49.475 130.445 49.785 131.245 ;
        RECT 49.955 131.075 51.075 131.245 ;
        RECT 49.955 130.615 50.215 131.075 ;
        RECT 50.385 130.445 50.640 130.905 ;
        RECT 50.815 130.615 51.075 131.075 ;
        RECT 51.245 130.445 51.530 131.315 ;
        RECT 51.955 130.445 52.235 131.115 ;
        RECT 52.405 130.785 52.705 131.335 ;
        RECT 53.635 131.165 53.885 132.535 ;
        RECT 54.060 132.175 54.335 132.995 ;
        RECT 54.505 132.355 54.835 132.825 ;
        RECT 55.005 132.525 55.175 132.995 ;
        RECT 55.345 132.355 55.675 132.825 ;
        RECT 55.845 132.525 56.015 132.995 ;
        RECT 56.185 132.355 56.515 132.825 ;
        RECT 56.685 132.525 56.855 132.995 ;
        RECT 57.025 132.355 57.355 132.825 ;
        RECT 57.525 132.525 57.810 132.995 ;
        RECT 59.115 132.615 60.005 132.785 ;
        RECT 54.505 132.175 58.025 132.355 ;
        RECT 54.110 131.805 55.770 132.005 ;
        RECT 56.090 131.805 57.455 132.005 ;
        RECT 57.625 131.635 58.025 132.175 ;
        RECT 59.115 132.060 59.665 132.445 ;
        RECT 59.835 131.890 60.005 132.615 ;
        RECT 52.905 130.445 53.235 131.165 ;
        RECT 53.425 130.615 53.885 131.165 ;
        RECT 54.060 131.415 56.095 131.625 ;
        RECT 54.060 130.615 54.335 131.415 ;
        RECT 54.505 130.445 54.835 131.245 ;
        RECT 55.005 130.615 55.175 131.415 ;
        RECT 55.345 130.445 55.595 131.245 ;
        RECT 55.765 130.785 56.095 131.415 ;
        RECT 56.265 131.335 58.025 131.635 ;
        RECT 59.115 131.820 60.005 131.890 ;
        RECT 60.175 132.290 60.395 132.775 ;
        RECT 60.565 132.455 60.815 132.995 ;
        RECT 60.985 132.345 61.245 132.825 ;
        RECT 60.175 131.865 60.505 132.290 ;
        RECT 59.115 131.795 60.010 131.820 ;
        RECT 59.115 131.780 60.020 131.795 ;
        RECT 59.115 131.765 60.025 131.780 ;
        RECT 59.115 131.760 60.035 131.765 ;
        RECT 59.115 131.750 60.040 131.760 ;
        RECT 59.115 131.740 60.045 131.750 ;
        RECT 59.115 131.735 60.055 131.740 ;
        RECT 59.115 131.725 60.065 131.735 ;
        RECT 59.115 131.720 60.075 131.725 ;
        RECT 56.265 130.955 56.435 131.335 ;
        RECT 56.605 130.785 56.935 131.145 ;
        RECT 57.105 130.955 57.275 131.335 ;
        RECT 59.115 131.270 59.375 131.720 ;
        RECT 59.740 131.715 60.075 131.720 ;
        RECT 59.740 131.710 60.090 131.715 ;
        RECT 59.740 131.700 60.105 131.710 ;
        RECT 59.740 131.695 60.130 131.700 ;
        RECT 60.675 131.695 60.905 132.090 ;
        RECT 59.740 131.690 60.905 131.695 ;
        RECT 59.770 131.655 60.905 131.690 ;
        RECT 59.805 131.630 60.905 131.655 ;
        RECT 59.835 131.600 60.905 131.630 ;
        RECT 59.855 131.570 60.905 131.600 ;
        RECT 59.875 131.540 60.905 131.570 ;
        RECT 59.945 131.530 60.905 131.540 ;
        RECT 59.970 131.520 60.905 131.530 ;
        RECT 59.990 131.505 60.905 131.520 ;
        RECT 60.010 131.490 60.905 131.505 ;
        RECT 60.015 131.480 60.800 131.490 ;
        RECT 60.030 131.445 60.800 131.480 ;
        RECT 57.445 130.785 57.860 131.165 ;
        RECT 59.545 131.125 59.875 131.370 ;
        RECT 60.045 131.195 60.800 131.445 ;
        RECT 61.075 131.315 61.245 132.345 ;
        RECT 59.545 131.100 59.730 131.125 ;
        RECT 55.765 130.615 57.860 130.785 ;
        RECT 59.115 131.000 59.730 131.100 ;
        RECT 59.115 130.445 59.720 131.000 ;
        RECT 59.895 130.615 60.375 130.955 ;
        RECT 60.545 130.445 60.800 130.990 ;
        RECT 60.970 130.615 61.245 131.315 ;
        RECT 61.415 132.255 61.800 132.825 ;
        RECT 61.970 132.535 62.295 132.995 ;
        RECT 62.815 132.365 63.095 132.825 ;
        RECT 61.415 131.585 61.695 132.255 ;
        RECT 61.970 132.195 63.095 132.365 ;
        RECT 61.970 132.085 62.420 132.195 ;
        RECT 61.865 131.755 62.420 132.085 ;
        RECT 63.285 132.025 63.685 132.825 ;
        RECT 64.085 132.535 64.355 132.995 ;
        RECT 64.525 132.365 64.810 132.825 ;
        RECT 61.415 130.615 61.800 131.585 ;
        RECT 61.970 131.295 62.420 131.755 ;
        RECT 62.590 131.465 63.685 132.025 ;
        RECT 61.970 131.075 63.095 131.295 ;
        RECT 61.970 130.445 62.295 130.905 ;
        RECT 62.815 130.615 63.095 131.075 ;
        RECT 63.285 130.615 63.685 131.465 ;
        RECT 63.855 132.195 64.810 132.365 ;
        RECT 65.145 132.340 65.475 132.775 ;
        RECT 65.645 132.385 65.815 132.995 ;
        RECT 65.095 132.255 65.475 132.340 ;
        RECT 65.985 132.255 66.315 132.780 ;
        RECT 66.575 132.465 66.785 132.995 ;
        RECT 67.060 132.545 67.845 132.715 ;
        RECT 68.015 132.545 68.420 132.715 ;
        RECT 65.095 132.215 65.320 132.255 ;
        RECT 63.855 131.295 64.065 132.195 ;
        RECT 64.235 131.465 64.925 132.025 ;
        RECT 65.095 131.635 65.265 132.215 ;
        RECT 65.985 132.085 66.185 132.255 ;
        RECT 67.060 132.085 67.230 132.545 ;
        RECT 65.435 131.755 66.185 132.085 ;
        RECT 66.355 131.755 67.230 132.085 ;
        RECT 65.095 131.585 65.310 131.635 ;
        RECT 65.095 131.505 65.485 131.585 ;
        RECT 63.855 131.075 64.810 131.295 ;
        RECT 64.085 130.445 64.355 130.905 ;
        RECT 64.525 130.615 64.810 131.075 ;
        RECT 65.155 130.660 65.485 131.505 ;
        RECT 65.995 131.550 66.185 131.755 ;
        RECT 65.655 130.445 65.825 131.455 ;
        RECT 65.995 131.175 66.890 131.550 ;
        RECT 65.995 130.615 66.335 131.175 ;
        RECT 66.565 130.445 66.880 130.945 ;
        RECT 67.060 130.915 67.230 131.755 ;
        RECT 67.400 132.045 67.865 132.375 ;
        RECT 68.250 132.315 68.420 132.545 ;
        RECT 68.600 132.495 68.970 132.995 ;
        RECT 69.290 132.545 69.965 132.715 ;
        RECT 70.160 132.545 70.495 132.715 ;
        RECT 67.400 131.085 67.720 132.045 ;
        RECT 68.250 132.015 69.080 132.315 ;
        RECT 67.890 131.115 68.080 131.835 ;
        RECT 68.250 130.945 68.420 132.015 ;
        RECT 68.880 131.985 69.080 132.015 ;
        RECT 68.590 131.765 68.760 131.835 ;
        RECT 69.290 131.765 69.460 132.545 ;
        RECT 70.325 132.405 70.495 132.545 ;
        RECT 70.665 132.535 70.915 132.995 ;
        RECT 68.590 131.595 69.460 131.765 ;
        RECT 69.630 132.125 70.155 132.345 ;
        RECT 70.325 132.275 70.550 132.405 ;
        RECT 68.590 131.505 69.100 131.595 ;
        RECT 67.060 130.745 67.945 130.915 ;
        RECT 68.170 130.615 68.420 130.945 ;
        RECT 68.590 130.445 68.760 131.245 ;
        RECT 68.930 130.890 69.100 131.505 ;
        RECT 69.630 131.425 69.800 132.125 ;
        RECT 69.270 131.060 69.800 131.425 ;
        RECT 69.970 131.360 70.210 131.955 ;
        RECT 70.380 131.170 70.550 132.275 ;
        RECT 70.720 131.415 71.000 132.365 ;
        RECT 70.245 131.040 70.550 131.170 ;
        RECT 68.930 130.720 70.035 130.890 ;
        RECT 70.245 130.615 70.495 131.040 ;
        RECT 70.665 130.445 70.930 130.905 ;
        RECT 71.170 130.615 71.355 132.735 ;
        RECT 71.525 132.615 71.855 132.995 ;
        RECT 72.025 132.445 72.195 132.735 ;
        RECT 71.530 132.275 72.195 132.445 ;
        RECT 72.455 132.320 72.715 132.825 ;
        RECT 72.895 132.615 73.225 132.995 ;
        RECT 73.405 132.445 73.575 132.825 ;
        RECT 71.530 131.285 71.760 132.275 ;
        RECT 71.930 131.455 72.280 132.105 ;
        RECT 72.455 131.520 72.625 132.320 ;
        RECT 72.910 132.275 73.575 132.445 ;
        RECT 72.910 132.020 73.080 132.275 ;
        RECT 74.295 132.270 74.585 132.995 ;
        RECT 74.845 132.445 75.015 132.735 ;
        RECT 75.185 132.615 75.515 132.995 ;
        RECT 74.845 132.275 75.510 132.445 ;
        RECT 72.795 131.690 73.080 132.020 ;
        RECT 73.315 131.725 73.645 132.095 ;
        RECT 72.910 131.545 73.080 131.690 ;
        RECT 71.530 131.115 72.195 131.285 ;
        RECT 71.525 130.445 71.855 130.945 ;
        RECT 72.025 130.615 72.195 131.115 ;
        RECT 72.455 130.615 72.725 131.520 ;
        RECT 72.910 131.375 73.575 131.545 ;
        RECT 72.895 130.445 73.225 131.205 ;
        RECT 73.405 130.615 73.575 131.375 ;
        RECT 74.295 130.445 74.585 131.610 ;
        RECT 74.760 131.455 75.110 132.105 ;
        RECT 75.280 131.285 75.510 132.275 ;
        RECT 74.845 131.115 75.510 131.285 ;
        RECT 74.845 130.615 75.015 131.115 ;
        RECT 75.185 130.445 75.515 130.945 ;
        RECT 75.685 130.615 75.870 132.735 ;
        RECT 76.125 132.535 76.375 132.995 ;
        RECT 76.545 132.545 76.880 132.715 ;
        RECT 77.075 132.545 77.750 132.715 ;
        RECT 76.545 132.405 76.715 132.545 ;
        RECT 76.040 131.415 76.320 132.365 ;
        RECT 76.490 132.275 76.715 132.405 ;
        RECT 76.490 131.170 76.660 132.275 ;
        RECT 76.885 132.125 77.410 132.345 ;
        RECT 76.830 131.360 77.070 131.955 ;
        RECT 77.240 131.425 77.410 132.125 ;
        RECT 77.580 131.765 77.750 132.545 ;
        RECT 78.070 132.495 78.440 132.995 ;
        RECT 78.620 132.545 79.025 132.715 ;
        RECT 79.195 132.545 79.980 132.715 ;
        RECT 78.620 132.315 78.790 132.545 ;
        RECT 77.960 132.015 78.790 132.315 ;
        RECT 79.175 132.045 79.640 132.375 ;
        RECT 77.960 131.985 78.160 132.015 ;
        RECT 78.280 131.765 78.450 131.835 ;
        RECT 77.580 131.595 78.450 131.765 ;
        RECT 77.940 131.505 78.450 131.595 ;
        RECT 76.490 131.040 76.795 131.170 ;
        RECT 77.240 131.060 77.770 131.425 ;
        RECT 76.110 130.445 76.375 130.905 ;
        RECT 76.545 130.615 76.795 131.040 ;
        RECT 77.940 130.890 78.110 131.505 ;
        RECT 77.005 130.720 78.110 130.890 ;
        RECT 78.280 130.445 78.450 131.245 ;
        RECT 78.620 130.945 78.790 132.015 ;
        RECT 78.960 131.115 79.150 131.835 ;
        RECT 79.320 131.085 79.640 132.045 ;
        RECT 79.810 132.085 79.980 132.545 ;
        RECT 80.255 132.465 80.465 132.995 ;
        RECT 80.725 132.255 81.055 132.780 ;
        RECT 81.225 132.385 81.395 132.995 ;
        RECT 81.565 132.340 81.895 132.775 ;
        RECT 82.205 132.445 82.375 132.735 ;
        RECT 82.545 132.615 82.875 132.995 ;
        RECT 81.565 132.255 81.945 132.340 ;
        RECT 82.205 132.275 82.870 132.445 ;
        RECT 80.855 132.085 81.055 132.255 ;
        RECT 81.720 132.215 81.945 132.255 ;
        RECT 79.810 131.755 80.685 132.085 ;
        RECT 80.855 131.755 81.605 132.085 ;
        RECT 78.620 130.615 78.870 130.945 ;
        RECT 79.810 130.915 79.980 131.755 ;
        RECT 80.855 131.550 81.045 131.755 ;
        RECT 81.775 131.635 81.945 132.215 ;
        RECT 81.730 131.585 81.945 131.635 ;
        RECT 80.150 131.175 81.045 131.550 ;
        RECT 81.555 131.505 81.945 131.585 ;
        RECT 79.095 130.745 79.980 130.915 ;
        RECT 80.160 130.445 80.475 130.945 ;
        RECT 80.705 130.615 81.045 131.175 ;
        RECT 81.215 130.445 81.385 131.455 ;
        RECT 81.555 130.660 81.885 131.505 ;
        RECT 82.120 131.455 82.470 132.105 ;
        RECT 82.640 131.285 82.870 132.275 ;
        RECT 82.205 131.115 82.870 131.285 ;
        RECT 82.205 130.615 82.375 131.115 ;
        RECT 82.545 130.445 82.875 130.945 ;
        RECT 83.045 130.615 83.230 132.735 ;
        RECT 83.485 132.535 83.735 132.995 ;
        RECT 83.905 132.545 84.240 132.715 ;
        RECT 84.435 132.545 85.110 132.715 ;
        RECT 83.905 132.405 84.075 132.545 ;
        RECT 83.400 131.415 83.680 132.365 ;
        RECT 83.850 132.275 84.075 132.405 ;
        RECT 83.850 131.170 84.020 132.275 ;
        RECT 84.245 132.125 84.770 132.345 ;
        RECT 84.190 131.360 84.430 131.955 ;
        RECT 84.600 131.425 84.770 132.125 ;
        RECT 84.940 131.765 85.110 132.545 ;
        RECT 85.430 132.495 85.800 132.995 ;
        RECT 85.980 132.545 86.385 132.715 ;
        RECT 86.555 132.545 87.340 132.715 ;
        RECT 85.980 132.315 86.150 132.545 ;
        RECT 85.320 132.015 86.150 132.315 ;
        RECT 86.535 132.045 87.000 132.375 ;
        RECT 85.320 131.985 85.520 132.015 ;
        RECT 85.640 131.765 85.810 131.835 ;
        RECT 84.940 131.595 85.810 131.765 ;
        RECT 85.300 131.505 85.810 131.595 ;
        RECT 83.850 131.040 84.155 131.170 ;
        RECT 84.600 131.060 85.130 131.425 ;
        RECT 83.470 130.445 83.735 130.905 ;
        RECT 83.905 130.615 84.155 131.040 ;
        RECT 85.300 130.890 85.470 131.505 ;
        RECT 84.365 130.720 85.470 130.890 ;
        RECT 85.640 130.445 85.810 131.245 ;
        RECT 85.980 130.945 86.150 132.015 ;
        RECT 86.320 131.115 86.510 131.835 ;
        RECT 86.680 131.085 87.000 132.045 ;
        RECT 87.170 132.085 87.340 132.545 ;
        RECT 87.615 132.465 87.825 132.995 ;
        RECT 88.085 132.255 88.415 132.780 ;
        RECT 88.585 132.385 88.755 132.995 ;
        RECT 88.925 132.340 89.255 132.775 ;
        RECT 88.925 132.255 89.305 132.340 ;
        RECT 88.215 132.085 88.415 132.255 ;
        RECT 89.080 132.215 89.305 132.255 ;
        RECT 87.170 131.755 88.045 132.085 ;
        RECT 88.215 131.755 88.965 132.085 ;
        RECT 85.980 130.615 86.230 130.945 ;
        RECT 87.170 130.915 87.340 131.755 ;
        RECT 88.215 131.550 88.405 131.755 ;
        RECT 89.135 131.635 89.305 132.215 ;
        RECT 89.090 131.585 89.305 131.635 ;
        RECT 87.510 131.175 88.405 131.550 ;
        RECT 88.915 131.505 89.305 131.585 ;
        RECT 89.480 132.255 89.735 132.825 ;
        RECT 89.905 132.595 90.235 132.995 ;
        RECT 90.660 132.460 91.190 132.825 ;
        RECT 90.660 132.425 90.835 132.460 ;
        RECT 89.905 132.255 90.835 132.425 ;
        RECT 89.480 131.585 89.650 132.255 ;
        RECT 89.905 132.085 90.075 132.255 ;
        RECT 89.820 131.755 90.075 132.085 ;
        RECT 90.300 131.755 90.495 132.085 ;
        RECT 86.455 130.745 87.340 130.915 ;
        RECT 87.520 130.445 87.835 130.945 ;
        RECT 88.065 130.615 88.405 131.175 ;
        RECT 88.575 130.445 88.745 131.455 ;
        RECT 88.915 130.660 89.245 131.505 ;
        RECT 89.480 130.615 89.815 131.585 ;
        RECT 89.985 130.445 90.155 131.585 ;
        RECT 90.325 130.785 90.495 131.755 ;
        RECT 90.665 131.125 90.835 132.255 ;
        RECT 91.005 131.465 91.175 132.265 ;
        RECT 91.380 131.975 91.655 132.825 ;
        RECT 91.375 131.805 91.655 131.975 ;
        RECT 91.380 131.665 91.655 131.805 ;
        RECT 91.825 131.465 92.015 132.825 ;
        RECT 92.195 132.460 92.705 132.995 ;
        RECT 92.925 132.185 93.170 132.790 ;
        RECT 94.080 132.255 94.335 132.825 ;
        RECT 94.505 132.595 94.835 132.995 ;
        RECT 95.260 132.460 95.790 132.825 ;
        RECT 95.260 132.425 95.435 132.460 ;
        RECT 94.505 132.255 95.435 132.425 ;
        RECT 92.215 132.015 93.445 132.185 ;
        RECT 91.005 131.295 92.015 131.465 ;
        RECT 92.185 131.450 92.935 131.640 ;
        RECT 90.665 130.955 91.790 131.125 ;
        RECT 92.185 130.785 92.355 131.450 ;
        RECT 93.105 131.205 93.445 132.015 ;
        RECT 90.325 130.615 92.355 130.785 ;
        RECT 92.525 130.445 92.695 131.205 ;
        RECT 92.930 130.795 93.445 131.205 ;
        RECT 94.080 131.585 94.250 132.255 ;
        RECT 94.505 132.085 94.675 132.255 ;
        RECT 94.420 131.755 94.675 132.085 ;
        RECT 94.900 131.755 95.095 132.085 ;
        RECT 94.080 130.615 94.415 131.585 ;
        RECT 94.585 130.445 94.755 131.585 ;
        RECT 94.925 130.785 95.095 131.755 ;
        RECT 95.265 131.125 95.435 132.255 ;
        RECT 95.605 131.465 95.775 132.265 ;
        RECT 95.980 131.975 96.255 132.825 ;
        RECT 95.975 131.805 96.255 131.975 ;
        RECT 95.980 131.665 96.255 131.805 ;
        RECT 96.425 131.465 96.615 132.825 ;
        RECT 96.795 132.460 97.305 132.995 ;
        RECT 97.525 132.185 97.770 132.790 ;
        RECT 98.675 132.195 98.985 132.995 ;
        RECT 99.190 132.195 99.885 132.825 ;
        RECT 100.055 132.270 100.345 132.995 ;
        RECT 100.565 132.340 100.895 132.775 ;
        RECT 101.065 132.385 101.235 132.995 ;
        RECT 100.515 132.255 100.895 132.340 ;
        RECT 101.405 132.255 101.735 132.780 ;
        RECT 101.995 132.465 102.205 132.995 ;
        RECT 102.480 132.545 103.265 132.715 ;
        RECT 103.435 132.545 103.840 132.715 ;
        RECT 100.515 132.215 100.740 132.255 ;
        RECT 96.815 132.015 98.045 132.185 ;
        RECT 99.190 132.145 99.365 132.195 ;
        RECT 95.605 131.295 96.615 131.465 ;
        RECT 96.785 131.450 97.535 131.640 ;
        RECT 95.265 130.955 96.390 131.125 ;
        RECT 96.785 130.785 96.955 131.450 ;
        RECT 97.705 131.205 98.045 132.015 ;
        RECT 98.685 131.755 99.020 132.025 ;
        RECT 99.190 131.595 99.360 132.145 ;
        RECT 99.530 131.755 99.865 132.005 ;
        RECT 100.515 131.635 100.685 132.215 ;
        RECT 101.405 132.085 101.605 132.255 ;
        RECT 102.480 132.085 102.650 132.545 ;
        RECT 100.855 131.755 101.605 132.085 ;
        RECT 101.775 131.755 102.650 132.085 ;
        RECT 94.925 130.615 96.955 130.785 ;
        RECT 97.125 130.445 97.295 131.205 ;
        RECT 97.530 130.795 98.045 131.205 ;
        RECT 98.675 130.445 98.955 131.585 ;
        RECT 99.125 130.615 99.455 131.595 ;
        RECT 99.625 130.445 99.885 131.585 ;
        RECT 100.055 130.445 100.345 131.610 ;
        RECT 100.515 131.585 100.730 131.635 ;
        RECT 100.515 131.505 100.905 131.585 ;
        RECT 100.575 130.660 100.905 131.505 ;
        RECT 101.415 131.550 101.605 131.755 ;
        RECT 101.075 130.445 101.245 131.455 ;
        RECT 101.415 131.175 102.310 131.550 ;
        RECT 101.415 130.615 101.755 131.175 ;
        RECT 101.985 130.445 102.300 130.945 ;
        RECT 102.480 130.915 102.650 131.755 ;
        RECT 102.820 132.045 103.285 132.375 ;
        RECT 103.670 132.315 103.840 132.545 ;
        RECT 104.020 132.495 104.390 132.995 ;
        RECT 104.710 132.545 105.385 132.715 ;
        RECT 105.580 132.545 105.915 132.715 ;
        RECT 102.820 131.085 103.140 132.045 ;
        RECT 103.670 132.015 104.500 132.315 ;
        RECT 103.310 131.115 103.500 131.835 ;
        RECT 103.670 130.945 103.840 132.015 ;
        RECT 104.300 131.985 104.500 132.015 ;
        RECT 104.010 131.765 104.180 131.835 ;
        RECT 104.710 131.765 104.880 132.545 ;
        RECT 105.745 132.405 105.915 132.545 ;
        RECT 106.085 132.535 106.335 132.995 ;
        RECT 104.010 131.595 104.880 131.765 ;
        RECT 105.050 132.125 105.575 132.345 ;
        RECT 105.745 132.275 105.970 132.405 ;
        RECT 104.010 131.505 104.520 131.595 ;
        RECT 102.480 130.745 103.365 130.915 ;
        RECT 103.590 130.615 103.840 130.945 ;
        RECT 104.010 130.445 104.180 131.245 ;
        RECT 104.350 130.890 104.520 131.505 ;
        RECT 105.050 131.425 105.220 132.125 ;
        RECT 104.690 131.060 105.220 131.425 ;
        RECT 105.390 131.360 105.630 131.955 ;
        RECT 105.800 131.170 105.970 132.275 ;
        RECT 106.140 131.415 106.420 132.365 ;
        RECT 105.665 131.040 105.970 131.170 ;
        RECT 104.350 130.720 105.455 130.890 ;
        RECT 105.665 130.615 105.915 131.040 ;
        RECT 106.085 130.445 106.350 130.905 ;
        RECT 106.590 130.615 106.775 132.735 ;
        RECT 106.945 132.615 107.275 132.995 ;
        RECT 107.445 132.445 107.615 132.735 ;
        RECT 106.950 132.275 107.615 132.445 ;
        RECT 107.965 132.445 108.135 132.735 ;
        RECT 108.305 132.615 108.635 132.995 ;
        RECT 107.965 132.275 108.630 132.445 ;
        RECT 106.950 131.285 107.180 132.275 ;
        RECT 107.350 131.455 107.700 132.105 ;
        RECT 107.880 131.455 108.230 132.105 ;
        RECT 108.400 131.285 108.630 132.275 ;
        RECT 106.950 131.115 107.615 131.285 ;
        RECT 106.945 130.445 107.275 130.945 ;
        RECT 107.445 130.615 107.615 131.115 ;
        RECT 107.965 131.115 108.630 131.285 ;
        RECT 107.965 130.615 108.135 131.115 ;
        RECT 108.305 130.445 108.635 130.945 ;
        RECT 108.805 130.615 108.990 132.735 ;
        RECT 109.245 132.535 109.495 132.995 ;
        RECT 109.665 132.545 110.000 132.715 ;
        RECT 110.195 132.545 110.870 132.715 ;
        RECT 109.665 132.405 109.835 132.545 ;
        RECT 109.160 131.415 109.440 132.365 ;
        RECT 109.610 132.275 109.835 132.405 ;
        RECT 109.610 131.170 109.780 132.275 ;
        RECT 110.005 132.125 110.530 132.345 ;
        RECT 109.950 131.360 110.190 131.955 ;
        RECT 110.360 131.425 110.530 132.125 ;
        RECT 110.700 131.765 110.870 132.545 ;
        RECT 111.190 132.495 111.560 132.995 ;
        RECT 111.740 132.545 112.145 132.715 ;
        RECT 112.315 132.545 113.100 132.715 ;
        RECT 111.740 132.315 111.910 132.545 ;
        RECT 111.080 132.015 111.910 132.315 ;
        RECT 112.295 132.045 112.760 132.375 ;
        RECT 111.080 131.985 111.280 132.015 ;
        RECT 111.400 131.765 111.570 131.835 ;
        RECT 110.700 131.595 111.570 131.765 ;
        RECT 111.060 131.505 111.570 131.595 ;
        RECT 109.610 131.040 109.915 131.170 ;
        RECT 110.360 131.060 110.890 131.425 ;
        RECT 109.230 130.445 109.495 130.905 ;
        RECT 109.665 130.615 109.915 131.040 ;
        RECT 111.060 130.890 111.230 131.505 ;
        RECT 110.125 130.720 111.230 130.890 ;
        RECT 111.400 130.445 111.570 131.245 ;
        RECT 111.740 130.945 111.910 132.015 ;
        RECT 112.080 131.115 112.270 131.835 ;
        RECT 112.440 131.085 112.760 132.045 ;
        RECT 112.930 132.085 113.100 132.545 ;
        RECT 113.375 132.465 113.585 132.995 ;
        RECT 113.845 132.255 114.175 132.780 ;
        RECT 114.345 132.385 114.515 132.995 ;
        RECT 114.685 132.340 115.015 132.775 ;
        RECT 115.265 132.605 119.025 132.825 ;
        RECT 114.685 132.255 115.065 132.340 ;
        RECT 113.975 132.085 114.175 132.255 ;
        RECT 114.840 132.215 115.065 132.255 ;
        RECT 112.930 131.755 113.805 132.085 ;
        RECT 113.975 131.755 114.725 132.085 ;
        RECT 111.740 130.615 111.990 130.945 ;
        RECT 112.930 130.915 113.100 131.755 ;
        RECT 113.975 131.550 114.165 131.755 ;
        RECT 114.895 131.635 115.065 132.215 ;
        RECT 114.850 131.585 115.065 131.635 ;
        RECT 113.270 131.175 114.165 131.550 ;
        RECT 114.675 131.505 115.065 131.585 ;
        RECT 115.235 132.260 118.555 132.435 ;
        RECT 112.215 130.745 113.100 130.915 ;
        RECT 113.280 130.445 113.595 130.945 ;
        RECT 113.825 130.615 114.165 131.175 ;
        RECT 114.335 130.445 114.505 131.455 ;
        RECT 114.675 130.660 115.005 131.505 ;
        RECT 115.235 131.295 115.405 132.260 ;
        RECT 115.575 131.635 115.795 132.085 ;
        RECT 116.050 131.805 117.400 132.005 ;
        RECT 117.570 131.635 118.215 132.085 ;
        RECT 115.575 131.465 118.215 131.635 ;
        RECT 118.385 131.635 118.555 132.260 ;
        RECT 118.725 132.345 119.025 132.605 ;
        RECT 119.195 132.525 119.365 132.995 ;
        RECT 119.535 132.355 119.865 132.825 ;
        RECT 120.035 132.525 120.205 132.995 ;
        RECT 120.375 132.355 120.705 132.825 ;
        RECT 120.875 132.525 121.045 132.995 ;
        RECT 119.535 132.345 120.705 132.355 ;
        RECT 121.215 132.355 121.545 132.825 ;
        RECT 121.715 132.525 121.885 132.995 ;
        RECT 122.055 132.355 122.385 132.825 ;
        RECT 121.215 132.345 122.385 132.355 ;
        RECT 118.725 132.175 122.385 132.345 ;
        RECT 123.055 132.495 123.355 132.825 ;
        RECT 123.525 132.515 123.800 132.995 ;
        RECT 118.905 131.835 119.235 132.005 ;
        RECT 118.935 131.635 119.235 131.835 ;
        RECT 119.415 131.805 120.825 132.005 ;
        RECT 121.095 131.805 122.425 132.005 ;
        RECT 121.095 131.635 121.360 131.805 ;
        RECT 118.385 131.465 118.765 131.635 ;
        RECT 118.935 131.465 121.445 131.635 ;
        RECT 118.595 131.295 118.765 131.465 ;
        RECT 121.675 131.295 121.925 131.635 ;
        RECT 115.235 131.125 117.255 131.295 ;
        RECT 116.165 130.955 116.415 131.125 ;
        RECT 117.005 130.955 117.255 131.125 ;
        RECT 117.425 131.125 118.425 131.295 ;
        RECT 118.595 131.125 120.665 131.295 ;
        RECT 115.295 130.445 115.575 130.955 ;
        RECT 115.745 130.785 115.995 130.945 ;
        RECT 116.585 130.785 116.835 130.955 ;
        RECT 117.425 130.785 117.675 131.125 ;
        RECT 118.255 130.955 118.425 131.125 ;
        RECT 119.575 130.955 119.825 131.125 ;
        RECT 120.415 130.955 120.665 131.125 ;
        RECT 120.835 131.125 121.925 131.295 ;
        RECT 115.745 130.615 117.675 130.785 ;
        RECT 117.845 130.445 118.085 130.955 ;
        RECT 118.255 130.615 118.555 130.955 ;
        RECT 118.725 130.445 118.945 130.955 ;
        RECT 119.115 130.785 119.405 130.955 ;
        RECT 119.995 130.785 120.245 130.955 ;
        RECT 120.835 130.785 121.085 131.125 ;
        RECT 119.115 130.615 121.085 130.785 ;
        RECT 121.255 130.445 121.505 130.955 ;
        RECT 121.675 130.615 121.925 131.125 ;
        RECT 122.095 130.445 122.345 131.635 ;
        RECT 123.055 131.585 123.225 132.495 ;
        RECT 123.980 132.345 124.275 132.735 ;
        RECT 124.445 132.515 124.700 132.995 ;
        RECT 124.875 132.345 125.135 132.735 ;
        RECT 125.305 132.515 125.585 132.995 ;
        RECT 123.395 131.755 123.745 132.325 ;
        RECT 123.980 132.175 125.630 132.345 ;
        RECT 125.815 132.270 126.105 132.995 ;
        RECT 126.390 132.365 126.675 132.825 ;
        RECT 126.845 132.535 127.115 132.995 ;
        RECT 126.390 132.195 127.345 132.365 ;
        RECT 123.915 131.835 125.055 132.005 ;
        RECT 123.915 131.585 124.085 131.835 ;
        RECT 125.225 131.665 125.630 132.175 ;
        RECT 123.055 131.415 124.085 131.585 ;
        RECT 124.875 131.495 125.630 131.665 ;
        RECT 123.055 130.615 123.365 131.415 ;
        RECT 124.875 131.245 125.135 131.495 ;
        RECT 123.535 130.445 123.845 131.245 ;
        RECT 124.015 131.075 125.135 131.245 ;
        RECT 124.015 130.615 124.275 131.075 ;
        RECT 124.445 130.445 124.700 130.905 ;
        RECT 124.875 130.615 125.135 131.075 ;
        RECT 125.305 130.445 125.590 131.315 ;
        RECT 125.815 130.445 126.105 131.610 ;
        RECT 126.275 131.465 126.965 132.025 ;
        RECT 127.135 131.295 127.345 132.195 ;
        RECT 126.390 131.075 127.345 131.295 ;
        RECT 127.515 132.025 127.915 132.825 ;
        RECT 128.105 132.365 128.385 132.825 ;
        RECT 128.905 132.535 129.230 132.995 ;
        RECT 128.105 132.195 129.230 132.365 ;
        RECT 129.400 132.255 129.785 132.825 ;
        RECT 128.780 132.085 129.230 132.195 ;
        RECT 127.515 131.465 128.610 132.025 ;
        RECT 128.780 131.755 129.335 132.085 ;
        RECT 126.390 130.615 126.675 131.075 ;
        RECT 126.845 130.445 127.115 130.905 ;
        RECT 127.515 130.615 127.915 131.465 ;
        RECT 128.780 131.295 129.230 131.755 ;
        RECT 129.505 131.585 129.785 132.255 ;
        RECT 130.415 132.195 130.725 132.995 ;
        RECT 130.930 132.195 131.625 132.825 ;
        RECT 131.795 132.355 132.135 132.760 ;
        RECT 132.305 132.525 132.475 132.995 ;
        RECT 132.645 132.355 132.895 132.760 ;
        RECT 130.930 132.145 131.105 132.195 ;
        RECT 131.795 132.175 132.895 132.355 ;
        RECT 133.065 132.390 133.315 132.760 ;
        RECT 133.485 132.515 133.930 132.685 ;
        RECT 134.100 132.655 134.320 132.700 ;
        RECT 130.425 131.755 130.760 132.025 ;
        RECT 130.930 131.595 131.100 132.145 ;
        RECT 133.065 132.005 133.235 132.390 ;
        RECT 131.270 131.755 131.605 132.005 ;
        RECT 128.105 131.075 129.230 131.295 ;
        RECT 128.105 130.615 128.385 131.075 ;
        RECT 128.905 130.445 129.230 130.905 ;
        RECT 129.400 130.615 129.785 131.585 ;
        RECT 130.415 130.445 130.695 131.585 ;
        RECT 130.865 130.615 131.195 131.595 ;
        RECT 131.365 130.445 131.625 131.585 ;
        RECT 131.795 131.435 132.140 132.005 ;
        RECT 132.310 131.755 132.870 132.005 ;
        RECT 133.040 131.835 133.235 132.005 ;
        RECT 131.795 130.445 132.140 131.265 ;
        RECT 132.310 130.655 132.485 131.755 ;
        RECT 133.040 131.585 133.210 131.835 ;
        RECT 133.485 131.725 133.655 132.515 ;
        RECT 134.100 132.485 134.325 132.655 ;
        RECT 134.100 132.345 134.320 132.485 ;
        RECT 133.825 132.175 134.320 132.345 ;
        RECT 134.600 132.330 134.770 132.995 ;
        RECT 134.965 132.255 135.305 132.825 ;
        RECT 133.825 131.980 134.000 132.175 ;
        RECT 134.170 131.805 134.620 132.005 ;
        RECT 132.655 131.195 133.210 131.585 ;
        RECT 133.380 131.585 133.655 131.725 ;
        RECT 134.790 131.635 134.960 132.085 ;
        RECT 133.380 131.365 134.395 131.585 ;
        RECT 134.565 131.465 134.960 131.635 ;
        RECT 134.565 131.195 134.735 131.465 ;
        RECT 135.130 131.285 135.305 132.255 ;
        RECT 132.655 131.025 134.735 131.195 ;
        RECT 132.655 130.790 132.985 131.025 ;
        RECT 133.275 130.445 133.675 130.845 ;
        RECT 134.545 130.445 134.875 130.845 ;
        RECT 135.045 130.615 135.305 131.285 ;
        RECT 135.475 132.235 136.185 132.825 ;
        RECT 136.695 132.465 137.025 132.825 ;
        RECT 137.225 132.635 137.555 132.995 ;
        RECT 137.725 132.465 138.055 132.825 ;
        RECT 136.695 132.255 138.055 132.465 ;
        RECT 138.435 132.365 138.765 132.725 ;
        RECT 139.385 132.535 139.635 132.995 ;
        RECT 139.805 132.535 140.365 132.825 ;
        RECT 135.475 131.265 135.680 132.235 ;
        RECT 138.435 132.175 139.825 132.365 ;
        RECT 139.655 132.085 139.825 132.175 ;
        RECT 135.850 131.465 136.180 132.005 ;
        RECT 136.355 131.755 136.850 132.085 ;
        RECT 137.170 131.755 137.545 132.085 ;
        RECT 137.755 131.755 138.065 132.085 ;
        RECT 138.250 131.755 138.925 132.005 ;
        RECT 139.145 131.755 139.485 132.005 ;
        RECT 139.655 131.755 139.945 132.085 ;
        RECT 136.355 131.465 136.680 131.755 ;
        RECT 136.875 131.265 137.205 131.485 ;
        RECT 135.475 131.035 137.205 131.265 ;
        RECT 135.475 130.615 136.175 131.035 ;
        RECT 136.375 130.445 136.705 130.805 ;
        RECT 136.875 130.635 137.205 131.035 ;
        RECT 137.375 130.830 137.545 131.755 ;
        RECT 137.725 130.445 138.055 131.505 ;
        RECT 138.250 131.395 138.515 131.755 ;
        RECT 139.655 131.505 139.825 131.755 ;
        RECT 138.885 131.335 139.825 131.505 ;
        RECT 138.435 130.445 138.715 131.115 ;
        RECT 138.885 130.785 139.185 131.335 ;
        RECT 140.115 131.165 140.365 132.535 ;
        RECT 140.535 132.245 141.745 132.995 ;
        RECT 142.080 132.485 142.320 132.995 ;
        RECT 142.500 132.485 142.780 132.815 ;
        RECT 143.010 132.485 143.225 132.995 ;
        RECT 140.535 131.705 141.055 132.245 ;
        RECT 141.225 131.535 141.745 132.075 ;
        RECT 141.975 131.755 142.330 132.315 ;
        RECT 142.500 131.585 142.670 132.485 ;
        RECT 142.840 131.755 143.105 132.315 ;
        RECT 143.395 132.255 144.010 132.825 ;
        RECT 143.355 131.585 143.525 132.085 ;
        RECT 139.385 130.445 139.715 131.165 ;
        RECT 139.905 130.615 140.365 131.165 ;
        RECT 140.535 130.445 141.745 131.535 ;
        RECT 142.100 131.415 143.525 131.585 ;
        RECT 142.100 131.240 142.490 131.415 ;
        RECT 142.975 130.445 143.305 131.245 ;
        RECT 143.695 131.235 144.010 132.255 ;
        RECT 144.215 132.225 146.805 132.995 ;
        RECT 147.065 132.445 147.235 132.825 ;
        RECT 147.415 132.615 147.745 132.995 ;
        RECT 147.065 132.275 147.730 132.445 ;
        RECT 147.925 132.320 148.185 132.825 ;
        RECT 144.215 131.705 145.425 132.225 ;
        RECT 145.595 131.535 146.805 132.055 ;
        RECT 146.995 131.725 147.325 132.095 ;
        RECT 147.560 132.020 147.730 132.275 ;
        RECT 147.560 131.690 147.845 132.020 ;
        RECT 147.560 131.545 147.730 131.690 ;
        RECT 143.475 130.615 144.010 131.235 ;
        RECT 144.215 130.445 146.805 131.535 ;
        RECT 147.065 131.375 147.730 131.545 ;
        RECT 148.015 131.520 148.185 132.320 ;
        RECT 148.355 132.225 150.945 132.995 ;
        RECT 151.575 132.270 151.865 132.995 ;
        RECT 152.035 132.225 155.545 132.995 ;
        RECT 155.715 132.245 156.925 132.995 ;
        RECT 148.355 131.705 149.565 132.225 ;
        RECT 149.735 131.535 150.945 132.055 ;
        RECT 152.035 131.705 153.685 132.225 ;
        RECT 147.065 130.615 147.235 131.375 ;
        RECT 147.415 130.445 147.745 131.205 ;
        RECT 147.915 130.615 148.185 131.520 ;
        RECT 148.355 130.445 150.945 131.535 ;
        RECT 151.575 130.445 151.865 131.610 ;
        RECT 153.855 131.535 155.545 132.055 ;
        RECT 152.035 130.445 155.545 131.535 ;
        RECT 155.715 131.535 156.235 132.075 ;
        RECT 156.405 131.705 156.925 132.245 ;
        RECT 155.715 130.445 156.925 131.535 ;
        RECT 22.690 130.275 157.010 130.445 ;
        RECT 22.775 129.185 23.985 130.275 ;
        RECT 22.775 128.475 23.295 129.015 ;
        RECT 23.465 128.645 23.985 129.185 ;
        RECT 24.615 129.135 25.000 130.105 ;
        RECT 25.170 129.815 25.495 130.275 ;
        RECT 26.015 129.645 26.295 130.105 ;
        RECT 25.170 129.425 26.295 129.645 ;
        RECT 22.775 127.725 23.985 128.475 ;
        RECT 24.615 128.465 24.895 129.135 ;
        RECT 25.170 128.965 25.620 129.425 ;
        RECT 26.485 129.255 26.885 130.105 ;
        RECT 27.285 129.815 27.555 130.275 ;
        RECT 27.725 129.645 28.010 130.105 ;
        RECT 25.065 128.635 25.620 128.965 ;
        RECT 25.790 128.695 26.885 129.255 ;
        RECT 25.170 128.525 25.620 128.635 ;
        RECT 24.615 127.895 25.000 128.465 ;
        RECT 25.170 128.355 26.295 128.525 ;
        RECT 25.170 127.725 25.495 128.185 ;
        RECT 26.015 127.895 26.295 128.355 ;
        RECT 26.485 127.895 26.885 128.695 ;
        RECT 27.055 129.425 28.010 129.645 ;
        RECT 28.385 129.605 28.555 130.105 ;
        RECT 28.725 129.775 29.055 130.275 ;
        RECT 28.385 129.435 29.050 129.605 ;
        RECT 27.055 128.525 27.265 129.425 ;
        RECT 27.435 128.695 28.125 129.255 ;
        RECT 28.300 128.615 28.650 129.265 ;
        RECT 27.055 128.355 28.010 128.525 ;
        RECT 28.820 128.445 29.050 129.435 ;
        RECT 27.285 127.725 27.555 128.185 ;
        RECT 27.725 127.895 28.010 128.355 ;
        RECT 28.385 128.275 29.050 128.445 ;
        RECT 28.385 127.985 28.555 128.275 ;
        RECT 28.725 127.725 29.055 128.105 ;
        RECT 29.225 127.985 29.410 130.105 ;
        RECT 29.650 129.815 29.915 130.275 ;
        RECT 30.085 129.680 30.335 130.105 ;
        RECT 30.545 129.830 31.650 130.000 ;
        RECT 30.030 129.550 30.335 129.680 ;
        RECT 29.580 128.355 29.860 129.305 ;
        RECT 30.030 128.445 30.200 129.550 ;
        RECT 30.370 128.765 30.610 129.360 ;
        RECT 30.780 129.295 31.310 129.660 ;
        RECT 30.780 128.595 30.950 129.295 ;
        RECT 31.480 129.215 31.650 129.830 ;
        RECT 31.820 129.475 31.990 130.275 ;
        RECT 32.160 129.775 32.410 130.105 ;
        RECT 32.635 129.805 33.520 129.975 ;
        RECT 31.480 129.125 31.990 129.215 ;
        RECT 30.030 128.315 30.255 128.445 ;
        RECT 30.425 128.375 30.950 128.595 ;
        RECT 31.120 128.955 31.990 129.125 ;
        RECT 29.665 127.725 29.915 128.185 ;
        RECT 30.085 128.175 30.255 128.315 ;
        RECT 31.120 128.175 31.290 128.955 ;
        RECT 31.820 128.885 31.990 128.955 ;
        RECT 31.500 128.705 31.700 128.735 ;
        RECT 32.160 128.705 32.330 129.775 ;
        RECT 32.500 128.885 32.690 129.605 ;
        RECT 31.500 128.405 32.330 128.705 ;
        RECT 32.860 128.675 33.180 129.635 ;
        RECT 30.085 128.005 30.420 128.175 ;
        RECT 30.615 128.005 31.290 128.175 ;
        RECT 31.610 127.725 31.980 128.225 ;
        RECT 32.160 128.175 32.330 128.405 ;
        RECT 32.715 128.345 33.180 128.675 ;
        RECT 33.350 128.965 33.520 129.805 ;
        RECT 33.700 129.775 34.015 130.275 ;
        RECT 34.245 129.545 34.585 130.105 ;
        RECT 33.690 129.170 34.585 129.545 ;
        RECT 34.755 129.265 34.925 130.275 ;
        RECT 34.395 128.965 34.585 129.170 ;
        RECT 35.095 129.215 35.425 130.060 ;
        RECT 35.095 129.135 35.485 129.215 ;
        RECT 35.270 129.085 35.485 129.135 ;
        RECT 35.655 129.110 35.945 130.275 ;
        RECT 36.320 129.305 36.650 130.105 ;
        RECT 36.820 129.475 37.150 130.275 ;
        RECT 37.450 129.305 37.780 130.105 ;
        RECT 38.425 129.475 38.675 130.275 ;
        RECT 36.320 129.135 38.755 129.305 ;
        RECT 38.945 129.135 39.115 130.275 ;
        RECT 39.285 129.135 39.625 130.105 ;
        RECT 40.265 129.465 40.560 130.275 ;
        RECT 33.350 128.635 34.225 128.965 ;
        RECT 34.395 128.635 35.145 128.965 ;
        RECT 33.350 128.175 33.520 128.635 ;
        RECT 34.395 128.465 34.595 128.635 ;
        RECT 35.315 128.505 35.485 129.085 ;
        RECT 36.115 128.715 36.465 128.965 ;
        RECT 36.650 128.505 36.820 129.135 ;
        RECT 36.990 128.715 37.320 128.915 ;
        RECT 37.490 128.715 37.820 128.915 ;
        RECT 37.990 128.715 38.410 128.915 ;
        RECT 38.585 128.885 38.755 129.135 ;
        RECT 38.585 128.715 39.280 128.885 ;
        RECT 35.260 128.465 35.485 128.505 ;
        RECT 32.160 128.005 32.565 128.175 ;
        RECT 32.735 128.005 33.520 128.175 ;
        RECT 33.795 127.725 34.005 128.255 ;
        RECT 34.265 127.940 34.595 128.465 ;
        RECT 35.105 128.380 35.485 128.465 ;
        RECT 34.765 127.725 34.935 128.335 ;
        RECT 35.105 127.945 35.435 128.380 ;
        RECT 35.655 127.725 35.945 128.450 ;
        RECT 36.320 127.895 36.820 128.505 ;
        RECT 37.450 128.375 38.675 128.545 ;
        RECT 39.450 128.525 39.625 129.135 ;
        RECT 40.740 128.965 40.985 130.105 ;
        RECT 41.160 129.465 41.420 130.275 ;
        RECT 42.020 130.270 48.295 130.275 ;
        RECT 41.600 128.965 41.850 130.100 ;
        RECT 42.020 129.475 42.280 130.270 ;
        RECT 42.450 129.375 42.710 130.100 ;
        RECT 42.880 129.545 43.140 130.270 ;
        RECT 43.310 129.375 43.570 130.100 ;
        RECT 43.740 129.545 44.000 130.270 ;
        RECT 44.170 129.375 44.430 130.100 ;
        RECT 44.600 129.545 44.860 130.270 ;
        RECT 45.030 129.375 45.290 130.100 ;
        RECT 45.460 129.545 45.705 130.270 ;
        RECT 45.875 129.375 46.135 130.100 ;
        RECT 46.320 129.545 46.565 130.270 ;
        RECT 46.735 129.375 46.995 130.100 ;
        RECT 47.180 129.545 47.425 130.270 ;
        RECT 47.595 129.375 47.855 130.100 ;
        RECT 48.040 129.545 48.295 130.270 ;
        RECT 42.450 129.360 47.855 129.375 ;
        RECT 48.465 129.360 48.755 130.100 ;
        RECT 48.925 129.530 49.195 130.275 ;
        RECT 49.560 129.815 49.730 130.275 ;
        RECT 49.900 129.645 50.230 130.105 ;
        RECT 49.455 129.475 50.230 129.645 ;
        RECT 50.400 129.475 50.570 130.275 ;
        RECT 51.805 129.815 52.015 130.275 ;
        RECT 52.505 129.685 53.005 130.105 ;
        RECT 42.450 129.135 49.195 129.360 ;
        RECT 37.450 127.895 37.780 128.375 ;
        RECT 37.950 127.725 38.175 128.185 ;
        RECT 38.345 127.895 38.675 128.375 ;
        RECT 38.865 127.725 39.115 128.525 ;
        RECT 39.285 127.895 39.625 128.525 ;
        RECT 40.255 128.405 40.570 128.965 ;
        RECT 40.740 128.715 47.860 128.965 ;
        RECT 40.255 127.725 40.560 128.235 ;
        RECT 40.740 127.905 40.990 128.715 ;
        RECT 41.160 127.725 41.420 128.250 ;
        RECT 41.600 127.905 41.850 128.715 ;
        RECT 48.030 128.545 49.195 129.135 ;
        RECT 42.450 128.375 49.195 128.545 ;
        RECT 49.455 128.465 49.885 129.475 ;
        RECT 51.155 129.305 51.515 129.480 ;
        RECT 50.055 129.135 51.515 129.305 ;
        RECT 50.055 128.635 50.225 129.135 ;
        RECT 42.020 127.725 42.280 128.285 ;
        RECT 42.450 127.920 42.710 128.375 ;
        RECT 42.880 127.725 43.140 128.205 ;
        RECT 43.310 127.920 43.570 128.375 ;
        RECT 43.740 127.725 44.000 128.205 ;
        RECT 44.170 127.920 44.430 128.375 ;
        RECT 44.600 127.725 44.845 128.205 ;
        RECT 45.015 127.920 45.290 128.375 ;
        RECT 45.460 127.725 45.705 128.205 ;
        RECT 45.875 127.920 46.135 128.375 ;
        RECT 46.315 127.725 46.565 128.205 ;
        RECT 46.735 127.920 46.995 128.375 ;
        RECT 47.175 127.725 47.425 128.205 ;
        RECT 47.595 127.920 47.855 128.375 ;
        RECT 48.035 127.725 48.295 128.205 ;
        RECT 48.465 127.920 48.725 128.375 ;
        RECT 49.455 128.295 50.150 128.465 ;
        RECT 50.395 128.405 50.805 128.965 ;
        RECT 48.895 127.725 49.195 128.205 ;
        RECT 49.480 127.725 49.810 128.125 ;
        RECT 49.980 128.025 50.150 128.295 ;
        RECT 50.975 128.235 51.155 129.135 ;
        RECT 51.325 128.575 51.520 128.965 ;
        RECT 51.325 128.405 51.525 128.575 ;
        RECT 51.755 128.305 51.995 129.630 ;
        RECT 52.165 129.475 53.005 129.685 ;
        RECT 52.165 128.465 52.335 129.475 ;
        RECT 52.505 129.055 52.905 129.305 ;
        RECT 53.195 129.255 53.395 130.045 ;
        RECT 53.075 129.085 53.395 129.255 ;
        RECT 53.565 129.095 53.885 130.275 ;
        RECT 54.145 129.605 54.315 130.105 ;
        RECT 54.485 129.775 54.815 130.275 ;
        RECT 54.145 129.435 54.810 129.605 ;
        RECT 52.505 128.635 52.675 129.055 ;
        RECT 53.075 128.885 53.255 129.085 ;
        RECT 52.890 128.715 53.255 128.885 ;
        RECT 53.425 128.715 53.885 128.915 ;
        RECT 54.060 128.615 54.410 129.265 ;
        RECT 52.855 128.465 53.885 128.505 ;
        RECT 52.165 128.285 52.515 128.465 ;
        RECT 52.685 128.335 53.885 128.465 ;
        RECT 54.580 128.445 54.810 129.435 ;
        RECT 50.320 127.725 50.635 128.235 ;
        RECT 50.865 127.895 51.155 128.235 ;
        RECT 51.325 127.725 51.565 128.235 ;
        RECT 52.685 128.115 53.015 128.335 ;
        RECT 51.755 127.935 53.015 128.115 ;
        RECT 53.205 127.725 53.375 128.165 ;
        RECT 53.545 127.920 53.885 128.335 ;
        RECT 54.145 128.275 54.810 128.445 ;
        RECT 54.145 127.985 54.315 128.275 ;
        RECT 54.485 127.725 54.815 128.105 ;
        RECT 54.985 127.985 55.170 130.105 ;
        RECT 55.410 129.815 55.675 130.275 ;
        RECT 55.845 129.680 56.095 130.105 ;
        RECT 56.305 129.830 57.410 130.000 ;
        RECT 55.790 129.550 56.095 129.680 ;
        RECT 55.340 128.355 55.620 129.305 ;
        RECT 55.790 128.445 55.960 129.550 ;
        RECT 56.130 128.765 56.370 129.360 ;
        RECT 56.540 129.295 57.070 129.660 ;
        RECT 56.540 128.595 56.710 129.295 ;
        RECT 57.240 129.215 57.410 129.830 ;
        RECT 57.580 129.475 57.750 130.275 ;
        RECT 57.920 129.775 58.170 130.105 ;
        RECT 58.395 129.805 59.280 129.975 ;
        RECT 57.240 129.125 57.750 129.215 ;
        RECT 55.790 128.315 56.015 128.445 ;
        RECT 56.185 128.375 56.710 128.595 ;
        RECT 56.880 128.955 57.750 129.125 ;
        RECT 55.425 127.725 55.675 128.185 ;
        RECT 55.845 128.175 56.015 128.315 ;
        RECT 56.880 128.175 57.050 128.955 ;
        RECT 57.580 128.885 57.750 128.955 ;
        RECT 57.260 128.705 57.460 128.735 ;
        RECT 57.920 128.705 58.090 129.775 ;
        RECT 58.260 128.885 58.450 129.605 ;
        RECT 57.260 128.405 58.090 128.705 ;
        RECT 58.620 128.675 58.940 129.635 ;
        RECT 55.845 128.005 56.180 128.175 ;
        RECT 56.375 128.005 57.050 128.175 ;
        RECT 57.370 127.725 57.740 128.225 ;
        RECT 57.920 128.175 58.090 128.405 ;
        RECT 58.475 128.345 58.940 128.675 ;
        RECT 59.110 128.965 59.280 129.805 ;
        RECT 59.460 129.775 59.775 130.275 ;
        RECT 60.005 129.545 60.345 130.105 ;
        RECT 59.450 129.170 60.345 129.545 ;
        RECT 60.515 129.265 60.685 130.275 ;
        RECT 60.155 128.965 60.345 129.170 ;
        RECT 60.855 129.215 61.185 130.060 ;
        RECT 60.855 129.135 61.245 129.215 ;
        RECT 61.030 129.085 61.245 129.135 ;
        RECT 61.415 129.110 61.705 130.275 ;
        RECT 59.110 128.635 59.985 128.965 ;
        RECT 60.155 128.635 60.905 128.965 ;
        RECT 59.110 128.175 59.280 128.635 ;
        RECT 60.155 128.465 60.355 128.635 ;
        RECT 61.075 128.505 61.245 129.085 ;
        RECT 61.020 128.465 61.245 128.505 ;
        RECT 57.920 128.005 58.325 128.175 ;
        RECT 58.495 128.005 59.280 128.175 ;
        RECT 59.555 127.725 59.765 128.255 ;
        RECT 60.025 127.940 60.355 128.465 ;
        RECT 60.865 128.380 61.245 128.465 ;
        RECT 60.525 127.725 60.695 128.335 ;
        RECT 60.865 127.945 61.195 128.380 ;
        RECT 61.415 127.725 61.705 128.450 ;
        RECT 62.345 127.905 62.605 130.095 ;
        RECT 62.775 129.545 63.115 130.275 ;
        RECT 63.295 129.365 63.565 130.095 ;
        RECT 62.795 129.145 63.565 129.365 ;
        RECT 63.745 129.385 63.975 130.095 ;
        RECT 64.145 129.565 64.475 130.275 ;
        RECT 64.645 129.385 64.905 130.095 ;
        RECT 65.185 129.605 65.355 130.105 ;
        RECT 65.525 129.775 65.855 130.275 ;
        RECT 65.185 129.435 65.850 129.605 ;
        RECT 63.745 129.145 64.905 129.385 ;
        RECT 62.795 128.475 63.085 129.145 ;
        RECT 63.265 128.655 63.730 128.965 ;
        RECT 63.910 128.655 64.435 128.965 ;
        RECT 62.795 128.275 64.025 128.475 ;
        RECT 62.865 127.725 63.535 128.095 ;
        RECT 63.715 127.905 64.025 128.275 ;
        RECT 64.205 128.015 64.435 128.655 ;
        RECT 64.615 128.635 64.915 128.965 ;
        RECT 65.100 128.615 65.450 129.265 ;
        RECT 64.615 127.725 64.905 128.455 ;
        RECT 65.620 128.445 65.850 129.435 ;
        RECT 65.185 128.275 65.850 128.445 ;
        RECT 65.185 127.985 65.355 128.275 ;
        RECT 65.525 127.725 65.855 128.105 ;
        RECT 66.025 127.985 66.210 130.105 ;
        RECT 66.450 129.815 66.715 130.275 ;
        RECT 66.885 129.680 67.135 130.105 ;
        RECT 67.345 129.830 68.450 130.000 ;
        RECT 66.830 129.550 67.135 129.680 ;
        RECT 66.380 128.355 66.660 129.305 ;
        RECT 66.830 128.445 67.000 129.550 ;
        RECT 67.170 128.765 67.410 129.360 ;
        RECT 67.580 129.295 68.110 129.660 ;
        RECT 67.580 128.595 67.750 129.295 ;
        RECT 68.280 129.215 68.450 129.830 ;
        RECT 68.620 129.475 68.790 130.275 ;
        RECT 68.960 129.775 69.210 130.105 ;
        RECT 69.435 129.805 70.320 129.975 ;
        RECT 68.280 129.125 68.790 129.215 ;
        RECT 66.830 128.315 67.055 128.445 ;
        RECT 67.225 128.375 67.750 128.595 ;
        RECT 67.920 128.955 68.790 129.125 ;
        RECT 66.465 127.725 66.715 128.185 ;
        RECT 66.885 128.175 67.055 128.315 ;
        RECT 67.920 128.175 68.090 128.955 ;
        RECT 68.620 128.885 68.790 128.955 ;
        RECT 68.300 128.705 68.500 128.735 ;
        RECT 68.960 128.705 69.130 129.775 ;
        RECT 69.300 128.885 69.490 129.605 ;
        RECT 68.300 128.405 69.130 128.705 ;
        RECT 69.660 128.675 69.980 129.635 ;
        RECT 66.885 128.005 67.220 128.175 ;
        RECT 67.415 128.005 68.090 128.175 ;
        RECT 68.410 127.725 68.780 128.225 ;
        RECT 68.960 128.175 69.130 128.405 ;
        RECT 69.515 128.345 69.980 128.675 ;
        RECT 70.150 128.965 70.320 129.805 ;
        RECT 70.500 129.775 70.815 130.275 ;
        RECT 71.045 129.545 71.385 130.105 ;
        RECT 70.490 129.170 71.385 129.545 ;
        RECT 71.555 129.265 71.725 130.275 ;
        RECT 71.195 128.965 71.385 129.170 ;
        RECT 71.895 129.215 72.225 130.060 ;
        RECT 71.895 129.135 72.285 129.215 ;
        RECT 72.070 129.085 72.285 129.135 ;
        RECT 70.150 128.635 71.025 128.965 ;
        RECT 71.195 128.635 71.945 128.965 ;
        RECT 70.150 128.175 70.320 128.635 ;
        RECT 71.195 128.465 71.395 128.635 ;
        RECT 72.115 128.505 72.285 129.085 ;
        RECT 72.060 128.465 72.285 128.505 ;
        RECT 68.960 128.005 69.365 128.175 ;
        RECT 69.535 128.005 70.320 128.175 ;
        RECT 70.595 127.725 70.805 128.255 ;
        RECT 71.065 127.940 71.395 128.465 ;
        RECT 71.905 128.380 72.285 128.465 ;
        RECT 72.455 129.135 72.840 130.105 ;
        RECT 73.010 129.815 73.335 130.275 ;
        RECT 73.855 129.645 74.135 130.105 ;
        RECT 73.010 129.425 74.135 129.645 ;
        RECT 72.455 128.465 72.735 129.135 ;
        RECT 73.010 128.965 73.460 129.425 ;
        RECT 74.325 129.255 74.725 130.105 ;
        RECT 75.125 129.815 75.395 130.275 ;
        RECT 75.565 129.645 75.850 130.105 ;
        RECT 72.905 128.635 73.460 128.965 ;
        RECT 73.630 128.695 74.725 129.255 ;
        RECT 73.010 128.525 73.460 128.635 ;
        RECT 71.565 127.725 71.735 128.335 ;
        RECT 71.905 127.945 72.235 128.380 ;
        RECT 72.455 127.895 72.840 128.465 ;
        RECT 73.010 128.355 74.135 128.525 ;
        RECT 73.010 127.725 73.335 128.185 ;
        RECT 73.855 127.895 74.135 128.355 ;
        RECT 74.325 127.895 74.725 128.695 ;
        RECT 74.895 129.425 75.850 129.645 ;
        RECT 74.895 128.525 75.105 129.425 ;
        RECT 75.275 128.695 75.965 129.255 ;
        RECT 76.135 129.185 77.805 130.275 ;
        RECT 74.895 128.355 75.850 128.525 ;
        RECT 75.125 127.725 75.395 128.185 ;
        RECT 75.565 127.895 75.850 128.355 ;
        RECT 76.135 128.495 76.885 129.015 ;
        RECT 77.055 128.665 77.805 129.185 ;
        RECT 78.435 129.295 78.755 130.105 ;
        RECT 78.925 129.465 79.175 130.275 ;
        RECT 79.345 129.935 80.475 130.105 ;
        RECT 79.345 129.295 79.595 129.935 ;
        RECT 78.435 129.085 79.595 129.295 ;
        RECT 78.830 128.705 79.270 128.915 ;
        RECT 79.765 128.535 80.015 129.765 ;
        RECT 80.185 129.530 80.475 129.935 ;
        RECT 80.185 129.085 80.440 129.530 ;
        RECT 80.745 129.255 80.915 130.100 ;
        RECT 81.125 129.785 81.375 130.275 ;
        RECT 81.260 129.595 81.475 129.605 ;
        RECT 81.255 129.425 81.475 129.595 ;
        RECT 80.610 129.085 80.915 129.255 ;
        RECT 80.610 128.885 80.780 129.085 ;
        RECT 81.260 128.915 81.475 129.425 ;
        RECT 81.655 129.185 83.325 130.275 ;
        RECT 80.225 128.715 80.780 128.885 ;
        RECT 80.565 128.535 80.780 128.715 ;
        RECT 80.950 128.705 81.475 128.915 ;
        RECT 76.135 127.725 77.805 128.495 ;
        RECT 78.435 127.725 78.715 128.535 ;
        RECT 78.885 128.365 80.055 128.535 ;
        RECT 78.885 127.895 79.215 128.365 ;
        RECT 79.385 127.725 79.555 128.195 ;
        RECT 79.725 127.895 80.055 128.365 ;
        RECT 80.225 127.725 80.395 128.535 ;
        RECT 80.565 128.365 80.915 128.535 ;
        RECT 81.655 128.495 82.405 129.015 ;
        RECT 82.575 128.665 83.325 129.185 ;
        RECT 83.495 129.200 83.765 130.105 ;
        RECT 83.935 129.515 84.265 130.275 ;
        RECT 84.445 129.345 84.615 130.105 ;
        RECT 85.075 129.605 85.355 130.275 ;
        RECT 80.745 128.085 80.915 128.365 ;
        RECT 81.125 127.725 81.380 128.485 ;
        RECT 81.655 127.725 83.325 128.495 ;
        RECT 83.495 128.400 83.665 129.200 ;
        RECT 83.950 129.175 84.615 129.345 ;
        RECT 85.525 129.385 85.825 129.935 ;
        RECT 86.025 129.555 86.355 130.275 ;
        RECT 86.545 129.555 87.005 130.105 ;
        RECT 83.950 129.030 84.120 129.175 ;
        RECT 83.835 128.700 84.120 129.030 ;
        RECT 83.950 128.445 84.120 128.700 ;
        RECT 84.355 128.625 84.685 128.995 ;
        RECT 84.890 128.965 85.155 129.325 ;
        RECT 85.525 129.215 86.465 129.385 ;
        RECT 86.295 128.965 86.465 129.215 ;
        RECT 84.890 128.715 85.565 128.965 ;
        RECT 85.785 128.715 86.125 128.965 ;
        RECT 86.295 128.635 86.585 128.965 ;
        RECT 86.295 128.545 86.465 128.635 ;
        RECT 83.495 127.895 83.755 128.400 ;
        RECT 83.950 128.275 84.615 128.445 ;
        RECT 83.935 127.725 84.265 128.105 ;
        RECT 84.445 127.895 84.615 128.275 ;
        RECT 85.075 128.355 86.465 128.545 ;
        RECT 85.075 127.995 85.405 128.355 ;
        RECT 86.755 128.185 87.005 129.555 ;
        RECT 87.175 129.110 87.465 130.275 ;
        RECT 87.635 129.305 87.945 130.105 ;
        RECT 88.115 129.475 88.425 130.275 ;
        RECT 88.595 129.645 88.855 130.105 ;
        RECT 89.025 129.815 89.280 130.275 ;
        RECT 89.455 129.645 89.715 130.105 ;
        RECT 88.595 129.475 89.715 129.645 ;
        RECT 87.635 129.135 88.665 129.305 ;
        RECT 86.025 127.725 86.275 128.185 ;
        RECT 86.445 127.895 87.005 128.185 ;
        RECT 87.175 127.725 87.465 128.450 ;
        RECT 87.635 128.225 87.805 129.135 ;
        RECT 87.975 128.395 88.325 128.965 ;
        RECT 88.495 128.885 88.665 129.135 ;
        RECT 89.455 129.225 89.715 129.475 ;
        RECT 89.885 129.405 90.170 130.275 ;
        RECT 91.515 129.605 91.795 130.275 ;
        RECT 91.965 129.385 92.265 129.935 ;
        RECT 92.465 129.555 92.795 130.275 ;
        RECT 92.985 129.555 93.445 130.105 ;
        RECT 93.675 129.765 93.955 130.275 ;
        RECT 94.125 129.935 96.055 130.105 ;
        RECT 94.125 129.775 94.375 129.935 ;
        RECT 94.965 129.765 95.215 129.935 ;
        RECT 94.545 129.595 94.795 129.765 ;
        RECT 95.385 129.595 95.635 129.765 ;
        RECT 89.455 129.055 90.210 129.225 ;
        RECT 88.495 128.715 89.635 128.885 ;
        RECT 89.805 128.545 90.210 129.055 ;
        RECT 91.330 128.965 91.595 129.325 ;
        RECT 91.965 129.215 92.905 129.385 ;
        RECT 92.735 128.965 92.905 129.215 ;
        RECT 91.330 128.715 92.005 128.965 ;
        RECT 92.225 128.715 92.565 128.965 ;
        RECT 92.735 128.635 93.025 128.965 ;
        RECT 92.735 128.545 92.905 128.635 ;
        RECT 88.560 128.375 90.210 128.545 ;
        RECT 87.635 127.895 87.935 128.225 ;
        RECT 88.105 127.725 88.380 128.205 ;
        RECT 88.560 127.985 88.855 128.375 ;
        RECT 89.025 127.725 89.280 128.205 ;
        RECT 89.455 127.985 89.715 128.375 ;
        RECT 91.515 128.355 92.905 128.545 ;
        RECT 89.885 127.725 90.165 128.205 ;
        RECT 91.515 127.995 91.845 128.355 ;
        RECT 93.195 128.185 93.445 129.555 ;
        RECT 93.615 129.425 95.635 129.595 ;
        RECT 95.805 129.595 96.055 129.935 ;
        RECT 96.225 129.765 96.465 130.275 ;
        RECT 96.635 129.765 96.935 130.105 ;
        RECT 97.105 129.765 97.325 130.275 ;
        RECT 97.495 129.935 99.465 130.105 ;
        RECT 97.495 129.765 97.785 129.935 ;
        RECT 98.375 129.765 98.625 129.935 ;
        RECT 96.635 129.595 96.805 129.765 ;
        RECT 97.955 129.595 98.205 129.765 ;
        RECT 98.795 129.595 99.045 129.765 ;
        RECT 95.805 129.425 96.805 129.595 ;
        RECT 96.975 129.425 99.045 129.595 ;
        RECT 99.215 129.595 99.465 129.935 ;
        RECT 99.635 129.765 99.885 130.275 ;
        RECT 100.055 129.595 100.305 130.105 ;
        RECT 99.215 129.425 100.305 129.595 ;
        RECT 93.615 128.460 93.785 129.425 ;
        RECT 96.975 129.255 97.145 129.425 ;
        RECT 93.955 129.085 96.595 129.255 ;
        RECT 93.955 128.635 94.175 129.085 ;
        RECT 94.430 128.715 95.780 128.915 ;
        RECT 95.950 128.635 96.595 129.085 ;
        RECT 96.765 129.085 97.145 129.255 ;
        RECT 97.315 129.085 99.825 129.255 ;
        RECT 100.055 129.085 100.305 129.425 ;
        RECT 100.475 129.085 100.725 130.275 ;
        RECT 100.975 129.840 106.320 130.275 ;
        RECT 96.765 128.460 96.935 129.085 ;
        RECT 97.315 128.885 97.615 129.085 ;
        RECT 99.475 128.915 99.740 129.085 ;
        RECT 97.285 128.715 97.615 128.885 ;
        RECT 97.795 128.715 99.205 128.915 ;
        RECT 99.475 128.715 100.805 128.915 ;
        RECT 93.615 128.285 96.935 128.460 ;
        RECT 97.105 128.375 100.765 128.545 ;
        RECT 92.465 127.725 92.715 128.185 ;
        RECT 92.885 127.895 93.445 128.185 ;
        RECT 97.105 128.115 97.405 128.375 ;
        RECT 97.915 128.365 99.085 128.375 ;
        RECT 93.645 127.895 97.405 128.115 ;
        RECT 97.575 127.725 97.745 128.195 ;
        RECT 97.915 127.895 98.245 128.365 ;
        RECT 98.415 127.725 98.585 128.195 ;
        RECT 98.755 127.895 99.085 128.365 ;
        RECT 99.595 128.365 100.765 128.375 ;
        RECT 99.255 127.725 99.425 128.195 ;
        RECT 99.595 127.895 99.925 128.365 ;
        RECT 100.095 127.725 100.265 128.195 ;
        RECT 100.435 127.895 100.765 128.365 ;
        RECT 102.560 128.270 102.900 129.100 ;
        RECT 104.380 128.590 104.730 129.840 ;
        RECT 106.495 129.185 107.705 130.275 ;
        RECT 106.495 128.475 107.015 129.015 ;
        RECT 107.185 128.645 107.705 129.185 ;
        RECT 107.880 129.135 108.215 130.105 ;
        RECT 108.385 129.135 108.555 130.275 ;
        RECT 108.725 129.935 110.755 130.105 ;
        RECT 100.975 127.725 106.320 128.270 ;
        RECT 106.495 127.725 107.705 128.475 ;
        RECT 107.880 128.465 108.050 129.135 ;
        RECT 108.725 128.965 108.895 129.935 ;
        RECT 108.220 128.635 108.475 128.965 ;
        RECT 108.700 128.635 108.895 128.965 ;
        RECT 109.065 129.595 110.190 129.765 ;
        RECT 108.305 128.465 108.475 128.635 ;
        RECT 109.065 128.465 109.235 129.595 ;
        RECT 107.880 127.895 108.135 128.465 ;
        RECT 108.305 128.295 109.235 128.465 ;
        RECT 109.405 129.255 110.415 129.425 ;
        RECT 109.405 128.455 109.575 129.255 ;
        RECT 109.780 128.915 110.055 129.055 ;
        RECT 109.775 128.745 110.055 128.915 ;
        RECT 109.060 128.260 109.235 128.295 ;
        RECT 108.305 127.725 108.635 128.125 ;
        RECT 109.060 127.895 109.590 128.260 ;
        RECT 109.780 127.895 110.055 128.745 ;
        RECT 110.225 127.895 110.415 129.255 ;
        RECT 110.585 129.270 110.755 129.935 ;
        RECT 110.925 129.515 111.095 130.275 ;
        RECT 111.330 129.515 111.845 129.925 ;
        RECT 110.585 129.080 111.335 129.270 ;
        RECT 111.505 128.705 111.845 129.515 ;
        RECT 112.935 129.110 113.225 130.275 ;
        RECT 113.395 129.185 115.065 130.275 ;
        RECT 115.290 129.405 115.575 130.275 ;
        RECT 115.745 129.645 116.005 130.105 ;
        RECT 116.180 129.815 116.435 130.275 ;
        RECT 116.605 129.645 116.865 130.105 ;
        RECT 115.745 129.475 116.865 129.645 ;
        RECT 117.035 129.475 117.345 130.275 ;
        RECT 115.745 129.225 116.005 129.475 ;
        RECT 117.515 129.305 117.825 130.105 ;
        RECT 110.615 128.535 111.845 128.705 ;
        RECT 110.595 127.725 111.105 128.260 ;
        RECT 111.325 127.930 111.570 128.535 ;
        RECT 113.395 128.495 114.145 129.015 ;
        RECT 114.315 128.665 115.065 129.185 ;
        RECT 115.250 129.055 116.005 129.225 ;
        RECT 116.795 129.135 117.825 129.305 ;
        RECT 118.055 129.215 118.385 130.060 ;
        RECT 118.555 129.265 118.725 130.275 ;
        RECT 118.895 129.545 119.235 130.105 ;
        RECT 119.465 129.775 119.780 130.275 ;
        RECT 119.960 129.805 120.845 129.975 ;
        RECT 115.250 128.545 115.655 129.055 ;
        RECT 116.795 128.885 116.965 129.135 ;
        RECT 115.825 128.715 116.965 128.885 ;
        RECT 112.935 127.725 113.225 128.450 ;
        RECT 113.395 127.725 115.065 128.495 ;
        RECT 115.250 128.375 116.900 128.545 ;
        RECT 117.135 128.395 117.485 128.965 ;
        RECT 115.295 127.725 115.575 128.205 ;
        RECT 115.745 127.985 116.005 128.375 ;
        RECT 116.180 127.725 116.435 128.205 ;
        RECT 116.605 127.985 116.900 128.375 ;
        RECT 117.655 128.225 117.825 129.135 ;
        RECT 117.995 129.135 118.385 129.215 ;
        RECT 118.895 129.170 119.790 129.545 ;
        RECT 117.995 129.085 118.210 129.135 ;
        RECT 117.995 128.505 118.165 129.085 ;
        RECT 118.895 128.965 119.085 129.170 ;
        RECT 119.960 128.965 120.130 129.805 ;
        RECT 121.070 129.775 121.320 130.105 ;
        RECT 118.335 128.635 119.085 128.965 ;
        RECT 119.255 128.635 120.130 128.965 ;
        RECT 117.995 128.465 118.220 128.505 ;
        RECT 118.885 128.465 119.085 128.635 ;
        RECT 117.995 128.380 118.375 128.465 ;
        RECT 117.080 127.725 117.355 128.205 ;
        RECT 117.525 127.895 117.825 128.225 ;
        RECT 118.045 127.945 118.375 128.380 ;
        RECT 118.545 127.725 118.715 128.335 ;
        RECT 118.885 127.940 119.215 128.465 ;
        RECT 119.475 127.725 119.685 128.255 ;
        RECT 119.960 128.175 120.130 128.635 ;
        RECT 120.300 128.675 120.620 129.635 ;
        RECT 120.790 128.885 120.980 129.605 ;
        RECT 121.150 128.705 121.320 129.775 ;
        RECT 121.490 129.475 121.660 130.275 ;
        RECT 121.830 129.830 122.935 130.000 ;
        RECT 121.830 129.215 122.000 129.830 ;
        RECT 123.145 129.680 123.395 130.105 ;
        RECT 123.565 129.815 123.830 130.275 ;
        RECT 122.170 129.295 122.700 129.660 ;
        RECT 123.145 129.550 123.450 129.680 ;
        RECT 121.490 129.125 122.000 129.215 ;
        RECT 121.490 128.955 122.360 129.125 ;
        RECT 121.490 128.885 121.660 128.955 ;
        RECT 121.780 128.705 121.980 128.735 ;
        RECT 120.300 128.345 120.765 128.675 ;
        RECT 121.150 128.405 121.980 128.705 ;
        RECT 121.150 128.175 121.320 128.405 ;
        RECT 119.960 128.005 120.745 128.175 ;
        RECT 120.915 128.005 121.320 128.175 ;
        RECT 121.500 127.725 121.870 128.225 ;
        RECT 122.190 128.175 122.360 128.955 ;
        RECT 122.530 128.595 122.700 129.295 ;
        RECT 122.870 128.765 123.110 129.360 ;
        RECT 122.530 128.375 123.055 128.595 ;
        RECT 123.280 128.445 123.450 129.550 ;
        RECT 123.225 128.315 123.450 128.445 ;
        RECT 123.620 128.355 123.900 129.305 ;
        RECT 123.225 128.175 123.395 128.315 ;
        RECT 122.190 128.005 122.865 128.175 ;
        RECT 123.060 128.005 123.395 128.175 ;
        RECT 123.565 127.725 123.815 128.185 ;
        RECT 124.070 127.985 124.255 130.105 ;
        RECT 124.425 129.775 124.755 130.275 ;
        RECT 124.925 129.605 125.095 130.105 ;
        RECT 126.295 129.765 126.595 130.275 ;
        RECT 126.765 129.765 127.145 129.935 ;
        RECT 127.725 129.765 128.355 130.275 ;
        RECT 124.430 129.435 125.095 129.605 ;
        RECT 126.765 129.595 126.935 129.765 ;
        RECT 128.525 129.595 128.855 130.105 ;
        RECT 129.025 129.765 129.325 130.275 ;
        RECT 124.430 128.445 124.660 129.435 ;
        RECT 126.275 129.395 126.935 129.595 ;
        RECT 127.105 129.425 129.325 129.595 ;
        RECT 124.830 128.615 125.180 129.265 ;
        RECT 126.275 128.465 126.445 129.395 ;
        RECT 127.105 129.225 127.275 129.425 ;
        RECT 126.615 129.055 127.275 129.225 ;
        RECT 127.445 129.085 128.985 129.255 ;
        RECT 126.615 128.635 126.785 129.055 ;
        RECT 127.445 128.885 127.615 129.085 ;
        RECT 127.015 128.715 127.615 128.885 ;
        RECT 127.785 128.715 128.480 128.915 ;
        RECT 128.740 128.635 128.985 129.085 ;
        RECT 127.105 128.465 128.015 128.545 ;
        RECT 124.430 128.275 125.095 128.445 ;
        RECT 124.425 127.725 124.755 128.105 ;
        RECT 124.925 127.985 125.095 128.275 ;
        RECT 126.275 127.985 126.595 128.465 ;
        RECT 126.765 128.375 128.015 128.465 ;
        RECT 126.765 128.295 127.275 128.375 ;
        RECT 126.765 127.895 126.995 128.295 ;
        RECT 127.165 127.725 127.515 128.115 ;
        RECT 127.685 127.895 128.015 128.375 ;
        RECT 128.185 127.725 128.355 128.545 ;
        RECT 129.155 128.465 129.325 129.425 ;
        RECT 129.495 129.185 131.165 130.275 ;
        RECT 128.860 127.920 129.325 128.465 ;
        RECT 129.495 128.495 130.245 129.015 ;
        RECT 130.415 128.665 131.165 129.185 ;
        RECT 131.335 129.135 131.720 130.105 ;
        RECT 131.890 129.815 132.215 130.275 ;
        RECT 132.735 129.645 133.015 130.105 ;
        RECT 131.890 129.425 133.015 129.645 ;
        RECT 129.495 127.725 131.165 128.495 ;
        RECT 131.335 128.465 131.615 129.135 ;
        RECT 131.890 128.965 132.340 129.425 ;
        RECT 133.205 129.255 133.605 130.105 ;
        RECT 134.005 129.815 134.275 130.275 ;
        RECT 134.445 129.645 134.730 130.105 ;
        RECT 131.785 128.635 132.340 128.965 ;
        RECT 132.510 128.695 133.605 129.255 ;
        RECT 131.890 128.525 132.340 128.635 ;
        RECT 131.335 127.895 131.720 128.465 ;
        RECT 131.890 128.355 133.015 128.525 ;
        RECT 131.890 127.725 132.215 128.185 ;
        RECT 132.735 127.895 133.015 128.355 ;
        RECT 133.205 127.895 133.605 128.695 ;
        RECT 133.775 129.425 134.730 129.645 ;
        RECT 133.775 128.525 133.985 129.425 ;
        RECT 134.155 128.695 134.845 129.255 ;
        RECT 135.015 129.135 135.285 130.105 ;
        RECT 135.495 129.475 135.775 130.275 ;
        RECT 135.955 129.725 137.150 130.055 ;
        RECT 136.280 129.305 136.700 129.555 ;
        RECT 135.455 129.135 136.700 129.305 ;
        RECT 133.775 128.355 134.730 128.525 ;
        RECT 134.005 127.725 134.275 128.185 ;
        RECT 134.445 127.895 134.730 128.355 ;
        RECT 135.015 128.400 135.185 129.135 ;
        RECT 135.455 128.965 135.625 129.135 ;
        RECT 136.925 128.965 137.095 129.525 ;
        RECT 137.345 129.135 137.600 130.275 ;
        RECT 138.695 129.110 138.985 130.275 ;
        RECT 139.215 129.135 139.425 130.275 ;
        RECT 139.595 129.125 139.925 130.105 ;
        RECT 140.095 129.135 140.325 130.275 ;
        RECT 140.535 129.135 140.795 130.275 ;
        RECT 140.965 129.125 141.295 130.105 ;
        RECT 141.465 129.135 141.745 130.275 ;
        RECT 141.915 129.135 142.195 130.275 ;
        RECT 142.365 129.125 142.695 130.105 ;
        RECT 142.865 129.135 143.125 130.275 ;
        RECT 143.295 129.720 143.900 130.275 ;
        RECT 144.075 129.765 144.555 130.105 ;
        RECT 144.725 129.730 144.980 130.275 ;
        RECT 143.295 129.620 143.910 129.720 ;
        RECT 143.725 129.595 143.910 129.620 ;
        RECT 135.395 128.635 135.625 128.965 ;
        RECT 136.355 128.635 137.095 128.965 ;
        RECT 137.265 128.715 137.600 128.965 ;
        RECT 135.455 128.465 135.625 128.635 ;
        RECT 136.845 128.545 137.095 128.635 ;
        RECT 135.015 128.055 135.285 128.400 ;
        RECT 135.455 128.295 136.195 128.465 ;
        RECT 136.845 128.375 137.580 128.545 ;
        RECT 135.475 127.725 135.855 128.125 ;
        RECT 136.025 127.945 136.195 128.295 ;
        RECT 136.365 127.725 137.100 128.205 ;
        RECT 137.270 127.905 137.580 128.375 ;
        RECT 138.695 127.725 138.985 128.450 ;
        RECT 139.215 127.725 139.425 128.545 ;
        RECT 139.595 128.525 139.845 129.125 ;
        RECT 140.015 128.715 140.345 128.965 ;
        RECT 140.555 128.715 140.890 128.965 ;
        RECT 139.595 127.895 139.925 128.525 ;
        RECT 140.095 127.725 140.325 128.545 ;
        RECT 141.060 128.525 141.230 129.125 ;
        RECT 141.400 128.695 141.735 128.965 ;
        RECT 141.925 128.695 142.260 128.965 ;
        RECT 142.430 128.525 142.600 129.125 ;
        RECT 143.295 129.000 143.555 129.450 ;
        RECT 143.725 129.350 144.055 129.595 ;
        RECT 144.225 129.275 144.980 129.525 ;
        RECT 145.150 129.405 145.425 130.105 ;
        RECT 144.210 129.240 144.980 129.275 ;
        RECT 144.195 129.230 144.980 129.240 ;
        RECT 144.190 129.215 145.085 129.230 ;
        RECT 144.170 129.200 145.085 129.215 ;
        RECT 144.150 129.190 145.085 129.200 ;
        RECT 144.125 129.180 145.085 129.190 ;
        RECT 144.055 129.150 145.085 129.180 ;
        RECT 144.035 129.120 145.085 129.150 ;
        RECT 144.015 129.090 145.085 129.120 ;
        RECT 143.985 129.065 145.085 129.090 ;
        RECT 143.950 129.030 145.085 129.065 ;
        RECT 143.920 129.025 145.085 129.030 ;
        RECT 143.920 129.020 144.310 129.025 ;
        RECT 143.920 129.010 144.285 129.020 ;
        RECT 143.920 129.005 144.270 129.010 ;
        RECT 143.920 129.000 144.255 129.005 ;
        RECT 143.295 128.995 144.255 129.000 ;
        RECT 143.295 128.985 144.245 128.995 ;
        RECT 143.295 128.980 144.235 128.985 ;
        RECT 143.295 128.970 144.225 128.980 ;
        RECT 142.770 128.715 143.105 128.965 ;
        RECT 143.295 128.960 144.220 128.970 ;
        RECT 143.295 128.955 144.215 128.960 ;
        RECT 143.295 128.940 144.205 128.955 ;
        RECT 143.295 128.925 144.200 128.940 ;
        RECT 143.295 128.900 144.190 128.925 ;
        RECT 143.295 128.830 144.185 128.900 ;
        RECT 140.535 127.895 141.230 128.525 ;
        RECT 141.435 127.725 141.745 128.525 ;
        RECT 141.915 127.725 142.225 128.525 ;
        RECT 142.430 127.895 143.125 128.525 ;
        RECT 143.295 128.275 143.845 128.660 ;
        RECT 144.015 128.105 144.185 128.830 ;
        RECT 143.295 127.935 144.185 128.105 ;
        RECT 144.355 128.430 144.685 128.855 ;
        RECT 144.855 128.630 145.085 129.025 ;
        RECT 144.355 128.405 144.605 128.430 ;
        RECT 144.355 127.945 144.575 128.405 ;
        RECT 145.255 128.375 145.425 129.405 ;
        RECT 145.780 129.305 146.170 129.480 ;
        RECT 146.655 129.475 146.985 130.275 ;
        RECT 147.155 129.485 147.690 130.105 ;
        RECT 145.780 129.135 147.205 129.305 ;
        RECT 145.655 128.405 146.010 128.965 ;
        RECT 144.745 127.725 144.995 128.265 ;
        RECT 145.165 127.895 145.425 128.375 ;
        RECT 146.180 128.235 146.350 129.135 ;
        RECT 146.520 128.405 146.785 128.965 ;
        RECT 147.035 128.635 147.205 129.135 ;
        RECT 147.375 128.465 147.690 129.485 ;
        RECT 147.955 129.215 148.285 130.060 ;
        RECT 148.455 129.265 148.625 130.275 ;
        RECT 148.795 129.545 149.135 130.105 ;
        RECT 149.365 129.775 149.680 130.275 ;
        RECT 149.860 129.805 150.745 129.975 ;
        RECT 145.760 127.725 146.000 128.235 ;
        RECT 146.180 127.905 146.460 128.235 ;
        RECT 146.690 127.725 146.905 128.235 ;
        RECT 147.075 127.895 147.690 128.465 ;
        RECT 147.895 129.135 148.285 129.215 ;
        RECT 148.795 129.170 149.690 129.545 ;
        RECT 147.895 129.085 148.110 129.135 ;
        RECT 147.895 128.505 148.065 129.085 ;
        RECT 148.795 128.965 148.985 129.170 ;
        RECT 149.860 128.965 150.030 129.805 ;
        RECT 150.970 129.775 151.220 130.105 ;
        RECT 148.235 128.635 148.985 128.965 ;
        RECT 149.155 128.635 150.030 128.965 ;
        RECT 147.895 128.465 148.120 128.505 ;
        RECT 148.785 128.465 148.985 128.635 ;
        RECT 147.895 128.380 148.275 128.465 ;
        RECT 147.945 127.945 148.275 128.380 ;
        RECT 148.445 127.725 148.615 128.335 ;
        RECT 148.785 127.940 149.115 128.465 ;
        RECT 149.375 127.725 149.585 128.255 ;
        RECT 149.860 128.175 150.030 128.635 ;
        RECT 150.200 128.675 150.520 129.635 ;
        RECT 150.690 128.885 150.880 129.605 ;
        RECT 151.050 128.705 151.220 129.775 ;
        RECT 151.390 129.475 151.560 130.275 ;
        RECT 151.730 129.830 152.835 130.000 ;
        RECT 151.730 129.215 151.900 129.830 ;
        RECT 153.045 129.680 153.295 130.105 ;
        RECT 153.465 129.815 153.730 130.275 ;
        RECT 152.070 129.295 152.600 129.660 ;
        RECT 153.045 129.550 153.350 129.680 ;
        RECT 151.390 129.125 151.900 129.215 ;
        RECT 151.390 128.955 152.260 129.125 ;
        RECT 151.390 128.885 151.560 128.955 ;
        RECT 151.680 128.705 151.880 128.735 ;
        RECT 150.200 128.345 150.665 128.675 ;
        RECT 151.050 128.405 151.880 128.705 ;
        RECT 151.050 128.175 151.220 128.405 ;
        RECT 149.860 128.005 150.645 128.175 ;
        RECT 150.815 128.005 151.220 128.175 ;
        RECT 151.400 127.725 151.770 128.225 ;
        RECT 152.090 128.175 152.260 128.955 ;
        RECT 152.430 128.595 152.600 129.295 ;
        RECT 152.770 128.765 153.010 129.360 ;
        RECT 152.430 128.375 152.955 128.595 ;
        RECT 153.180 128.445 153.350 129.550 ;
        RECT 153.125 128.315 153.350 128.445 ;
        RECT 153.520 128.355 153.800 129.305 ;
        RECT 153.125 128.175 153.295 128.315 ;
        RECT 152.090 128.005 152.765 128.175 ;
        RECT 152.960 128.005 153.295 128.175 ;
        RECT 153.465 127.725 153.715 128.185 ;
        RECT 153.970 127.985 154.155 130.105 ;
        RECT 154.325 129.775 154.655 130.275 ;
        RECT 154.825 129.605 154.995 130.105 ;
        RECT 154.330 129.435 154.995 129.605 ;
        RECT 154.330 128.445 154.560 129.435 ;
        RECT 154.730 128.615 155.080 129.265 ;
        RECT 155.715 129.185 156.925 130.275 ;
        RECT 155.715 128.645 156.235 129.185 ;
        RECT 156.405 128.475 156.925 129.015 ;
        RECT 154.330 128.275 154.995 128.445 ;
        RECT 154.325 127.725 154.655 128.105 ;
        RECT 154.825 127.985 154.995 128.275 ;
        RECT 155.715 127.725 156.925 128.475 ;
        RECT 22.690 127.555 157.010 127.725 ;
        RECT 22.775 126.805 23.985 127.555 ;
        RECT 24.245 127.005 24.415 127.295 ;
        RECT 24.585 127.175 24.915 127.555 ;
        RECT 24.245 126.835 24.910 127.005 ;
        RECT 22.775 126.265 23.295 126.805 ;
        RECT 23.465 126.095 23.985 126.635 ;
        RECT 22.775 125.005 23.985 126.095 ;
        RECT 24.160 126.015 24.510 126.665 ;
        RECT 24.680 125.845 24.910 126.835 ;
        RECT 24.245 125.675 24.910 125.845 ;
        RECT 24.245 125.175 24.415 125.675 ;
        RECT 24.585 125.005 24.915 125.505 ;
        RECT 25.085 125.175 25.270 127.295 ;
        RECT 25.525 127.095 25.775 127.555 ;
        RECT 25.945 127.105 26.280 127.275 ;
        RECT 26.475 127.105 27.150 127.275 ;
        RECT 25.945 126.965 26.115 127.105 ;
        RECT 25.440 125.975 25.720 126.925 ;
        RECT 25.890 126.835 26.115 126.965 ;
        RECT 25.890 125.730 26.060 126.835 ;
        RECT 26.285 126.685 26.810 126.905 ;
        RECT 26.230 125.920 26.470 126.515 ;
        RECT 26.640 125.985 26.810 126.685 ;
        RECT 26.980 126.325 27.150 127.105 ;
        RECT 27.470 127.055 27.840 127.555 ;
        RECT 28.020 127.105 28.425 127.275 ;
        RECT 28.595 127.105 29.380 127.275 ;
        RECT 28.020 126.875 28.190 127.105 ;
        RECT 27.360 126.575 28.190 126.875 ;
        RECT 28.575 126.605 29.040 126.935 ;
        RECT 27.360 126.545 27.560 126.575 ;
        RECT 27.680 126.325 27.850 126.395 ;
        RECT 26.980 126.155 27.850 126.325 ;
        RECT 27.340 126.065 27.850 126.155 ;
        RECT 25.890 125.600 26.195 125.730 ;
        RECT 26.640 125.620 27.170 125.985 ;
        RECT 25.510 125.005 25.775 125.465 ;
        RECT 25.945 125.175 26.195 125.600 ;
        RECT 27.340 125.450 27.510 126.065 ;
        RECT 26.405 125.280 27.510 125.450 ;
        RECT 27.680 125.005 27.850 125.805 ;
        RECT 28.020 125.505 28.190 126.575 ;
        RECT 28.360 125.675 28.550 126.395 ;
        RECT 28.720 125.645 29.040 126.605 ;
        RECT 29.210 126.645 29.380 127.105 ;
        RECT 29.655 127.025 29.865 127.555 ;
        RECT 30.125 126.815 30.455 127.340 ;
        RECT 30.625 126.945 30.795 127.555 ;
        RECT 30.965 126.900 31.295 127.335 ;
        RECT 30.965 126.815 31.345 126.900 ;
        RECT 30.255 126.645 30.455 126.815 ;
        RECT 31.120 126.775 31.345 126.815 ;
        RECT 29.210 126.315 30.085 126.645 ;
        RECT 30.255 126.315 31.005 126.645 ;
        RECT 28.020 125.175 28.270 125.505 ;
        RECT 29.210 125.475 29.380 126.315 ;
        RECT 30.255 126.110 30.445 126.315 ;
        RECT 31.175 126.195 31.345 126.775 ;
        RECT 31.515 126.805 32.725 127.555 ;
        RECT 31.515 126.265 32.035 126.805 ;
        RECT 33.100 126.775 33.600 127.385 ;
        RECT 31.130 126.145 31.345 126.195 ;
        RECT 29.550 125.735 30.445 126.110 ;
        RECT 30.955 126.065 31.345 126.145 ;
        RECT 32.205 126.095 32.725 126.635 ;
        RECT 32.895 126.315 33.245 126.565 ;
        RECT 33.430 126.145 33.600 126.775 ;
        RECT 34.230 126.905 34.560 127.385 ;
        RECT 34.730 127.095 34.955 127.555 ;
        RECT 35.125 126.905 35.455 127.385 ;
        RECT 34.230 126.735 35.455 126.905 ;
        RECT 35.645 126.755 35.895 127.555 ;
        RECT 36.065 126.755 36.405 127.385 ;
        RECT 36.690 126.925 36.975 127.385 ;
        RECT 37.145 127.095 37.415 127.555 ;
        RECT 36.690 126.755 37.645 126.925 ;
        RECT 33.770 126.365 34.100 126.565 ;
        RECT 34.270 126.365 34.600 126.565 ;
        RECT 34.770 126.365 35.190 126.565 ;
        RECT 35.365 126.395 36.060 126.565 ;
        RECT 35.365 126.145 35.535 126.395 ;
        RECT 36.230 126.195 36.405 126.755 ;
        RECT 36.175 126.145 36.405 126.195 ;
        RECT 28.495 125.305 29.380 125.475 ;
        RECT 29.560 125.005 29.875 125.505 ;
        RECT 30.105 125.175 30.445 125.735 ;
        RECT 30.615 125.005 30.785 126.015 ;
        RECT 30.955 125.220 31.285 126.065 ;
        RECT 31.515 125.005 32.725 126.095 ;
        RECT 33.100 125.975 35.535 126.145 ;
        RECT 33.100 125.175 33.430 125.975 ;
        RECT 33.600 125.005 33.930 125.805 ;
        RECT 34.230 125.175 34.560 125.975 ;
        RECT 35.205 125.005 35.455 125.805 ;
        RECT 35.725 125.005 35.895 126.145 ;
        RECT 36.065 125.175 36.405 126.145 ;
        RECT 36.575 126.025 37.265 126.585 ;
        RECT 37.435 125.855 37.645 126.755 ;
        RECT 36.690 125.635 37.645 125.855 ;
        RECT 37.815 126.585 38.215 127.385 ;
        RECT 38.405 126.925 38.685 127.385 ;
        RECT 39.205 127.095 39.530 127.555 ;
        RECT 38.405 126.755 39.530 126.925 ;
        RECT 39.700 126.815 40.085 127.385 ;
        RECT 39.080 126.645 39.530 126.755 ;
        RECT 37.815 126.025 38.910 126.585 ;
        RECT 39.080 126.315 39.635 126.645 ;
        RECT 36.690 125.175 36.975 125.635 ;
        RECT 37.145 125.005 37.415 125.465 ;
        RECT 37.815 125.175 38.215 126.025 ;
        RECT 39.080 125.855 39.530 126.315 ;
        RECT 39.805 126.145 40.085 126.815 ;
        RECT 38.405 125.635 39.530 125.855 ;
        RECT 38.405 125.175 38.685 125.635 ;
        RECT 39.205 125.005 39.530 125.465 ;
        RECT 39.700 125.175 40.085 126.145 ;
        RECT 40.255 126.815 40.640 127.385 ;
        RECT 40.810 127.095 41.135 127.555 ;
        RECT 41.655 126.925 41.935 127.385 ;
        RECT 40.255 126.145 40.535 126.815 ;
        RECT 40.810 126.755 41.935 126.925 ;
        RECT 40.810 126.645 41.260 126.755 ;
        RECT 40.705 126.315 41.260 126.645 ;
        RECT 42.125 126.585 42.525 127.385 ;
        RECT 42.925 127.095 43.195 127.555 ;
        RECT 43.365 126.925 43.650 127.385 ;
        RECT 40.255 125.175 40.640 126.145 ;
        RECT 40.810 125.855 41.260 126.315 ;
        RECT 41.430 126.025 42.525 126.585 ;
        RECT 40.810 125.635 41.935 125.855 ;
        RECT 40.810 125.005 41.135 125.465 ;
        RECT 41.655 125.175 41.935 125.635 ;
        RECT 42.125 125.175 42.525 126.025 ;
        RECT 42.695 126.755 43.650 126.925 ;
        RECT 44.970 126.925 45.255 127.385 ;
        RECT 45.425 127.095 45.695 127.555 ;
        RECT 44.970 126.755 45.925 126.925 ;
        RECT 42.695 125.855 42.905 126.755 ;
        RECT 43.075 126.025 43.765 126.585 ;
        RECT 44.855 126.025 45.545 126.585 ;
        RECT 45.715 125.855 45.925 126.755 ;
        RECT 42.695 125.635 43.650 125.855 ;
        RECT 42.925 125.005 43.195 125.465 ;
        RECT 43.365 125.175 43.650 125.635 ;
        RECT 44.970 125.635 45.925 125.855 ;
        RECT 46.095 126.585 46.495 127.385 ;
        RECT 46.685 126.925 46.965 127.385 ;
        RECT 47.485 127.095 47.810 127.555 ;
        RECT 46.685 126.755 47.810 126.925 ;
        RECT 47.980 126.815 48.365 127.385 ;
        RECT 48.535 126.830 48.825 127.555 ;
        RECT 47.360 126.645 47.810 126.755 ;
        RECT 46.095 126.025 47.190 126.585 ;
        RECT 47.360 126.315 47.915 126.645 ;
        RECT 44.970 125.175 45.255 125.635 ;
        RECT 45.425 125.005 45.695 125.465 ;
        RECT 46.095 125.175 46.495 126.025 ;
        RECT 47.360 125.855 47.810 126.315 ;
        RECT 48.085 126.145 48.365 126.815 ;
        RECT 49.455 126.815 49.840 127.385 ;
        RECT 50.010 127.095 50.335 127.555 ;
        RECT 50.855 126.925 51.135 127.385 ;
        RECT 46.685 125.635 47.810 125.855 ;
        RECT 46.685 125.175 46.965 125.635 ;
        RECT 47.485 125.005 47.810 125.465 ;
        RECT 47.980 125.175 48.365 126.145 ;
        RECT 48.535 125.005 48.825 126.170 ;
        RECT 49.455 126.145 49.735 126.815 ;
        RECT 50.010 126.755 51.135 126.925 ;
        RECT 50.010 126.645 50.460 126.755 ;
        RECT 49.905 126.315 50.460 126.645 ;
        RECT 51.325 126.585 51.725 127.385 ;
        RECT 52.125 127.095 52.395 127.555 ;
        RECT 52.565 126.925 52.850 127.385 ;
        RECT 49.455 125.175 49.840 126.145 ;
        RECT 50.010 125.855 50.460 126.315 ;
        RECT 50.630 126.025 51.725 126.585 ;
        RECT 50.010 125.635 51.135 125.855 ;
        RECT 50.010 125.005 50.335 125.465 ;
        RECT 50.855 125.175 51.135 125.635 ;
        RECT 51.325 125.175 51.725 126.025 ;
        RECT 51.895 126.755 52.850 126.925 ;
        RECT 53.685 127.005 53.855 127.295 ;
        RECT 54.025 127.175 54.355 127.555 ;
        RECT 53.685 126.835 54.350 127.005 ;
        RECT 51.895 125.855 52.105 126.755 ;
        RECT 52.275 126.025 52.965 126.585 ;
        RECT 53.600 126.015 53.950 126.665 ;
        RECT 51.895 125.635 52.850 125.855 ;
        RECT 54.120 125.845 54.350 126.835 ;
        RECT 52.125 125.005 52.395 125.465 ;
        RECT 52.565 125.175 52.850 125.635 ;
        RECT 53.685 125.675 54.350 125.845 ;
        RECT 53.685 125.175 53.855 125.675 ;
        RECT 54.025 125.005 54.355 125.505 ;
        RECT 54.525 125.175 54.710 127.295 ;
        RECT 54.965 127.095 55.215 127.555 ;
        RECT 55.385 127.105 55.720 127.275 ;
        RECT 55.915 127.105 56.590 127.275 ;
        RECT 55.385 126.965 55.555 127.105 ;
        RECT 54.880 125.975 55.160 126.925 ;
        RECT 55.330 126.835 55.555 126.965 ;
        RECT 55.330 125.730 55.500 126.835 ;
        RECT 55.725 126.685 56.250 126.905 ;
        RECT 55.670 125.920 55.910 126.515 ;
        RECT 56.080 125.985 56.250 126.685 ;
        RECT 56.420 126.325 56.590 127.105 ;
        RECT 56.910 127.055 57.280 127.555 ;
        RECT 57.460 127.105 57.865 127.275 ;
        RECT 58.035 127.105 58.820 127.275 ;
        RECT 57.460 126.875 57.630 127.105 ;
        RECT 56.800 126.575 57.630 126.875 ;
        RECT 58.015 126.605 58.480 126.935 ;
        RECT 56.800 126.545 57.000 126.575 ;
        RECT 57.120 126.325 57.290 126.395 ;
        RECT 56.420 126.155 57.290 126.325 ;
        RECT 56.780 126.065 57.290 126.155 ;
        RECT 55.330 125.600 55.635 125.730 ;
        RECT 56.080 125.620 56.610 125.985 ;
        RECT 54.950 125.005 55.215 125.465 ;
        RECT 55.385 125.175 55.635 125.600 ;
        RECT 56.780 125.450 56.950 126.065 ;
        RECT 55.845 125.280 56.950 125.450 ;
        RECT 57.120 125.005 57.290 125.805 ;
        RECT 57.460 125.505 57.630 126.575 ;
        RECT 57.800 125.675 57.990 126.395 ;
        RECT 58.160 125.645 58.480 126.605 ;
        RECT 58.650 126.645 58.820 127.105 ;
        RECT 59.095 127.025 59.305 127.555 ;
        RECT 59.565 126.815 59.895 127.340 ;
        RECT 60.065 126.945 60.235 127.555 ;
        RECT 60.405 126.900 60.735 127.335 ;
        RECT 60.405 126.815 60.785 126.900 ;
        RECT 59.695 126.645 59.895 126.815 ;
        RECT 60.560 126.775 60.785 126.815 ;
        RECT 58.650 126.315 59.525 126.645 ;
        RECT 59.695 126.315 60.445 126.645 ;
        RECT 57.460 125.175 57.710 125.505 ;
        RECT 58.650 125.475 58.820 126.315 ;
        RECT 59.695 126.110 59.885 126.315 ;
        RECT 60.615 126.195 60.785 126.775 ;
        RECT 60.570 126.145 60.785 126.195 ;
        RECT 58.990 125.735 59.885 126.110 ;
        RECT 60.395 126.065 60.785 126.145 ;
        RECT 57.935 125.305 58.820 125.475 ;
        RECT 59.000 125.005 59.315 125.505 ;
        RECT 59.545 125.175 59.885 125.735 ;
        RECT 60.055 125.005 60.225 126.015 ;
        RECT 60.395 125.220 60.725 126.065 ;
        RECT 61.425 125.185 61.685 127.375 ;
        RECT 61.945 127.185 62.615 127.555 ;
        RECT 62.795 127.005 63.105 127.375 ;
        RECT 61.875 126.805 63.105 127.005 ;
        RECT 61.875 126.135 62.165 126.805 ;
        RECT 63.285 126.625 63.515 127.265 ;
        RECT 63.695 126.825 63.985 127.555 ;
        RECT 64.175 126.905 64.435 127.385 ;
        RECT 64.605 127.015 64.855 127.555 ;
        RECT 62.345 126.315 62.810 126.625 ;
        RECT 62.990 126.315 63.515 126.625 ;
        RECT 63.695 126.315 63.995 126.645 ;
        RECT 61.875 125.915 62.645 126.135 ;
        RECT 61.855 125.005 62.195 125.735 ;
        RECT 62.375 125.185 62.645 125.915 ;
        RECT 62.825 125.895 63.985 126.135 ;
        RECT 62.825 125.185 63.055 125.895 ;
        RECT 63.225 125.005 63.555 125.715 ;
        RECT 63.725 125.185 63.985 125.895 ;
        RECT 64.175 125.875 64.345 126.905 ;
        RECT 65.025 126.875 65.245 127.335 ;
        RECT 64.995 126.850 65.245 126.875 ;
        RECT 64.515 126.255 64.745 126.650 ;
        RECT 64.915 126.425 65.245 126.850 ;
        RECT 65.415 127.175 66.305 127.345 ;
        RECT 65.415 126.450 65.585 127.175 ;
        RECT 65.755 126.620 66.305 127.005 ;
        RECT 65.415 126.380 66.305 126.450 ;
        RECT 65.410 126.355 66.305 126.380 ;
        RECT 65.400 126.340 66.305 126.355 ;
        RECT 65.395 126.325 66.305 126.340 ;
        RECT 65.385 126.320 66.305 126.325 ;
        RECT 65.380 126.310 66.305 126.320 ;
        RECT 65.375 126.300 66.305 126.310 ;
        RECT 65.365 126.295 66.305 126.300 ;
        RECT 65.355 126.285 66.305 126.295 ;
        RECT 65.345 126.280 66.305 126.285 ;
        RECT 65.345 126.275 65.680 126.280 ;
        RECT 65.330 126.270 65.680 126.275 ;
        RECT 65.315 126.260 65.680 126.270 ;
        RECT 65.290 126.255 65.680 126.260 ;
        RECT 64.515 126.250 65.680 126.255 ;
        RECT 64.515 126.215 65.650 126.250 ;
        RECT 64.515 126.190 65.615 126.215 ;
        RECT 64.515 126.160 65.585 126.190 ;
        RECT 64.515 126.130 65.565 126.160 ;
        RECT 64.515 126.100 65.545 126.130 ;
        RECT 64.515 126.090 65.475 126.100 ;
        RECT 64.515 126.080 65.450 126.090 ;
        RECT 64.515 126.065 65.430 126.080 ;
        RECT 64.515 126.050 65.410 126.065 ;
        RECT 64.620 126.040 65.405 126.050 ;
        RECT 64.620 126.005 65.390 126.040 ;
        RECT 64.175 125.175 64.450 125.875 ;
        RECT 64.620 125.755 65.375 126.005 ;
        RECT 65.545 125.685 65.875 125.930 ;
        RECT 66.045 125.830 66.305 126.280 ;
        RECT 65.690 125.660 65.875 125.685 ;
        RECT 65.690 125.560 66.305 125.660 ;
        RECT 64.620 125.005 64.875 125.550 ;
        RECT 65.045 125.175 65.525 125.515 ;
        RECT 65.700 125.005 66.305 125.560 ;
        RECT 66.945 125.185 67.205 127.375 ;
        RECT 67.465 127.185 68.135 127.555 ;
        RECT 68.315 127.005 68.625 127.375 ;
        RECT 67.395 126.805 68.625 127.005 ;
        RECT 67.395 126.135 67.685 126.805 ;
        RECT 68.805 126.625 69.035 127.265 ;
        RECT 69.215 126.825 69.505 127.555 ;
        RECT 69.695 126.905 69.955 127.385 ;
        RECT 70.125 127.015 70.375 127.555 ;
        RECT 67.865 126.315 68.330 126.625 ;
        RECT 68.510 126.315 69.035 126.625 ;
        RECT 69.215 126.315 69.515 126.645 ;
        RECT 67.395 125.915 68.165 126.135 ;
        RECT 67.375 125.005 67.715 125.735 ;
        RECT 67.895 125.185 68.165 125.915 ;
        RECT 68.345 125.895 69.505 126.135 ;
        RECT 68.345 125.185 68.575 125.895 ;
        RECT 68.745 125.005 69.075 125.715 ;
        RECT 69.245 125.185 69.505 125.895 ;
        RECT 69.695 125.875 69.865 126.905 ;
        RECT 70.545 126.850 70.765 127.335 ;
        RECT 70.035 126.255 70.265 126.650 ;
        RECT 70.435 126.425 70.765 126.850 ;
        RECT 70.935 127.175 71.825 127.345 ;
        RECT 70.935 126.450 71.105 127.175 ;
        RECT 71.275 126.620 71.825 127.005 ;
        RECT 72.035 126.735 72.265 127.555 ;
        RECT 72.435 126.755 72.765 127.385 ;
        RECT 70.935 126.380 71.825 126.450 ;
        RECT 70.930 126.355 71.825 126.380 ;
        RECT 70.920 126.340 71.825 126.355 ;
        RECT 70.915 126.325 71.825 126.340 ;
        RECT 70.905 126.320 71.825 126.325 ;
        RECT 70.900 126.310 71.825 126.320 ;
        RECT 72.015 126.315 72.345 126.565 ;
        RECT 70.895 126.300 71.825 126.310 ;
        RECT 70.885 126.295 71.825 126.300 ;
        RECT 70.875 126.285 71.825 126.295 ;
        RECT 70.865 126.280 71.825 126.285 ;
        RECT 70.865 126.275 71.200 126.280 ;
        RECT 70.850 126.270 71.200 126.275 ;
        RECT 70.835 126.260 71.200 126.270 ;
        RECT 70.810 126.255 71.200 126.260 ;
        RECT 70.035 126.250 71.200 126.255 ;
        RECT 70.035 126.215 71.170 126.250 ;
        RECT 70.035 126.190 71.135 126.215 ;
        RECT 70.035 126.160 71.105 126.190 ;
        RECT 70.035 126.130 71.085 126.160 ;
        RECT 70.035 126.100 71.065 126.130 ;
        RECT 70.035 126.090 70.995 126.100 ;
        RECT 70.035 126.080 70.970 126.090 ;
        RECT 70.035 126.065 70.950 126.080 ;
        RECT 70.035 126.050 70.930 126.065 ;
        RECT 70.140 126.040 70.925 126.050 ;
        RECT 70.140 126.005 70.910 126.040 ;
        RECT 69.695 125.175 69.970 125.875 ;
        RECT 70.140 125.755 70.895 126.005 ;
        RECT 71.065 125.685 71.395 125.930 ;
        RECT 71.565 125.830 71.825 126.280 ;
        RECT 72.515 126.155 72.765 126.755 ;
        RECT 72.935 126.735 73.145 127.555 ;
        RECT 74.295 126.830 74.585 127.555 ;
        RECT 74.870 126.925 75.155 127.385 ;
        RECT 75.325 127.095 75.595 127.555 ;
        RECT 74.870 126.755 75.825 126.925 ;
        RECT 71.210 125.660 71.395 125.685 ;
        RECT 71.210 125.560 71.825 125.660 ;
        RECT 70.140 125.005 70.395 125.550 ;
        RECT 70.565 125.175 71.045 125.515 ;
        RECT 71.220 125.005 71.825 125.560 ;
        RECT 72.035 125.005 72.265 126.145 ;
        RECT 72.435 125.175 72.765 126.155 ;
        RECT 72.935 125.005 73.145 126.145 ;
        RECT 74.295 125.005 74.585 126.170 ;
        RECT 74.755 126.025 75.445 126.585 ;
        RECT 75.615 125.855 75.825 126.755 ;
        RECT 74.870 125.635 75.825 125.855 ;
        RECT 75.995 126.585 76.395 127.385 ;
        RECT 76.585 126.925 76.865 127.385 ;
        RECT 77.385 127.095 77.710 127.555 ;
        RECT 76.585 126.755 77.710 126.925 ;
        RECT 77.880 126.815 78.265 127.385 ;
        RECT 77.260 126.645 77.710 126.755 ;
        RECT 75.995 126.025 77.090 126.585 ;
        RECT 77.260 126.315 77.815 126.645 ;
        RECT 74.870 125.175 75.155 125.635 ;
        RECT 75.325 125.005 75.595 125.465 ;
        RECT 75.995 125.175 76.395 126.025 ;
        RECT 77.260 125.855 77.710 126.315 ;
        RECT 77.985 126.145 78.265 126.815 ;
        RECT 79.630 126.745 79.875 127.350 ;
        RECT 80.095 127.020 80.605 127.555 ;
        RECT 76.585 125.635 77.710 125.855 ;
        RECT 76.585 125.175 76.865 125.635 ;
        RECT 77.385 125.005 77.710 125.465 ;
        RECT 77.880 125.175 78.265 126.145 ;
        RECT 79.355 126.575 80.585 126.745 ;
        RECT 79.355 125.765 79.695 126.575 ;
        RECT 79.865 126.010 80.615 126.200 ;
        RECT 79.355 125.355 79.870 125.765 ;
        RECT 80.105 125.005 80.275 125.765 ;
        RECT 80.445 125.345 80.615 126.010 ;
        RECT 80.785 126.025 80.975 127.385 ;
        RECT 81.145 126.875 81.420 127.385 ;
        RECT 81.610 127.020 82.140 127.385 ;
        RECT 82.565 127.155 82.895 127.555 ;
        RECT 81.965 126.985 82.140 127.020 ;
        RECT 81.145 126.705 81.425 126.875 ;
        RECT 81.145 126.225 81.420 126.705 ;
        RECT 81.625 126.025 81.795 126.825 ;
        RECT 80.785 125.855 81.795 126.025 ;
        RECT 81.965 126.815 82.895 126.985 ;
        RECT 83.065 126.815 83.320 127.385 ;
        RECT 81.965 125.685 82.135 126.815 ;
        RECT 82.725 126.645 82.895 126.815 ;
        RECT 81.010 125.515 82.135 125.685 ;
        RECT 82.305 126.315 82.500 126.645 ;
        RECT 82.725 126.315 82.980 126.645 ;
        RECT 82.305 125.345 82.475 126.315 ;
        RECT 83.150 126.145 83.320 126.815 ;
        RECT 83.495 126.785 87.005 127.555 ;
        RECT 88.185 127.005 88.355 127.385 ;
        RECT 88.535 127.175 88.865 127.555 ;
        RECT 88.185 126.835 88.850 127.005 ;
        RECT 89.045 126.880 89.305 127.385 ;
        RECT 83.495 126.265 85.145 126.785 ;
        RECT 80.445 125.175 82.475 125.345 ;
        RECT 82.645 125.005 82.815 126.145 ;
        RECT 82.985 125.175 83.320 126.145 ;
        RECT 85.315 126.095 87.005 126.615 ;
        RECT 88.115 126.285 88.445 126.655 ;
        RECT 88.680 126.580 88.850 126.835 ;
        RECT 88.680 126.250 88.965 126.580 ;
        RECT 88.680 126.105 88.850 126.250 ;
        RECT 83.495 125.005 87.005 126.095 ;
        RECT 88.185 125.935 88.850 126.105 ;
        RECT 89.135 126.080 89.305 126.880 ;
        RECT 89.565 127.005 89.735 127.295 ;
        RECT 89.905 127.175 90.235 127.555 ;
        RECT 89.565 126.835 90.230 127.005 ;
        RECT 88.185 125.175 88.355 125.935 ;
        RECT 88.535 125.005 88.865 125.765 ;
        RECT 89.035 125.175 89.305 126.080 ;
        RECT 89.480 126.015 89.830 126.665 ;
        RECT 90.000 125.845 90.230 126.835 ;
        RECT 89.565 125.675 90.230 125.845 ;
        RECT 89.565 125.175 89.735 125.675 ;
        RECT 89.905 125.005 90.235 125.505 ;
        RECT 90.405 125.175 90.590 127.295 ;
        RECT 90.845 127.095 91.095 127.555 ;
        RECT 91.265 127.105 91.600 127.275 ;
        RECT 91.795 127.105 92.470 127.275 ;
        RECT 91.265 126.965 91.435 127.105 ;
        RECT 90.760 125.975 91.040 126.925 ;
        RECT 91.210 126.835 91.435 126.965 ;
        RECT 91.210 125.730 91.380 126.835 ;
        RECT 91.605 126.685 92.130 126.905 ;
        RECT 91.550 125.920 91.790 126.515 ;
        RECT 91.960 125.985 92.130 126.685 ;
        RECT 92.300 126.325 92.470 127.105 ;
        RECT 92.790 127.055 93.160 127.555 ;
        RECT 93.340 127.105 93.745 127.275 ;
        RECT 93.915 127.105 94.700 127.275 ;
        RECT 93.340 126.875 93.510 127.105 ;
        RECT 92.680 126.575 93.510 126.875 ;
        RECT 93.895 126.605 94.360 126.935 ;
        RECT 92.680 126.545 92.880 126.575 ;
        RECT 93.000 126.325 93.170 126.395 ;
        RECT 92.300 126.155 93.170 126.325 ;
        RECT 92.660 126.065 93.170 126.155 ;
        RECT 91.210 125.600 91.515 125.730 ;
        RECT 91.960 125.620 92.490 125.985 ;
        RECT 90.830 125.005 91.095 125.465 ;
        RECT 91.265 125.175 91.515 125.600 ;
        RECT 92.660 125.450 92.830 126.065 ;
        RECT 91.725 125.280 92.830 125.450 ;
        RECT 93.000 125.005 93.170 125.805 ;
        RECT 93.340 125.505 93.510 126.575 ;
        RECT 93.680 125.675 93.870 126.395 ;
        RECT 94.040 125.645 94.360 126.605 ;
        RECT 94.530 126.645 94.700 127.105 ;
        RECT 94.975 127.025 95.185 127.555 ;
        RECT 95.445 126.815 95.775 127.340 ;
        RECT 95.945 126.945 96.115 127.555 ;
        RECT 96.285 126.900 96.615 127.335 ;
        RECT 96.285 126.815 96.665 126.900 ;
        RECT 95.575 126.645 95.775 126.815 ;
        RECT 96.440 126.775 96.665 126.815 ;
        RECT 94.530 126.315 95.405 126.645 ;
        RECT 95.575 126.315 96.325 126.645 ;
        RECT 93.340 125.175 93.590 125.505 ;
        RECT 94.530 125.475 94.700 126.315 ;
        RECT 95.575 126.110 95.765 126.315 ;
        RECT 96.495 126.195 96.665 126.775 ;
        RECT 96.835 126.785 99.425 127.555 ;
        RECT 100.055 126.830 100.345 127.555 ;
        RECT 100.515 126.785 102.185 127.555 ;
        RECT 102.355 127.095 102.915 127.385 ;
        RECT 103.085 127.095 103.335 127.555 ;
        RECT 96.835 126.265 98.045 126.785 ;
        RECT 96.450 126.145 96.665 126.195 ;
        RECT 94.870 125.735 95.765 126.110 ;
        RECT 96.275 126.065 96.665 126.145 ;
        RECT 98.215 126.095 99.425 126.615 ;
        RECT 100.515 126.265 101.265 126.785 ;
        RECT 93.815 125.305 94.700 125.475 ;
        RECT 94.880 125.005 95.195 125.505 ;
        RECT 95.425 125.175 95.765 125.735 ;
        RECT 95.935 125.005 96.105 126.015 ;
        RECT 96.275 125.220 96.605 126.065 ;
        RECT 96.835 125.005 99.425 126.095 ;
        RECT 100.055 125.005 100.345 126.170 ;
        RECT 101.435 126.095 102.185 126.615 ;
        RECT 100.515 125.005 102.185 126.095 ;
        RECT 102.355 125.725 102.605 127.095 ;
        RECT 103.955 126.925 104.285 127.285 ;
        RECT 102.895 126.735 104.285 126.925 ;
        RECT 104.655 126.785 107.245 127.555 ;
        RECT 107.445 127.165 111.205 127.385 ;
        RECT 107.415 126.820 110.735 126.995 ;
        RECT 102.895 126.645 103.065 126.735 ;
        RECT 102.775 126.315 103.065 126.645 ;
        RECT 103.235 126.315 103.575 126.565 ;
        RECT 103.795 126.315 104.470 126.565 ;
        RECT 102.895 126.065 103.065 126.315 ;
        RECT 102.895 125.895 103.835 126.065 ;
        RECT 104.205 125.955 104.470 126.315 ;
        RECT 104.655 126.265 105.865 126.785 ;
        RECT 106.035 126.095 107.245 126.615 ;
        RECT 102.355 125.175 102.815 125.725 ;
        RECT 103.005 125.005 103.335 125.725 ;
        RECT 103.535 125.345 103.835 125.895 ;
        RECT 104.005 125.005 104.285 125.675 ;
        RECT 104.655 125.005 107.245 126.095 ;
        RECT 107.415 125.855 107.585 126.820 ;
        RECT 107.755 126.195 107.975 126.645 ;
        RECT 108.230 126.365 109.580 126.565 ;
        RECT 109.750 126.195 110.395 126.645 ;
        RECT 107.755 126.025 110.395 126.195 ;
        RECT 110.565 126.195 110.735 126.820 ;
        RECT 110.905 126.905 111.205 127.165 ;
        RECT 111.375 127.085 111.545 127.555 ;
        RECT 111.715 126.915 112.045 127.385 ;
        RECT 112.215 127.085 112.385 127.555 ;
        RECT 112.555 126.915 112.885 127.385 ;
        RECT 113.055 127.085 113.225 127.555 ;
        RECT 111.715 126.905 112.885 126.915 ;
        RECT 113.395 126.915 113.725 127.385 ;
        RECT 113.895 127.085 114.065 127.555 ;
        RECT 114.235 126.915 114.565 127.385 ;
        RECT 113.395 126.905 114.565 126.915 ;
        RECT 110.905 126.735 114.565 126.905 ;
        RECT 114.775 126.785 117.365 127.555 ;
        RECT 117.540 127.025 117.830 127.375 ;
        RECT 118.025 127.195 118.355 127.555 ;
        RECT 118.525 127.025 118.755 127.330 ;
        RECT 117.540 126.855 118.755 127.025 ;
        RECT 111.085 126.395 111.415 126.565 ;
        RECT 111.115 126.195 111.415 126.395 ;
        RECT 111.595 126.365 113.005 126.565 ;
        RECT 113.275 126.365 114.605 126.565 ;
        RECT 113.275 126.195 113.540 126.365 ;
        RECT 114.775 126.265 115.985 126.785 ;
        RECT 118.945 126.685 119.115 127.250 ;
        RECT 110.565 126.025 110.945 126.195 ;
        RECT 111.115 126.025 113.540 126.195 ;
        RECT 110.775 125.855 110.945 126.025 ;
        RECT 113.855 125.855 114.105 126.195 ;
        RECT 107.415 125.685 109.435 125.855 ;
        RECT 108.345 125.515 108.595 125.685 ;
        RECT 109.185 125.515 109.435 125.685 ;
        RECT 109.605 125.685 110.605 125.855 ;
        RECT 110.775 125.685 112.845 125.855 ;
        RECT 107.475 125.005 107.755 125.515 ;
        RECT 107.925 125.345 108.175 125.505 ;
        RECT 108.765 125.345 109.015 125.515 ;
        RECT 109.605 125.345 109.855 125.685 ;
        RECT 110.435 125.515 110.605 125.685 ;
        RECT 111.755 125.515 112.005 125.685 ;
        RECT 112.595 125.515 112.845 125.685 ;
        RECT 113.015 125.685 114.105 125.855 ;
        RECT 107.925 125.175 109.855 125.345 ;
        RECT 110.025 125.005 110.265 125.515 ;
        RECT 110.435 125.175 110.735 125.515 ;
        RECT 110.905 125.005 111.125 125.515 ;
        RECT 111.295 125.345 111.585 125.515 ;
        RECT 112.175 125.345 112.425 125.515 ;
        RECT 113.015 125.345 113.265 125.685 ;
        RECT 111.295 125.175 113.265 125.345 ;
        RECT 113.435 125.005 113.685 125.515 ;
        RECT 113.855 125.175 114.105 125.685 ;
        RECT 114.275 125.005 114.525 126.195 ;
        RECT 116.155 126.095 117.365 126.615 ;
        RECT 117.600 126.535 117.860 126.645 ;
        RECT 117.595 126.365 117.860 126.535 ;
        RECT 117.600 126.315 117.860 126.365 ;
        RECT 118.040 126.315 118.425 126.645 ;
        RECT 118.595 126.515 119.115 126.685 ;
        RECT 119.375 127.055 119.675 127.385 ;
        RECT 119.845 127.075 120.120 127.555 ;
        RECT 114.775 125.005 117.365 126.095 ;
        RECT 117.540 125.005 117.860 126.145 ;
        RECT 118.040 125.265 118.235 126.315 ;
        RECT 118.595 126.135 118.765 126.515 ;
        RECT 118.415 125.855 118.765 126.135 ;
        RECT 118.955 125.985 119.200 126.345 ;
        RECT 119.375 126.145 119.545 127.055 ;
        RECT 120.300 126.905 120.595 127.295 ;
        RECT 120.765 127.075 121.020 127.555 ;
        RECT 121.195 126.905 121.455 127.295 ;
        RECT 121.625 127.075 121.905 127.555 ;
        RECT 122.380 127.095 122.725 127.270 ;
        RECT 119.715 126.315 120.065 126.885 ;
        RECT 120.300 126.735 121.950 126.905 ;
        RECT 120.235 126.395 121.375 126.565 ;
        RECT 120.235 126.145 120.405 126.395 ;
        RECT 121.545 126.225 121.950 126.735 ;
        RECT 122.150 126.315 122.375 126.915 ;
        RECT 119.375 125.975 120.405 126.145 ;
        RECT 121.195 126.055 121.950 126.225 ;
        RECT 122.545 126.130 122.725 127.095 ;
        RECT 122.905 126.745 123.115 127.555 ;
        RECT 123.285 126.915 123.615 127.385 ;
        RECT 123.785 127.085 124.170 127.555 ;
        RECT 123.285 126.745 124.265 126.915 ;
        RECT 123.010 126.315 123.375 126.575 ;
        RECT 123.585 126.395 123.915 126.565 ;
        RECT 123.585 126.130 123.755 126.395 ;
        RECT 118.415 125.175 118.745 125.855 ;
        RECT 118.945 125.005 119.200 125.805 ;
        RECT 119.375 125.175 119.685 125.975 ;
        RECT 121.195 125.805 121.455 126.055 ;
        RECT 122.465 125.960 123.755 126.130 ;
        RECT 119.855 125.005 120.165 125.805 ;
        RECT 120.335 125.635 121.455 125.805 ;
        RECT 120.335 125.175 120.595 125.635 ;
        RECT 120.765 125.005 121.020 125.465 ;
        RECT 121.195 125.175 121.455 125.635 ;
        RECT 121.625 125.005 121.910 125.875 ;
        RECT 122.465 125.735 122.725 125.960 ;
        RECT 124.085 125.790 124.265 126.745 ;
        RECT 124.435 126.805 125.645 127.555 ;
        RECT 125.815 126.830 126.105 127.555 ;
        RECT 126.275 127.055 126.535 127.385 ;
        RECT 126.705 127.195 127.035 127.555 ;
        RECT 127.290 127.175 128.590 127.385 ;
        RECT 124.435 126.265 124.955 126.805 ;
        RECT 125.125 126.095 125.645 126.635 ;
        RECT 122.925 125.005 123.255 125.785 ;
        RECT 123.705 125.175 124.265 125.790 ;
        RECT 124.435 125.005 125.645 126.095 ;
        RECT 125.815 125.005 126.105 126.170 ;
        RECT 126.275 125.855 126.445 127.055 ;
        RECT 127.290 127.025 127.460 127.175 ;
        RECT 126.705 126.900 127.460 127.025 ;
        RECT 126.615 126.855 127.460 126.900 ;
        RECT 126.615 126.735 126.885 126.855 ;
        RECT 126.615 126.160 126.785 126.735 ;
        RECT 127.015 126.295 127.425 126.600 ;
        RECT 127.715 126.565 127.925 126.965 ;
        RECT 127.595 126.355 127.925 126.565 ;
        RECT 128.170 126.565 128.390 126.965 ;
        RECT 128.865 126.790 129.320 127.555 ;
        RECT 129.495 127.055 129.795 127.385 ;
        RECT 129.965 127.075 130.240 127.555 ;
        RECT 128.170 126.355 128.645 126.565 ;
        RECT 128.835 126.365 129.325 126.565 ;
        RECT 126.615 126.125 126.815 126.160 ;
        RECT 128.145 126.125 129.320 126.185 ;
        RECT 126.615 126.015 129.320 126.125 ;
        RECT 126.675 125.955 128.475 126.015 ;
        RECT 128.145 125.925 128.475 125.955 ;
        RECT 126.275 125.175 126.535 125.855 ;
        RECT 126.705 125.005 126.955 125.785 ;
        RECT 127.205 125.755 128.040 125.765 ;
        RECT 128.630 125.755 128.815 125.845 ;
        RECT 127.205 125.555 128.815 125.755 ;
        RECT 127.205 125.175 127.455 125.555 ;
        RECT 128.585 125.515 128.815 125.555 ;
        RECT 129.065 125.395 129.320 126.015 ;
        RECT 127.625 125.005 127.980 125.385 ;
        RECT 128.985 125.175 129.320 125.395 ;
        RECT 129.495 126.145 129.665 127.055 ;
        RECT 130.420 126.905 130.715 127.295 ;
        RECT 130.885 127.075 131.140 127.555 ;
        RECT 131.315 126.905 131.575 127.295 ;
        RECT 131.745 127.075 132.025 127.555 ;
        RECT 132.255 126.970 132.565 127.385 ;
        RECT 132.760 127.175 133.090 127.555 ;
        RECT 133.260 127.215 134.665 127.385 ;
        RECT 133.260 126.985 133.430 127.215 ;
        RECT 129.835 126.315 130.185 126.885 ;
        RECT 130.420 126.735 132.070 126.905 ;
        RECT 130.355 126.395 131.495 126.565 ;
        RECT 130.355 126.145 130.525 126.395 ;
        RECT 131.665 126.225 132.070 126.735 ;
        RECT 129.495 125.975 130.525 126.145 ;
        RECT 131.315 126.055 132.070 126.225 ;
        RECT 129.495 125.175 129.805 125.975 ;
        RECT 131.315 125.805 131.575 126.055 ;
        RECT 129.975 125.005 130.285 125.805 ;
        RECT 130.455 125.635 131.575 125.805 ;
        RECT 130.455 125.175 130.715 125.635 ;
        RECT 130.885 125.005 131.140 125.465 ;
        RECT 131.315 125.175 131.575 125.635 ;
        RECT 131.745 125.005 132.030 125.875 ;
        RECT 132.255 125.855 132.425 126.970 ;
        RECT 132.735 126.815 133.430 126.985 ;
        RECT 134.495 126.985 134.665 127.215 ;
        RECT 134.935 127.155 135.265 127.555 ;
        RECT 135.505 126.985 135.675 127.385 ;
        RECT 132.735 126.645 132.905 126.815 ;
        RECT 132.595 126.315 132.905 126.645 ;
        RECT 133.075 126.315 133.410 126.645 ;
        RECT 133.680 126.315 133.875 126.890 ;
        RECT 134.135 126.645 134.325 126.875 ;
        RECT 134.495 126.815 135.675 126.985 ;
        RECT 135.975 126.735 136.205 127.555 ;
        RECT 136.375 126.755 136.705 127.385 ;
        RECT 134.135 126.315 134.480 126.645 ;
        RECT 134.790 126.315 135.265 126.645 ;
        RECT 135.520 126.315 135.705 126.645 ;
        RECT 135.955 126.315 136.285 126.565 ;
        RECT 132.735 126.145 132.905 126.315 ;
        RECT 136.455 126.155 136.705 126.755 ;
        RECT 136.875 126.735 137.085 127.555 ;
        RECT 137.315 126.785 140.825 127.555 ;
        RECT 141.455 126.835 141.795 127.345 ;
        RECT 137.315 126.265 138.965 126.785 ;
        RECT 132.735 125.975 135.675 126.145 ;
        RECT 132.255 125.215 132.595 125.855 ;
        RECT 133.185 125.635 134.745 125.805 ;
        RECT 132.765 125.005 133.010 125.465 ;
        RECT 133.185 125.175 133.435 125.635 ;
        RECT 133.625 125.005 134.295 125.385 ;
        RECT 134.495 125.175 134.745 125.635 ;
        RECT 135.505 125.175 135.675 125.975 ;
        RECT 135.975 125.005 136.205 126.145 ;
        RECT 136.375 125.175 136.705 126.155 ;
        RECT 136.875 125.005 137.085 126.145 ;
        RECT 139.135 126.095 140.825 126.615 ;
        RECT 137.315 125.005 140.825 126.095 ;
        RECT 141.455 125.435 141.715 126.835 ;
        RECT 141.965 126.755 142.235 127.555 ;
        RECT 141.890 126.315 142.220 126.565 ;
        RECT 142.415 126.315 142.695 127.285 ;
        RECT 142.875 126.315 143.175 127.285 ;
        RECT 143.355 126.315 143.705 127.280 ;
        RECT 143.925 127.055 144.420 127.385 ;
        RECT 141.905 126.145 142.220 126.315 ;
        RECT 143.925 126.145 144.095 127.055 ;
        RECT 141.905 125.975 144.095 126.145 ;
        RECT 141.455 125.175 141.795 125.435 ;
        RECT 141.965 125.005 142.295 125.805 ;
        RECT 142.760 125.175 143.010 125.975 ;
        RECT 143.195 125.005 143.525 125.725 ;
        RECT 143.745 125.175 143.995 125.975 ;
        RECT 144.265 125.565 144.505 126.875 ;
        RECT 144.675 126.735 144.935 127.555 ;
        RECT 145.105 126.735 145.435 127.155 ;
        RECT 145.615 127.070 146.405 127.335 ;
        RECT 145.185 126.645 145.435 126.735 ;
        RECT 144.675 125.685 145.015 126.565 ;
        RECT 145.185 126.395 145.980 126.645 ;
        RECT 144.165 125.005 144.500 125.385 ;
        RECT 144.675 125.005 144.935 125.515 ;
        RECT 145.185 125.175 145.355 126.395 ;
        RECT 146.150 126.215 146.405 127.070 ;
        RECT 146.575 126.915 146.775 127.335 ;
        RECT 146.965 127.095 147.295 127.555 ;
        RECT 146.575 126.395 146.985 126.915 ;
        RECT 147.465 126.905 147.725 127.385 ;
        RECT 147.895 127.175 148.785 127.345 ;
        RECT 147.155 126.215 147.385 126.645 ;
        RECT 145.595 126.045 147.385 126.215 ;
        RECT 145.595 125.680 145.845 126.045 ;
        RECT 146.015 125.685 146.345 125.875 ;
        RECT 146.565 125.750 147.280 126.045 ;
        RECT 147.555 125.875 147.725 126.905 ;
        RECT 147.895 126.620 148.445 127.005 ;
        RECT 148.615 126.450 148.785 127.175 ;
        RECT 146.015 125.510 146.210 125.685 ;
        RECT 145.595 125.005 146.210 125.510 ;
        RECT 146.380 125.175 146.855 125.515 ;
        RECT 147.025 125.005 147.240 125.550 ;
        RECT 147.450 125.175 147.725 125.875 ;
        RECT 147.895 126.380 148.785 126.450 ;
        RECT 148.955 126.850 149.175 127.335 ;
        RECT 149.345 127.015 149.595 127.555 ;
        RECT 149.765 126.905 150.025 127.385 ;
        RECT 148.955 126.425 149.285 126.850 ;
        RECT 147.895 126.355 148.790 126.380 ;
        RECT 147.895 126.340 148.800 126.355 ;
        RECT 147.895 126.325 148.805 126.340 ;
        RECT 147.895 126.320 148.815 126.325 ;
        RECT 147.895 126.310 148.820 126.320 ;
        RECT 147.895 126.300 148.825 126.310 ;
        RECT 147.895 126.295 148.835 126.300 ;
        RECT 147.895 126.285 148.845 126.295 ;
        RECT 147.895 126.280 148.855 126.285 ;
        RECT 147.895 125.830 148.155 126.280 ;
        RECT 148.520 126.275 148.855 126.280 ;
        RECT 148.520 126.270 148.870 126.275 ;
        RECT 148.520 126.260 148.885 126.270 ;
        RECT 148.520 126.255 148.910 126.260 ;
        RECT 149.455 126.255 149.685 126.650 ;
        RECT 148.520 126.250 149.685 126.255 ;
        RECT 148.550 126.215 149.685 126.250 ;
        RECT 148.585 126.190 149.685 126.215 ;
        RECT 148.615 126.160 149.685 126.190 ;
        RECT 148.635 126.130 149.685 126.160 ;
        RECT 148.655 126.100 149.685 126.130 ;
        RECT 148.725 126.090 149.685 126.100 ;
        RECT 148.750 126.080 149.685 126.090 ;
        RECT 148.770 126.065 149.685 126.080 ;
        RECT 148.790 126.050 149.685 126.065 ;
        RECT 148.795 126.040 149.580 126.050 ;
        RECT 148.810 126.005 149.580 126.040 ;
        RECT 148.325 125.685 148.655 125.930 ;
        RECT 148.825 125.755 149.580 126.005 ;
        RECT 149.855 125.875 150.025 126.905 ;
        RECT 150.285 127.005 150.455 127.385 ;
        RECT 150.635 127.175 150.965 127.555 ;
        RECT 150.285 126.835 150.950 127.005 ;
        RECT 151.145 126.880 151.405 127.385 ;
        RECT 150.215 126.285 150.545 126.655 ;
        RECT 150.780 126.580 150.950 126.835 ;
        RECT 150.780 126.250 151.065 126.580 ;
        RECT 150.780 126.105 150.950 126.250 ;
        RECT 148.325 125.660 148.510 125.685 ;
        RECT 147.895 125.560 148.510 125.660 ;
        RECT 147.895 125.005 148.500 125.560 ;
        RECT 148.675 125.175 149.155 125.515 ;
        RECT 149.325 125.005 149.580 125.550 ;
        RECT 149.750 125.175 150.025 125.875 ;
        RECT 150.285 125.935 150.950 126.105 ;
        RECT 151.235 126.080 151.405 126.880 ;
        RECT 151.575 126.830 151.865 127.555 ;
        RECT 152.035 126.880 152.295 127.385 ;
        RECT 152.475 127.175 152.805 127.555 ;
        RECT 152.985 127.005 153.155 127.385 ;
        RECT 150.285 125.175 150.455 125.935 ;
        RECT 150.635 125.005 150.965 125.765 ;
        RECT 151.135 125.175 151.405 126.080 ;
        RECT 151.575 125.005 151.865 126.170 ;
        RECT 152.035 126.080 152.205 126.880 ;
        RECT 152.490 126.835 153.155 127.005 ;
        RECT 152.490 126.580 152.660 126.835 ;
        RECT 153.415 126.785 155.085 127.555 ;
        RECT 155.715 126.805 156.925 127.555 ;
        RECT 152.375 126.250 152.660 126.580 ;
        RECT 152.895 126.285 153.225 126.655 ;
        RECT 153.415 126.265 154.165 126.785 ;
        RECT 152.490 126.105 152.660 126.250 ;
        RECT 152.035 125.175 152.305 126.080 ;
        RECT 152.490 125.935 153.155 126.105 ;
        RECT 154.335 126.095 155.085 126.615 ;
        RECT 152.475 125.005 152.805 125.765 ;
        RECT 152.985 125.175 153.155 125.935 ;
        RECT 153.415 125.005 155.085 126.095 ;
        RECT 155.715 126.095 156.235 126.635 ;
        RECT 156.405 126.265 156.925 126.805 ;
        RECT 155.715 125.005 156.925 126.095 ;
        RECT 22.690 124.835 157.010 125.005 ;
        RECT 22.775 123.745 23.985 124.835 ;
        RECT 22.775 123.035 23.295 123.575 ;
        RECT 23.465 123.205 23.985 123.745 ;
        RECT 25.260 123.865 25.650 124.040 ;
        RECT 26.135 124.035 26.465 124.835 ;
        RECT 26.635 124.045 27.170 124.665 ;
        RECT 25.260 123.695 26.685 123.865 ;
        RECT 22.775 122.285 23.985 123.035 ;
        RECT 25.135 122.965 25.490 123.525 ;
        RECT 25.660 122.795 25.830 123.695 ;
        RECT 26.000 122.965 26.265 123.525 ;
        RECT 26.515 123.195 26.685 123.695 ;
        RECT 26.855 123.025 27.170 124.045 ;
        RECT 27.490 124.205 27.775 124.665 ;
        RECT 27.945 124.375 28.215 124.835 ;
        RECT 27.490 123.985 28.445 124.205 ;
        RECT 27.375 123.255 28.065 123.815 ;
        RECT 28.235 123.085 28.445 123.985 ;
        RECT 25.240 122.285 25.480 122.795 ;
        RECT 25.660 122.465 25.940 122.795 ;
        RECT 26.170 122.285 26.385 122.795 ;
        RECT 26.555 122.455 27.170 123.025 ;
        RECT 27.490 122.915 28.445 123.085 ;
        RECT 28.615 123.815 29.015 124.665 ;
        RECT 29.205 124.205 29.485 124.665 ;
        RECT 30.005 124.375 30.330 124.835 ;
        RECT 29.205 123.985 30.330 124.205 ;
        RECT 28.615 123.255 29.710 123.815 ;
        RECT 29.880 123.525 30.330 123.985 ;
        RECT 30.500 123.695 30.885 124.665 ;
        RECT 27.490 122.455 27.775 122.915 ;
        RECT 27.945 122.285 28.215 122.745 ;
        RECT 28.615 122.455 29.015 123.255 ;
        RECT 29.880 123.195 30.435 123.525 ;
        RECT 29.880 123.085 30.330 123.195 ;
        RECT 29.205 122.915 30.330 123.085 ;
        RECT 30.605 123.025 30.885 123.695 ;
        RECT 29.205 122.455 29.485 122.915 ;
        RECT 30.005 122.285 30.330 122.745 ;
        RECT 30.500 122.455 30.885 123.025 ;
        RECT 31.055 123.695 31.440 124.665 ;
        RECT 31.610 124.375 31.935 124.835 ;
        RECT 32.455 124.205 32.735 124.665 ;
        RECT 31.610 123.985 32.735 124.205 ;
        RECT 31.055 123.025 31.335 123.695 ;
        RECT 31.610 123.525 32.060 123.985 ;
        RECT 32.925 123.815 33.325 124.665 ;
        RECT 33.725 124.375 33.995 124.835 ;
        RECT 34.165 124.205 34.450 124.665 ;
        RECT 31.505 123.195 32.060 123.525 ;
        RECT 32.230 123.255 33.325 123.815 ;
        RECT 31.610 123.085 32.060 123.195 ;
        RECT 31.055 122.455 31.440 123.025 ;
        RECT 31.610 122.915 32.735 123.085 ;
        RECT 31.610 122.285 31.935 122.745 ;
        RECT 32.455 122.455 32.735 122.915 ;
        RECT 32.925 122.455 33.325 123.255 ;
        RECT 33.495 123.985 34.450 124.205 ;
        RECT 33.495 123.085 33.705 123.985 ;
        RECT 33.875 123.255 34.565 123.815 ;
        RECT 35.655 123.670 35.945 124.835 ;
        RECT 36.175 123.775 36.505 124.620 ;
        RECT 36.675 123.825 36.845 124.835 ;
        RECT 37.015 124.105 37.355 124.665 ;
        RECT 37.585 124.335 37.900 124.835 ;
        RECT 38.080 124.365 38.965 124.535 ;
        RECT 36.115 123.695 36.505 123.775 ;
        RECT 37.015 123.730 37.910 124.105 ;
        RECT 36.115 123.645 36.330 123.695 ;
        RECT 33.495 122.915 34.450 123.085 ;
        RECT 36.115 123.065 36.285 123.645 ;
        RECT 37.015 123.525 37.205 123.730 ;
        RECT 38.080 123.525 38.250 124.365 ;
        RECT 39.190 124.335 39.440 124.665 ;
        RECT 36.455 123.195 37.205 123.525 ;
        RECT 37.375 123.195 38.250 123.525 ;
        RECT 36.115 123.025 36.340 123.065 ;
        RECT 37.005 123.025 37.205 123.195 ;
        RECT 33.725 122.285 33.995 122.745 ;
        RECT 34.165 122.455 34.450 122.915 ;
        RECT 35.655 122.285 35.945 123.010 ;
        RECT 36.115 122.940 36.495 123.025 ;
        RECT 36.165 122.505 36.495 122.940 ;
        RECT 36.665 122.285 36.835 122.895 ;
        RECT 37.005 122.500 37.335 123.025 ;
        RECT 37.595 122.285 37.805 122.815 ;
        RECT 38.080 122.735 38.250 123.195 ;
        RECT 38.420 123.235 38.740 124.195 ;
        RECT 38.910 123.445 39.100 124.165 ;
        RECT 39.270 123.265 39.440 124.335 ;
        RECT 39.610 124.035 39.780 124.835 ;
        RECT 39.950 124.390 41.055 124.560 ;
        RECT 39.950 123.775 40.120 124.390 ;
        RECT 41.265 124.240 41.515 124.665 ;
        RECT 41.685 124.375 41.950 124.835 ;
        RECT 40.290 123.855 40.820 124.220 ;
        RECT 41.265 124.110 41.570 124.240 ;
        RECT 39.610 123.685 40.120 123.775 ;
        RECT 39.610 123.515 40.480 123.685 ;
        RECT 39.610 123.445 39.780 123.515 ;
        RECT 39.900 123.265 40.100 123.295 ;
        RECT 38.420 122.905 38.885 123.235 ;
        RECT 39.270 122.965 40.100 123.265 ;
        RECT 39.270 122.735 39.440 122.965 ;
        RECT 38.080 122.565 38.865 122.735 ;
        RECT 39.035 122.565 39.440 122.735 ;
        RECT 39.620 122.285 39.990 122.785 ;
        RECT 40.310 122.735 40.480 123.515 ;
        RECT 40.650 123.155 40.820 123.855 ;
        RECT 40.990 123.325 41.230 123.920 ;
        RECT 40.650 122.935 41.175 123.155 ;
        RECT 41.400 123.005 41.570 124.110 ;
        RECT 41.345 122.875 41.570 123.005 ;
        RECT 41.740 122.915 42.020 123.865 ;
        RECT 41.345 122.735 41.515 122.875 ;
        RECT 40.310 122.565 40.985 122.735 ;
        RECT 41.180 122.565 41.515 122.735 ;
        RECT 41.685 122.285 41.935 122.745 ;
        RECT 42.190 122.545 42.375 124.665 ;
        RECT 42.545 124.335 42.875 124.835 ;
        RECT 43.045 124.165 43.215 124.665 ;
        RECT 42.550 123.995 43.215 124.165 ;
        RECT 42.550 123.005 42.780 123.995 ;
        RECT 42.950 123.175 43.300 123.825 ;
        RECT 43.995 123.775 44.325 124.620 ;
        RECT 44.495 123.825 44.665 124.835 ;
        RECT 44.835 124.105 45.175 124.665 ;
        RECT 45.405 124.335 45.720 124.835 ;
        RECT 45.900 124.365 46.785 124.535 ;
        RECT 43.935 123.695 44.325 123.775 ;
        RECT 44.835 123.730 45.730 124.105 ;
        RECT 43.935 123.645 44.150 123.695 ;
        RECT 43.935 123.065 44.105 123.645 ;
        RECT 44.835 123.525 45.025 123.730 ;
        RECT 45.900 123.525 46.070 124.365 ;
        RECT 47.010 124.335 47.260 124.665 ;
        RECT 44.275 123.195 45.025 123.525 ;
        RECT 45.195 123.195 46.070 123.525 ;
        RECT 43.935 123.025 44.160 123.065 ;
        RECT 44.825 123.025 45.025 123.195 ;
        RECT 42.550 122.835 43.215 123.005 ;
        RECT 43.935 122.940 44.315 123.025 ;
        RECT 42.545 122.285 42.875 122.665 ;
        RECT 43.045 122.545 43.215 122.835 ;
        RECT 43.985 122.505 44.315 122.940 ;
        RECT 44.485 122.285 44.655 122.895 ;
        RECT 44.825 122.500 45.155 123.025 ;
        RECT 45.415 122.285 45.625 122.815 ;
        RECT 45.900 122.735 46.070 123.195 ;
        RECT 46.240 123.235 46.560 124.195 ;
        RECT 46.730 123.445 46.920 124.165 ;
        RECT 47.090 123.265 47.260 124.335 ;
        RECT 47.430 124.035 47.600 124.835 ;
        RECT 47.770 124.390 48.875 124.560 ;
        RECT 47.770 123.775 47.940 124.390 ;
        RECT 49.085 124.240 49.335 124.665 ;
        RECT 49.505 124.375 49.770 124.835 ;
        RECT 48.110 123.855 48.640 124.220 ;
        RECT 49.085 124.110 49.390 124.240 ;
        RECT 47.430 123.685 47.940 123.775 ;
        RECT 47.430 123.515 48.300 123.685 ;
        RECT 47.430 123.445 47.600 123.515 ;
        RECT 47.720 123.265 47.920 123.295 ;
        RECT 46.240 122.905 46.705 123.235 ;
        RECT 47.090 122.965 47.920 123.265 ;
        RECT 47.090 122.735 47.260 122.965 ;
        RECT 45.900 122.565 46.685 122.735 ;
        RECT 46.855 122.565 47.260 122.735 ;
        RECT 47.440 122.285 47.810 122.785 ;
        RECT 48.130 122.735 48.300 123.515 ;
        RECT 48.470 123.155 48.640 123.855 ;
        RECT 48.810 123.325 49.050 123.920 ;
        RECT 48.470 122.935 48.995 123.155 ;
        RECT 49.220 123.005 49.390 124.110 ;
        RECT 49.165 122.875 49.390 123.005 ;
        RECT 49.560 122.915 49.840 123.865 ;
        RECT 49.165 122.735 49.335 122.875 ;
        RECT 48.130 122.565 48.805 122.735 ;
        RECT 49.000 122.565 49.335 122.735 ;
        RECT 49.505 122.285 49.755 122.745 ;
        RECT 50.010 122.545 50.195 124.665 ;
        RECT 50.365 124.335 50.695 124.835 ;
        RECT 50.865 124.165 51.035 124.665 ;
        RECT 50.370 123.995 51.035 124.165 ;
        RECT 50.370 123.005 50.600 123.995 ;
        RECT 51.480 123.865 51.870 124.040 ;
        RECT 52.355 124.035 52.685 124.835 ;
        RECT 52.855 124.045 53.390 124.665 ;
        RECT 50.770 123.175 51.120 123.825 ;
        RECT 51.480 123.695 52.905 123.865 ;
        RECT 50.370 122.835 51.035 123.005 ;
        RECT 51.355 122.965 51.710 123.525 ;
        RECT 50.365 122.285 50.695 122.665 ;
        RECT 50.865 122.545 51.035 122.835 ;
        RECT 51.880 122.795 52.050 123.695 ;
        RECT 52.220 122.965 52.485 123.525 ;
        RECT 52.735 123.195 52.905 123.695 ;
        RECT 53.075 123.025 53.390 124.045 ;
        RECT 53.605 124.225 53.935 124.655 ;
        RECT 54.115 124.395 54.310 124.835 ;
        RECT 54.480 124.225 54.810 124.655 ;
        RECT 53.605 124.055 54.810 124.225 ;
        RECT 53.605 123.725 54.500 124.055 ;
        RECT 54.980 123.885 55.255 124.655 ;
        RECT 54.670 123.695 55.255 123.885 ;
        RECT 55.440 123.695 55.760 124.835 ;
        RECT 53.610 123.195 53.905 123.525 ;
        RECT 54.085 123.195 54.500 123.525 ;
        RECT 51.460 122.285 51.700 122.795 ;
        RECT 51.880 122.465 52.160 122.795 ;
        RECT 52.390 122.285 52.605 122.795 ;
        RECT 52.775 122.455 53.390 123.025 ;
        RECT 53.605 122.285 53.905 123.015 ;
        RECT 54.085 122.575 54.315 123.195 ;
        RECT 54.670 123.025 54.845 123.695 ;
        RECT 55.940 123.525 56.135 124.575 ;
        RECT 56.315 123.985 56.645 124.665 ;
        RECT 56.845 124.035 57.100 124.835 ;
        RECT 56.315 123.705 56.665 123.985 ;
        RECT 54.515 122.845 54.845 123.025 ;
        RECT 55.015 122.875 55.255 123.525 ;
        RECT 55.500 123.475 55.760 123.525 ;
        RECT 55.495 123.305 55.760 123.475 ;
        RECT 55.500 123.195 55.760 123.305 ;
        RECT 55.940 123.195 56.325 123.525 ;
        RECT 56.495 123.325 56.665 123.705 ;
        RECT 56.855 123.495 57.100 123.855 ;
        RECT 57.275 123.745 60.785 124.835 ;
        RECT 56.495 123.155 57.015 123.325 ;
        RECT 54.515 122.465 54.740 122.845 ;
        RECT 55.440 122.815 56.655 122.985 ;
        RECT 54.910 122.285 55.240 122.675 ;
        RECT 55.440 122.465 55.730 122.815 ;
        RECT 55.925 122.285 56.255 122.645 ;
        RECT 56.425 122.510 56.655 122.815 ;
        RECT 56.845 122.590 57.015 123.155 ;
        RECT 57.275 123.055 58.925 123.575 ;
        RECT 59.095 123.225 60.785 123.745 ;
        RECT 61.415 123.670 61.705 124.835 ;
        RECT 61.875 123.745 64.465 124.835 ;
        RECT 65.105 124.025 65.400 124.835 ;
        RECT 61.875 123.055 63.085 123.575 ;
        RECT 63.255 123.225 64.465 123.745 ;
        RECT 65.580 123.525 65.825 124.665 ;
        RECT 66.000 124.025 66.260 124.835 ;
        RECT 66.860 124.830 73.135 124.835 ;
        RECT 66.440 123.525 66.690 124.660 ;
        RECT 66.860 124.035 67.120 124.830 ;
        RECT 67.290 123.935 67.550 124.660 ;
        RECT 67.720 124.105 67.980 124.830 ;
        RECT 68.150 123.935 68.410 124.660 ;
        RECT 68.580 124.105 68.840 124.830 ;
        RECT 69.010 123.935 69.270 124.660 ;
        RECT 69.440 124.105 69.700 124.830 ;
        RECT 69.870 123.935 70.130 124.660 ;
        RECT 70.300 124.105 70.545 124.830 ;
        RECT 70.715 123.935 70.975 124.660 ;
        RECT 71.160 124.105 71.405 124.830 ;
        RECT 71.575 123.935 71.835 124.660 ;
        RECT 72.020 124.105 72.265 124.830 ;
        RECT 72.435 123.935 72.695 124.660 ;
        RECT 72.880 124.105 73.135 124.830 ;
        RECT 67.290 123.920 72.695 123.935 ;
        RECT 73.305 123.920 73.595 124.660 ;
        RECT 73.765 124.090 74.035 124.835 ;
        RECT 67.290 123.695 74.035 123.920 ;
        RECT 74.295 123.745 75.965 124.835 ;
        RECT 76.225 124.165 76.395 124.665 ;
        RECT 76.565 124.335 76.895 124.835 ;
        RECT 76.225 123.995 76.890 124.165 ;
        RECT 57.275 122.285 60.785 123.055 ;
        RECT 61.415 122.285 61.705 123.010 ;
        RECT 61.875 122.285 64.465 123.055 ;
        RECT 65.095 122.965 65.410 123.525 ;
        RECT 65.580 123.275 72.700 123.525 ;
        RECT 65.095 122.285 65.400 122.795 ;
        RECT 65.580 122.465 65.830 123.275 ;
        RECT 66.000 122.285 66.260 122.810 ;
        RECT 66.440 122.465 66.690 123.275 ;
        RECT 72.870 123.105 74.035 123.695 ;
        RECT 67.290 122.935 74.035 123.105 ;
        RECT 74.295 123.055 75.045 123.575 ;
        RECT 75.215 123.225 75.965 123.745 ;
        RECT 76.140 123.175 76.490 123.825 ;
        RECT 66.860 122.285 67.120 122.845 ;
        RECT 67.290 122.480 67.550 122.935 ;
        RECT 67.720 122.285 67.980 122.765 ;
        RECT 68.150 122.480 68.410 122.935 ;
        RECT 68.580 122.285 68.840 122.765 ;
        RECT 69.010 122.480 69.270 122.935 ;
        RECT 69.440 122.285 69.685 122.765 ;
        RECT 69.855 122.480 70.130 122.935 ;
        RECT 70.300 122.285 70.545 122.765 ;
        RECT 70.715 122.480 70.975 122.935 ;
        RECT 71.155 122.285 71.405 122.765 ;
        RECT 71.575 122.480 71.835 122.935 ;
        RECT 72.015 122.285 72.265 122.765 ;
        RECT 72.435 122.480 72.695 122.935 ;
        RECT 72.875 122.285 73.135 122.765 ;
        RECT 73.305 122.480 73.565 122.935 ;
        RECT 73.735 122.285 74.035 122.765 ;
        RECT 74.295 122.285 75.965 123.055 ;
        RECT 76.660 123.005 76.890 123.995 ;
        RECT 76.225 122.835 76.890 123.005 ;
        RECT 76.225 122.545 76.395 122.835 ;
        RECT 76.565 122.285 76.895 122.665 ;
        RECT 77.065 122.545 77.250 124.665 ;
        RECT 77.490 124.375 77.755 124.835 ;
        RECT 77.925 124.240 78.175 124.665 ;
        RECT 78.385 124.390 79.490 124.560 ;
        RECT 77.870 124.110 78.175 124.240 ;
        RECT 77.420 122.915 77.700 123.865 ;
        RECT 77.870 123.005 78.040 124.110 ;
        RECT 78.210 123.325 78.450 123.920 ;
        RECT 78.620 123.855 79.150 124.220 ;
        RECT 78.620 123.155 78.790 123.855 ;
        RECT 79.320 123.775 79.490 124.390 ;
        RECT 79.660 124.035 79.830 124.835 ;
        RECT 80.000 124.335 80.250 124.665 ;
        RECT 80.475 124.365 81.360 124.535 ;
        RECT 79.320 123.685 79.830 123.775 ;
        RECT 77.870 122.875 78.095 123.005 ;
        RECT 78.265 122.935 78.790 123.155 ;
        RECT 78.960 123.515 79.830 123.685 ;
        RECT 77.505 122.285 77.755 122.745 ;
        RECT 77.925 122.735 78.095 122.875 ;
        RECT 78.960 122.735 79.130 123.515 ;
        RECT 79.660 123.445 79.830 123.515 ;
        RECT 79.340 123.265 79.540 123.295 ;
        RECT 80.000 123.265 80.170 124.335 ;
        RECT 80.340 123.445 80.530 124.165 ;
        RECT 79.340 122.965 80.170 123.265 ;
        RECT 80.700 123.235 81.020 124.195 ;
        RECT 77.925 122.565 78.260 122.735 ;
        RECT 78.455 122.565 79.130 122.735 ;
        RECT 79.450 122.285 79.820 122.785 ;
        RECT 80.000 122.735 80.170 122.965 ;
        RECT 80.555 122.905 81.020 123.235 ;
        RECT 81.190 123.525 81.360 124.365 ;
        RECT 81.540 124.335 81.855 124.835 ;
        RECT 82.085 124.105 82.425 124.665 ;
        RECT 81.530 123.730 82.425 124.105 ;
        RECT 82.595 123.825 82.765 124.835 ;
        RECT 82.235 123.525 82.425 123.730 ;
        RECT 82.935 123.775 83.265 124.620 ;
        RECT 83.495 124.115 83.955 124.665 ;
        RECT 84.145 124.115 84.475 124.835 ;
        RECT 82.935 123.695 83.325 123.775 ;
        RECT 83.110 123.645 83.325 123.695 ;
        RECT 81.190 123.195 82.065 123.525 ;
        RECT 82.235 123.195 82.985 123.525 ;
        RECT 81.190 122.735 81.360 123.195 ;
        RECT 82.235 123.025 82.435 123.195 ;
        RECT 83.155 123.065 83.325 123.645 ;
        RECT 83.100 123.025 83.325 123.065 ;
        RECT 80.000 122.565 80.405 122.735 ;
        RECT 80.575 122.565 81.360 122.735 ;
        RECT 81.635 122.285 81.845 122.815 ;
        RECT 82.105 122.500 82.435 123.025 ;
        RECT 82.945 122.940 83.325 123.025 ;
        RECT 82.605 122.285 82.775 122.895 ;
        RECT 82.945 122.505 83.275 122.940 ;
        RECT 83.495 122.745 83.745 124.115 ;
        RECT 84.675 123.945 84.975 124.495 ;
        RECT 85.145 124.165 85.425 124.835 ;
        RECT 84.035 123.775 84.975 123.945 ;
        RECT 84.035 123.525 84.205 123.775 ;
        RECT 85.345 123.525 85.610 123.885 ;
        RECT 85.795 123.745 87.005 124.835 ;
        RECT 83.915 123.195 84.205 123.525 ;
        RECT 84.375 123.275 84.715 123.525 ;
        RECT 84.935 123.275 85.610 123.525 ;
        RECT 84.035 123.105 84.205 123.195 ;
        RECT 84.035 122.915 85.425 123.105 ;
        RECT 83.495 122.455 84.055 122.745 ;
        RECT 84.225 122.285 84.475 122.745 ;
        RECT 85.095 122.555 85.425 122.915 ;
        RECT 85.795 123.035 86.315 123.575 ;
        RECT 86.485 123.205 87.005 123.745 ;
        RECT 87.175 123.670 87.465 124.835 ;
        RECT 87.835 124.165 88.115 124.835 ;
        RECT 88.285 123.945 88.585 124.495 ;
        RECT 88.785 124.115 89.115 124.835 ;
        RECT 89.305 124.115 89.765 124.665 ;
        RECT 87.650 123.525 87.915 123.885 ;
        RECT 88.285 123.775 89.225 123.945 ;
        RECT 89.055 123.525 89.225 123.775 ;
        RECT 87.650 123.275 88.325 123.525 ;
        RECT 88.545 123.275 88.885 123.525 ;
        RECT 89.055 123.195 89.345 123.525 ;
        RECT 89.055 123.105 89.225 123.195 ;
        RECT 85.795 122.285 87.005 123.035 ;
        RECT 87.175 122.285 87.465 123.010 ;
        RECT 87.835 122.915 89.225 123.105 ;
        RECT 87.835 122.555 88.165 122.915 ;
        RECT 89.515 122.745 89.765 124.115 ;
        RECT 89.935 123.745 91.605 124.835 ;
        RECT 88.785 122.285 89.035 122.745 ;
        RECT 89.205 122.455 89.765 122.745 ;
        RECT 89.935 123.055 90.685 123.575 ;
        RECT 90.855 123.225 91.605 123.745 ;
        RECT 91.775 123.760 92.045 124.665 ;
        RECT 92.215 124.075 92.545 124.835 ;
        RECT 92.725 123.905 92.895 124.665 ;
        RECT 93.355 124.165 93.635 124.835 ;
        RECT 89.935 122.285 91.605 123.055 ;
        RECT 91.775 122.960 91.945 123.760 ;
        RECT 92.230 123.735 92.895 123.905 ;
        RECT 93.805 123.945 94.105 124.495 ;
        RECT 94.305 124.115 94.635 124.835 ;
        RECT 94.825 124.115 95.285 124.665 ;
        RECT 92.230 123.590 92.400 123.735 ;
        RECT 92.115 123.260 92.400 123.590 ;
        RECT 92.230 123.005 92.400 123.260 ;
        RECT 92.635 123.185 92.965 123.555 ;
        RECT 93.170 123.525 93.435 123.885 ;
        RECT 93.805 123.775 94.745 123.945 ;
        RECT 94.575 123.525 94.745 123.775 ;
        RECT 93.170 123.275 93.845 123.525 ;
        RECT 94.065 123.275 94.405 123.525 ;
        RECT 94.575 123.195 94.865 123.525 ;
        RECT 94.575 123.105 94.745 123.195 ;
        RECT 91.775 122.455 92.035 122.960 ;
        RECT 92.230 122.835 92.895 123.005 ;
        RECT 92.215 122.285 92.545 122.665 ;
        RECT 92.725 122.455 92.895 122.835 ;
        RECT 93.355 122.915 94.745 123.105 ;
        RECT 93.355 122.555 93.685 122.915 ;
        RECT 95.035 122.745 95.285 124.115 ;
        RECT 95.455 123.745 97.125 124.835 ;
        RECT 94.305 122.285 94.555 122.745 ;
        RECT 94.725 122.455 95.285 122.745 ;
        RECT 95.455 123.055 96.205 123.575 ;
        RECT 96.375 123.225 97.125 123.745 ;
        RECT 97.385 123.905 97.555 124.665 ;
        RECT 97.735 124.075 98.065 124.835 ;
        RECT 97.385 123.735 98.050 123.905 ;
        RECT 98.235 123.760 98.505 124.665 ;
        RECT 98.765 124.165 98.935 124.665 ;
        RECT 99.105 124.335 99.435 124.835 ;
        RECT 98.765 123.995 99.430 124.165 ;
        RECT 97.880 123.590 98.050 123.735 ;
        RECT 97.315 123.185 97.645 123.555 ;
        RECT 97.880 123.260 98.165 123.590 ;
        RECT 95.455 122.285 97.125 123.055 ;
        RECT 97.880 123.005 98.050 123.260 ;
        RECT 97.385 122.835 98.050 123.005 ;
        RECT 98.335 122.960 98.505 123.760 ;
        RECT 98.680 123.175 99.030 123.825 ;
        RECT 99.200 123.005 99.430 123.995 ;
        RECT 97.385 122.455 97.555 122.835 ;
        RECT 97.735 122.285 98.065 122.665 ;
        RECT 98.245 122.455 98.505 122.960 ;
        RECT 98.765 122.835 99.430 123.005 ;
        RECT 98.765 122.545 98.935 122.835 ;
        RECT 99.105 122.285 99.435 122.665 ;
        RECT 99.605 122.545 99.790 124.665 ;
        RECT 100.030 124.375 100.295 124.835 ;
        RECT 100.465 124.240 100.715 124.665 ;
        RECT 100.925 124.390 102.030 124.560 ;
        RECT 100.410 124.110 100.715 124.240 ;
        RECT 99.960 122.915 100.240 123.865 ;
        RECT 100.410 123.005 100.580 124.110 ;
        RECT 100.750 123.325 100.990 123.920 ;
        RECT 101.160 123.855 101.690 124.220 ;
        RECT 101.160 123.155 101.330 123.855 ;
        RECT 101.860 123.775 102.030 124.390 ;
        RECT 102.200 124.035 102.370 124.835 ;
        RECT 102.540 124.335 102.790 124.665 ;
        RECT 103.015 124.365 103.900 124.535 ;
        RECT 101.860 123.685 102.370 123.775 ;
        RECT 100.410 122.875 100.635 123.005 ;
        RECT 100.805 122.935 101.330 123.155 ;
        RECT 101.500 123.515 102.370 123.685 ;
        RECT 100.045 122.285 100.295 122.745 ;
        RECT 100.465 122.735 100.635 122.875 ;
        RECT 101.500 122.735 101.670 123.515 ;
        RECT 102.200 123.445 102.370 123.515 ;
        RECT 101.880 123.265 102.080 123.295 ;
        RECT 102.540 123.265 102.710 124.335 ;
        RECT 102.880 123.445 103.070 124.165 ;
        RECT 101.880 122.965 102.710 123.265 ;
        RECT 103.240 123.235 103.560 124.195 ;
        RECT 100.465 122.565 100.800 122.735 ;
        RECT 100.995 122.565 101.670 122.735 ;
        RECT 101.990 122.285 102.360 122.785 ;
        RECT 102.540 122.735 102.710 122.965 ;
        RECT 103.095 122.905 103.560 123.235 ;
        RECT 103.730 123.525 103.900 124.365 ;
        RECT 104.080 124.335 104.395 124.835 ;
        RECT 104.625 124.105 104.965 124.665 ;
        RECT 104.070 123.730 104.965 124.105 ;
        RECT 105.135 123.825 105.305 124.835 ;
        RECT 104.775 123.525 104.965 123.730 ;
        RECT 105.475 123.775 105.805 124.620 ;
        RECT 105.475 123.695 105.865 123.775 ;
        RECT 105.650 123.645 105.865 123.695 ;
        RECT 103.730 123.195 104.605 123.525 ;
        RECT 104.775 123.195 105.525 123.525 ;
        RECT 103.730 122.735 103.900 123.195 ;
        RECT 104.775 123.025 104.975 123.195 ;
        RECT 105.695 123.065 105.865 123.645 ;
        RECT 105.640 123.025 105.865 123.065 ;
        RECT 102.540 122.565 102.945 122.735 ;
        RECT 103.115 122.565 103.900 122.735 ;
        RECT 104.175 122.285 104.385 122.815 ;
        RECT 104.645 122.500 104.975 123.025 ;
        RECT 105.485 122.940 105.865 123.025 ;
        RECT 106.035 123.760 106.305 124.665 ;
        RECT 106.475 124.075 106.805 124.835 ;
        RECT 106.985 123.905 107.155 124.665 ;
        RECT 106.035 122.960 106.205 123.760 ;
        RECT 106.490 123.735 107.155 123.905 ;
        RECT 106.490 123.590 106.660 123.735 ;
        RECT 106.375 123.260 106.660 123.590 ;
        RECT 107.420 123.695 107.755 124.665 ;
        RECT 107.925 123.695 108.095 124.835 ;
        RECT 108.265 124.495 110.295 124.665 ;
        RECT 106.490 123.005 106.660 123.260 ;
        RECT 106.895 123.185 107.225 123.555 ;
        RECT 107.420 123.025 107.590 123.695 ;
        RECT 108.265 123.525 108.435 124.495 ;
        RECT 107.760 123.195 108.015 123.525 ;
        RECT 108.240 123.195 108.435 123.525 ;
        RECT 108.605 124.155 109.730 124.325 ;
        RECT 107.845 123.025 108.015 123.195 ;
        RECT 108.605 123.025 108.775 124.155 ;
        RECT 105.145 122.285 105.315 122.895 ;
        RECT 105.485 122.505 105.815 122.940 ;
        RECT 106.035 122.455 106.295 122.960 ;
        RECT 106.490 122.835 107.155 123.005 ;
        RECT 106.475 122.285 106.805 122.665 ;
        RECT 106.985 122.455 107.155 122.835 ;
        RECT 107.420 122.455 107.675 123.025 ;
        RECT 107.845 122.855 108.775 123.025 ;
        RECT 108.945 123.815 109.955 123.985 ;
        RECT 108.945 123.015 109.115 123.815 ;
        RECT 108.600 122.820 108.775 122.855 ;
        RECT 107.845 122.285 108.175 122.685 ;
        RECT 108.600 122.455 109.130 122.820 ;
        RECT 109.320 122.795 109.595 123.615 ;
        RECT 109.315 122.625 109.595 122.795 ;
        RECT 109.320 122.455 109.595 122.625 ;
        RECT 109.765 122.455 109.955 123.815 ;
        RECT 110.125 123.830 110.295 124.495 ;
        RECT 110.465 124.075 110.635 124.835 ;
        RECT 110.870 124.075 111.385 124.485 ;
        RECT 110.125 123.640 110.875 123.830 ;
        RECT 111.045 123.265 111.385 124.075 ;
        RECT 111.555 123.745 112.765 124.835 ;
        RECT 110.155 123.095 111.385 123.265 ;
        RECT 110.135 122.285 110.645 122.820 ;
        RECT 110.865 122.490 111.110 123.095 ;
        RECT 111.555 123.035 112.075 123.575 ;
        RECT 112.245 123.205 112.765 123.745 ;
        RECT 112.935 123.670 113.225 124.835 ;
        RECT 113.395 123.745 116.905 124.835 ;
        RECT 118.005 124.025 118.300 124.835 ;
        RECT 113.395 123.055 115.045 123.575 ;
        RECT 115.215 123.225 116.905 123.745 ;
        RECT 118.480 123.525 118.725 124.665 ;
        RECT 118.900 124.025 119.160 124.835 ;
        RECT 119.760 124.830 126.035 124.835 ;
        RECT 119.340 123.525 119.590 124.660 ;
        RECT 119.760 124.035 120.020 124.830 ;
        RECT 120.190 123.935 120.450 124.660 ;
        RECT 120.620 124.105 120.880 124.830 ;
        RECT 121.050 123.935 121.310 124.660 ;
        RECT 121.480 124.105 121.740 124.830 ;
        RECT 121.910 123.935 122.170 124.660 ;
        RECT 122.340 124.105 122.600 124.830 ;
        RECT 122.770 123.935 123.030 124.660 ;
        RECT 123.200 124.105 123.445 124.830 ;
        RECT 123.615 123.935 123.875 124.660 ;
        RECT 124.060 124.105 124.305 124.830 ;
        RECT 124.475 123.935 124.735 124.660 ;
        RECT 124.920 124.105 125.165 124.830 ;
        RECT 125.335 123.935 125.595 124.660 ;
        RECT 125.780 124.105 126.035 124.830 ;
        RECT 120.190 123.920 125.595 123.935 ;
        RECT 126.205 123.920 126.495 124.660 ;
        RECT 126.665 124.090 126.935 124.835 ;
        RECT 127.285 124.165 127.455 124.665 ;
        RECT 127.625 124.335 127.955 124.835 ;
        RECT 127.285 123.995 127.950 124.165 ;
        RECT 120.190 123.695 126.935 123.920 ;
        RECT 111.555 122.285 112.765 123.035 ;
        RECT 112.935 122.285 113.225 123.010 ;
        RECT 113.395 122.285 116.905 123.055 ;
        RECT 117.995 122.965 118.310 123.525 ;
        RECT 118.480 123.275 125.600 123.525 ;
        RECT 117.995 122.285 118.300 122.795 ;
        RECT 118.480 122.465 118.730 123.275 ;
        RECT 118.900 122.285 119.160 122.810 ;
        RECT 119.340 122.465 119.590 123.275 ;
        RECT 125.770 123.105 126.935 123.695 ;
        RECT 127.200 123.175 127.550 123.825 ;
        RECT 120.190 122.935 126.935 123.105 ;
        RECT 127.720 123.005 127.950 123.995 ;
        RECT 119.760 122.285 120.020 122.845 ;
        RECT 120.190 122.480 120.450 122.935 ;
        RECT 120.620 122.285 120.880 122.765 ;
        RECT 121.050 122.480 121.310 122.935 ;
        RECT 121.480 122.285 121.740 122.765 ;
        RECT 121.910 122.480 122.170 122.935 ;
        RECT 122.340 122.285 122.585 122.765 ;
        RECT 122.755 122.480 123.030 122.935 ;
        RECT 123.200 122.285 123.445 122.765 ;
        RECT 123.615 122.480 123.875 122.935 ;
        RECT 124.055 122.285 124.305 122.765 ;
        RECT 124.475 122.480 124.735 122.935 ;
        RECT 124.915 122.285 125.165 122.765 ;
        RECT 125.335 122.480 125.595 122.935 ;
        RECT 125.775 122.285 126.035 122.765 ;
        RECT 126.205 122.480 126.465 122.935 ;
        RECT 127.285 122.835 127.950 123.005 ;
        RECT 126.635 122.285 126.935 122.765 ;
        RECT 127.285 122.545 127.455 122.835 ;
        RECT 127.625 122.285 127.955 122.665 ;
        RECT 128.125 122.545 128.310 124.665 ;
        RECT 128.550 124.375 128.815 124.835 ;
        RECT 128.985 124.240 129.235 124.665 ;
        RECT 129.445 124.390 130.550 124.560 ;
        RECT 128.930 124.110 129.235 124.240 ;
        RECT 128.480 122.915 128.760 123.865 ;
        RECT 128.930 123.005 129.100 124.110 ;
        RECT 129.270 123.325 129.510 123.920 ;
        RECT 129.680 123.855 130.210 124.220 ;
        RECT 129.680 123.155 129.850 123.855 ;
        RECT 130.380 123.775 130.550 124.390 ;
        RECT 130.720 124.035 130.890 124.835 ;
        RECT 131.060 124.335 131.310 124.665 ;
        RECT 131.535 124.365 132.420 124.535 ;
        RECT 130.380 123.685 130.890 123.775 ;
        RECT 128.930 122.875 129.155 123.005 ;
        RECT 129.325 122.935 129.850 123.155 ;
        RECT 130.020 123.515 130.890 123.685 ;
        RECT 128.565 122.285 128.815 122.745 ;
        RECT 128.985 122.735 129.155 122.875 ;
        RECT 130.020 122.735 130.190 123.515 ;
        RECT 130.720 123.445 130.890 123.515 ;
        RECT 130.400 123.265 130.600 123.295 ;
        RECT 131.060 123.265 131.230 124.335 ;
        RECT 131.400 123.445 131.590 124.165 ;
        RECT 130.400 122.965 131.230 123.265 ;
        RECT 131.760 123.235 132.080 124.195 ;
        RECT 128.985 122.565 129.320 122.735 ;
        RECT 129.515 122.565 130.190 122.735 ;
        RECT 130.510 122.285 130.880 122.785 ;
        RECT 131.060 122.735 131.230 122.965 ;
        RECT 131.615 122.905 132.080 123.235 ;
        RECT 132.250 123.525 132.420 124.365 ;
        RECT 132.600 124.335 132.915 124.835 ;
        RECT 133.145 124.105 133.485 124.665 ;
        RECT 132.590 123.730 133.485 124.105 ;
        RECT 133.655 123.825 133.825 124.835 ;
        RECT 133.295 123.525 133.485 123.730 ;
        RECT 133.995 123.775 134.325 124.620 ;
        RECT 133.995 123.695 134.385 123.775 ;
        RECT 134.170 123.645 134.385 123.695 ;
        RECT 132.250 123.195 133.125 123.525 ;
        RECT 133.295 123.195 134.045 123.525 ;
        RECT 132.250 122.735 132.420 123.195 ;
        RECT 133.295 123.025 133.495 123.195 ;
        RECT 134.215 123.065 134.385 123.645 ;
        RECT 134.160 123.025 134.385 123.065 ;
        RECT 131.060 122.565 131.465 122.735 ;
        RECT 131.635 122.565 132.420 122.735 ;
        RECT 132.695 122.285 132.905 122.815 ;
        RECT 133.165 122.500 133.495 123.025 ;
        RECT 134.005 122.940 134.385 123.025 ;
        RECT 134.555 123.695 134.940 124.665 ;
        RECT 135.110 124.375 135.435 124.835 ;
        RECT 135.955 124.205 136.235 124.665 ;
        RECT 135.110 123.985 136.235 124.205 ;
        RECT 134.555 123.025 134.835 123.695 ;
        RECT 135.110 123.525 135.560 123.985 ;
        RECT 136.425 123.815 136.825 124.665 ;
        RECT 137.225 124.375 137.495 124.835 ;
        RECT 137.665 124.205 137.950 124.665 ;
        RECT 135.005 123.195 135.560 123.525 ;
        RECT 135.730 123.255 136.825 123.815 ;
        RECT 135.110 123.085 135.560 123.195 ;
        RECT 133.665 122.285 133.835 122.895 ;
        RECT 134.005 122.505 134.335 122.940 ;
        RECT 134.555 122.455 134.940 123.025 ;
        RECT 135.110 122.915 136.235 123.085 ;
        RECT 135.110 122.285 135.435 122.745 ;
        RECT 135.955 122.455 136.235 122.915 ;
        RECT 136.425 122.455 136.825 123.255 ;
        RECT 136.995 123.985 137.950 124.205 ;
        RECT 136.995 123.085 137.205 123.985 ;
        RECT 137.375 123.255 138.065 123.815 ;
        RECT 138.695 123.670 138.985 124.835 ;
        RECT 139.155 123.725 139.415 124.665 ;
        RECT 139.585 124.435 139.915 124.835 ;
        RECT 141.060 124.570 141.315 124.665 ;
        RECT 140.175 124.400 141.315 124.570 ;
        RECT 141.485 124.455 141.815 124.625 ;
        RECT 140.175 124.175 140.345 124.400 ;
        RECT 139.585 124.005 140.345 124.175 ;
        RECT 141.060 124.265 141.315 124.400 ;
        RECT 136.995 122.915 137.950 123.085 ;
        RECT 139.155 123.010 139.330 123.725 ;
        RECT 139.585 123.525 139.755 124.005 ;
        RECT 140.610 123.915 140.780 124.105 ;
        RECT 141.060 124.095 141.470 124.265 ;
        RECT 139.500 123.195 139.755 123.525 ;
        RECT 139.980 123.195 140.310 123.815 ;
        RECT 140.610 123.745 141.130 123.915 ;
        RECT 140.480 123.195 140.770 123.575 ;
        RECT 140.960 123.025 141.130 123.745 ;
        RECT 137.225 122.285 137.495 122.745 ;
        RECT 137.665 122.455 137.950 122.915 ;
        RECT 138.695 122.285 138.985 123.010 ;
        RECT 139.155 122.455 139.415 123.010 ;
        RECT 140.250 122.855 141.130 123.025 ;
        RECT 141.300 123.070 141.470 124.095 ;
        RECT 141.645 124.205 141.815 124.455 ;
        RECT 141.985 124.375 142.235 124.835 ;
        RECT 142.405 124.205 142.585 124.665 ;
        RECT 141.645 124.035 142.585 124.205 ;
        RECT 141.670 123.555 142.150 123.855 ;
        RECT 141.300 122.900 141.650 123.070 ;
        RECT 141.890 122.965 142.150 123.555 ;
        RECT 142.350 122.965 142.610 123.855 ;
        RECT 142.835 123.695 143.110 124.665 ;
        RECT 143.320 124.035 143.600 124.835 ;
        RECT 143.770 124.325 145.385 124.655 ;
        RECT 143.770 123.985 144.945 124.155 ;
        RECT 143.770 123.865 143.940 123.985 ;
        RECT 143.280 123.695 143.940 123.865 ;
        RECT 139.585 122.285 140.015 122.730 ;
        RECT 140.250 122.455 140.420 122.855 ;
        RECT 140.590 122.285 141.310 122.685 ;
        RECT 141.480 122.455 141.650 122.900 ;
        RECT 142.835 122.960 143.005 123.695 ;
        RECT 143.280 123.525 143.450 123.695 ;
        RECT 144.200 123.525 144.445 123.815 ;
        RECT 144.615 123.695 144.945 123.985 ;
        RECT 145.205 123.525 145.375 124.085 ;
        RECT 145.625 123.695 145.885 124.835 ;
        RECT 146.095 123.695 146.325 124.835 ;
        RECT 146.495 123.685 146.825 124.665 ;
        RECT 146.995 123.695 147.205 124.835 ;
        RECT 147.955 123.775 148.285 124.620 ;
        RECT 148.455 123.825 148.625 124.835 ;
        RECT 148.795 124.105 149.135 124.665 ;
        RECT 149.365 124.335 149.680 124.835 ;
        RECT 149.860 124.365 150.745 124.535 ;
        RECT 147.895 123.695 148.285 123.775 ;
        RECT 148.795 123.730 149.690 124.105 ;
        RECT 143.175 123.195 143.450 123.525 ;
        RECT 143.620 123.195 144.445 123.525 ;
        RECT 144.660 123.195 145.375 123.525 ;
        RECT 145.545 123.275 145.880 123.525 ;
        RECT 146.075 123.275 146.405 123.525 ;
        RECT 143.280 123.025 143.450 123.195 ;
        RECT 145.125 123.105 145.375 123.195 ;
        RECT 142.225 122.285 142.625 122.795 ;
        RECT 142.835 122.615 143.110 122.960 ;
        RECT 143.280 122.855 144.945 123.025 ;
        RECT 143.300 122.285 143.675 122.685 ;
        RECT 143.845 122.505 144.015 122.855 ;
        RECT 144.185 122.285 144.515 122.685 ;
        RECT 144.685 122.455 144.945 122.855 ;
        RECT 145.125 122.685 145.455 123.105 ;
        RECT 145.625 122.285 145.885 123.105 ;
        RECT 146.095 122.285 146.325 123.105 ;
        RECT 146.575 123.085 146.825 123.685 ;
        RECT 147.895 123.645 148.110 123.695 ;
        RECT 146.495 122.455 146.825 123.085 ;
        RECT 146.995 122.285 147.205 123.105 ;
        RECT 147.895 123.065 148.065 123.645 ;
        RECT 148.795 123.525 148.985 123.730 ;
        RECT 149.860 123.525 150.030 124.365 ;
        RECT 150.970 124.335 151.220 124.665 ;
        RECT 148.235 123.195 148.985 123.525 ;
        RECT 149.155 123.195 150.030 123.525 ;
        RECT 147.895 123.025 148.120 123.065 ;
        RECT 148.785 123.025 148.985 123.195 ;
        RECT 147.895 122.940 148.275 123.025 ;
        RECT 147.945 122.505 148.275 122.940 ;
        RECT 148.445 122.285 148.615 122.895 ;
        RECT 148.785 122.500 149.115 123.025 ;
        RECT 149.375 122.285 149.585 122.815 ;
        RECT 149.860 122.735 150.030 123.195 ;
        RECT 150.200 123.235 150.520 124.195 ;
        RECT 150.690 123.445 150.880 124.165 ;
        RECT 151.050 123.265 151.220 124.335 ;
        RECT 151.390 124.035 151.560 124.835 ;
        RECT 151.730 124.390 152.835 124.560 ;
        RECT 151.730 123.775 151.900 124.390 ;
        RECT 153.045 124.240 153.295 124.665 ;
        RECT 153.465 124.375 153.730 124.835 ;
        RECT 152.070 123.855 152.600 124.220 ;
        RECT 153.045 124.110 153.350 124.240 ;
        RECT 151.390 123.685 151.900 123.775 ;
        RECT 151.390 123.515 152.260 123.685 ;
        RECT 151.390 123.445 151.560 123.515 ;
        RECT 151.680 123.265 151.880 123.295 ;
        RECT 150.200 122.905 150.665 123.235 ;
        RECT 151.050 122.965 151.880 123.265 ;
        RECT 151.050 122.735 151.220 122.965 ;
        RECT 149.860 122.565 150.645 122.735 ;
        RECT 150.815 122.565 151.220 122.735 ;
        RECT 151.400 122.285 151.770 122.785 ;
        RECT 152.090 122.735 152.260 123.515 ;
        RECT 152.430 123.155 152.600 123.855 ;
        RECT 152.770 123.325 153.010 123.920 ;
        RECT 152.430 122.935 152.955 123.155 ;
        RECT 153.180 123.005 153.350 124.110 ;
        RECT 153.125 122.875 153.350 123.005 ;
        RECT 153.520 122.915 153.800 123.865 ;
        RECT 153.125 122.735 153.295 122.875 ;
        RECT 152.090 122.565 152.765 122.735 ;
        RECT 152.960 122.565 153.295 122.735 ;
        RECT 153.465 122.285 153.715 122.745 ;
        RECT 153.970 122.545 154.155 124.665 ;
        RECT 154.325 124.335 154.655 124.835 ;
        RECT 154.825 124.165 154.995 124.665 ;
        RECT 154.330 123.995 154.995 124.165 ;
        RECT 154.330 123.005 154.560 123.995 ;
        RECT 154.730 123.175 155.080 123.825 ;
        RECT 155.715 123.745 156.925 124.835 ;
        RECT 155.715 123.205 156.235 123.745 ;
        RECT 156.405 123.035 156.925 123.575 ;
        RECT 154.330 122.835 154.995 123.005 ;
        RECT 154.325 122.285 154.655 122.665 ;
        RECT 154.825 122.545 154.995 122.835 ;
        RECT 155.715 122.285 156.925 123.035 ;
        RECT 22.690 122.115 157.010 122.285 ;
        RECT 22.775 121.365 23.985 122.115 ;
        RECT 24.205 121.460 24.535 121.895 ;
        RECT 24.705 121.505 24.875 122.115 ;
        RECT 24.155 121.375 24.535 121.460 ;
        RECT 25.045 121.375 25.375 121.900 ;
        RECT 25.635 121.585 25.845 122.115 ;
        RECT 26.120 121.665 26.905 121.835 ;
        RECT 27.075 121.665 27.480 121.835 ;
        RECT 22.775 120.825 23.295 121.365 ;
        RECT 24.155 121.335 24.380 121.375 ;
        RECT 23.465 120.655 23.985 121.195 ;
        RECT 22.775 119.565 23.985 120.655 ;
        RECT 24.155 120.755 24.325 121.335 ;
        RECT 25.045 121.205 25.245 121.375 ;
        RECT 26.120 121.205 26.290 121.665 ;
        RECT 24.495 120.875 25.245 121.205 ;
        RECT 25.415 120.875 26.290 121.205 ;
        RECT 24.155 120.705 24.370 120.755 ;
        RECT 24.155 120.625 24.545 120.705 ;
        RECT 24.215 119.780 24.545 120.625 ;
        RECT 25.055 120.670 25.245 120.875 ;
        RECT 24.715 119.565 24.885 120.575 ;
        RECT 25.055 120.295 25.950 120.670 ;
        RECT 25.055 119.735 25.395 120.295 ;
        RECT 25.625 119.565 25.940 120.065 ;
        RECT 26.120 120.035 26.290 120.875 ;
        RECT 26.460 121.165 26.925 121.495 ;
        RECT 27.310 121.435 27.480 121.665 ;
        RECT 27.660 121.615 28.030 122.115 ;
        RECT 28.350 121.665 29.025 121.835 ;
        RECT 29.220 121.665 29.555 121.835 ;
        RECT 26.460 120.205 26.780 121.165 ;
        RECT 27.310 121.135 28.140 121.435 ;
        RECT 26.950 120.235 27.140 120.955 ;
        RECT 27.310 120.065 27.480 121.135 ;
        RECT 27.940 121.105 28.140 121.135 ;
        RECT 27.650 120.885 27.820 120.955 ;
        RECT 28.350 120.885 28.520 121.665 ;
        RECT 29.385 121.525 29.555 121.665 ;
        RECT 29.725 121.655 29.975 122.115 ;
        RECT 27.650 120.715 28.520 120.885 ;
        RECT 28.690 121.245 29.215 121.465 ;
        RECT 29.385 121.395 29.610 121.525 ;
        RECT 27.650 120.625 28.160 120.715 ;
        RECT 26.120 119.865 27.005 120.035 ;
        RECT 27.230 119.735 27.480 120.065 ;
        RECT 27.650 119.565 27.820 120.365 ;
        RECT 27.990 120.010 28.160 120.625 ;
        RECT 28.690 120.545 28.860 121.245 ;
        RECT 28.330 120.180 28.860 120.545 ;
        RECT 29.030 120.480 29.270 121.075 ;
        RECT 29.440 120.290 29.610 121.395 ;
        RECT 29.780 120.535 30.060 121.485 ;
        RECT 29.305 120.160 29.610 120.290 ;
        RECT 27.990 119.840 29.095 120.010 ;
        RECT 29.305 119.735 29.555 120.160 ;
        RECT 29.725 119.565 29.990 120.025 ;
        RECT 30.230 119.735 30.415 121.855 ;
        RECT 30.585 121.735 30.915 122.115 ;
        RECT 31.085 121.565 31.255 121.855 ;
        RECT 30.590 121.395 31.255 121.565 ;
        RECT 30.590 120.405 30.820 121.395 ;
        RECT 31.720 121.335 32.220 121.945 ;
        RECT 30.990 120.575 31.340 121.225 ;
        RECT 31.515 120.875 31.865 121.125 ;
        RECT 32.050 120.705 32.220 121.335 ;
        RECT 32.850 121.465 33.180 121.945 ;
        RECT 33.350 121.655 33.575 122.115 ;
        RECT 33.745 121.465 34.075 121.945 ;
        RECT 32.850 121.295 34.075 121.465 ;
        RECT 34.265 121.315 34.515 122.115 ;
        RECT 34.685 121.315 35.025 121.945 ;
        RECT 35.200 121.715 35.535 122.115 ;
        RECT 35.705 121.545 35.910 121.945 ;
        RECT 36.120 121.635 36.395 122.115 ;
        RECT 36.605 121.615 36.865 121.945 ;
        RECT 37.045 121.615 37.375 122.115 ;
        RECT 32.390 120.925 32.720 121.125 ;
        RECT 32.890 120.925 33.220 121.125 ;
        RECT 33.390 120.925 33.810 121.125 ;
        RECT 33.985 120.955 34.680 121.125 ;
        RECT 33.985 120.705 34.155 120.955 ;
        RECT 34.850 120.705 35.025 121.315 ;
        RECT 31.720 120.535 34.155 120.705 ;
        RECT 30.590 120.235 31.255 120.405 ;
        RECT 30.585 119.565 30.915 120.065 ;
        RECT 31.085 119.735 31.255 120.235 ;
        RECT 31.720 119.735 32.050 120.535 ;
        RECT 32.220 119.565 32.550 120.365 ;
        RECT 32.850 119.735 33.180 120.535 ;
        RECT 33.825 119.565 34.075 120.365 ;
        RECT 34.345 119.565 34.515 120.705 ;
        RECT 34.685 119.735 35.025 120.705 ;
        RECT 35.225 121.375 35.910 121.545 ;
        RECT 35.225 120.345 35.565 121.375 ;
        RECT 35.735 120.705 35.985 121.205 ;
        RECT 36.165 120.875 36.525 121.455 ;
        RECT 36.695 120.705 36.865 121.615 ;
        RECT 37.575 121.545 37.745 121.895 ;
        RECT 37.945 121.715 38.275 122.115 ;
        RECT 38.445 121.545 38.615 121.895 ;
        RECT 38.785 121.715 39.165 122.115 ;
        RECT 37.040 120.875 37.390 121.445 ;
        RECT 37.575 121.375 39.185 121.545 ;
        RECT 39.355 121.440 39.625 121.785 ;
        RECT 39.015 121.205 39.185 121.375 ;
        RECT 35.735 120.535 36.865 120.705 ;
        RECT 35.225 120.170 35.890 120.345 ;
        RECT 35.200 119.565 35.535 119.990 ;
        RECT 35.705 119.765 35.890 120.170 ;
        RECT 36.095 119.565 36.425 120.345 ;
        RECT 36.595 119.765 36.865 120.535 ;
        RECT 37.040 120.415 37.360 120.705 ;
        RECT 37.560 120.585 38.270 121.205 ;
        RECT 38.440 120.875 38.845 121.205 ;
        RECT 39.015 120.875 39.285 121.205 ;
        RECT 39.015 120.705 39.185 120.875 ;
        RECT 39.455 120.705 39.625 121.440 ;
        RECT 38.460 120.535 39.185 120.705 ;
        RECT 38.460 120.415 38.630 120.535 ;
        RECT 37.040 120.245 38.630 120.415 ;
        RECT 37.040 119.785 38.695 120.075 ;
        RECT 38.865 119.565 39.145 120.365 ;
        RECT 39.355 119.735 39.625 120.705 ;
        RECT 39.795 121.375 40.235 121.935 ;
        RECT 40.405 121.375 40.855 122.115 ;
        RECT 41.025 121.545 41.195 121.945 ;
        RECT 41.365 121.715 41.785 122.115 ;
        RECT 41.955 121.545 42.185 121.945 ;
        RECT 41.025 121.375 42.185 121.545 ;
        RECT 42.355 121.375 42.845 121.945 ;
        RECT 39.795 120.365 40.105 121.375 ;
        RECT 40.275 120.755 40.445 121.205 ;
        RECT 40.615 120.925 41.005 121.205 ;
        RECT 41.190 120.875 41.435 121.205 ;
        RECT 40.275 120.585 41.065 120.755 ;
        RECT 39.795 119.735 40.235 120.365 ;
        RECT 40.410 119.565 40.725 120.415 ;
        RECT 40.895 119.905 41.065 120.585 ;
        RECT 41.235 120.075 41.435 120.875 ;
        RECT 41.635 120.075 41.885 121.205 ;
        RECT 42.100 120.875 42.505 121.205 ;
        RECT 42.675 120.705 42.845 121.375 ;
        RECT 43.290 121.305 43.535 121.910 ;
        RECT 43.755 121.580 44.265 122.115 ;
        RECT 42.075 120.535 42.845 120.705 ;
        RECT 43.015 121.135 44.245 121.305 ;
        RECT 42.075 119.905 42.325 120.535 ;
        RECT 40.895 119.735 42.325 119.905 ;
        RECT 42.505 119.565 42.835 120.365 ;
        RECT 43.015 120.325 43.355 121.135 ;
        RECT 43.525 120.570 44.275 120.760 ;
        RECT 43.015 119.915 43.530 120.325 ;
        RECT 43.765 119.565 43.935 120.325 ;
        RECT 44.105 119.905 44.275 120.570 ;
        RECT 44.445 120.585 44.635 121.945 ;
        RECT 44.805 121.435 45.080 121.945 ;
        RECT 45.270 121.580 45.800 121.945 ;
        RECT 46.225 121.715 46.555 122.115 ;
        RECT 45.625 121.545 45.800 121.580 ;
        RECT 44.805 121.265 45.085 121.435 ;
        RECT 44.805 120.785 45.080 121.265 ;
        RECT 45.285 120.585 45.455 121.385 ;
        RECT 44.445 120.415 45.455 120.585 ;
        RECT 45.625 121.375 46.555 121.545 ;
        RECT 46.725 121.375 46.980 121.945 ;
        RECT 45.625 120.245 45.795 121.375 ;
        RECT 46.385 121.205 46.555 121.375 ;
        RECT 44.670 120.075 45.795 120.245 ;
        RECT 45.965 120.875 46.160 121.205 ;
        RECT 46.385 120.875 46.640 121.205 ;
        RECT 45.965 119.905 46.135 120.875 ;
        RECT 46.810 120.705 46.980 121.375 ;
        RECT 47.155 121.365 48.365 122.115 ;
        RECT 48.535 121.390 48.825 122.115 ;
        RECT 49.545 121.565 49.715 121.855 ;
        RECT 49.885 121.735 50.215 122.115 ;
        RECT 49.545 121.395 50.210 121.565 ;
        RECT 47.155 120.825 47.675 121.365 ;
        RECT 44.105 119.735 46.135 119.905 ;
        RECT 46.305 119.565 46.475 120.705 ;
        RECT 46.645 119.735 46.980 120.705 ;
        RECT 47.845 120.655 48.365 121.195 ;
        RECT 47.155 119.565 48.365 120.655 ;
        RECT 48.535 119.565 48.825 120.730 ;
        RECT 49.460 120.575 49.810 121.225 ;
        RECT 49.980 120.405 50.210 121.395 ;
        RECT 49.545 120.235 50.210 120.405 ;
        RECT 49.545 119.735 49.715 120.235 ;
        RECT 49.885 119.565 50.215 120.065 ;
        RECT 50.385 119.735 50.570 121.855 ;
        RECT 50.825 121.655 51.075 122.115 ;
        RECT 51.245 121.665 51.580 121.835 ;
        RECT 51.775 121.665 52.450 121.835 ;
        RECT 51.245 121.525 51.415 121.665 ;
        RECT 50.740 120.535 51.020 121.485 ;
        RECT 51.190 121.395 51.415 121.525 ;
        RECT 51.190 120.290 51.360 121.395 ;
        RECT 51.585 121.245 52.110 121.465 ;
        RECT 51.530 120.480 51.770 121.075 ;
        RECT 51.940 120.545 52.110 121.245 ;
        RECT 52.280 120.885 52.450 121.665 ;
        RECT 52.770 121.615 53.140 122.115 ;
        RECT 53.320 121.665 53.725 121.835 ;
        RECT 53.895 121.665 54.680 121.835 ;
        RECT 53.320 121.435 53.490 121.665 ;
        RECT 52.660 121.135 53.490 121.435 ;
        RECT 53.875 121.165 54.340 121.495 ;
        RECT 52.660 121.105 52.860 121.135 ;
        RECT 52.980 120.885 53.150 120.955 ;
        RECT 52.280 120.715 53.150 120.885 ;
        RECT 52.640 120.625 53.150 120.715 ;
        RECT 51.190 120.160 51.495 120.290 ;
        RECT 51.940 120.180 52.470 120.545 ;
        RECT 50.810 119.565 51.075 120.025 ;
        RECT 51.245 119.735 51.495 120.160 ;
        RECT 52.640 120.010 52.810 120.625 ;
        RECT 51.705 119.840 52.810 120.010 ;
        RECT 52.980 119.565 53.150 120.365 ;
        RECT 53.320 120.065 53.490 121.135 ;
        RECT 53.660 120.235 53.850 120.955 ;
        RECT 54.020 120.205 54.340 121.165 ;
        RECT 54.510 121.205 54.680 121.665 ;
        RECT 54.955 121.585 55.165 122.115 ;
        RECT 55.425 121.375 55.755 121.900 ;
        RECT 55.925 121.505 56.095 122.115 ;
        RECT 56.265 121.460 56.595 121.895 ;
        RECT 56.265 121.375 56.645 121.460 ;
        RECT 55.555 121.205 55.755 121.375 ;
        RECT 56.420 121.335 56.645 121.375 ;
        RECT 54.510 120.875 55.385 121.205 ;
        RECT 55.555 120.875 56.305 121.205 ;
        RECT 53.320 119.735 53.570 120.065 ;
        RECT 54.510 120.035 54.680 120.875 ;
        RECT 55.555 120.670 55.745 120.875 ;
        RECT 56.475 120.755 56.645 121.335 ;
        RECT 56.430 120.705 56.645 120.755 ;
        RECT 54.850 120.295 55.745 120.670 ;
        RECT 56.255 120.625 56.645 120.705 ;
        RECT 56.815 121.375 57.200 121.945 ;
        RECT 57.370 121.655 57.695 122.115 ;
        RECT 58.215 121.485 58.495 121.945 ;
        RECT 56.815 120.705 57.095 121.375 ;
        RECT 57.370 121.315 58.495 121.485 ;
        RECT 57.370 121.205 57.820 121.315 ;
        RECT 57.265 120.875 57.820 121.205 ;
        RECT 58.685 121.145 59.085 121.945 ;
        RECT 59.485 121.655 59.755 122.115 ;
        RECT 59.925 121.485 60.210 121.945 ;
        RECT 53.795 119.865 54.680 120.035 ;
        RECT 54.860 119.565 55.175 120.065 ;
        RECT 55.405 119.735 55.745 120.295 ;
        RECT 55.915 119.565 56.085 120.575 ;
        RECT 56.255 119.780 56.585 120.625 ;
        RECT 56.815 119.735 57.200 120.705 ;
        RECT 57.370 120.415 57.820 120.875 ;
        RECT 57.990 120.585 59.085 121.145 ;
        RECT 57.370 120.195 58.495 120.415 ;
        RECT 57.370 119.565 57.695 120.025 ;
        RECT 58.215 119.735 58.495 120.195 ;
        RECT 58.685 119.735 59.085 120.585 ;
        RECT 59.255 121.315 60.210 121.485 ;
        RECT 60.495 121.375 60.960 121.920 ;
        RECT 59.255 120.415 59.465 121.315 ;
        RECT 59.635 120.585 60.325 121.145 ;
        RECT 60.495 120.415 60.665 121.375 ;
        RECT 61.465 121.295 61.635 122.115 ;
        RECT 61.805 121.465 62.135 121.945 ;
        RECT 62.305 121.725 62.655 122.115 ;
        RECT 62.825 121.545 63.055 121.945 ;
        RECT 62.545 121.465 63.055 121.545 ;
        RECT 61.805 121.375 63.055 121.465 ;
        RECT 63.225 121.375 63.545 121.855 ;
        RECT 61.805 121.295 62.715 121.375 ;
        RECT 60.835 120.755 61.080 121.205 ;
        RECT 61.340 120.925 62.035 121.125 ;
        RECT 62.205 120.955 62.805 121.125 ;
        RECT 62.205 120.755 62.375 120.955 ;
        RECT 63.035 120.785 63.205 121.205 ;
        RECT 60.835 120.585 62.375 120.755 ;
        RECT 62.545 120.615 63.205 120.785 ;
        RECT 62.545 120.415 62.715 120.615 ;
        RECT 63.375 120.445 63.545 121.375 ;
        RECT 63.715 121.345 66.305 122.115 ;
        RECT 66.985 121.460 67.315 121.895 ;
        RECT 67.485 121.505 67.655 122.115 ;
        RECT 66.935 121.375 67.315 121.460 ;
        RECT 67.825 121.375 68.155 121.900 ;
        RECT 68.415 121.585 68.625 122.115 ;
        RECT 68.900 121.665 69.685 121.835 ;
        RECT 69.855 121.665 70.260 121.835 ;
        RECT 63.715 120.825 64.925 121.345 ;
        RECT 66.935 121.335 67.160 121.375 ;
        RECT 65.095 120.655 66.305 121.175 ;
        RECT 59.255 120.195 60.210 120.415 ;
        RECT 60.495 120.245 62.715 120.415 ;
        RECT 62.885 120.245 63.545 120.445 ;
        RECT 59.485 119.565 59.755 120.025 ;
        RECT 59.925 119.735 60.210 120.195 ;
        RECT 60.495 119.565 60.795 120.075 ;
        RECT 60.965 119.735 61.295 120.245 ;
        RECT 62.885 120.075 63.055 120.245 ;
        RECT 61.465 119.565 62.095 120.075 ;
        RECT 62.675 119.905 63.055 120.075 ;
        RECT 63.225 119.565 63.525 120.075 ;
        RECT 63.715 119.565 66.305 120.655 ;
        RECT 66.935 120.755 67.105 121.335 ;
        RECT 67.825 121.205 68.025 121.375 ;
        RECT 68.900 121.205 69.070 121.665 ;
        RECT 67.275 120.875 68.025 121.205 ;
        RECT 68.195 120.875 69.070 121.205 ;
        RECT 66.935 120.705 67.150 120.755 ;
        RECT 66.935 120.625 67.325 120.705 ;
        RECT 66.995 119.780 67.325 120.625 ;
        RECT 67.835 120.670 68.025 120.875 ;
        RECT 67.495 119.565 67.665 120.575 ;
        RECT 67.835 120.295 68.730 120.670 ;
        RECT 67.835 119.735 68.175 120.295 ;
        RECT 68.405 119.565 68.720 120.065 ;
        RECT 68.900 120.035 69.070 120.875 ;
        RECT 69.240 121.165 69.705 121.495 ;
        RECT 70.090 121.435 70.260 121.665 ;
        RECT 70.440 121.615 70.810 122.115 ;
        RECT 71.130 121.665 71.805 121.835 ;
        RECT 72.000 121.665 72.335 121.835 ;
        RECT 69.240 120.205 69.560 121.165 ;
        RECT 70.090 121.135 70.920 121.435 ;
        RECT 69.730 120.235 69.920 120.955 ;
        RECT 70.090 120.065 70.260 121.135 ;
        RECT 70.720 121.105 70.920 121.135 ;
        RECT 70.430 120.885 70.600 120.955 ;
        RECT 71.130 120.885 71.300 121.665 ;
        RECT 72.165 121.525 72.335 121.665 ;
        RECT 72.505 121.655 72.755 122.115 ;
        RECT 70.430 120.715 71.300 120.885 ;
        RECT 71.470 121.245 71.995 121.465 ;
        RECT 72.165 121.395 72.390 121.525 ;
        RECT 70.430 120.625 70.940 120.715 ;
        RECT 68.900 119.865 69.785 120.035 ;
        RECT 70.010 119.735 70.260 120.065 ;
        RECT 70.430 119.565 70.600 120.365 ;
        RECT 70.770 120.010 70.940 120.625 ;
        RECT 71.470 120.545 71.640 121.245 ;
        RECT 71.110 120.180 71.640 120.545 ;
        RECT 71.810 120.480 72.050 121.075 ;
        RECT 72.220 120.290 72.390 121.395 ;
        RECT 72.560 120.535 72.840 121.485 ;
        RECT 72.085 120.160 72.390 120.290 ;
        RECT 70.770 119.840 71.875 120.010 ;
        RECT 72.085 119.735 72.335 120.160 ;
        RECT 72.505 119.565 72.770 120.025 ;
        RECT 73.010 119.735 73.195 121.855 ;
        RECT 73.365 121.735 73.695 122.115 ;
        RECT 73.865 121.565 74.035 121.855 ;
        RECT 73.370 121.395 74.035 121.565 ;
        RECT 73.370 120.405 73.600 121.395 ;
        RECT 74.295 121.390 74.585 122.115 ;
        RECT 74.755 121.375 75.140 121.945 ;
        RECT 75.310 121.655 75.635 122.115 ;
        RECT 76.155 121.485 76.435 121.945 ;
        RECT 73.770 120.575 74.120 121.225 ;
        RECT 73.370 120.235 74.035 120.405 ;
        RECT 73.365 119.565 73.695 120.065 ;
        RECT 73.865 119.735 74.035 120.235 ;
        RECT 74.295 119.565 74.585 120.730 ;
        RECT 74.755 120.705 75.035 121.375 ;
        RECT 75.310 121.315 76.435 121.485 ;
        RECT 75.310 121.205 75.760 121.315 ;
        RECT 75.205 120.875 75.760 121.205 ;
        RECT 76.625 121.145 77.025 121.945 ;
        RECT 77.425 121.655 77.695 122.115 ;
        RECT 77.865 121.485 78.150 121.945 ;
        RECT 74.755 119.735 75.140 120.705 ;
        RECT 75.310 120.415 75.760 120.875 ;
        RECT 75.930 120.585 77.025 121.145 ;
        RECT 75.310 120.195 76.435 120.415 ;
        RECT 75.310 119.565 75.635 120.025 ;
        RECT 76.155 119.735 76.435 120.195 ;
        RECT 76.625 119.735 77.025 120.585 ;
        RECT 77.195 121.315 78.150 121.485 ;
        RECT 77.195 120.415 77.405 121.315 ;
        RECT 77.575 120.585 78.265 121.145 ;
        RECT 77.195 120.195 78.150 120.415 ;
        RECT 77.425 119.565 77.695 120.025 ;
        RECT 77.865 119.735 78.150 120.195 ;
        RECT 78.445 119.745 78.705 121.935 ;
        RECT 78.965 121.745 79.635 122.115 ;
        RECT 79.815 121.565 80.125 121.935 ;
        RECT 78.895 121.365 80.125 121.565 ;
        RECT 78.895 120.695 79.185 121.365 ;
        RECT 80.305 121.185 80.535 121.825 ;
        RECT 80.715 121.385 81.005 122.115 ;
        RECT 81.195 121.440 81.455 121.945 ;
        RECT 81.635 121.735 81.965 122.115 ;
        RECT 82.145 121.565 82.315 121.945 ;
        RECT 79.365 120.875 79.830 121.185 ;
        RECT 80.010 120.875 80.535 121.185 ;
        RECT 80.715 120.875 81.015 121.205 ;
        RECT 78.895 120.475 79.665 120.695 ;
        RECT 78.875 119.565 79.215 120.295 ;
        RECT 79.395 119.745 79.665 120.475 ;
        RECT 79.845 120.455 81.005 120.695 ;
        RECT 79.845 119.745 80.075 120.455 ;
        RECT 80.245 119.565 80.575 120.275 ;
        RECT 80.745 119.745 81.005 120.455 ;
        RECT 81.195 120.640 81.365 121.440 ;
        RECT 81.650 121.395 82.315 121.565 ;
        RECT 82.665 121.565 82.835 121.855 ;
        RECT 83.005 121.735 83.335 122.115 ;
        RECT 82.665 121.395 83.330 121.565 ;
        RECT 81.650 121.140 81.820 121.395 ;
        RECT 81.535 120.810 81.820 121.140 ;
        RECT 82.055 120.845 82.385 121.215 ;
        RECT 81.650 120.665 81.820 120.810 ;
        RECT 81.195 119.735 81.465 120.640 ;
        RECT 81.650 120.495 82.315 120.665 ;
        RECT 82.580 120.575 82.930 121.225 ;
        RECT 81.635 119.565 81.965 120.325 ;
        RECT 82.145 119.735 82.315 120.495 ;
        RECT 83.100 120.405 83.330 121.395 ;
        RECT 82.665 120.235 83.330 120.405 ;
        RECT 82.665 119.735 82.835 120.235 ;
        RECT 83.005 119.565 83.335 120.065 ;
        RECT 83.505 119.735 83.690 121.855 ;
        RECT 83.945 121.655 84.195 122.115 ;
        RECT 84.365 121.665 84.700 121.835 ;
        RECT 84.895 121.665 85.570 121.835 ;
        RECT 84.365 121.525 84.535 121.665 ;
        RECT 83.860 120.535 84.140 121.485 ;
        RECT 84.310 121.395 84.535 121.525 ;
        RECT 84.310 120.290 84.480 121.395 ;
        RECT 84.705 121.245 85.230 121.465 ;
        RECT 84.650 120.480 84.890 121.075 ;
        RECT 85.060 120.545 85.230 121.245 ;
        RECT 85.400 120.885 85.570 121.665 ;
        RECT 85.890 121.615 86.260 122.115 ;
        RECT 86.440 121.665 86.845 121.835 ;
        RECT 87.015 121.665 87.800 121.835 ;
        RECT 86.440 121.435 86.610 121.665 ;
        RECT 85.780 121.135 86.610 121.435 ;
        RECT 86.995 121.165 87.460 121.495 ;
        RECT 85.780 121.105 85.980 121.135 ;
        RECT 86.100 120.885 86.270 120.955 ;
        RECT 85.400 120.715 86.270 120.885 ;
        RECT 85.760 120.625 86.270 120.715 ;
        RECT 84.310 120.160 84.615 120.290 ;
        RECT 85.060 120.180 85.590 120.545 ;
        RECT 83.930 119.565 84.195 120.025 ;
        RECT 84.365 119.735 84.615 120.160 ;
        RECT 85.760 120.010 85.930 120.625 ;
        RECT 84.825 119.840 85.930 120.010 ;
        RECT 86.100 119.565 86.270 120.365 ;
        RECT 86.440 120.065 86.610 121.135 ;
        RECT 86.780 120.235 86.970 120.955 ;
        RECT 87.140 120.205 87.460 121.165 ;
        RECT 87.630 121.205 87.800 121.665 ;
        RECT 88.075 121.585 88.285 122.115 ;
        RECT 88.545 121.375 88.875 121.900 ;
        RECT 89.045 121.505 89.215 122.115 ;
        RECT 89.385 121.460 89.715 121.895 ;
        RECT 90.025 121.565 90.195 121.855 ;
        RECT 90.365 121.735 90.695 122.115 ;
        RECT 89.385 121.375 89.765 121.460 ;
        RECT 90.025 121.395 90.690 121.565 ;
        RECT 88.675 121.205 88.875 121.375 ;
        RECT 89.540 121.335 89.765 121.375 ;
        RECT 87.630 120.875 88.505 121.205 ;
        RECT 88.675 120.875 89.425 121.205 ;
        RECT 86.440 119.735 86.690 120.065 ;
        RECT 87.630 120.035 87.800 120.875 ;
        RECT 88.675 120.670 88.865 120.875 ;
        RECT 89.595 120.755 89.765 121.335 ;
        RECT 89.550 120.705 89.765 120.755 ;
        RECT 87.970 120.295 88.865 120.670 ;
        RECT 89.375 120.625 89.765 120.705 ;
        RECT 86.915 119.865 87.800 120.035 ;
        RECT 87.980 119.565 88.295 120.065 ;
        RECT 88.525 119.735 88.865 120.295 ;
        RECT 89.035 119.565 89.205 120.575 ;
        RECT 89.375 119.780 89.705 120.625 ;
        RECT 89.940 120.575 90.290 121.225 ;
        RECT 90.460 120.405 90.690 121.395 ;
        RECT 90.025 120.235 90.690 120.405 ;
        RECT 90.025 119.735 90.195 120.235 ;
        RECT 90.365 119.565 90.695 120.065 ;
        RECT 90.865 119.735 91.050 121.855 ;
        RECT 91.305 121.655 91.555 122.115 ;
        RECT 91.725 121.665 92.060 121.835 ;
        RECT 92.255 121.665 92.930 121.835 ;
        RECT 91.725 121.525 91.895 121.665 ;
        RECT 91.220 120.535 91.500 121.485 ;
        RECT 91.670 121.395 91.895 121.525 ;
        RECT 91.670 120.290 91.840 121.395 ;
        RECT 92.065 121.245 92.590 121.465 ;
        RECT 92.010 120.480 92.250 121.075 ;
        RECT 92.420 120.545 92.590 121.245 ;
        RECT 92.760 120.885 92.930 121.665 ;
        RECT 93.250 121.615 93.620 122.115 ;
        RECT 93.800 121.665 94.205 121.835 ;
        RECT 94.375 121.665 95.160 121.835 ;
        RECT 93.800 121.435 93.970 121.665 ;
        RECT 93.140 121.135 93.970 121.435 ;
        RECT 94.355 121.165 94.820 121.495 ;
        RECT 93.140 121.105 93.340 121.135 ;
        RECT 93.460 120.885 93.630 120.955 ;
        RECT 92.760 120.715 93.630 120.885 ;
        RECT 93.120 120.625 93.630 120.715 ;
        RECT 91.670 120.160 91.975 120.290 ;
        RECT 92.420 120.180 92.950 120.545 ;
        RECT 91.290 119.565 91.555 120.025 ;
        RECT 91.725 119.735 91.975 120.160 ;
        RECT 93.120 120.010 93.290 120.625 ;
        RECT 92.185 119.840 93.290 120.010 ;
        RECT 93.460 119.565 93.630 120.365 ;
        RECT 93.800 120.065 93.970 121.135 ;
        RECT 94.140 120.235 94.330 120.955 ;
        RECT 94.500 120.205 94.820 121.165 ;
        RECT 94.990 121.205 95.160 121.665 ;
        RECT 95.435 121.585 95.645 122.115 ;
        RECT 95.905 121.375 96.235 121.900 ;
        RECT 96.405 121.505 96.575 122.115 ;
        RECT 96.745 121.460 97.075 121.895 ;
        RECT 97.245 121.600 97.415 122.115 ;
        RECT 96.745 121.375 97.125 121.460 ;
        RECT 96.035 121.205 96.235 121.375 ;
        RECT 96.900 121.335 97.125 121.375 ;
        RECT 94.990 120.875 95.865 121.205 ;
        RECT 96.035 120.875 96.785 121.205 ;
        RECT 93.800 119.735 94.050 120.065 ;
        RECT 94.990 120.035 95.160 120.875 ;
        RECT 96.035 120.670 96.225 120.875 ;
        RECT 96.955 120.755 97.125 121.335 ;
        RECT 97.755 121.345 99.425 122.115 ;
        RECT 100.055 121.390 100.345 122.115 ;
        RECT 100.520 121.375 100.775 121.945 ;
        RECT 100.945 121.715 101.275 122.115 ;
        RECT 101.700 121.580 102.230 121.945 ;
        RECT 102.420 121.775 102.695 121.945 ;
        RECT 102.415 121.605 102.695 121.775 ;
        RECT 101.700 121.545 101.875 121.580 ;
        RECT 100.945 121.375 101.875 121.545 ;
        RECT 97.755 120.825 98.505 121.345 ;
        RECT 96.910 120.705 97.125 120.755 ;
        RECT 95.330 120.295 96.225 120.670 ;
        RECT 96.735 120.625 97.125 120.705 ;
        RECT 98.675 120.655 99.425 121.175 ;
        RECT 94.275 119.865 95.160 120.035 ;
        RECT 95.340 119.565 95.655 120.065 ;
        RECT 95.885 119.735 96.225 120.295 ;
        RECT 96.395 119.565 96.565 120.575 ;
        RECT 96.735 119.780 97.065 120.625 ;
        RECT 97.235 119.565 97.405 120.480 ;
        RECT 97.755 119.565 99.425 120.655 ;
        RECT 100.055 119.565 100.345 120.730 ;
        RECT 100.520 120.705 100.690 121.375 ;
        RECT 100.945 121.205 101.115 121.375 ;
        RECT 100.860 120.875 101.115 121.205 ;
        RECT 101.340 120.875 101.535 121.205 ;
        RECT 100.520 119.735 100.855 120.705 ;
        RECT 101.025 119.565 101.195 120.705 ;
        RECT 101.365 119.905 101.535 120.875 ;
        RECT 101.705 120.245 101.875 121.375 ;
        RECT 102.045 120.585 102.215 121.385 ;
        RECT 102.420 120.785 102.695 121.605 ;
        RECT 102.865 120.585 103.055 121.945 ;
        RECT 103.235 121.580 103.745 122.115 ;
        RECT 103.965 121.305 104.210 121.910 ;
        RECT 105.205 121.565 105.375 121.855 ;
        RECT 105.545 121.735 105.875 122.115 ;
        RECT 105.205 121.395 105.870 121.565 ;
        RECT 103.255 121.135 104.485 121.305 ;
        RECT 102.045 120.415 103.055 120.585 ;
        RECT 103.225 120.570 103.975 120.760 ;
        RECT 101.705 120.075 102.830 120.245 ;
        RECT 103.225 119.905 103.395 120.570 ;
        RECT 104.145 120.325 104.485 121.135 ;
        RECT 105.120 120.575 105.470 121.225 ;
        RECT 105.640 120.405 105.870 121.395 ;
        RECT 101.365 119.735 103.395 119.905 ;
        RECT 103.565 119.565 103.735 120.325 ;
        RECT 103.970 119.915 104.485 120.325 ;
        RECT 105.205 120.235 105.870 120.405 ;
        RECT 105.205 119.735 105.375 120.235 ;
        RECT 105.545 119.565 105.875 120.065 ;
        RECT 106.045 119.735 106.230 121.855 ;
        RECT 106.485 121.655 106.735 122.115 ;
        RECT 106.905 121.665 107.240 121.835 ;
        RECT 107.435 121.665 108.110 121.835 ;
        RECT 106.905 121.525 107.075 121.665 ;
        RECT 106.400 120.535 106.680 121.485 ;
        RECT 106.850 121.395 107.075 121.525 ;
        RECT 106.850 120.290 107.020 121.395 ;
        RECT 107.245 121.245 107.770 121.465 ;
        RECT 107.190 120.480 107.430 121.075 ;
        RECT 107.600 120.545 107.770 121.245 ;
        RECT 107.940 120.885 108.110 121.665 ;
        RECT 108.430 121.615 108.800 122.115 ;
        RECT 108.980 121.665 109.385 121.835 ;
        RECT 109.555 121.665 110.340 121.835 ;
        RECT 108.980 121.435 109.150 121.665 ;
        RECT 108.320 121.135 109.150 121.435 ;
        RECT 109.535 121.165 110.000 121.495 ;
        RECT 108.320 121.105 108.520 121.135 ;
        RECT 108.640 120.885 108.810 120.955 ;
        RECT 107.940 120.715 108.810 120.885 ;
        RECT 108.300 120.625 108.810 120.715 ;
        RECT 106.850 120.160 107.155 120.290 ;
        RECT 107.600 120.180 108.130 120.545 ;
        RECT 106.470 119.565 106.735 120.025 ;
        RECT 106.905 119.735 107.155 120.160 ;
        RECT 108.300 120.010 108.470 120.625 ;
        RECT 107.365 119.840 108.470 120.010 ;
        RECT 108.640 119.565 108.810 120.365 ;
        RECT 108.980 120.065 109.150 121.135 ;
        RECT 109.320 120.235 109.510 120.955 ;
        RECT 109.680 120.205 110.000 121.165 ;
        RECT 110.170 121.205 110.340 121.665 ;
        RECT 110.615 121.585 110.825 122.115 ;
        RECT 111.085 121.375 111.415 121.900 ;
        RECT 111.585 121.505 111.755 122.115 ;
        RECT 111.925 121.460 112.255 121.895 ;
        RECT 111.925 121.375 112.305 121.460 ;
        RECT 111.215 121.205 111.415 121.375 ;
        RECT 112.080 121.335 112.305 121.375 ;
        RECT 110.170 120.875 111.045 121.205 ;
        RECT 111.215 120.875 111.965 121.205 ;
        RECT 108.980 119.735 109.230 120.065 ;
        RECT 110.170 120.035 110.340 120.875 ;
        RECT 111.215 120.670 111.405 120.875 ;
        RECT 112.135 120.755 112.305 121.335 ;
        RECT 112.475 121.365 113.685 122.115 ;
        RECT 113.905 121.460 114.235 121.895 ;
        RECT 114.405 121.505 114.575 122.115 ;
        RECT 113.855 121.375 114.235 121.460 ;
        RECT 114.745 121.375 115.075 121.900 ;
        RECT 115.335 121.585 115.545 122.115 ;
        RECT 115.820 121.665 116.605 121.835 ;
        RECT 116.775 121.665 117.180 121.835 ;
        RECT 112.475 120.825 112.995 121.365 ;
        RECT 113.855 121.335 114.080 121.375 ;
        RECT 112.090 120.705 112.305 120.755 ;
        RECT 110.510 120.295 111.405 120.670 ;
        RECT 111.915 120.625 112.305 120.705 ;
        RECT 113.165 120.655 113.685 121.195 ;
        RECT 109.455 119.865 110.340 120.035 ;
        RECT 110.520 119.565 110.835 120.065 ;
        RECT 111.065 119.735 111.405 120.295 ;
        RECT 111.575 119.565 111.745 120.575 ;
        RECT 111.915 119.780 112.245 120.625 ;
        RECT 112.475 119.565 113.685 120.655 ;
        RECT 113.855 120.755 114.025 121.335 ;
        RECT 114.745 121.205 114.945 121.375 ;
        RECT 115.820 121.205 115.990 121.665 ;
        RECT 114.195 120.875 114.945 121.205 ;
        RECT 115.115 120.875 115.990 121.205 ;
        RECT 113.855 120.705 114.070 120.755 ;
        RECT 113.855 120.625 114.245 120.705 ;
        RECT 113.915 119.780 114.245 120.625 ;
        RECT 114.755 120.670 114.945 120.875 ;
        RECT 114.415 119.565 114.585 120.575 ;
        RECT 114.755 120.295 115.650 120.670 ;
        RECT 114.755 119.735 115.095 120.295 ;
        RECT 115.325 119.565 115.640 120.065 ;
        RECT 115.820 120.035 115.990 120.875 ;
        RECT 116.160 121.165 116.625 121.495 ;
        RECT 117.010 121.435 117.180 121.665 ;
        RECT 117.360 121.615 117.730 122.115 ;
        RECT 118.050 121.665 118.725 121.835 ;
        RECT 118.920 121.665 119.255 121.835 ;
        RECT 116.160 120.205 116.480 121.165 ;
        RECT 117.010 121.135 117.840 121.435 ;
        RECT 116.650 120.235 116.840 120.955 ;
        RECT 117.010 120.065 117.180 121.135 ;
        RECT 117.640 121.105 117.840 121.135 ;
        RECT 117.350 120.885 117.520 120.955 ;
        RECT 118.050 120.885 118.220 121.665 ;
        RECT 119.085 121.525 119.255 121.665 ;
        RECT 119.425 121.655 119.675 122.115 ;
        RECT 117.350 120.715 118.220 120.885 ;
        RECT 118.390 121.245 118.915 121.465 ;
        RECT 119.085 121.395 119.310 121.525 ;
        RECT 117.350 120.625 117.860 120.715 ;
        RECT 115.820 119.865 116.705 120.035 ;
        RECT 116.930 119.735 117.180 120.065 ;
        RECT 117.350 119.565 117.520 120.365 ;
        RECT 117.690 120.010 117.860 120.625 ;
        RECT 118.390 120.545 118.560 121.245 ;
        RECT 118.030 120.180 118.560 120.545 ;
        RECT 118.730 120.480 118.970 121.075 ;
        RECT 119.140 120.290 119.310 121.395 ;
        RECT 119.480 120.535 119.760 121.485 ;
        RECT 119.005 120.160 119.310 120.290 ;
        RECT 117.690 119.840 118.795 120.010 ;
        RECT 119.005 119.735 119.255 120.160 ;
        RECT 119.425 119.565 119.690 120.025 ;
        RECT 119.930 119.735 120.115 121.855 ;
        RECT 120.285 121.735 120.615 122.115 ;
        RECT 120.785 121.565 120.955 121.855 ;
        RECT 120.290 121.395 120.955 121.565 ;
        RECT 122.135 121.615 122.395 121.945 ;
        RECT 122.565 121.755 122.895 122.115 ;
        RECT 123.150 121.735 124.450 121.945 ;
        RECT 122.135 121.605 122.365 121.615 ;
        RECT 120.290 120.405 120.520 121.395 ;
        RECT 120.690 120.575 121.040 121.225 ;
        RECT 122.135 120.415 122.305 121.605 ;
        RECT 123.150 121.585 123.320 121.735 ;
        RECT 122.565 121.460 123.320 121.585 ;
        RECT 122.475 121.415 123.320 121.460 ;
        RECT 122.475 121.295 122.745 121.415 ;
        RECT 122.475 120.720 122.645 121.295 ;
        RECT 122.875 120.855 123.285 121.160 ;
        RECT 123.575 121.125 123.785 121.525 ;
        RECT 123.455 120.915 123.785 121.125 ;
        RECT 124.030 121.125 124.250 121.525 ;
        RECT 124.725 121.350 125.180 122.115 ;
        RECT 125.815 121.390 126.105 122.115 ;
        RECT 126.365 121.565 126.535 121.855 ;
        RECT 126.705 121.735 127.035 122.115 ;
        RECT 126.365 121.395 127.030 121.565 ;
        RECT 124.030 120.915 124.505 121.125 ;
        RECT 124.695 120.925 125.185 121.125 ;
        RECT 122.475 120.685 122.675 120.720 ;
        RECT 124.005 120.685 125.180 120.745 ;
        RECT 122.475 120.575 125.180 120.685 ;
        RECT 122.535 120.515 124.335 120.575 ;
        RECT 124.005 120.485 124.335 120.515 ;
        RECT 120.290 120.235 120.955 120.405 ;
        RECT 120.285 119.565 120.615 120.065 ;
        RECT 120.785 119.735 120.955 120.235 ;
        RECT 122.135 119.735 122.395 120.415 ;
        RECT 122.565 119.565 122.815 120.345 ;
        RECT 123.065 120.315 123.900 120.325 ;
        RECT 124.490 120.315 124.675 120.405 ;
        RECT 123.065 120.115 124.675 120.315 ;
        RECT 123.065 119.735 123.315 120.115 ;
        RECT 124.445 120.075 124.675 120.115 ;
        RECT 124.925 119.955 125.180 120.575 ;
        RECT 123.485 119.565 123.840 119.945 ;
        RECT 124.845 119.735 125.180 119.955 ;
        RECT 125.815 119.565 126.105 120.730 ;
        RECT 126.280 120.575 126.630 121.225 ;
        RECT 126.800 120.405 127.030 121.395 ;
        RECT 126.365 120.235 127.030 120.405 ;
        RECT 126.365 119.735 126.535 120.235 ;
        RECT 126.705 119.565 127.035 120.065 ;
        RECT 127.205 119.735 127.390 121.855 ;
        RECT 127.645 121.655 127.895 122.115 ;
        RECT 128.065 121.665 128.400 121.835 ;
        RECT 128.595 121.665 129.270 121.835 ;
        RECT 128.065 121.525 128.235 121.665 ;
        RECT 127.560 120.535 127.840 121.485 ;
        RECT 128.010 121.395 128.235 121.525 ;
        RECT 128.010 120.290 128.180 121.395 ;
        RECT 128.405 121.245 128.930 121.465 ;
        RECT 128.350 120.480 128.590 121.075 ;
        RECT 128.760 120.545 128.930 121.245 ;
        RECT 129.100 120.885 129.270 121.665 ;
        RECT 129.590 121.615 129.960 122.115 ;
        RECT 130.140 121.665 130.545 121.835 ;
        RECT 130.715 121.665 131.500 121.835 ;
        RECT 130.140 121.435 130.310 121.665 ;
        RECT 129.480 121.135 130.310 121.435 ;
        RECT 130.695 121.165 131.160 121.495 ;
        RECT 129.480 121.105 129.680 121.135 ;
        RECT 129.800 120.885 129.970 120.955 ;
        RECT 129.100 120.715 129.970 120.885 ;
        RECT 129.460 120.625 129.970 120.715 ;
        RECT 128.010 120.160 128.315 120.290 ;
        RECT 128.760 120.180 129.290 120.545 ;
        RECT 127.630 119.565 127.895 120.025 ;
        RECT 128.065 119.735 128.315 120.160 ;
        RECT 129.460 120.010 129.630 120.625 ;
        RECT 128.525 119.840 129.630 120.010 ;
        RECT 129.800 119.565 129.970 120.365 ;
        RECT 130.140 120.065 130.310 121.135 ;
        RECT 130.480 120.235 130.670 120.955 ;
        RECT 130.840 120.205 131.160 121.165 ;
        RECT 131.330 121.205 131.500 121.665 ;
        RECT 131.775 121.585 131.985 122.115 ;
        RECT 132.245 121.375 132.575 121.900 ;
        RECT 132.745 121.505 132.915 122.115 ;
        RECT 133.085 121.460 133.415 121.895 ;
        RECT 133.085 121.375 133.465 121.460 ;
        RECT 132.375 121.205 132.575 121.375 ;
        RECT 133.240 121.335 133.465 121.375 ;
        RECT 131.330 120.875 132.205 121.205 ;
        RECT 132.375 120.875 133.125 121.205 ;
        RECT 130.140 119.735 130.390 120.065 ;
        RECT 131.330 120.035 131.500 120.875 ;
        RECT 132.375 120.670 132.565 120.875 ;
        RECT 133.295 120.755 133.465 121.335 ;
        RECT 133.250 120.705 133.465 120.755 ;
        RECT 131.670 120.295 132.565 120.670 ;
        RECT 133.075 120.625 133.465 120.705 ;
        RECT 133.645 121.390 133.975 121.900 ;
        RECT 134.145 121.715 134.475 122.115 ;
        RECT 135.525 121.545 135.855 121.885 ;
        RECT 136.025 121.715 136.355 122.115 ;
        RECT 133.645 120.625 133.835 121.390 ;
        RECT 134.145 121.375 136.510 121.545 ;
        RECT 134.145 121.205 134.315 121.375 ;
        RECT 134.005 120.875 134.315 121.205 ;
        RECT 134.485 120.875 134.790 121.205 ;
        RECT 130.615 119.865 131.500 120.035 ;
        RECT 131.680 119.565 131.995 120.065 ;
        RECT 132.225 119.735 132.565 120.295 ;
        RECT 132.735 119.565 132.905 120.575 ;
        RECT 133.075 119.780 133.405 120.625 ;
        RECT 133.645 119.775 133.975 120.625 ;
        RECT 134.145 119.565 134.395 120.705 ;
        RECT 134.575 120.545 134.790 120.875 ;
        RECT 134.965 120.545 135.250 121.205 ;
        RECT 135.445 120.545 135.710 121.205 ;
        RECT 135.925 120.545 136.170 121.205 ;
        RECT 136.340 120.375 136.510 121.375 ;
        RECT 134.585 120.205 135.875 120.375 ;
        RECT 134.585 119.785 134.835 120.205 ;
        RECT 135.065 119.565 135.395 120.035 ;
        RECT 135.625 119.785 135.875 120.205 ;
        RECT 136.055 120.205 136.510 120.375 ;
        RECT 136.860 120.515 137.195 121.935 ;
        RECT 137.375 121.745 138.120 122.115 ;
        RECT 138.685 121.575 138.940 121.935 ;
        RECT 139.120 121.745 139.450 122.115 ;
        RECT 139.630 121.575 139.855 121.935 ;
        RECT 137.370 121.385 139.855 121.575 ;
        RECT 137.370 120.695 137.595 121.385 ;
        RECT 140.095 121.305 140.335 122.115 ;
        RECT 140.505 121.305 140.835 121.945 ;
        RECT 141.005 121.305 141.275 122.115 ;
        RECT 141.455 121.655 142.015 121.945 ;
        RECT 142.185 121.655 142.435 122.115 ;
        RECT 137.795 120.875 138.075 121.205 ;
        RECT 138.255 120.875 138.830 121.205 ;
        RECT 139.010 120.875 139.445 121.205 ;
        RECT 139.625 120.875 139.895 121.205 ;
        RECT 140.075 120.875 140.425 121.125 ;
        RECT 140.595 120.705 140.765 121.305 ;
        RECT 140.935 120.875 141.285 121.125 ;
        RECT 137.370 120.515 139.865 120.695 ;
        RECT 136.055 119.775 136.385 120.205 ;
        RECT 136.860 119.745 137.125 120.515 ;
        RECT 137.295 119.565 137.625 120.285 ;
        RECT 137.815 120.105 139.005 120.335 ;
        RECT 137.815 119.745 138.075 120.105 ;
        RECT 138.245 119.565 138.575 119.935 ;
        RECT 138.745 119.745 139.005 120.105 ;
        RECT 139.575 119.745 139.865 120.515 ;
        RECT 140.085 120.535 140.765 120.705 ;
        RECT 140.085 119.750 140.415 120.535 ;
        RECT 140.945 119.565 141.275 120.705 ;
        RECT 141.455 120.285 141.705 121.655 ;
        RECT 143.055 121.485 143.385 121.845 ;
        RECT 141.995 121.295 143.385 121.485 ;
        RECT 144.265 121.460 144.595 121.895 ;
        RECT 144.765 121.505 144.935 122.115 ;
        RECT 144.215 121.375 144.595 121.460 ;
        RECT 145.105 121.375 145.435 121.900 ;
        RECT 145.695 121.585 145.905 122.115 ;
        RECT 146.180 121.665 146.965 121.835 ;
        RECT 147.135 121.665 147.540 121.835 ;
        RECT 144.215 121.335 144.440 121.375 ;
        RECT 141.995 121.205 142.165 121.295 ;
        RECT 141.875 120.875 142.165 121.205 ;
        RECT 142.335 120.875 142.675 121.125 ;
        RECT 142.895 120.875 143.570 121.125 ;
        RECT 141.995 120.625 142.165 120.875 ;
        RECT 141.995 120.455 142.935 120.625 ;
        RECT 143.305 120.515 143.570 120.875 ;
        RECT 144.215 120.755 144.385 121.335 ;
        RECT 145.105 121.205 145.305 121.375 ;
        RECT 146.180 121.205 146.350 121.665 ;
        RECT 144.555 120.875 145.305 121.205 ;
        RECT 145.475 120.875 146.350 121.205 ;
        RECT 144.215 120.705 144.430 120.755 ;
        RECT 144.215 120.625 144.605 120.705 ;
        RECT 141.455 119.735 141.915 120.285 ;
        RECT 142.105 119.565 142.435 120.285 ;
        RECT 142.635 119.905 142.935 120.455 ;
        RECT 143.105 119.565 143.385 120.235 ;
        RECT 144.275 119.780 144.605 120.625 ;
        RECT 145.115 120.670 145.305 120.875 ;
        RECT 144.775 119.565 144.945 120.575 ;
        RECT 145.115 120.295 146.010 120.670 ;
        RECT 145.115 119.735 145.455 120.295 ;
        RECT 145.685 119.565 146.000 120.065 ;
        RECT 146.180 120.035 146.350 120.875 ;
        RECT 146.520 121.165 146.985 121.495 ;
        RECT 147.370 121.435 147.540 121.665 ;
        RECT 147.720 121.615 148.090 122.115 ;
        RECT 148.410 121.665 149.085 121.835 ;
        RECT 149.280 121.665 149.615 121.835 ;
        RECT 146.520 120.205 146.840 121.165 ;
        RECT 147.370 121.135 148.200 121.435 ;
        RECT 147.010 120.235 147.200 120.955 ;
        RECT 147.370 120.065 147.540 121.135 ;
        RECT 148.000 121.105 148.200 121.135 ;
        RECT 147.710 120.885 147.880 120.955 ;
        RECT 148.410 120.885 148.580 121.665 ;
        RECT 149.445 121.525 149.615 121.665 ;
        RECT 149.785 121.655 150.035 122.115 ;
        RECT 147.710 120.715 148.580 120.885 ;
        RECT 148.750 121.245 149.275 121.465 ;
        RECT 149.445 121.395 149.670 121.525 ;
        RECT 147.710 120.625 148.220 120.715 ;
        RECT 146.180 119.865 147.065 120.035 ;
        RECT 147.290 119.735 147.540 120.065 ;
        RECT 147.710 119.565 147.880 120.365 ;
        RECT 148.050 120.010 148.220 120.625 ;
        RECT 148.750 120.545 148.920 121.245 ;
        RECT 148.390 120.180 148.920 120.545 ;
        RECT 149.090 120.480 149.330 121.075 ;
        RECT 149.500 120.290 149.670 121.395 ;
        RECT 149.840 120.535 150.120 121.485 ;
        RECT 149.365 120.160 149.670 120.290 ;
        RECT 148.050 119.840 149.155 120.010 ;
        RECT 149.365 119.735 149.615 120.160 ;
        RECT 149.785 119.565 150.050 120.025 ;
        RECT 150.290 119.735 150.475 121.855 ;
        RECT 150.645 121.735 150.975 122.115 ;
        RECT 151.145 121.565 151.315 121.855 ;
        RECT 150.650 121.395 151.315 121.565 ;
        RECT 150.650 120.405 150.880 121.395 ;
        RECT 151.575 121.390 151.865 122.115 ;
        RECT 152.035 121.345 155.545 122.115 ;
        RECT 155.715 121.365 156.925 122.115 ;
        RECT 151.050 120.575 151.400 121.225 ;
        RECT 152.035 120.825 153.685 121.345 ;
        RECT 150.650 120.235 151.315 120.405 ;
        RECT 150.645 119.565 150.975 120.065 ;
        RECT 151.145 119.735 151.315 120.235 ;
        RECT 151.575 119.565 151.865 120.730 ;
        RECT 153.855 120.655 155.545 121.175 ;
        RECT 152.035 119.565 155.545 120.655 ;
        RECT 155.715 120.655 156.235 121.195 ;
        RECT 156.405 120.825 156.925 121.365 ;
        RECT 155.715 119.565 156.925 120.655 ;
        RECT 22.690 119.395 157.010 119.565 ;
        RECT 22.775 118.305 23.985 119.395 ;
        RECT 24.155 118.305 25.825 119.395 ;
        RECT 22.775 117.595 23.295 118.135 ;
        RECT 23.465 117.765 23.985 118.305 ;
        RECT 24.155 117.615 24.905 118.135 ;
        RECT 25.075 117.785 25.825 118.305 ;
        RECT 26.180 118.425 26.570 118.600 ;
        RECT 27.055 118.595 27.385 119.395 ;
        RECT 27.555 118.605 28.090 119.225 ;
        RECT 26.180 118.255 27.605 118.425 ;
        RECT 22.775 116.845 23.985 117.595 ;
        RECT 24.155 116.845 25.825 117.615 ;
        RECT 26.055 117.525 26.410 118.085 ;
        RECT 26.580 117.355 26.750 118.255 ;
        RECT 26.920 117.525 27.185 118.085 ;
        RECT 27.435 117.755 27.605 118.255 ;
        RECT 27.775 117.585 28.090 118.605 ;
        RECT 28.355 118.335 28.685 119.180 ;
        RECT 28.855 118.385 29.025 119.395 ;
        RECT 29.195 118.665 29.535 119.225 ;
        RECT 29.765 118.895 30.080 119.395 ;
        RECT 30.260 118.925 31.145 119.095 ;
        RECT 26.160 116.845 26.400 117.355 ;
        RECT 26.580 117.025 26.860 117.355 ;
        RECT 27.090 116.845 27.305 117.355 ;
        RECT 27.475 117.015 28.090 117.585 ;
        RECT 28.295 118.255 28.685 118.335 ;
        RECT 29.195 118.290 30.090 118.665 ;
        RECT 28.295 118.205 28.510 118.255 ;
        RECT 28.295 117.625 28.465 118.205 ;
        RECT 29.195 118.085 29.385 118.290 ;
        RECT 30.260 118.085 30.430 118.925 ;
        RECT 31.370 118.895 31.620 119.225 ;
        RECT 28.635 117.755 29.385 118.085 ;
        RECT 29.555 117.755 30.430 118.085 ;
        RECT 28.295 117.585 28.520 117.625 ;
        RECT 29.185 117.585 29.385 117.755 ;
        RECT 28.295 117.500 28.675 117.585 ;
        RECT 28.345 117.065 28.675 117.500 ;
        RECT 28.845 116.845 29.015 117.455 ;
        RECT 29.185 117.060 29.515 117.585 ;
        RECT 29.775 116.845 29.985 117.375 ;
        RECT 30.260 117.295 30.430 117.755 ;
        RECT 30.600 117.795 30.920 118.755 ;
        RECT 31.090 118.005 31.280 118.725 ;
        RECT 31.450 117.825 31.620 118.895 ;
        RECT 31.790 118.595 31.960 119.395 ;
        RECT 32.130 118.950 33.235 119.120 ;
        RECT 32.130 118.335 32.300 118.950 ;
        RECT 33.445 118.800 33.695 119.225 ;
        RECT 33.865 118.935 34.130 119.395 ;
        RECT 32.470 118.415 33.000 118.780 ;
        RECT 33.445 118.670 33.750 118.800 ;
        RECT 31.790 118.245 32.300 118.335 ;
        RECT 31.790 118.075 32.660 118.245 ;
        RECT 31.790 118.005 31.960 118.075 ;
        RECT 32.080 117.825 32.280 117.855 ;
        RECT 30.600 117.465 31.065 117.795 ;
        RECT 31.450 117.525 32.280 117.825 ;
        RECT 31.450 117.295 31.620 117.525 ;
        RECT 30.260 117.125 31.045 117.295 ;
        RECT 31.215 117.125 31.620 117.295 ;
        RECT 31.800 116.845 32.170 117.345 ;
        RECT 32.490 117.295 32.660 118.075 ;
        RECT 32.830 117.715 33.000 118.415 ;
        RECT 33.170 117.885 33.410 118.480 ;
        RECT 32.830 117.495 33.355 117.715 ;
        RECT 33.580 117.565 33.750 118.670 ;
        RECT 33.525 117.435 33.750 117.565 ;
        RECT 33.920 117.475 34.200 118.425 ;
        RECT 33.525 117.295 33.695 117.435 ;
        RECT 32.490 117.125 33.165 117.295 ;
        RECT 33.360 117.125 33.695 117.295 ;
        RECT 33.865 116.845 34.115 117.305 ;
        RECT 34.370 117.105 34.555 119.225 ;
        RECT 34.725 118.895 35.055 119.395 ;
        RECT 35.225 118.725 35.395 119.225 ;
        RECT 34.730 118.555 35.395 118.725 ;
        RECT 34.730 117.565 34.960 118.555 ;
        RECT 35.130 117.735 35.480 118.385 ;
        RECT 35.655 118.230 35.945 119.395 ;
        RECT 36.115 118.255 36.500 119.225 ;
        RECT 36.670 118.935 36.995 119.395 ;
        RECT 37.515 118.765 37.795 119.225 ;
        RECT 36.670 118.545 37.795 118.765 ;
        RECT 36.115 117.585 36.395 118.255 ;
        RECT 36.670 118.085 37.120 118.545 ;
        RECT 37.985 118.375 38.385 119.225 ;
        RECT 38.785 118.935 39.055 119.395 ;
        RECT 39.225 118.765 39.510 119.225 ;
        RECT 36.565 117.755 37.120 118.085 ;
        RECT 37.290 117.815 38.385 118.375 ;
        RECT 36.670 117.645 37.120 117.755 ;
        RECT 34.730 117.395 35.395 117.565 ;
        RECT 34.725 116.845 35.055 117.225 ;
        RECT 35.225 117.105 35.395 117.395 ;
        RECT 35.655 116.845 35.945 117.570 ;
        RECT 36.115 117.015 36.500 117.585 ;
        RECT 36.670 117.475 37.795 117.645 ;
        RECT 36.670 116.845 36.995 117.305 ;
        RECT 37.515 117.015 37.795 117.475 ;
        RECT 37.985 117.015 38.385 117.815 ;
        RECT 38.555 118.545 39.510 118.765 ;
        RECT 38.555 117.645 38.765 118.545 ;
        RECT 38.935 117.815 39.625 118.375 ;
        RECT 39.795 118.255 40.135 119.225 ;
        RECT 40.305 118.255 40.475 119.395 ;
        RECT 40.745 118.595 40.995 119.395 ;
        RECT 41.640 118.425 41.970 119.225 ;
        RECT 42.270 118.595 42.600 119.395 ;
        RECT 42.770 118.425 43.100 119.225 ;
        RECT 40.665 118.255 43.100 118.425 ;
        RECT 43.475 118.255 43.860 119.225 ;
        RECT 44.030 118.935 44.355 119.395 ;
        RECT 44.875 118.765 45.155 119.225 ;
        RECT 44.030 118.545 45.155 118.765 ;
        RECT 39.795 117.645 39.970 118.255 ;
        RECT 40.665 118.005 40.835 118.255 ;
        RECT 40.140 117.835 40.835 118.005 ;
        RECT 41.010 117.835 41.430 118.035 ;
        RECT 41.600 117.835 41.930 118.035 ;
        RECT 42.100 117.835 42.430 118.035 ;
        RECT 38.555 117.475 39.510 117.645 ;
        RECT 38.785 116.845 39.055 117.305 ;
        RECT 39.225 117.015 39.510 117.475 ;
        RECT 39.795 117.015 40.135 117.645 ;
        RECT 40.305 116.845 40.555 117.645 ;
        RECT 40.745 117.495 41.970 117.665 ;
        RECT 40.745 117.015 41.075 117.495 ;
        RECT 41.245 116.845 41.470 117.305 ;
        RECT 41.640 117.015 41.970 117.495 ;
        RECT 42.600 117.625 42.770 118.255 ;
        RECT 42.955 117.835 43.305 118.085 ;
        RECT 42.600 117.015 43.100 117.625 ;
        RECT 43.475 117.585 43.755 118.255 ;
        RECT 44.030 118.085 44.480 118.545 ;
        RECT 45.345 118.375 45.745 119.225 ;
        RECT 46.145 118.935 46.415 119.395 ;
        RECT 46.585 118.765 46.870 119.225 ;
        RECT 43.925 117.755 44.480 118.085 ;
        RECT 44.650 117.815 45.745 118.375 ;
        RECT 44.030 117.645 44.480 117.755 ;
        RECT 43.475 117.015 43.860 117.585 ;
        RECT 44.030 117.475 45.155 117.645 ;
        RECT 44.030 116.845 44.355 117.305 ;
        RECT 44.875 117.015 45.155 117.475 ;
        RECT 45.345 117.015 45.745 117.815 ;
        RECT 45.915 118.545 46.870 118.765 ;
        RECT 45.915 117.645 46.125 118.545 ;
        RECT 48.280 118.425 48.610 119.225 ;
        RECT 48.780 118.595 49.110 119.395 ;
        RECT 49.410 118.425 49.740 119.225 ;
        RECT 50.385 118.595 50.635 119.395 ;
        RECT 46.295 117.815 46.985 118.375 ;
        RECT 48.280 118.255 50.715 118.425 ;
        RECT 50.905 118.255 51.075 119.395 ;
        RECT 51.245 118.255 51.585 119.225 ;
        RECT 51.870 118.765 52.155 119.225 ;
        RECT 52.325 118.935 52.595 119.395 ;
        RECT 51.870 118.545 52.825 118.765 ;
        RECT 48.075 117.835 48.425 118.085 ;
        RECT 45.915 117.475 46.870 117.645 ;
        RECT 48.610 117.625 48.780 118.255 ;
        RECT 48.950 117.835 49.280 118.035 ;
        RECT 49.450 117.835 49.780 118.035 ;
        RECT 49.950 117.835 50.370 118.035 ;
        RECT 50.545 118.005 50.715 118.255 ;
        RECT 50.545 117.835 51.240 118.005 ;
        RECT 46.145 116.845 46.415 117.305 ;
        RECT 46.585 117.015 46.870 117.475 ;
        RECT 48.280 117.015 48.780 117.625 ;
        RECT 49.410 117.495 50.635 117.665 ;
        RECT 51.410 117.645 51.585 118.255 ;
        RECT 51.755 117.815 52.445 118.375 ;
        RECT 52.615 117.645 52.825 118.545 ;
        RECT 49.410 117.015 49.740 117.495 ;
        RECT 49.910 116.845 50.135 117.305 ;
        RECT 50.305 117.015 50.635 117.495 ;
        RECT 50.825 116.845 51.075 117.645 ;
        RECT 51.245 117.015 51.585 117.645 ;
        RECT 51.870 117.475 52.825 117.645 ;
        RECT 52.995 118.375 53.395 119.225 ;
        RECT 53.585 118.765 53.865 119.225 ;
        RECT 54.385 118.935 54.710 119.395 ;
        RECT 53.585 118.545 54.710 118.765 ;
        RECT 52.995 117.815 54.090 118.375 ;
        RECT 54.260 118.085 54.710 118.545 ;
        RECT 54.880 118.255 55.265 119.225 ;
        RECT 51.870 117.015 52.155 117.475 ;
        RECT 52.325 116.845 52.595 117.305 ;
        RECT 52.995 117.015 53.395 117.815 ;
        RECT 54.260 117.755 54.815 118.085 ;
        RECT 54.260 117.645 54.710 117.755 ;
        RECT 53.585 117.475 54.710 117.645 ;
        RECT 54.985 117.585 55.265 118.255 ;
        RECT 53.585 117.015 53.865 117.475 ;
        RECT 54.385 116.845 54.710 117.305 ;
        RECT 54.880 117.015 55.265 117.585 ;
        RECT 55.470 118.605 56.005 119.225 ;
        RECT 55.470 117.585 55.785 118.605 ;
        RECT 56.175 118.595 56.505 119.395 ;
        RECT 56.990 118.425 57.380 118.600 ;
        RECT 55.955 118.255 57.380 118.425 ;
        RECT 57.735 118.255 58.005 119.225 ;
        RECT 58.215 118.595 58.495 119.395 ;
        RECT 58.675 118.845 59.870 119.175 ;
        RECT 59.000 118.425 59.420 118.675 ;
        RECT 58.175 118.255 59.420 118.425 ;
        RECT 55.955 117.755 56.125 118.255 ;
        RECT 55.470 117.015 56.085 117.585 ;
        RECT 56.375 117.525 56.640 118.085 ;
        RECT 56.810 117.355 56.980 118.255 ;
        RECT 57.150 117.525 57.505 118.085 ;
        RECT 57.735 117.520 57.905 118.255 ;
        RECT 58.175 118.085 58.345 118.255 ;
        RECT 59.645 118.085 59.815 118.645 ;
        RECT 60.065 118.255 60.320 119.395 ;
        RECT 61.415 118.230 61.705 119.395 ;
        RECT 61.875 118.305 65.385 119.395 ;
        RECT 58.115 117.755 58.345 118.085 ;
        RECT 59.075 117.755 59.815 118.085 ;
        RECT 59.985 117.835 60.320 118.085 ;
        RECT 58.175 117.585 58.345 117.755 ;
        RECT 59.565 117.665 59.815 117.755 ;
        RECT 56.255 116.845 56.470 117.355 ;
        RECT 56.700 117.025 56.980 117.355 ;
        RECT 57.160 116.845 57.400 117.355 ;
        RECT 57.735 117.175 58.005 117.520 ;
        RECT 58.175 117.415 58.915 117.585 ;
        RECT 59.565 117.495 60.300 117.665 ;
        RECT 61.875 117.615 63.525 118.135 ;
        RECT 63.695 117.785 65.385 118.305 ;
        RECT 66.020 118.255 66.355 119.225 ;
        RECT 66.525 118.255 66.695 119.395 ;
        RECT 66.865 119.055 68.895 119.225 ;
        RECT 58.195 116.845 58.575 117.245 ;
        RECT 58.745 117.065 58.915 117.415 ;
        RECT 59.085 116.845 59.820 117.325 ;
        RECT 59.990 117.025 60.300 117.495 ;
        RECT 61.415 116.845 61.705 117.570 ;
        RECT 61.875 116.845 65.385 117.615 ;
        RECT 66.020 117.585 66.190 118.255 ;
        RECT 66.865 118.085 67.035 119.055 ;
        RECT 66.360 117.755 66.615 118.085 ;
        RECT 66.840 117.755 67.035 118.085 ;
        RECT 67.205 118.715 68.330 118.885 ;
        RECT 66.445 117.585 66.615 117.755 ;
        RECT 67.205 117.585 67.375 118.715 ;
        RECT 66.020 117.015 66.275 117.585 ;
        RECT 66.445 117.415 67.375 117.585 ;
        RECT 67.545 118.375 68.555 118.545 ;
        RECT 67.545 117.575 67.715 118.375 ;
        RECT 67.920 117.695 68.195 118.175 ;
        RECT 67.915 117.525 68.195 117.695 ;
        RECT 67.200 117.380 67.375 117.415 ;
        RECT 66.445 116.845 66.775 117.245 ;
        RECT 67.200 117.015 67.730 117.380 ;
        RECT 67.920 117.015 68.195 117.525 ;
        RECT 68.365 117.015 68.555 118.375 ;
        RECT 68.725 118.390 68.895 119.055 ;
        RECT 69.065 118.635 69.235 119.395 ;
        RECT 69.470 118.635 69.985 119.045 ;
        RECT 68.725 118.200 69.475 118.390 ;
        RECT 69.645 117.825 69.985 118.635 ;
        RECT 70.215 118.255 70.425 119.395 ;
        RECT 68.755 117.655 69.985 117.825 ;
        RECT 70.595 118.245 70.925 119.225 ;
        RECT 71.095 118.255 71.325 119.395 ;
        RECT 71.535 118.960 76.880 119.395 ;
        RECT 68.735 116.845 69.245 117.380 ;
        RECT 69.465 117.050 69.710 117.655 ;
        RECT 70.215 116.845 70.425 117.665 ;
        RECT 70.595 117.645 70.845 118.245 ;
        RECT 71.015 117.835 71.345 118.085 ;
        RECT 70.595 117.015 70.925 117.645 ;
        RECT 71.095 116.845 71.325 117.665 ;
        RECT 73.120 117.390 73.460 118.220 ;
        RECT 74.940 117.710 75.290 118.960 ;
        RECT 77.515 118.840 78.120 119.395 ;
        RECT 78.295 118.885 78.775 119.225 ;
        RECT 78.945 118.850 79.200 119.395 ;
        RECT 77.515 118.740 78.130 118.840 ;
        RECT 77.945 118.715 78.130 118.740 ;
        RECT 77.515 118.120 77.775 118.570 ;
        RECT 77.945 118.470 78.275 118.715 ;
        RECT 78.445 118.395 79.200 118.645 ;
        RECT 79.370 118.525 79.645 119.225 ;
        RECT 78.430 118.360 79.200 118.395 ;
        RECT 78.415 118.350 79.200 118.360 ;
        RECT 78.410 118.335 79.305 118.350 ;
        RECT 78.390 118.320 79.305 118.335 ;
        RECT 78.370 118.310 79.305 118.320 ;
        RECT 78.345 118.300 79.305 118.310 ;
        RECT 78.275 118.270 79.305 118.300 ;
        RECT 78.255 118.240 79.305 118.270 ;
        RECT 78.235 118.210 79.305 118.240 ;
        RECT 78.205 118.185 79.305 118.210 ;
        RECT 78.170 118.150 79.305 118.185 ;
        RECT 78.140 118.145 79.305 118.150 ;
        RECT 78.140 118.140 78.530 118.145 ;
        RECT 78.140 118.130 78.505 118.140 ;
        RECT 78.140 118.125 78.490 118.130 ;
        RECT 78.140 118.120 78.475 118.125 ;
        RECT 77.515 118.115 78.475 118.120 ;
        RECT 77.515 118.105 78.465 118.115 ;
        RECT 77.515 118.100 78.455 118.105 ;
        RECT 77.515 118.090 78.445 118.100 ;
        RECT 77.515 118.080 78.440 118.090 ;
        RECT 77.515 118.075 78.435 118.080 ;
        RECT 77.515 118.060 78.425 118.075 ;
        RECT 77.515 118.045 78.420 118.060 ;
        RECT 77.515 118.020 78.410 118.045 ;
        RECT 77.515 117.950 78.405 118.020 ;
        RECT 77.515 117.395 78.065 117.780 ;
        RECT 71.535 116.845 76.880 117.390 ;
        RECT 78.235 117.225 78.405 117.950 ;
        RECT 77.515 117.055 78.405 117.225 ;
        RECT 78.575 117.550 78.905 117.975 ;
        RECT 79.075 117.750 79.305 118.145 ;
        RECT 78.575 117.065 78.795 117.550 ;
        RECT 79.475 117.495 79.645 118.525 ;
        RECT 78.965 116.845 79.215 117.385 ;
        RECT 79.385 117.015 79.645 117.495 ;
        RECT 79.815 118.320 80.085 119.225 ;
        RECT 80.255 118.635 80.585 119.395 ;
        RECT 80.765 118.465 80.935 119.225 ;
        RECT 79.815 117.520 79.985 118.320 ;
        RECT 80.270 118.295 80.935 118.465 ;
        RECT 81.655 118.675 82.115 119.225 ;
        RECT 82.305 118.675 82.635 119.395 ;
        RECT 80.270 118.150 80.440 118.295 ;
        RECT 80.155 117.820 80.440 118.150 ;
        RECT 80.270 117.565 80.440 117.820 ;
        RECT 80.675 117.745 81.005 118.115 ;
        RECT 79.815 117.015 80.075 117.520 ;
        RECT 80.270 117.395 80.935 117.565 ;
        RECT 80.255 116.845 80.585 117.225 ;
        RECT 80.765 117.015 80.935 117.395 ;
        RECT 81.655 117.305 81.905 118.675 ;
        RECT 82.835 118.505 83.135 119.055 ;
        RECT 83.305 118.725 83.585 119.395 ;
        RECT 82.195 118.335 83.135 118.505 ;
        RECT 82.195 118.085 82.365 118.335 ;
        RECT 83.505 118.085 83.770 118.445 ;
        RECT 82.075 117.755 82.365 118.085 ;
        RECT 82.535 117.835 82.875 118.085 ;
        RECT 83.095 117.835 83.770 118.085 ;
        RECT 83.955 118.320 84.225 119.225 ;
        RECT 84.395 118.635 84.725 119.395 ;
        RECT 84.905 118.465 85.075 119.225 ;
        RECT 82.195 117.665 82.365 117.755 ;
        RECT 82.195 117.475 83.585 117.665 ;
        RECT 81.655 117.015 82.215 117.305 ;
        RECT 82.385 116.845 82.635 117.305 ;
        RECT 83.255 117.115 83.585 117.475 ;
        RECT 83.955 117.520 84.125 118.320 ;
        RECT 84.410 118.295 85.075 118.465 ;
        RECT 85.335 118.305 87.005 119.395 ;
        RECT 84.410 118.150 84.580 118.295 ;
        RECT 84.295 117.820 84.580 118.150 ;
        RECT 84.410 117.565 84.580 117.820 ;
        RECT 84.815 117.745 85.145 118.115 ;
        RECT 85.335 117.615 86.085 118.135 ;
        RECT 86.255 117.785 87.005 118.305 ;
        RECT 87.175 118.230 87.465 119.395 ;
        RECT 87.640 118.255 87.975 119.225 ;
        RECT 88.145 118.255 88.315 119.395 ;
        RECT 88.485 119.055 90.515 119.225 ;
        RECT 83.955 117.015 84.215 117.520 ;
        RECT 84.410 117.395 85.075 117.565 ;
        RECT 84.395 116.845 84.725 117.225 ;
        RECT 84.905 117.015 85.075 117.395 ;
        RECT 85.335 116.845 87.005 117.615 ;
        RECT 87.640 117.585 87.810 118.255 ;
        RECT 88.485 118.085 88.655 119.055 ;
        RECT 87.980 117.755 88.235 118.085 ;
        RECT 88.460 117.755 88.655 118.085 ;
        RECT 88.825 118.715 89.950 118.885 ;
        RECT 88.065 117.585 88.235 117.755 ;
        RECT 88.825 117.585 88.995 118.715 ;
        RECT 87.175 116.845 87.465 117.570 ;
        RECT 87.640 117.015 87.895 117.585 ;
        RECT 88.065 117.415 88.995 117.585 ;
        RECT 89.165 118.375 90.175 118.545 ;
        RECT 89.165 117.575 89.335 118.375 ;
        RECT 89.540 117.695 89.815 118.175 ;
        RECT 89.535 117.525 89.815 117.695 ;
        RECT 88.820 117.380 88.995 117.415 ;
        RECT 88.065 116.845 88.395 117.245 ;
        RECT 88.820 117.015 89.350 117.380 ;
        RECT 89.540 117.015 89.815 117.525 ;
        RECT 89.985 117.015 90.175 118.375 ;
        RECT 90.345 118.390 90.515 119.055 ;
        RECT 90.685 118.635 90.855 119.395 ;
        RECT 91.090 118.635 91.605 119.045 ;
        RECT 90.345 118.200 91.095 118.390 ;
        RECT 91.265 117.825 91.605 118.635 ;
        RECT 90.375 117.655 91.605 117.825 ;
        RECT 92.700 118.255 93.035 119.225 ;
        RECT 93.205 118.255 93.375 119.395 ;
        RECT 93.545 119.055 95.575 119.225 ;
        RECT 90.355 116.845 90.865 117.380 ;
        RECT 91.085 117.050 91.330 117.655 ;
        RECT 92.700 117.585 92.870 118.255 ;
        RECT 93.545 118.085 93.715 119.055 ;
        RECT 93.040 117.755 93.295 118.085 ;
        RECT 93.520 117.755 93.715 118.085 ;
        RECT 93.885 118.715 95.010 118.885 ;
        RECT 93.125 117.585 93.295 117.755 ;
        RECT 93.885 117.585 94.055 118.715 ;
        RECT 92.700 117.015 92.955 117.585 ;
        RECT 93.125 117.415 94.055 117.585 ;
        RECT 94.225 118.375 95.235 118.545 ;
        RECT 94.225 117.575 94.395 118.375 ;
        RECT 94.600 118.035 94.875 118.175 ;
        RECT 94.595 117.865 94.875 118.035 ;
        RECT 93.880 117.380 94.055 117.415 ;
        RECT 93.125 116.845 93.455 117.245 ;
        RECT 93.880 117.015 94.410 117.380 ;
        RECT 94.600 117.015 94.875 117.865 ;
        RECT 95.045 117.015 95.235 118.375 ;
        RECT 95.405 118.390 95.575 119.055 ;
        RECT 95.745 118.635 95.915 119.395 ;
        RECT 96.150 118.635 96.665 119.045 ;
        RECT 95.405 118.200 96.155 118.390 ;
        RECT 96.325 117.825 96.665 118.635 ;
        RECT 96.835 118.305 98.505 119.395 ;
        RECT 95.435 117.655 96.665 117.825 ;
        RECT 95.415 116.845 95.925 117.380 ;
        RECT 96.145 117.050 96.390 117.655 ;
        RECT 96.835 117.615 97.585 118.135 ;
        RECT 97.755 117.785 98.505 118.305 ;
        RECT 99.140 118.255 99.475 119.225 ;
        RECT 99.645 118.255 99.815 119.395 ;
        RECT 99.985 119.055 102.015 119.225 ;
        RECT 96.835 116.845 98.505 117.615 ;
        RECT 99.140 117.585 99.310 118.255 ;
        RECT 99.985 118.085 100.155 119.055 ;
        RECT 99.480 117.755 99.735 118.085 ;
        RECT 99.960 117.755 100.155 118.085 ;
        RECT 100.325 118.715 101.450 118.885 ;
        RECT 99.565 117.585 99.735 117.755 ;
        RECT 100.325 117.585 100.495 118.715 ;
        RECT 99.140 117.015 99.395 117.585 ;
        RECT 99.565 117.415 100.495 117.585 ;
        RECT 100.665 118.375 101.675 118.545 ;
        RECT 100.665 117.575 100.835 118.375 ;
        RECT 101.040 118.035 101.315 118.175 ;
        RECT 101.035 117.865 101.315 118.035 ;
        RECT 100.320 117.380 100.495 117.415 ;
        RECT 99.565 116.845 99.895 117.245 ;
        RECT 100.320 117.015 100.850 117.380 ;
        RECT 101.040 117.015 101.315 117.865 ;
        RECT 101.485 117.015 101.675 118.375 ;
        RECT 101.845 118.390 102.015 119.055 ;
        RECT 102.185 118.635 102.355 119.395 ;
        RECT 102.590 118.635 103.105 119.045 ;
        RECT 103.275 118.960 108.620 119.395 ;
        RECT 101.845 118.200 102.595 118.390 ;
        RECT 102.765 117.825 103.105 118.635 ;
        RECT 101.875 117.655 103.105 117.825 ;
        RECT 101.855 116.845 102.365 117.380 ;
        RECT 102.585 117.050 102.830 117.655 ;
        RECT 104.860 117.390 105.200 118.220 ;
        RECT 106.680 117.710 107.030 118.960 ;
        RECT 108.795 118.305 110.465 119.395 ;
        RECT 108.795 117.615 109.545 118.135 ;
        RECT 109.715 117.785 110.465 118.305 ;
        RECT 110.635 118.675 111.095 119.225 ;
        RECT 111.285 118.675 111.615 119.395 ;
        RECT 103.275 116.845 108.620 117.390 ;
        RECT 108.795 116.845 110.465 117.615 ;
        RECT 110.635 117.305 110.885 118.675 ;
        RECT 111.815 118.505 112.115 119.055 ;
        RECT 112.285 118.725 112.565 119.395 ;
        RECT 111.175 118.335 112.115 118.505 ;
        RECT 111.175 118.085 111.345 118.335 ;
        RECT 112.485 118.085 112.750 118.445 ;
        RECT 112.935 118.230 113.225 119.395 ;
        RECT 113.405 118.415 113.735 119.225 ;
        RECT 113.905 118.595 114.145 119.395 ;
        RECT 113.405 118.245 114.120 118.415 ;
        RECT 111.055 117.755 111.345 118.085 ;
        RECT 111.515 117.835 111.855 118.085 ;
        RECT 112.075 117.835 112.750 118.085 ;
        RECT 113.400 117.835 113.780 118.075 ;
        RECT 113.950 118.005 114.120 118.245 ;
        RECT 114.325 118.375 114.495 119.225 ;
        RECT 114.665 118.595 114.995 119.395 ;
        RECT 115.165 118.375 115.335 119.225 ;
        RECT 114.325 118.205 115.335 118.375 ;
        RECT 115.505 118.245 115.835 119.395 ;
        RECT 116.270 118.765 116.555 119.225 ;
        RECT 116.725 118.935 116.995 119.395 ;
        RECT 116.270 118.545 117.225 118.765 ;
        RECT 113.950 117.835 114.450 118.005 ;
        RECT 111.175 117.665 111.345 117.755 ;
        RECT 113.950 117.665 114.120 117.835 ;
        RECT 114.840 117.695 115.335 118.205 ;
        RECT 116.155 117.815 116.845 118.375 ;
        RECT 114.835 117.665 115.335 117.695 ;
        RECT 111.175 117.475 112.565 117.665 ;
        RECT 110.635 117.015 111.195 117.305 ;
        RECT 111.365 116.845 111.615 117.305 ;
        RECT 112.235 117.115 112.565 117.475 ;
        RECT 112.935 116.845 113.225 117.570 ;
        RECT 113.485 117.495 114.120 117.665 ;
        RECT 114.325 117.495 115.335 117.665 ;
        RECT 117.015 117.645 117.225 118.545 ;
        RECT 113.485 117.015 113.655 117.495 ;
        RECT 113.835 116.845 114.075 117.325 ;
        RECT 114.325 117.015 114.495 117.495 ;
        RECT 114.665 116.845 114.995 117.325 ;
        RECT 115.165 117.015 115.335 117.495 ;
        RECT 115.505 116.845 115.835 117.645 ;
        RECT 116.270 117.475 117.225 117.645 ;
        RECT 117.395 118.375 117.795 119.225 ;
        RECT 117.985 118.765 118.265 119.225 ;
        RECT 118.785 118.935 119.110 119.395 ;
        RECT 117.985 118.545 119.110 118.765 ;
        RECT 117.395 117.815 118.490 118.375 ;
        RECT 118.660 118.085 119.110 118.545 ;
        RECT 119.280 118.255 119.665 119.225 ;
        RECT 116.270 117.015 116.555 117.475 ;
        RECT 116.725 116.845 116.995 117.305 ;
        RECT 117.395 117.015 117.795 117.815 ;
        RECT 118.660 117.755 119.215 118.085 ;
        RECT 118.660 117.645 119.110 117.755 ;
        RECT 117.985 117.475 119.110 117.645 ;
        RECT 119.385 117.585 119.665 118.255 ;
        RECT 117.985 117.015 118.265 117.475 ;
        RECT 118.785 116.845 119.110 117.305 ;
        RECT 119.280 117.015 119.665 117.585 ;
        RECT 119.845 117.025 120.105 119.215 ;
        RECT 120.275 118.665 120.615 119.395 ;
        RECT 120.795 118.485 121.065 119.215 ;
        RECT 120.295 118.265 121.065 118.485 ;
        RECT 121.245 118.505 121.475 119.215 ;
        RECT 121.645 118.685 121.975 119.395 ;
        RECT 122.145 118.505 122.405 119.215 ;
        RECT 121.245 118.265 122.405 118.505 ;
        RECT 122.595 118.320 122.865 119.225 ;
        RECT 123.035 118.635 123.365 119.395 ;
        RECT 123.545 118.465 123.715 119.225 ;
        RECT 120.295 117.595 120.585 118.265 ;
        RECT 120.765 117.775 121.230 118.085 ;
        RECT 121.410 117.775 121.935 118.085 ;
        RECT 120.295 117.395 121.525 117.595 ;
        RECT 120.365 116.845 121.035 117.215 ;
        RECT 121.215 117.025 121.525 117.395 ;
        RECT 121.705 117.135 121.935 117.775 ;
        RECT 122.115 117.755 122.415 118.085 ;
        RECT 122.115 116.845 122.405 117.575 ;
        RECT 122.595 117.520 122.765 118.320 ;
        RECT 123.050 118.295 123.715 118.465 ;
        RECT 124.440 119.005 124.775 119.225 ;
        RECT 125.780 119.015 126.135 119.395 ;
        RECT 124.440 118.385 124.695 119.005 ;
        RECT 124.945 118.845 125.175 118.885 ;
        RECT 126.305 118.845 126.555 119.225 ;
        RECT 124.945 118.645 126.555 118.845 ;
        RECT 124.945 118.555 125.130 118.645 ;
        RECT 125.720 118.635 126.555 118.645 ;
        RECT 126.805 118.615 127.055 119.395 ;
        RECT 127.225 118.545 127.485 119.225 ;
        RECT 125.285 118.445 125.615 118.475 ;
        RECT 125.285 118.385 127.085 118.445 ;
        RECT 123.050 118.150 123.220 118.295 ;
        RECT 124.440 118.275 127.145 118.385 ;
        RECT 124.440 118.215 125.615 118.275 ;
        RECT 126.945 118.240 127.145 118.275 ;
        RECT 122.935 117.820 123.220 118.150 ;
        RECT 123.050 117.565 123.220 117.820 ;
        RECT 123.455 117.745 123.785 118.115 ;
        RECT 124.435 117.835 124.925 118.035 ;
        RECT 125.115 117.835 125.590 118.045 ;
        RECT 122.595 117.015 122.855 117.520 ;
        RECT 123.050 117.395 123.715 117.565 ;
        RECT 123.035 116.845 123.365 117.225 ;
        RECT 123.545 117.015 123.715 117.395 ;
        RECT 124.440 116.845 124.895 117.610 ;
        RECT 125.370 117.435 125.590 117.835 ;
        RECT 125.835 117.835 126.165 118.045 ;
        RECT 125.835 117.435 126.045 117.835 ;
        RECT 126.335 117.800 126.745 118.105 ;
        RECT 126.975 117.665 127.145 118.240 ;
        RECT 126.875 117.545 127.145 117.665 ;
        RECT 126.300 117.500 127.145 117.545 ;
        RECT 126.300 117.375 127.055 117.500 ;
        RECT 126.300 117.225 126.470 117.375 ;
        RECT 127.315 117.355 127.485 118.545 ;
        RECT 127.655 118.305 128.865 119.395 ;
        RECT 127.255 117.345 127.485 117.355 ;
        RECT 125.170 117.015 126.470 117.225 ;
        RECT 126.725 116.845 127.055 117.205 ;
        RECT 127.225 117.015 127.485 117.345 ;
        RECT 127.655 117.595 128.175 118.135 ;
        RECT 128.345 117.765 128.865 118.305 ;
        RECT 129.035 118.255 129.420 119.225 ;
        RECT 129.590 118.935 129.915 119.395 ;
        RECT 130.435 118.765 130.715 119.225 ;
        RECT 129.590 118.545 130.715 118.765 ;
        RECT 127.655 116.845 128.865 117.595 ;
        RECT 129.035 117.585 129.315 118.255 ;
        RECT 129.590 118.085 130.040 118.545 ;
        RECT 130.905 118.375 131.305 119.225 ;
        RECT 131.705 118.935 131.975 119.395 ;
        RECT 132.145 118.765 132.430 119.225 ;
        RECT 129.485 117.755 130.040 118.085 ;
        RECT 130.210 117.815 131.305 118.375 ;
        RECT 129.590 117.645 130.040 117.755 ;
        RECT 129.035 117.015 129.420 117.585 ;
        RECT 129.590 117.475 130.715 117.645 ;
        RECT 129.590 116.845 129.915 117.305 ;
        RECT 130.435 117.015 130.715 117.475 ;
        RECT 130.905 117.015 131.305 117.815 ;
        RECT 131.475 118.545 132.430 118.765 ;
        RECT 132.715 118.545 132.975 119.225 ;
        RECT 133.145 118.615 133.395 119.395 ;
        RECT 133.645 118.845 133.895 119.225 ;
        RECT 134.065 119.015 134.420 119.395 ;
        RECT 135.425 119.005 135.760 119.225 ;
        RECT 135.025 118.845 135.255 118.885 ;
        RECT 133.645 118.645 135.255 118.845 ;
        RECT 133.645 118.635 134.480 118.645 ;
        RECT 135.070 118.555 135.255 118.645 ;
        RECT 131.475 117.645 131.685 118.545 ;
        RECT 131.855 117.815 132.545 118.375 ;
        RECT 131.475 117.475 132.430 117.645 ;
        RECT 131.705 116.845 131.975 117.305 ;
        RECT 132.145 117.015 132.430 117.475 ;
        RECT 132.715 117.355 132.885 118.545 ;
        RECT 134.585 118.445 134.915 118.475 ;
        RECT 133.115 118.385 134.915 118.445 ;
        RECT 135.505 118.385 135.760 119.005 ;
        RECT 133.055 118.275 135.760 118.385 ;
        RECT 133.055 118.240 133.255 118.275 ;
        RECT 133.055 117.665 133.225 118.240 ;
        RECT 134.585 118.215 135.760 118.275 ;
        RECT 135.970 118.605 136.505 119.225 ;
        RECT 133.455 117.800 133.865 118.105 ;
        RECT 134.035 117.835 134.365 118.045 ;
        RECT 133.055 117.545 133.325 117.665 ;
        RECT 133.055 117.500 133.900 117.545 ;
        RECT 133.145 117.375 133.900 117.500 ;
        RECT 134.155 117.435 134.365 117.835 ;
        RECT 134.610 117.835 135.085 118.045 ;
        RECT 135.275 117.835 135.765 118.035 ;
        RECT 134.610 117.435 134.830 117.835 ;
        RECT 132.715 117.345 132.945 117.355 ;
        RECT 132.715 117.015 132.975 117.345 ;
        RECT 133.730 117.225 133.900 117.375 ;
        RECT 133.145 116.845 133.475 117.205 ;
        RECT 133.730 117.015 135.030 117.225 ;
        RECT 135.305 116.845 135.760 117.610 ;
        RECT 135.970 117.585 136.285 118.605 ;
        RECT 136.675 118.595 137.005 119.395 ;
        RECT 137.490 118.425 137.880 118.600 ;
        RECT 136.455 118.255 137.880 118.425 ;
        RECT 136.455 117.755 136.625 118.255 ;
        RECT 135.970 117.015 136.585 117.585 ;
        RECT 136.875 117.525 137.140 118.085 ;
        RECT 137.310 117.355 137.480 118.255 ;
        RECT 138.695 118.230 138.985 119.395 ;
        RECT 139.155 118.255 139.415 119.395 ;
        RECT 139.585 118.245 139.915 119.225 ;
        RECT 140.085 118.255 140.365 119.395 ;
        RECT 140.535 118.885 140.795 119.395 ;
        RECT 139.675 118.205 139.850 118.245 ;
        RECT 137.650 117.525 138.005 118.085 ;
        RECT 139.175 117.835 139.510 118.085 ;
        RECT 139.680 117.645 139.850 118.205 ;
        RECT 140.020 117.815 140.355 118.085 ;
        RECT 140.535 117.835 140.875 118.715 ;
        RECT 141.045 118.005 141.215 119.225 ;
        RECT 141.455 118.890 142.070 119.395 ;
        RECT 141.455 118.355 141.705 118.720 ;
        RECT 141.875 118.715 142.070 118.890 ;
        RECT 142.240 118.885 142.715 119.225 ;
        RECT 142.885 118.850 143.100 119.395 ;
        RECT 141.875 118.525 142.205 118.715 ;
        RECT 142.425 118.355 143.140 118.650 ;
        RECT 143.310 118.525 143.585 119.225 ;
        RECT 141.455 118.185 143.245 118.355 ;
        RECT 141.045 117.755 141.840 118.005 ;
        RECT 141.045 117.665 141.295 117.755 ;
        RECT 136.755 116.845 136.970 117.355 ;
        RECT 137.200 117.025 137.480 117.355 ;
        RECT 137.660 116.845 137.900 117.355 ;
        RECT 138.695 116.845 138.985 117.570 ;
        RECT 139.155 117.015 139.850 117.645 ;
        RECT 140.055 116.845 140.365 117.645 ;
        RECT 140.535 116.845 140.795 117.665 ;
        RECT 140.965 117.245 141.295 117.665 ;
        RECT 142.010 117.330 142.265 118.185 ;
        RECT 141.475 117.065 142.265 117.330 ;
        RECT 142.435 117.485 142.845 118.005 ;
        RECT 143.015 117.755 143.245 118.185 ;
        RECT 143.415 117.495 143.585 118.525 ;
        RECT 142.435 117.065 142.635 117.485 ;
        RECT 142.825 116.845 143.155 117.305 ;
        RECT 143.325 117.015 143.585 117.495 ;
        RECT 143.755 118.255 144.140 119.225 ;
        RECT 144.310 118.935 144.635 119.395 ;
        RECT 145.155 118.765 145.435 119.225 ;
        RECT 144.310 118.545 145.435 118.765 ;
        RECT 143.755 117.585 144.035 118.255 ;
        RECT 144.310 118.085 144.760 118.545 ;
        RECT 145.625 118.375 146.025 119.225 ;
        RECT 146.425 118.935 146.695 119.395 ;
        RECT 146.865 118.765 147.150 119.225 ;
        RECT 144.205 117.755 144.760 118.085 ;
        RECT 144.930 117.815 146.025 118.375 ;
        RECT 144.310 117.645 144.760 117.755 ;
        RECT 143.755 117.015 144.140 117.585 ;
        RECT 144.310 117.475 145.435 117.645 ;
        RECT 144.310 116.845 144.635 117.305 ;
        RECT 145.155 117.015 145.435 117.475 ;
        RECT 145.625 117.015 146.025 117.815 ;
        RECT 146.195 118.545 147.150 118.765 ;
        RECT 146.195 117.645 146.405 118.545 ;
        RECT 146.575 117.815 147.265 118.375 ;
        RECT 147.495 118.335 147.825 119.180 ;
        RECT 147.995 118.385 148.165 119.395 ;
        RECT 148.335 118.665 148.675 119.225 ;
        RECT 148.905 118.895 149.220 119.395 ;
        RECT 149.400 118.925 150.285 119.095 ;
        RECT 147.435 118.255 147.825 118.335 ;
        RECT 148.335 118.290 149.230 118.665 ;
        RECT 147.435 118.205 147.650 118.255 ;
        RECT 146.195 117.475 147.150 117.645 ;
        RECT 147.435 117.625 147.605 118.205 ;
        RECT 148.335 118.085 148.525 118.290 ;
        RECT 149.400 118.085 149.570 118.925 ;
        RECT 150.510 118.895 150.760 119.225 ;
        RECT 147.775 117.755 148.525 118.085 ;
        RECT 148.695 117.755 149.570 118.085 ;
        RECT 147.435 117.585 147.660 117.625 ;
        RECT 148.325 117.585 148.525 117.755 ;
        RECT 147.435 117.500 147.815 117.585 ;
        RECT 146.425 116.845 146.695 117.305 ;
        RECT 146.865 117.015 147.150 117.475 ;
        RECT 147.485 117.065 147.815 117.500 ;
        RECT 147.985 116.845 148.155 117.455 ;
        RECT 148.325 117.060 148.655 117.585 ;
        RECT 148.915 116.845 149.125 117.375 ;
        RECT 149.400 117.295 149.570 117.755 ;
        RECT 149.740 117.795 150.060 118.755 ;
        RECT 150.230 118.005 150.420 118.725 ;
        RECT 150.590 117.825 150.760 118.895 ;
        RECT 150.930 118.595 151.100 119.395 ;
        RECT 151.270 118.950 152.375 119.120 ;
        RECT 151.270 118.335 151.440 118.950 ;
        RECT 152.585 118.800 152.835 119.225 ;
        RECT 153.005 118.935 153.270 119.395 ;
        RECT 151.610 118.415 152.140 118.780 ;
        RECT 152.585 118.670 152.890 118.800 ;
        RECT 150.930 118.245 151.440 118.335 ;
        RECT 150.930 118.075 151.800 118.245 ;
        RECT 150.930 118.005 151.100 118.075 ;
        RECT 151.220 117.825 151.420 117.855 ;
        RECT 149.740 117.465 150.205 117.795 ;
        RECT 150.590 117.525 151.420 117.825 ;
        RECT 150.590 117.295 150.760 117.525 ;
        RECT 149.400 117.125 150.185 117.295 ;
        RECT 150.355 117.125 150.760 117.295 ;
        RECT 150.940 116.845 151.310 117.345 ;
        RECT 151.630 117.295 151.800 118.075 ;
        RECT 151.970 117.715 152.140 118.415 ;
        RECT 152.310 117.885 152.550 118.480 ;
        RECT 151.970 117.495 152.495 117.715 ;
        RECT 152.720 117.565 152.890 118.670 ;
        RECT 152.665 117.435 152.890 117.565 ;
        RECT 153.060 117.475 153.340 118.425 ;
        RECT 152.665 117.295 152.835 117.435 ;
        RECT 151.630 117.125 152.305 117.295 ;
        RECT 152.500 117.125 152.835 117.295 ;
        RECT 153.005 116.845 153.255 117.305 ;
        RECT 153.510 117.105 153.695 119.225 ;
        RECT 153.865 118.895 154.195 119.395 ;
        RECT 154.365 118.725 154.535 119.225 ;
        RECT 153.870 118.555 154.535 118.725 ;
        RECT 153.870 117.565 154.100 118.555 ;
        RECT 154.270 117.735 154.620 118.385 ;
        RECT 155.715 118.305 156.925 119.395 ;
        RECT 155.715 117.765 156.235 118.305 ;
        RECT 156.405 117.595 156.925 118.135 ;
        RECT 153.870 117.395 154.535 117.565 ;
        RECT 153.865 116.845 154.195 117.225 ;
        RECT 154.365 117.105 154.535 117.395 ;
        RECT 155.715 116.845 156.925 117.595 ;
        RECT 22.690 116.675 157.010 116.845 ;
        RECT 22.775 115.925 23.985 116.675 ;
        RECT 25.240 116.165 25.480 116.675 ;
        RECT 25.660 116.165 25.940 116.495 ;
        RECT 26.170 116.165 26.385 116.675 ;
        RECT 22.775 115.385 23.295 115.925 ;
        RECT 23.465 115.215 23.985 115.755 ;
        RECT 25.135 115.435 25.490 115.995 ;
        RECT 25.660 115.265 25.830 116.165 ;
        RECT 26.000 115.435 26.265 115.995 ;
        RECT 26.555 115.935 27.170 116.505 ;
        RECT 26.515 115.265 26.685 115.765 ;
        RECT 22.775 114.125 23.985 115.215 ;
        RECT 25.260 115.095 26.685 115.265 ;
        RECT 25.260 114.920 25.650 115.095 ;
        RECT 26.135 114.125 26.465 114.925 ;
        RECT 26.855 114.915 27.170 115.935 ;
        RECT 27.580 115.895 28.080 116.505 ;
        RECT 27.375 115.435 27.725 115.685 ;
        RECT 27.910 115.265 28.080 115.895 ;
        RECT 28.710 116.025 29.040 116.505 ;
        RECT 29.210 116.215 29.435 116.675 ;
        RECT 29.605 116.025 29.935 116.505 ;
        RECT 28.710 115.855 29.935 116.025 ;
        RECT 30.125 115.875 30.375 116.675 ;
        RECT 30.545 115.875 30.885 116.505 ;
        RECT 31.170 116.045 31.455 116.505 ;
        RECT 31.625 116.215 31.895 116.675 ;
        RECT 31.170 115.875 32.125 116.045 ;
        RECT 28.250 115.485 28.580 115.685 ;
        RECT 28.750 115.485 29.080 115.685 ;
        RECT 29.250 115.485 29.670 115.685 ;
        RECT 29.845 115.515 30.540 115.685 ;
        RECT 29.845 115.265 30.015 115.515 ;
        RECT 30.710 115.315 30.885 115.875 ;
        RECT 30.655 115.265 30.885 115.315 ;
        RECT 26.635 114.295 27.170 114.915 ;
        RECT 27.580 115.095 30.015 115.265 ;
        RECT 27.580 114.295 27.910 115.095 ;
        RECT 28.080 114.125 28.410 114.925 ;
        RECT 28.710 114.295 29.040 115.095 ;
        RECT 29.685 114.125 29.935 114.925 ;
        RECT 30.205 114.125 30.375 115.265 ;
        RECT 30.545 114.295 30.885 115.265 ;
        RECT 31.055 115.145 31.745 115.705 ;
        RECT 31.915 114.975 32.125 115.875 ;
        RECT 31.170 114.755 32.125 114.975 ;
        RECT 32.295 115.705 32.695 116.505 ;
        RECT 32.885 116.045 33.165 116.505 ;
        RECT 33.685 116.215 34.010 116.675 ;
        RECT 32.885 115.875 34.010 116.045 ;
        RECT 34.180 115.935 34.565 116.505 ;
        RECT 34.745 116.175 35.075 116.675 ;
        RECT 35.275 116.105 35.445 116.455 ;
        RECT 35.645 116.275 35.975 116.675 ;
        RECT 36.145 116.105 36.315 116.455 ;
        RECT 36.485 116.275 36.865 116.675 ;
        RECT 33.560 115.765 34.010 115.875 ;
        RECT 32.295 115.145 33.390 115.705 ;
        RECT 33.560 115.435 34.115 115.765 ;
        RECT 31.170 114.295 31.455 114.755 ;
        RECT 31.625 114.125 31.895 114.585 ;
        RECT 32.295 114.295 32.695 115.145 ;
        RECT 33.560 114.975 34.010 115.435 ;
        RECT 34.285 115.265 34.565 115.935 ;
        RECT 34.740 115.435 35.090 116.005 ;
        RECT 35.275 115.935 36.885 116.105 ;
        RECT 37.055 116.000 37.325 116.345 ;
        RECT 36.715 115.765 36.885 115.935 ;
        RECT 32.885 114.755 34.010 114.975 ;
        RECT 32.885 114.295 33.165 114.755 ;
        RECT 33.685 114.125 34.010 114.585 ;
        RECT 34.180 114.295 34.565 115.265 ;
        RECT 34.740 114.975 35.060 115.265 ;
        RECT 35.260 115.145 35.970 115.765 ;
        RECT 36.140 115.435 36.545 115.765 ;
        RECT 36.715 115.435 36.985 115.765 ;
        RECT 36.715 115.265 36.885 115.435 ;
        RECT 37.155 115.265 37.325 116.000 ;
        RECT 37.585 116.125 37.755 116.415 ;
        RECT 37.925 116.295 38.255 116.675 ;
        RECT 37.585 115.955 38.250 116.125 ;
        RECT 36.160 115.095 36.885 115.265 ;
        RECT 36.160 114.975 36.330 115.095 ;
        RECT 34.740 114.805 36.330 114.975 ;
        RECT 34.740 114.345 36.395 114.635 ;
        RECT 36.565 114.125 36.845 114.925 ;
        RECT 37.055 114.295 37.325 115.265 ;
        RECT 37.500 115.135 37.850 115.785 ;
        RECT 38.020 114.965 38.250 115.955 ;
        RECT 37.585 114.795 38.250 114.965 ;
        RECT 37.585 114.295 37.755 114.795 ;
        RECT 37.925 114.125 38.255 114.625 ;
        RECT 38.425 114.295 38.610 116.415 ;
        RECT 38.865 116.215 39.115 116.675 ;
        RECT 39.285 116.225 39.620 116.395 ;
        RECT 39.815 116.225 40.490 116.395 ;
        RECT 39.285 116.085 39.455 116.225 ;
        RECT 38.780 115.095 39.060 116.045 ;
        RECT 39.230 115.955 39.455 116.085 ;
        RECT 39.230 114.850 39.400 115.955 ;
        RECT 39.625 115.805 40.150 116.025 ;
        RECT 39.570 115.040 39.810 115.635 ;
        RECT 39.980 115.105 40.150 115.805 ;
        RECT 40.320 115.445 40.490 116.225 ;
        RECT 40.810 116.175 41.180 116.675 ;
        RECT 41.360 116.225 41.765 116.395 ;
        RECT 41.935 116.225 42.720 116.395 ;
        RECT 41.360 115.995 41.530 116.225 ;
        RECT 40.700 115.695 41.530 115.995 ;
        RECT 41.915 115.725 42.380 116.055 ;
        RECT 40.700 115.665 40.900 115.695 ;
        RECT 41.020 115.445 41.190 115.515 ;
        RECT 40.320 115.275 41.190 115.445 ;
        RECT 40.680 115.185 41.190 115.275 ;
        RECT 39.230 114.720 39.535 114.850 ;
        RECT 39.980 114.740 40.510 115.105 ;
        RECT 38.850 114.125 39.115 114.585 ;
        RECT 39.285 114.295 39.535 114.720 ;
        RECT 40.680 114.570 40.850 115.185 ;
        RECT 39.745 114.400 40.850 114.570 ;
        RECT 41.020 114.125 41.190 114.925 ;
        RECT 41.360 114.625 41.530 115.695 ;
        RECT 41.700 114.795 41.890 115.515 ;
        RECT 42.060 114.765 42.380 115.725 ;
        RECT 42.550 115.765 42.720 116.225 ;
        RECT 42.995 116.145 43.205 116.675 ;
        RECT 43.465 115.935 43.795 116.460 ;
        RECT 43.965 116.065 44.135 116.675 ;
        RECT 44.305 116.020 44.635 116.455 ;
        RECT 44.305 115.935 44.685 116.020 ;
        RECT 43.595 115.765 43.795 115.935 ;
        RECT 44.460 115.895 44.685 115.935 ;
        RECT 45.060 115.895 45.560 116.505 ;
        RECT 42.550 115.435 43.425 115.765 ;
        RECT 43.595 115.435 44.345 115.765 ;
        RECT 41.360 114.295 41.610 114.625 ;
        RECT 42.550 114.595 42.720 115.435 ;
        RECT 43.595 115.230 43.785 115.435 ;
        RECT 44.515 115.315 44.685 115.895 ;
        RECT 44.855 115.435 45.205 115.685 ;
        RECT 44.470 115.265 44.685 115.315 ;
        RECT 45.390 115.265 45.560 115.895 ;
        RECT 46.190 116.025 46.520 116.505 ;
        RECT 46.690 116.215 46.915 116.675 ;
        RECT 47.085 116.025 47.415 116.505 ;
        RECT 46.190 115.855 47.415 116.025 ;
        RECT 47.605 115.875 47.855 116.675 ;
        RECT 48.025 115.875 48.365 116.505 ;
        RECT 48.535 115.950 48.825 116.675 ;
        RECT 48.135 115.825 48.365 115.875 ;
        RECT 45.730 115.485 46.060 115.685 ;
        RECT 46.230 115.485 46.560 115.685 ;
        RECT 46.730 115.485 47.150 115.685 ;
        RECT 47.325 115.515 48.020 115.685 ;
        RECT 47.325 115.265 47.495 115.515 ;
        RECT 48.190 115.265 48.365 115.825 ;
        RECT 48.995 115.905 50.665 116.675 ;
        RECT 50.885 116.020 51.215 116.455 ;
        RECT 51.385 116.065 51.555 116.675 ;
        RECT 50.835 115.935 51.215 116.020 ;
        RECT 51.725 115.935 52.055 116.460 ;
        RECT 52.315 116.145 52.525 116.675 ;
        RECT 52.800 116.225 53.585 116.395 ;
        RECT 53.755 116.225 54.160 116.395 ;
        RECT 48.995 115.385 49.745 115.905 ;
        RECT 50.835 115.895 51.060 115.935 ;
        RECT 42.890 114.855 43.785 115.230 ;
        RECT 44.295 115.185 44.685 115.265 ;
        RECT 41.835 114.425 42.720 114.595 ;
        RECT 42.900 114.125 43.215 114.625 ;
        RECT 43.445 114.295 43.785 114.855 ;
        RECT 43.955 114.125 44.125 115.135 ;
        RECT 44.295 114.340 44.625 115.185 ;
        RECT 45.060 115.095 47.495 115.265 ;
        RECT 45.060 114.295 45.390 115.095 ;
        RECT 45.560 114.125 45.890 114.925 ;
        RECT 46.190 114.295 46.520 115.095 ;
        RECT 47.165 114.125 47.415 114.925 ;
        RECT 47.685 114.125 47.855 115.265 ;
        RECT 48.025 114.295 48.365 115.265 ;
        RECT 48.535 114.125 48.825 115.290 ;
        RECT 49.915 115.215 50.665 115.735 ;
        RECT 48.995 114.125 50.665 115.215 ;
        RECT 50.835 115.315 51.005 115.895 ;
        RECT 51.725 115.765 51.925 115.935 ;
        RECT 52.800 115.765 52.970 116.225 ;
        RECT 51.175 115.435 51.925 115.765 ;
        RECT 52.095 115.435 52.970 115.765 ;
        RECT 50.835 115.265 51.050 115.315 ;
        RECT 50.835 115.185 51.225 115.265 ;
        RECT 50.895 114.340 51.225 115.185 ;
        RECT 51.735 115.230 51.925 115.435 ;
        RECT 51.395 114.125 51.565 115.135 ;
        RECT 51.735 114.855 52.630 115.230 ;
        RECT 51.735 114.295 52.075 114.855 ;
        RECT 52.305 114.125 52.620 114.625 ;
        RECT 52.800 114.595 52.970 115.435 ;
        RECT 53.140 115.725 53.605 116.055 ;
        RECT 53.990 115.995 54.160 116.225 ;
        RECT 54.340 116.175 54.710 116.675 ;
        RECT 55.030 116.225 55.705 116.395 ;
        RECT 55.900 116.225 56.235 116.395 ;
        RECT 53.140 114.765 53.460 115.725 ;
        RECT 53.990 115.695 54.820 115.995 ;
        RECT 53.630 114.795 53.820 115.515 ;
        RECT 53.990 114.625 54.160 115.695 ;
        RECT 54.620 115.665 54.820 115.695 ;
        RECT 54.330 115.445 54.500 115.515 ;
        RECT 55.030 115.445 55.200 116.225 ;
        RECT 56.065 116.085 56.235 116.225 ;
        RECT 56.405 116.215 56.655 116.675 ;
        RECT 54.330 115.275 55.200 115.445 ;
        RECT 55.370 115.805 55.895 116.025 ;
        RECT 56.065 115.955 56.290 116.085 ;
        RECT 54.330 115.185 54.840 115.275 ;
        RECT 52.800 114.425 53.685 114.595 ;
        RECT 53.910 114.295 54.160 114.625 ;
        RECT 54.330 114.125 54.500 114.925 ;
        RECT 54.670 114.570 54.840 115.185 ;
        RECT 55.370 115.105 55.540 115.805 ;
        RECT 55.010 114.740 55.540 115.105 ;
        RECT 55.710 115.040 55.950 115.635 ;
        RECT 56.120 114.850 56.290 115.955 ;
        RECT 56.460 115.095 56.740 116.045 ;
        RECT 55.985 114.720 56.290 114.850 ;
        RECT 54.670 114.400 55.775 114.570 ;
        RECT 55.985 114.295 56.235 114.720 ;
        RECT 56.405 114.125 56.670 114.585 ;
        RECT 56.910 114.295 57.095 116.415 ;
        RECT 57.265 116.295 57.595 116.675 ;
        RECT 57.765 116.125 57.935 116.415 ;
        RECT 57.270 115.955 57.935 116.125 ;
        RECT 57.270 114.965 57.500 115.955 ;
        RECT 58.235 115.855 58.465 116.675 ;
        RECT 58.635 115.875 58.965 116.505 ;
        RECT 57.670 115.135 58.020 115.785 ;
        RECT 58.215 115.435 58.545 115.685 ;
        RECT 58.715 115.275 58.965 115.875 ;
        RECT 59.135 115.855 59.345 116.675 ;
        RECT 59.575 115.905 61.245 116.675 ;
        RECT 59.575 115.385 60.325 115.905 ;
        RECT 61.430 115.895 61.725 116.675 ;
        RECT 62.285 116.145 62.630 116.505 ;
        RECT 63.090 116.315 63.420 116.675 ;
        RECT 63.625 116.145 63.945 116.505 ;
        RECT 62.285 115.975 63.945 116.145 ;
        RECT 57.270 114.795 57.935 114.965 ;
        RECT 57.265 114.125 57.595 114.625 ;
        RECT 57.765 114.295 57.935 114.795 ;
        RECT 58.235 114.125 58.465 115.265 ;
        RECT 58.635 114.295 58.965 115.275 ;
        RECT 59.135 114.125 59.345 115.265 ;
        RECT 60.495 115.215 61.245 115.735 ;
        RECT 59.575 114.125 61.245 115.215 ;
        RECT 61.475 115.265 61.975 115.725 ;
        RECT 62.145 115.435 62.755 115.765 ;
        RECT 62.935 115.515 63.265 115.685 ;
        RECT 62.935 115.265 63.260 115.515 ;
        RECT 61.475 115.085 63.260 115.265 ;
        RECT 61.440 114.735 63.475 114.905 ;
        RECT 61.440 114.655 62.550 114.735 ;
        RECT 61.440 114.295 61.700 114.655 ;
        RECT 61.870 114.125 62.200 114.485 ;
        RECT 62.380 114.295 62.550 114.655 ;
        RECT 62.805 114.125 62.975 114.565 ;
        RECT 63.145 114.475 63.475 114.735 ;
        RECT 63.645 114.645 63.945 115.975 ;
        RECT 64.125 115.935 64.455 116.675 ;
        RECT 65.095 115.855 65.355 116.675 ;
        RECT 65.525 115.855 65.855 116.275 ;
        RECT 66.035 116.105 66.295 116.505 ;
        RECT 66.465 116.275 66.795 116.675 ;
        RECT 66.965 116.105 67.135 116.455 ;
        RECT 67.305 116.275 67.680 116.675 ;
        RECT 66.035 115.935 67.700 116.105 ;
        RECT 67.870 116.000 68.145 116.345 ;
        RECT 65.605 115.765 65.855 115.855 ;
        RECT 67.530 115.765 67.700 115.935 ;
        RECT 64.130 115.135 64.405 115.765 ;
        RECT 65.100 115.435 65.435 115.685 ;
        RECT 65.605 115.435 66.320 115.765 ;
        RECT 66.535 115.435 67.360 115.765 ;
        RECT 67.530 115.435 67.805 115.765 ;
        RECT 64.115 114.475 64.420 114.965 ;
        RECT 63.145 114.295 64.420 114.475 ;
        RECT 65.095 114.125 65.355 115.265 ;
        RECT 65.605 114.875 65.775 115.435 ;
        RECT 66.035 114.975 66.365 115.265 ;
        RECT 66.535 115.145 66.780 115.435 ;
        RECT 67.530 115.265 67.700 115.435 ;
        RECT 67.975 115.265 68.145 116.000 ;
        RECT 69.050 115.865 69.295 116.470 ;
        RECT 69.515 116.140 70.025 116.675 ;
        RECT 67.040 115.095 67.700 115.265 ;
        RECT 67.040 114.975 67.210 115.095 ;
        RECT 66.035 114.805 67.210 114.975 ;
        RECT 65.595 114.305 67.210 114.635 ;
        RECT 67.380 114.125 67.660 114.925 ;
        RECT 67.870 114.295 68.145 115.265 ;
        RECT 68.775 115.695 70.005 115.865 ;
        RECT 68.775 114.885 69.115 115.695 ;
        RECT 69.285 115.130 70.035 115.320 ;
        RECT 68.775 114.475 69.290 114.885 ;
        RECT 69.525 114.125 69.695 114.885 ;
        RECT 69.865 114.465 70.035 115.130 ;
        RECT 70.205 115.145 70.395 116.505 ;
        RECT 70.565 116.335 70.840 116.505 ;
        RECT 70.565 116.165 70.845 116.335 ;
        RECT 70.565 115.345 70.840 116.165 ;
        RECT 71.030 116.140 71.560 116.505 ;
        RECT 71.985 116.275 72.315 116.675 ;
        RECT 71.385 116.105 71.560 116.140 ;
        RECT 71.045 115.145 71.215 115.945 ;
        RECT 70.205 114.975 71.215 115.145 ;
        RECT 71.385 115.935 72.315 116.105 ;
        RECT 72.485 115.935 72.740 116.505 ;
        RECT 71.385 114.805 71.555 115.935 ;
        RECT 72.145 115.765 72.315 115.935 ;
        RECT 70.430 114.635 71.555 114.805 ;
        RECT 71.725 115.435 71.920 115.765 ;
        RECT 72.145 115.435 72.400 115.765 ;
        RECT 71.725 114.465 71.895 115.435 ;
        RECT 72.570 115.265 72.740 115.935 ;
        RECT 69.865 114.295 71.895 114.465 ;
        RECT 72.065 114.125 72.235 115.265 ;
        RECT 72.405 114.295 72.740 115.265 ;
        RECT 72.915 116.000 73.175 116.505 ;
        RECT 73.355 116.295 73.685 116.675 ;
        RECT 73.865 116.125 74.035 116.505 ;
        RECT 72.915 115.200 73.085 116.000 ;
        RECT 73.370 115.955 74.035 116.125 ;
        RECT 73.370 115.700 73.540 115.955 ;
        RECT 74.295 115.950 74.585 116.675 ;
        RECT 75.305 116.125 75.475 116.415 ;
        RECT 75.645 116.295 75.975 116.675 ;
        RECT 75.305 115.955 75.970 116.125 ;
        RECT 73.255 115.370 73.540 115.700 ;
        RECT 73.775 115.405 74.105 115.775 ;
        RECT 73.370 115.225 73.540 115.370 ;
        RECT 72.915 114.295 73.185 115.200 ;
        RECT 73.370 115.055 74.035 115.225 ;
        RECT 73.355 114.125 73.685 114.885 ;
        RECT 73.865 114.295 74.035 115.055 ;
        RECT 74.295 114.125 74.585 115.290 ;
        RECT 75.220 115.135 75.570 115.785 ;
        RECT 75.740 114.965 75.970 115.955 ;
        RECT 75.305 114.795 75.970 114.965 ;
        RECT 75.305 114.295 75.475 114.795 ;
        RECT 75.645 114.125 75.975 114.625 ;
        RECT 76.145 114.295 76.330 116.415 ;
        RECT 76.585 116.215 76.835 116.675 ;
        RECT 77.005 116.225 77.340 116.395 ;
        RECT 77.535 116.225 78.210 116.395 ;
        RECT 77.005 116.085 77.175 116.225 ;
        RECT 76.500 115.095 76.780 116.045 ;
        RECT 76.950 115.955 77.175 116.085 ;
        RECT 76.950 114.850 77.120 115.955 ;
        RECT 77.345 115.805 77.870 116.025 ;
        RECT 77.290 115.040 77.530 115.635 ;
        RECT 77.700 115.105 77.870 115.805 ;
        RECT 78.040 115.445 78.210 116.225 ;
        RECT 78.530 116.175 78.900 116.675 ;
        RECT 79.080 116.225 79.485 116.395 ;
        RECT 79.655 116.225 80.440 116.395 ;
        RECT 79.080 115.995 79.250 116.225 ;
        RECT 78.420 115.695 79.250 115.995 ;
        RECT 79.635 115.725 80.100 116.055 ;
        RECT 78.420 115.665 78.620 115.695 ;
        RECT 78.740 115.445 78.910 115.515 ;
        RECT 78.040 115.275 78.910 115.445 ;
        RECT 78.400 115.185 78.910 115.275 ;
        RECT 76.950 114.720 77.255 114.850 ;
        RECT 77.700 114.740 78.230 115.105 ;
        RECT 76.570 114.125 76.835 114.585 ;
        RECT 77.005 114.295 77.255 114.720 ;
        RECT 78.400 114.570 78.570 115.185 ;
        RECT 77.465 114.400 78.570 114.570 ;
        RECT 78.740 114.125 78.910 114.925 ;
        RECT 79.080 114.625 79.250 115.695 ;
        RECT 79.420 114.795 79.610 115.515 ;
        RECT 79.780 114.765 80.100 115.725 ;
        RECT 80.270 115.765 80.440 116.225 ;
        RECT 80.715 116.145 80.925 116.675 ;
        RECT 81.185 115.935 81.515 116.460 ;
        RECT 81.685 116.065 81.855 116.675 ;
        RECT 82.025 116.020 82.355 116.455 ;
        RECT 83.495 116.165 83.800 116.675 ;
        RECT 82.025 115.935 82.405 116.020 ;
        RECT 81.315 115.765 81.515 115.935 ;
        RECT 82.180 115.895 82.405 115.935 ;
        RECT 80.270 115.435 81.145 115.765 ;
        RECT 81.315 115.435 82.065 115.765 ;
        RECT 79.080 114.295 79.330 114.625 ;
        RECT 80.270 114.595 80.440 115.435 ;
        RECT 81.315 115.230 81.505 115.435 ;
        RECT 82.235 115.315 82.405 115.895 ;
        RECT 83.495 115.435 83.810 115.995 ;
        RECT 83.980 115.685 84.230 116.495 ;
        RECT 84.400 116.150 84.660 116.675 ;
        RECT 84.840 115.685 85.090 116.495 ;
        RECT 85.260 116.115 85.520 116.675 ;
        RECT 85.690 116.025 85.950 116.480 ;
        RECT 86.120 116.195 86.380 116.675 ;
        RECT 86.550 116.025 86.810 116.480 ;
        RECT 86.980 116.195 87.240 116.675 ;
        RECT 87.410 116.025 87.670 116.480 ;
        RECT 87.840 116.195 88.085 116.675 ;
        RECT 88.255 116.025 88.530 116.480 ;
        RECT 88.700 116.195 88.945 116.675 ;
        RECT 89.115 116.025 89.375 116.480 ;
        RECT 89.555 116.195 89.805 116.675 ;
        RECT 89.975 116.025 90.235 116.480 ;
        RECT 90.415 116.195 90.665 116.675 ;
        RECT 90.835 116.025 91.095 116.480 ;
        RECT 91.275 116.195 91.535 116.675 ;
        RECT 91.705 116.025 91.965 116.480 ;
        RECT 92.135 116.195 92.435 116.675 ;
        RECT 85.690 115.995 92.435 116.025 ;
        RECT 85.690 115.855 92.465 115.995 ;
        RECT 92.715 115.865 92.955 116.675 ;
        RECT 93.125 115.865 93.455 116.505 ;
        RECT 93.625 115.865 93.895 116.675 ;
        RECT 94.075 115.905 95.745 116.675 ;
        RECT 96.465 116.125 96.635 116.505 ;
        RECT 96.815 116.295 97.145 116.675 ;
        RECT 96.465 115.955 97.130 116.125 ;
        RECT 97.325 116.000 97.585 116.505 ;
        RECT 91.270 115.825 92.465 115.855 ;
        RECT 83.980 115.435 91.100 115.685 ;
        RECT 82.190 115.265 82.405 115.315 ;
        RECT 80.610 114.855 81.505 115.230 ;
        RECT 82.015 115.185 82.405 115.265 ;
        RECT 79.555 114.425 80.440 114.595 ;
        RECT 80.620 114.125 80.935 114.625 ;
        RECT 81.165 114.295 81.505 114.855 ;
        RECT 81.675 114.125 81.845 115.135 ;
        RECT 82.015 114.340 82.345 115.185 ;
        RECT 83.505 114.125 83.800 114.935 ;
        RECT 83.980 114.295 84.225 115.435 ;
        RECT 84.400 114.125 84.660 114.935 ;
        RECT 84.840 114.300 85.090 115.435 ;
        RECT 91.270 115.265 92.435 115.825 ;
        RECT 92.695 115.435 93.045 115.685 ;
        RECT 93.215 115.265 93.385 115.865 ;
        RECT 93.555 115.435 93.905 115.685 ;
        RECT 94.075 115.385 94.825 115.905 ;
        RECT 85.690 115.040 92.435 115.265 ;
        RECT 92.705 115.095 93.385 115.265 ;
        RECT 85.690 115.025 91.095 115.040 ;
        RECT 85.260 114.130 85.520 114.925 ;
        RECT 85.690 114.300 85.950 115.025 ;
        RECT 86.120 114.130 86.380 114.855 ;
        RECT 86.550 114.300 86.810 115.025 ;
        RECT 86.980 114.130 87.240 114.855 ;
        RECT 87.410 114.300 87.670 115.025 ;
        RECT 87.840 114.130 88.100 114.855 ;
        RECT 88.270 114.300 88.530 115.025 ;
        RECT 88.700 114.130 88.945 114.855 ;
        RECT 89.115 114.300 89.375 115.025 ;
        RECT 89.560 114.130 89.805 114.855 ;
        RECT 89.975 114.300 90.235 115.025 ;
        RECT 90.420 114.130 90.665 114.855 ;
        RECT 90.835 114.300 91.095 115.025 ;
        RECT 91.280 114.130 91.535 114.855 ;
        RECT 91.705 114.300 91.995 115.040 ;
        RECT 85.260 114.125 91.535 114.130 ;
        RECT 92.165 114.125 92.435 114.870 ;
        RECT 92.705 114.310 93.035 115.095 ;
        RECT 93.565 114.125 93.895 115.265 ;
        RECT 94.995 115.215 95.745 115.735 ;
        RECT 96.395 115.405 96.725 115.775 ;
        RECT 96.960 115.700 97.130 115.955 ;
        RECT 96.960 115.370 97.245 115.700 ;
        RECT 96.960 115.225 97.130 115.370 ;
        RECT 94.075 114.125 95.745 115.215 ;
        RECT 96.465 115.055 97.130 115.225 ;
        RECT 97.415 115.200 97.585 116.000 ;
        RECT 97.955 116.045 98.285 116.405 ;
        RECT 98.905 116.215 99.155 116.675 ;
        RECT 99.325 116.215 99.885 116.505 ;
        RECT 97.955 115.855 99.345 116.045 ;
        RECT 99.175 115.765 99.345 115.855 ;
        RECT 96.465 114.295 96.635 115.055 ;
        RECT 96.815 114.125 97.145 114.885 ;
        RECT 97.315 114.295 97.585 115.200 ;
        RECT 97.770 115.435 98.445 115.685 ;
        RECT 98.665 115.435 99.005 115.685 ;
        RECT 99.175 115.435 99.465 115.765 ;
        RECT 97.770 115.075 98.035 115.435 ;
        RECT 99.175 115.185 99.345 115.435 ;
        RECT 98.405 115.015 99.345 115.185 ;
        RECT 97.955 114.125 98.235 114.795 ;
        RECT 98.405 114.465 98.705 115.015 ;
        RECT 99.635 114.845 99.885 116.215 ;
        RECT 100.055 115.950 100.345 116.675 ;
        RECT 100.565 116.020 100.895 116.455 ;
        RECT 101.065 116.065 101.235 116.675 ;
        RECT 100.515 115.935 100.895 116.020 ;
        RECT 101.405 115.935 101.735 116.460 ;
        RECT 101.995 116.145 102.205 116.675 ;
        RECT 102.480 116.225 103.265 116.395 ;
        RECT 103.435 116.225 103.840 116.395 ;
        RECT 100.515 115.895 100.740 115.935 ;
        RECT 100.515 115.315 100.685 115.895 ;
        RECT 101.405 115.765 101.605 115.935 ;
        RECT 102.480 115.765 102.650 116.225 ;
        RECT 100.855 115.435 101.605 115.765 ;
        RECT 101.775 115.435 102.650 115.765 ;
        RECT 98.905 114.125 99.235 114.845 ;
        RECT 99.425 114.295 99.885 114.845 ;
        RECT 100.055 114.125 100.345 115.290 ;
        RECT 100.515 115.265 100.730 115.315 ;
        RECT 100.515 115.185 100.905 115.265 ;
        RECT 100.575 114.340 100.905 115.185 ;
        RECT 101.415 115.230 101.605 115.435 ;
        RECT 101.075 114.125 101.245 115.135 ;
        RECT 101.415 114.855 102.310 115.230 ;
        RECT 101.415 114.295 101.755 114.855 ;
        RECT 101.985 114.125 102.300 114.625 ;
        RECT 102.480 114.595 102.650 115.435 ;
        RECT 102.820 115.725 103.285 116.055 ;
        RECT 103.670 115.995 103.840 116.225 ;
        RECT 104.020 116.175 104.390 116.675 ;
        RECT 104.710 116.225 105.385 116.395 ;
        RECT 105.580 116.225 105.915 116.395 ;
        RECT 102.820 114.765 103.140 115.725 ;
        RECT 103.670 115.695 104.500 115.995 ;
        RECT 103.310 114.795 103.500 115.515 ;
        RECT 103.670 114.625 103.840 115.695 ;
        RECT 104.300 115.665 104.500 115.695 ;
        RECT 104.010 115.445 104.180 115.515 ;
        RECT 104.710 115.445 104.880 116.225 ;
        RECT 105.745 116.085 105.915 116.225 ;
        RECT 106.085 116.215 106.335 116.675 ;
        RECT 104.010 115.275 104.880 115.445 ;
        RECT 105.050 115.805 105.575 116.025 ;
        RECT 105.745 115.955 105.970 116.085 ;
        RECT 104.010 115.185 104.520 115.275 ;
        RECT 102.480 114.425 103.365 114.595 ;
        RECT 103.590 114.295 103.840 114.625 ;
        RECT 104.010 114.125 104.180 114.925 ;
        RECT 104.350 114.570 104.520 115.185 ;
        RECT 105.050 115.105 105.220 115.805 ;
        RECT 104.690 114.740 105.220 115.105 ;
        RECT 105.390 115.040 105.630 115.635 ;
        RECT 105.800 114.850 105.970 115.955 ;
        RECT 106.140 115.095 106.420 116.045 ;
        RECT 105.665 114.720 105.970 114.850 ;
        RECT 104.350 114.400 105.455 114.570 ;
        RECT 105.665 114.295 105.915 114.720 ;
        RECT 106.085 114.125 106.350 114.585 ;
        RECT 106.590 114.295 106.775 116.415 ;
        RECT 106.945 116.295 107.275 116.675 ;
        RECT 107.445 116.125 107.615 116.415 ;
        RECT 106.950 115.955 107.615 116.125 ;
        RECT 108.425 116.125 108.595 116.415 ;
        RECT 108.765 116.295 109.095 116.675 ;
        RECT 108.425 115.955 109.090 116.125 ;
        RECT 106.950 114.965 107.180 115.955 ;
        RECT 107.350 115.135 107.700 115.785 ;
        RECT 108.340 115.135 108.690 115.785 ;
        RECT 108.860 114.965 109.090 115.955 ;
        RECT 106.950 114.795 107.615 114.965 ;
        RECT 106.945 114.125 107.275 114.625 ;
        RECT 107.445 114.295 107.615 114.795 ;
        RECT 108.425 114.795 109.090 114.965 ;
        RECT 108.425 114.295 108.595 114.795 ;
        RECT 108.765 114.125 109.095 114.625 ;
        RECT 109.265 114.295 109.450 116.415 ;
        RECT 109.705 116.215 109.955 116.675 ;
        RECT 110.125 116.225 110.460 116.395 ;
        RECT 110.655 116.225 111.330 116.395 ;
        RECT 110.125 116.085 110.295 116.225 ;
        RECT 109.620 115.095 109.900 116.045 ;
        RECT 110.070 115.955 110.295 116.085 ;
        RECT 110.070 114.850 110.240 115.955 ;
        RECT 110.465 115.805 110.990 116.025 ;
        RECT 110.410 115.040 110.650 115.635 ;
        RECT 110.820 115.105 110.990 115.805 ;
        RECT 111.160 115.445 111.330 116.225 ;
        RECT 111.650 116.175 112.020 116.675 ;
        RECT 112.200 116.225 112.605 116.395 ;
        RECT 112.775 116.225 113.560 116.395 ;
        RECT 112.200 115.995 112.370 116.225 ;
        RECT 111.540 115.695 112.370 115.995 ;
        RECT 112.755 115.725 113.220 116.055 ;
        RECT 111.540 115.665 111.740 115.695 ;
        RECT 111.860 115.445 112.030 115.515 ;
        RECT 111.160 115.275 112.030 115.445 ;
        RECT 111.520 115.185 112.030 115.275 ;
        RECT 110.070 114.720 110.375 114.850 ;
        RECT 110.820 114.740 111.350 115.105 ;
        RECT 109.690 114.125 109.955 114.585 ;
        RECT 110.125 114.295 110.375 114.720 ;
        RECT 111.520 114.570 111.690 115.185 ;
        RECT 110.585 114.400 111.690 114.570 ;
        RECT 111.860 114.125 112.030 114.925 ;
        RECT 112.200 114.625 112.370 115.695 ;
        RECT 112.540 114.795 112.730 115.515 ;
        RECT 112.900 114.765 113.220 115.725 ;
        RECT 113.390 115.765 113.560 116.225 ;
        RECT 113.835 116.145 114.045 116.675 ;
        RECT 114.305 115.935 114.635 116.460 ;
        RECT 114.805 116.065 114.975 116.675 ;
        RECT 115.145 116.020 115.475 116.455 ;
        RECT 115.145 115.935 115.525 116.020 ;
        RECT 114.435 115.765 114.635 115.935 ;
        RECT 115.300 115.895 115.525 115.935 ;
        RECT 113.390 115.435 114.265 115.765 ;
        RECT 114.435 115.435 115.185 115.765 ;
        RECT 112.200 114.295 112.450 114.625 ;
        RECT 113.390 114.595 113.560 115.435 ;
        RECT 114.435 115.230 114.625 115.435 ;
        RECT 115.355 115.315 115.525 115.895 ;
        RECT 115.310 115.265 115.525 115.315 ;
        RECT 113.730 114.855 114.625 115.230 ;
        RECT 115.135 115.185 115.525 115.265 ;
        RECT 115.700 115.935 115.955 116.505 ;
        RECT 116.125 116.275 116.455 116.675 ;
        RECT 116.880 116.140 117.410 116.505 ;
        RECT 116.880 116.105 117.055 116.140 ;
        RECT 116.125 115.935 117.055 116.105 ;
        RECT 115.700 115.265 115.870 115.935 ;
        RECT 116.125 115.765 116.295 115.935 ;
        RECT 116.040 115.435 116.295 115.765 ;
        RECT 116.520 115.435 116.715 115.765 ;
        RECT 112.675 114.425 113.560 114.595 ;
        RECT 113.740 114.125 114.055 114.625 ;
        RECT 114.285 114.295 114.625 114.855 ;
        RECT 114.795 114.125 114.965 115.135 ;
        RECT 115.135 114.340 115.465 115.185 ;
        RECT 115.700 114.295 116.035 115.265 ;
        RECT 116.205 114.125 116.375 115.265 ;
        RECT 116.545 114.465 116.715 115.435 ;
        RECT 116.885 114.805 117.055 115.935 ;
        RECT 117.225 115.145 117.395 115.945 ;
        RECT 117.600 115.655 117.875 116.505 ;
        RECT 117.595 115.485 117.875 115.655 ;
        RECT 117.600 115.345 117.875 115.485 ;
        RECT 118.045 115.145 118.235 116.505 ;
        RECT 118.415 116.140 118.925 116.675 ;
        RECT 119.145 115.865 119.390 116.470 ;
        RECT 120.110 115.865 120.355 116.470 ;
        RECT 120.575 116.140 121.085 116.675 ;
        RECT 118.435 115.695 119.665 115.865 ;
        RECT 117.225 114.975 118.235 115.145 ;
        RECT 118.405 115.130 119.155 115.320 ;
        RECT 116.885 114.635 118.010 114.805 ;
        RECT 118.405 114.465 118.575 115.130 ;
        RECT 119.325 114.885 119.665 115.695 ;
        RECT 116.545 114.295 118.575 114.465 ;
        RECT 118.745 114.125 118.915 114.885 ;
        RECT 119.150 114.475 119.665 114.885 ;
        RECT 119.835 115.695 121.065 115.865 ;
        RECT 119.835 114.885 120.175 115.695 ;
        RECT 120.345 115.130 121.095 115.320 ;
        RECT 119.835 114.475 120.350 114.885 ;
        RECT 120.585 114.125 120.755 114.885 ;
        RECT 120.925 114.465 121.095 115.130 ;
        RECT 121.265 115.145 121.455 116.505 ;
        RECT 121.625 115.655 121.900 116.505 ;
        RECT 122.090 116.140 122.620 116.505 ;
        RECT 123.045 116.275 123.375 116.675 ;
        RECT 122.445 116.105 122.620 116.140 ;
        RECT 121.625 115.485 121.905 115.655 ;
        RECT 121.625 115.345 121.900 115.485 ;
        RECT 122.105 115.145 122.275 115.945 ;
        RECT 121.265 114.975 122.275 115.145 ;
        RECT 122.445 115.935 123.375 116.105 ;
        RECT 123.545 115.935 123.800 116.505 ;
        RECT 122.445 114.805 122.615 115.935 ;
        RECT 123.205 115.765 123.375 115.935 ;
        RECT 121.490 114.635 122.615 114.805 ;
        RECT 122.785 115.435 122.980 115.765 ;
        RECT 123.205 115.435 123.460 115.765 ;
        RECT 122.785 114.465 122.955 115.435 ;
        RECT 123.630 115.265 123.800 115.935 ;
        RECT 123.975 115.905 125.645 116.675 ;
        RECT 125.815 115.950 126.105 116.675 ;
        RECT 126.365 116.125 126.535 116.415 ;
        RECT 126.705 116.295 127.035 116.675 ;
        RECT 126.365 115.955 127.030 116.125 ;
        RECT 123.975 115.385 124.725 115.905 ;
        RECT 120.925 114.295 122.955 114.465 ;
        RECT 123.125 114.125 123.295 115.265 ;
        RECT 123.465 114.295 123.800 115.265 ;
        RECT 124.895 115.215 125.645 115.735 ;
        RECT 123.975 114.125 125.645 115.215 ;
        RECT 125.815 114.125 126.105 115.290 ;
        RECT 126.280 115.135 126.630 115.785 ;
        RECT 126.800 114.965 127.030 115.955 ;
        RECT 126.365 114.795 127.030 114.965 ;
        RECT 126.365 114.295 126.535 114.795 ;
        RECT 126.705 114.125 127.035 114.625 ;
        RECT 127.205 114.295 127.390 116.415 ;
        RECT 127.645 116.215 127.895 116.675 ;
        RECT 128.065 116.225 128.400 116.395 ;
        RECT 128.595 116.225 129.270 116.395 ;
        RECT 128.065 116.085 128.235 116.225 ;
        RECT 127.560 115.095 127.840 116.045 ;
        RECT 128.010 115.955 128.235 116.085 ;
        RECT 128.010 114.850 128.180 115.955 ;
        RECT 128.405 115.805 128.930 116.025 ;
        RECT 128.350 115.040 128.590 115.635 ;
        RECT 128.760 115.105 128.930 115.805 ;
        RECT 129.100 115.445 129.270 116.225 ;
        RECT 129.590 116.175 129.960 116.675 ;
        RECT 130.140 116.225 130.545 116.395 ;
        RECT 130.715 116.225 131.500 116.395 ;
        RECT 130.140 115.995 130.310 116.225 ;
        RECT 129.480 115.695 130.310 115.995 ;
        RECT 130.695 115.725 131.160 116.055 ;
        RECT 129.480 115.665 129.680 115.695 ;
        RECT 129.800 115.445 129.970 115.515 ;
        RECT 129.100 115.275 129.970 115.445 ;
        RECT 129.460 115.185 129.970 115.275 ;
        RECT 128.010 114.720 128.315 114.850 ;
        RECT 128.760 114.740 129.290 115.105 ;
        RECT 127.630 114.125 127.895 114.585 ;
        RECT 128.065 114.295 128.315 114.720 ;
        RECT 129.460 114.570 129.630 115.185 ;
        RECT 128.525 114.400 129.630 114.570 ;
        RECT 129.800 114.125 129.970 114.925 ;
        RECT 130.140 114.625 130.310 115.695 ;
        RECT 130.480 114.795 130.670 115.515 ;
        RECT 130.840 114.765 131.160 115.725 ;
        RECT 131.330 115.765 131.500 116.225 ;
        RECT 131.775 116.145 131.985 116.675 ;
        RECT 132.245 115.935 132.575 116.460 ;
        RECT 132.745 116.065 132.915 116.675 ;
        RECT 133.085 116.020 133.415 116.455 ;
        RECT 133.750 116.045 134.035 116.505 ;
        RECT 134.205 116.215 134.475 116.675 ;
        RECT 133.085 115.935 133.465 116.020 ;
        RECT 132.375 115.765 132.575 115.935 ;
        RECT 133.240 115.895 133.465 115.935 ;
        RECT 131.330 115.435 132.205 115.765 ;
        RECT 132.375 115.435 133.125 115.765 ;
        RECT 130.140 114.295 130.390 114.625 ;
        RECT 131.330 114.595 131.500 115.435 ;
        RECT 132.375 115.230 132.565 115.435 ;
        RECT 133.295 115.315 133.465 115.895 ;
        RECT 133.750 115.875 134.705 116.045 ;
        RECT 133.250 115.265 133.465 115.315 ;
        RECT 131.670 114.855 132.565 115.230 ;
        RECT 133.075 115.185 133.465 115.265 ;
        RECT 130.615 114.425 131.500 114.595 ;
        RECT 131.680 114.125 131.995 114.625 ;
        RECT 132.225 114.295 132.565 114.855 ;
        RECT 132.735 114.125 132.905 115.135 ;
        RECT 133.075 114.340 133.405 115.185 ;
        RECT 133.635 115.145 134.325 115.705 ;
        RECT 134.495 114.975 134.705 115.875 ;
        RECT 133.750 114.755 134.705 114.975 ;
        RECT 134.875 115.705 135.275 116.505 ;
        RECT 135.465 116.045 135.745 116.505 ;
        RECT 136.265 116.215 136.590 116.675 ;
        RECT 135.465 115.875 136.590 116.045 ;
        RECT 136.760 115.935 137.145 116.505 ;
        RECT 137.595 116.045 137.975 116.495 ;
        RECT 136.140 115.765 136.590 115.875 ;
        RECT 134.875 115.145 135.970 115.705 ;
        RECT 136.140 115.435 136.695 115.765 ;
        RECT 133.750 114.295 134.035 114.755 ;
        RECT 134.205 114.125 134.475 114.585 ;
        RECT 134.875 114.295 135.275 115.145 ;
        RECT 136.140 114.975 136.590 115.435 ;
        RECT 136.865 115.265 137.145 115.935 ;
        RECT 135.465 114.755 136.590 114.975 ;
        RECT 135.465 114.295 135.745 114.755 ;
        RECT 136.265 114.125 136.590 114.585 ;
        RECT 136.760 114.295 137.145 115.265 ;
        RECT 137.335 115.095 137.565 115.785 ;
        RECT 137.745 115.595 137.975 116.045 ;
        RECT 138.155 115.895 138.385 116.675 ;
        RECT 138.565 115.965 138.995 116.495 ;
        RECT 138.565 115.715 138.810 115.965 ;
        RECT 139.175 115.765 139.385 116.385 ;
        RECT 139.555 115.945 139.885 116.675 ;
        RECT 140.075 115.935 140.460 116.505 ;
        RECT 140.630 116.215 140.955 116.675 ;
        RECT 141.475 116.045 141.755 116.505 ;
        RECT 137.745 114.915 138.085 115.595 ;
        RECT 137.325 114.715 138.085 114.915 ;
        RECT 138.275 115.415 138.810 115.715 ;
        RECT 138.990 115.415 139.385 115.765 ;
        RECT 139.580 115.415 139.870 115.765 ;
        RECT 137.325 114.325 137.585 114.715 ;
        RECT 137.755 114.125 138.085 114.535 ;
        RECT 138.275 114.305 138.605 115.415 ;
        RECT 140.075 115.265 140.355 115.935 ;
        RECT 140.630 115.875 141.755 116.045 ;
        RECT 140.630 115.765 141.080 115.875 ;
        RECT 140.525 115.435 141.080 115.765 ;
        RECT 141.945 115.705 142.345 116.505 ;
        RECT 142.745 116.215 143.015 116.675 ;
        RECT 143.185 116.045 143.470 116.505 ;
        RECT 138.775 115.035 139.815 115.235 ;
        RECT 138.775 114.305 138.965 115.035 ;
        RECT 139.135 114.125 139.465 114.855 ;
        RECT 139.645 114.305 139.815 115.035 ;
        RECT 140.075 114.295 140.460 115.265 ;
        RECT 140.630 114.975 141.080 115.435 ;
        RECT 141.250 115.145 142.345 115.705 ;
        RECT 140.630 114.755 141.755 114.975 ;
        RECT 140.630 114.125 140.955 114.585 ;
        RECT 141.475 114.295 141.755 114.755 ;
        RECT 141.945 114.295 142.345 115.145 ;
        RECT 142.515 115.875 143.470 116.045 ;
        RECT 144.305 116.125 144.475 116.415 ;
        RECT 144.645 116.295 144.975 116.675 ;
        RECT 144.305 115.955 144.970 116.125 ;
        RECT 142.515 114.975 142.725 115.875 ;
        RECT 142.895 115.145 143.585 115.705 ;
        RECT 144.220 115.135 144.570 115.785 ;
        RECT 142.515 114.755 143.470 114.975 ;
        RECT 144.740 114.965 144.970 115.955 ;
        RECT 142.745 114.125 143.015 114.585 ;
        RECT 143.185 114.295 143.470 114.755 ;
        RECT 144.305 114.795 144.970 114.965 ;
        RECT 144.305 114.295 144.475 114.795 ;
        RECT 144.645 114.125 144.975 114.625 ;
        RECT 145.145 114.295 145.330 116.415 ;
        RECT 145.585 116.215 145.835 116.675 ;
        RECT 146.005 116.225 146.340 116.395 ;
        RECT 146.535 116.225 147.210 116.395 ;
        RECT 146.005 116.085 146.175 116.225 ;
        RECT 145.500 115.095 145.780 116.045 ;
        RECT 145.950 115.955 146.175 116.085 ;
        RECT 145.950 114.850 146.120 115.955 ;
        RECT 146.345 115.805 146.870 116.025 ;
        RECT 146.290 115.040 146.530 115.635 ;
        RECT 146.700 115.105 146.870 115.805 ;
        RECT 147.040 115.445 147.210 116.225 ;
        RECT 147.530 116.175 147.900 116.675 ;
        RECT 148.080 116.225 148.485 116.395 ;
        RECT 148.655 116.225 149.440 116.395 ;
        RECT 148.080 115.995 148.250 116.225 ;
        RECT 147.420 115.695 148.250 115.995 ;
        RECT 148.635 115.725 149.100 116.055 ;
        RECT 147.420 115.665 147.620 115.695 ;
        RECT 147.740 115.445 147.910 115.515 ;
        RECT 147.040 115.275 147.910 115.445 ;
        RECT 147.400 115.185 147.910 115.275 ;
        RECT 145.950 114.720 146.255 114.850 ;
        RECT 146.700 114.740 147.230 115.105 ;
        RECT 145.570 114.125 145.835 114.585 ;
        RECT 146.005 114.295 146.255 114.720 ;
        RECT 147.400 114.570 147.570 115.185 ;
        RECT 146.465 114.400 147.570 114.570 ;
        RECT 147.740 114.125 147.910 114.925 ;
        RECT 148.080 114.625 148.250 115.695 ;
        RECT 148.420 114.795 148.610 115.515 ;
        RECT 148.780 114.765 149.100 115.725 ;
        RECT 149.270 115.765 149.440 116.225 ;
        RECT 149.715 116.145 149.925 116.675 ;
        RECT 150.185 115.935 150.515 116.460 ;
        RECT 150.685 116.065 150.855 116.675 ;
        RECT 151.025 116.020 151.355 116.455 ;
        RECT 151.025 115.935 151.405 116.020 ;
        RECT 151.575 115.950 151.865 116.675 ;
        RECT 152.125 116.125 152.295 116.505 ;
        RECT 152.475 116.295 152.805 116.675 ;
        RECT 152.125 115.955 152.790 116.125 ;
        RECT 152.985 116.000 153.245 116.505 ;
        RECT 150.315 115.765 150.515 115.935 ;
        RECT 151.180 115.895 151.405 115.935 ;
        RECT 149.270 115.435 150.145 115.765 ;
        RECT 150.315 115.435 151.065 115.765 ;
        RECT 148.080 114.295 148.330 114.625 ;
        RECT 149.270 114.595 149.440 115.435 ;
        RECT 150.315 115.230 150.505 115.435 ;
        RECT 151.235 115.315 151.405 115.895 ;
        RECT 152.055 115.405 152.385 115.775 ;
        RECT 152.620 115.700 152.790 115.955 ;
        RECT 151.190 115.265 151.405 115.315 ;
        RECT 152.620 115.370 152.905 115.700 ;
        RECT 149.610 114.855 150.505 115.230 ;
        RECT 151.015 115.185 151.405 115.265 ;
        RECT 148.555 114.425 149.440 114.595 ;
        RECT 149.620 114.125 149.935 114.625 ;
        RECT 150.165 114.295 150.505 114.855 ;
        RECT 150.675 114.125 150.845 115.135 ;
        RECT 151.015 114.340 151.345 115.185 ;
        RECT 151.575 114.125 151.865 115.290 ;
        RECT 152.620 115.225 152.790 115.370 ;
        RECT 152.125 115.055 152.790 115.225 ;
        RECT 153.075 115.200 153.245 116.000 ;
        RECT 153.415 115.905 155.085 116.675 ;
        RECT 155.715 115.925 156.925 116.675 ;
        RECT 153.415 115.385 154.165 115.905 ;
        RECT 154.335 115.215 155.085 115.735 ;
        RECT 152.125 114.295 152.295 115.055 ;
        RECT 152.475 114.125 152.805 114.885 ;
        RECT 152.975 114.295 153.245 115.200 ;
        RECT 153.415 114.125 155.085 115.215 ;
        RECT 155.715 115.215 156.235 115.755 ;
        RECT 156.405 115.385 156.925 115.925 ;
        RECT 155.715 114.125 156.925 115.215 ;
        RECT 22.690 113.955 157.010 114.125 ;
        RECT 22.775 112.865 23.985 113.955 ;
        RECT 22.775 112.155 23.295 112.695 ;
        RECT 23.465 112.325 23.985 112.865 ;
        RECT 25.110 113.165 25.645 113.785 ;
        RECT 22.775 111.405 23.985 112.155 ;
        RECT 25.110 112.145 25.425 113.165 ;
        RECT 25.815 113.155 26.145 113.955 ;
        RECT 26.630 112.985 27.020 113.160 ;
        RECT 25.595 112.815 27.020 112.985 ;
        RECT 27.375 112.815 27.715 113.785 ;
        RECT 27.885 112.815 28.055 113.955 ;
        RECT 28.325 113.155 28.575 113.955 ;
        RECT 29.220 112.985 29.550 113.785 ;
        RECT 29.850 113.155 30.180 113.955 ;
        RECT 30.350 112.985 30.680 113.785 ;
        RECT 28.245 112.815 30.680 112.985 ;
        RECT 31.055 112.815 31.440 113.785 ;
        RECT 31.610 113.495 31.935 113.955 ;
        RECT 32.455 113.325 32.735 113.785 ;
        RECT 31.610 113.105 32.735 113.325 ;
        RECT 25.595 112.315 25.765 112.815 ;
        RECT 25.110 111.575 25.725 112.145 ;
        RECT 26.015 112.085 26.280 112.645 ;
        RECT 26.450 111.915 26.620 112.815 ;
        RECT 26.790 112.085 27.145 112.645 ;
        RECT 27.375 112.205 27.550 112.815 ;
        RECT 28.245 112.565 28.415 112.815 ;
        RECT 27.720 112.395 28.415 112.565 ;
        RECT 28.590 112.395 29.010 112.595 ;
        RECT 29.180 112.395 29.510 112.595 ;
        RECT 29.680 112.395 30.010 112.595 ;
        RECT 25.895 111.405 26.110 111.915 ;
        RECT 26.340 111.585 26.620 111.915 ;
        RECT 26.800 111.405 27.040 111.915 ;
        RECT 27.375 111.575 27.715 112.205 ;
        RECT 27.885 111.405 28.135 112.205 ;
        RECT 28.325 112.055 29.550 112.225 ;
        RECT 28.325 111.575 28.655 112.055 ;
        RECT 28.825 111.405 29.050 111.865 ;
        RECT 29.220 111.575 29.550 112.055 ;
        RECT 30.180 112.185 30.350 112.815 ;
        RECT 30.535 112.395 30.885 112.645 ;
        RECT 30.180 111.575 30.680 112.185 ;
        RECT 31.055 112.145 31.335 112.815 ;
        RECT 31.610 112.645 32.060 113.105 ;
        RECT 32.925 112.935 33.325 113.785 ;
        RECT 33.725 113.495 33.995 113.955 ;
        RECT 34.165 113.325 34.450 113.785 ;
        RECT 31.505 112.315 32.060 112.645 ;
        RECT 32.230 112.375 33.325 112.935 ;
        RECT 31.610 112.205 32.060 112.315 ;
        RECT 31.055 111.575 31.440 112.145 ;
        RECT 31.610 112.035 32.735 112.205 ;
        RECT 31.610 111.405 31.935 111.865 ;
        RECT 32.455 111.575 32.735 112.035 ;
        RECT 32.925 111.575 33.325 112.375 ;
        RECT 33.495 113.105 34.450 113.325 ;
        RECT 33.495 112.205 33.705 113.105 ;
        RECT 33.875 112.375 34.565 112.935 ;
        RECT 35.655 112.790 35.945 113.955 ;
        RECT 36.115 112.865 37.325 113.955 ;
        RECT 33.495 112.035 34.450 112.205 ;
        RECT 36.115 112.155 36.635 112.695 ;
        RECT 36.805 112.325 37.325 112.865 ;
        RECT 37.495 112.815 37.880 113.785 ;
        RECT 38.050 113.495 38.375 113.955 ;
        RECT 38.895 113.325 39.175 113.785 ;
        RECT 38.050 113.105 39.175 113.325 ;
        RECT 33.725 111.405 33.995 111.865 ;
        RECT 34.165 111.575 34.450 112.035 ;
        RECT 35.655 111.405 35.945 112.130 ;
        RECT 36.115 111.405 37.325 112.155 ;
        RECT 37.495 112.145 37.775 112.815 ;
        RECT 38.050 112.645 38.500 113.105 ;
        RECT 39.365 112.935 39.765 113.785 ;
        RECT 40.165 113.495 40.435 113.955 ;
        RECT 40.605 113.325 40.890 113.785 ;
        RECT 37.945 112.315 38.500 112.645 ;
        RECT 38.670 112.375 39.765 112.935 ;
        RECT 38.050 112.205 38.500 112.315 ;
        RECT 37.495 111.575 37.880 112.145 ;
        RECT 38.050 112.035 39.175 112.205 ;
        RECT 38.050 111.405 38.375 111.865 ;
        RECT 38.895 111.575 39.175 112.035 ;
        RECT 39.365 111.575 39.765 112.375 ;
        RECT 39.935 113.105 40.890 113.325 ;
        RECT 39.935 112.205 40.145 113.105 ;
        RECT 40.315 112.375 41.005 112.935 ;
        RECT 41.180 112.805 41.440 113.955 ;
        RECT 41.615 112.880 41.870 113.785 ;
        RECT 42.040 113.195 42.370 113.955 ;
        RECT 42.585 113.025 42.755 113.785 ;
        RECT 43.130 113.325 43.415 113.785 ;
        RECT 43.585 113.495 43.855 113.955 ;
        RECT 43.130 113.105 44.085 113.325 ;
        RECT 39.935 112.035 40.890 112.205 ;
        RECT 40.165 111.405 40.435 111.865 ;
        RECT 40.605 111.575 40.890 112.035 ;
        RECT 41.180 111.405 41.440 112.245 ;
        RECT 41.615 112.150 41.785 112.880 ;
        RECT 42.040 112.855 42.755 113.025 ;
        RECT 42.040 112.645 42.210 112.855 ;
        RECT 41.955 112.315 42.210 112.645 ;
        RECT 41.615 111.575 41.870 112.150 ;
        RECT 42.040 112.125 42.210 112.315 ;
        RECT 42.490 112.305 42.845 112.675 ;
        RECT 43.015 112.375 43.705 112.935 ;
        RECT 43.875 112.205 44.085 113.105 ;
        RECT 42.040 111.955 42.755 112.125 ;
        RECT 42.040 111.405 42.370 111.785 ;
        RECT 42.585 111.575 42.755 111.955 ;
        RECT 43.130 112.035 44.085 112.205 ;
        RECT 44.255 112.935 44.655 113.785 ;
        RECT 44.845 113.325 45.125 113.785 ;
        RECT 45.645 113.495 45.970 113.955 ;
        RECT 44.845 113.105 45.970 113.325 ;
        RECT 44.255 112.375 45.350 112.935 ;
        RECT 45.520 112.645 45.970 113.105 ;
        RECT 46.140 112.815 46.525 113.785 ;
        RECT 46.785 113.285 46.955 113.785 ;
        RECT 47.125 113.455 47.455 113.955 ;
        RECT 46.785 113.115 47.450 113.285 ;
        RECT 43.130 111.575 43.415 112.035 ;
        RECT 43.585 111.405 43.855 111.865 ;
        RECT 44.255 111.575 44.655 112.375 ;
        RECT 45.520 112.315 46.075 112.645 ;
        RECT 45.520 112.205 45.970 112.315 ;
        RECT 44.845 112.035 45.970 112.205 ;
        RECT 46.245 112.145 46.525 112.815 ;
        RECT 46.700 112.295 47.050 112.945 ;
        RECT 44.845 111.575 45.125 112.035 ;
        RECT 45.645 111.405 45.970 111.865 ;
        RECT 46.140 111.575 46.525 112.145 ;
        RECT 47.220 112.125 47.450 113.115 ;
        RECT 46.785 111.955 47.450 112.125 ;
        RECT 46.785 111.665 46.955 111.955 ;
        RECT 47.125 111.405 47.455 111.785 ;
        RECT 47.625 111.665 47.810 113.785 ;
        RECT 48.050 113.495 48.315 113.955 ;
        RECT 48.485 113.360 48.735 113.785 ;
        RECT 48.945 113.510 50.050 113.680 ;
        RECT 48.430 113.230 48.735 113.360 ;
        RECT 47.980 112.035 48.260 112.985 ;
        RECT 48.430 112.125 48.600 113.230 ;
        RECT 48.770 112.445 49.010 113.040 ;
        RECT 49.180 112.975 49.710 113.340 ;
        RECT 49.180 112.275 49.350 112.975 ;
        RECT 49.880 112.895 50.050 113.510 ;
        RECT 50.220 113.155 50.390 113.955 ;
        RECT 50.560 113.455 50.810 113.785 ;
        RECT 51.035 113.485 51.920 113.655 ;
        RECT 49.880 112.805 50.390 112.895 ;
        RECT 48.430 111.995 48.655 112.125 ;
        RECT 48.825 112.055 49.350 112.275 ;
        RECT 49.520 112.635 50.390 112.805 ;
        RECT 48.065 111.405 48.315 111.865 ;
        RECT 48.485 111.855 48.655 111.995 ;
        RECT 49.520 111.855 49.690 112.635 ;
        RECT 50.220 112.565 50.390 112.635 ;
        RECT 49.900 112.385 50.100 112.415 ;
        RECT 50.560 112.385 50.730 113.455 ;
        RECT 50.900 112.565 51.090 113.285 ;
        RECT 49.900 112.085 50.730 112.385 ;
        RECT 51.260 112.355 51.580 113.315 ;
        RECT 48.485 111.685 48.820 111.855 ;
        RECT 49.015 111.685 49.690 111.855 ;
        RECT 50.010 111.405 50.380 111.905 ;
        RECT 50.560 111.855 50.730 112.085 ;
        RECT 51.115 112.025 51.580 112.355 ;
        RECT 51.750 112.645 51.920 113.485 ;
        RECT 52.100 113.455 52.415 113.955 ;
        RECT 52.645 113.225 52.985 113.785 ;
        RECT 52.090 112.850 52.985 113.225 ;
        RECT 53.155 112.945 53.325 113.955 ;
        RECT 52.795 112.645 52.985 112.850 ;
        RECT 53.495 112.895 53.825 113.740 ;
        RECT 54.145 113.285 54.315 113.785 ;
        RECT 54.485 113.455 54.815 113.955 ;
        RECT 54.145 113.115 54.810 113.285 ;
        RECT 53.495 112.815 53.885 112.895 ;
        RECT 53.670 112.765 53.885 112.815 ;
        RECT 51.750 112.315 52.625 112.645 ;
        RECT 52.795 112.315 53.545 112.645 ;
        RECT 51.750 111.855 51.920 112.315 ;
        RECT 52.795 112.145 52.995 112.315 ;
        RECT 53.715 112.185 53.885 112.765 ;
        RECT 54.060 112.295 54.410 112.945 ;
        RECT 53.660 112.145 53.885 112.185 ;
        RECT 50.560 111.685 50.965 111.855 ;
        RECT 51.135 111.685 51.920 111.855 ;
        RECT 52.195 111.405 52.405 111.935 ;
        RECT 52.665 111.620 52.995 112.145 ;
        RECT 53.505 112.060 53.885 112.145 ;
        RECT 54.580 112.125 54.810 113.115 ;
        RECT 53.165 111.405 53.335 112.015 ;
        RECT 53.505 111.625 53.835 112.060 ;
        RECT 54.145 111.955 54.810 112.125 ;
        RECT 54.145 111.665 54.315 111.955 ;
        RECT 54.485 111.405 54.815 111.785 ;
        RECT 54.985 111.665 55.170 113.785 ;
        RECT 55.410 113.495 55.675 113.955 ;
        RECT 55.845 113.360 56.095 113.785 ;
        RECT 56.305 113.510 57.410 113.680 ;
        RECT 55.790 113.230 56.095 113.360 ;
        RECT 55.340 112.035 55.620 112.985 ;
        RECT 55.790 112.125 55.960 113.230 ;
        RECT 56.130 112.445 56.370 113.040 ;
        RECT 56.540 112.975 57.070 113.340 ;
        RECT 56.540 112.275 56.710 112.975 ;
        RECT 57.240 112.895 57.410 113.510 ;
        RECT 57.580 113.155 57.750 113.955 ;
        RECT 57.920 113.455 58.170 113.785 ;
        RECT 58.395 113.485 59.280 113.655 ;
        RECT 57.240 112.805 57.750 112.895 ;
        RECT 55.790 111.995 56.015 112.125 ;
        RECT 56.185 112.055 56.710 112.275 ;
        RECT 56.880 112.635 57.750 112.805 ;
        RECT 55.425 111.405 55.675 111.865 ;
        RECT 55.845 111.855 56.015 111.995 ;
        RECT 56.880 111.855 57.050 112.635 ;
        RECT 57.580 112.565 57.750 112.635 ;
        RECT 57.260 112.385 57.460 112.415 ;
        RECT 57.920 112.385 58.090 113.455 ;
        RECT 58.260 112.565 58.450 113.285 ;
        RECT 57.260 112.085 58.090 112.385 ;
        RECT 58.620 112.355 58.940 113.315 ;
        RECT 55.845 111.685 56.180 111.855 ;
        RECT 56.375 111.685 57.050 111.855 ;
        RECT 57.370 111.405 57.740 111.905 ;
        RECT 57.920 111.855 58.090 112.085 ;
        RECT 58.475 112.025 58.940 112.355 ;
        RECT 59.110 112.645 59.280 113.485 ;
        RECT 59.460 113.455 59.775 113.955 ;
        RECT 60.005 113.225 60.345 113.785 ;
        RECT 59.450 112.850 60.345 113.225 ;
        RECT 60.515 112.945 60.685 113.955 ;
        RECT 60.155 112.645 60.345 112.850 ;
        RECT 60.855 112.895 61.185 113.740 ;
        RECT 60.855 112.815 61.245 112.895 ;
        RECT 61.030 112.765 61.245 112.815 ;
        RECT 61.415 112.790 61.705 113.955 ;
        RECT 61.875 112.815 62.215 113.785 ;
        RECT 62.385 112.815 62.555 113.955 ;
        RECT 62.825 113.155 63.075 113.955 ;
        RECT 63.720 112.985 64.050 113.785 ;
        RECT 64.350 113.155 64.680 113.955 ;
        RECT 64.850 112.985 65.180 113.785 ;
        RECT 62.745 112.815 65.180 112.985 ;
        RECT 65.555 112.815 65.940 113.785 ;
        RECT 66.110 113.495 66.435 113.955 ;
        RECT 66.955 113.325 67.235 113.785 ;
        RECT 66.110 113.105 67.235 113.325 ;
        RECT 59.110 112.315 59.985 112.645 ;
        RECT 60.155 112.315 60.905 112.645 ;
        RECT 59.110 111.855 59.280 112.315 ;
        RECT 60.155 112.145 60.355 112.315 ;
        RECT 61.075 112.185 61.245 112.765 ;
        RECT 61.020 112.145 61.245 112.185 ;
        RECT 57.920 111.685 58.325 111.855 ;
        RECT 58.495 111.685 59.280 111.855 ;
        RECT 59.555 111.405 59.765 111.935 ;
        RECT 60.025 111.620 60.355 112.145 ;
        RECT 60.865 112.060 61.245 112.145 ;
        RECT 61.875 112.205 62.050 112.815 ;
        RECT 62.745 112.565 62.915 112.815 ;
        RECT 62.220 112.395 62.915 112.565 ;
        RECT 63.090 112.395 63.510 112.595 ;
        RECT 63.680 112.395 64.010 112.595 ;
        RECT 64.180 112.395 64.510 112.595 ;
        RECT 60.525 111.405 60.695 112.015 ;
        RECT 60.865 111.625 61.195 112.060 ;
        RECT 61.415 111.405 61.705 112.130 ;
        RECT 61.875 111.575 62.215 112.205 ;
        RECT 62.385 111.405 62.635 112.205 ;
        RECT 62.825 112.055 64.050 112.225 ;
        RECT 62.825 111.575 63.155 112.055 ;
        RECT 63.325 111.405 63.550 111.865 ;
        RECT 63.720 111.575 64.050 112.055 ;
        RECT 64.680 112.185 64.850 112.815 ;
        RECT 65.035 112.395 65.385 112.645 ;
        RECT 64.680 111.575 65.180 112.185 ;
        RECT 65.555 112.145 65.835 112.815 ;
        RECT 66.110 112.645 66.560 113.105 ;
        RECT 67.425 112.935 67.825 113.785 ;
        RECT 68.225 113.495 68.495 113.955 ;
        RECT 68.665 113.325 68.950 113.785 ;
        RECT 66.005 112.315 66.560 112.645 ;
        RECT 66.730 112.375 67.825 112.935 ;
        RECT 66.110 112.205 66.560 112.315 ;
        RECT 65.555 111.575 65.940 112.145 ;
        RECT 66.110 112.035 67.235 112.205 ;
        RECT 66.110 111.405 66.435 111.865 ;
        RECT 66.955 111.575 67.235 112.035 ;
        RECT 67.425 111.575 67.825 112.375 ;
        RECT 67.995 113.105 68.950 113.325 ;
        RECT 69.785 113.285 69.955 113.785 ;
        RECT 70.125 113.455 70.455 113.955 ;
        RECT 69.785 113.115 70.450 113.285 ;
        RECT 67.995 112.205 68.205 113.105 ;
        RECT 68.375 112.375 69.065 112.935 ;
        RECT 69.700 112.295 70.050 112.945 ;
        RECT 67.995 112.035 68.950 112.205 ;
        RECT 70.220 112.125 70.450 113.115 ;
        RECT 68.225 111.405 68.495 111.865 ;
        RECT 68.665 111.575 68.950 112.035 ;
        RECT 69.785 111.955 70.450 112.125 ;
        RECT 69.785 111.665 69.955 111.955 ;
        RECT 70.125 111.405 70.455 111.785 ;
        RECT 70.625 111.665 70.810 113.785 ;
        RECT 71.050 113.495 71.315 113.955 ;
        RECT 71.485 113.360 71.735 113.785 ;
        RECT 71.945 113.510 73.050 113.680 ;
        RECT 71.430 113.230 71.735 113.360 ;
        RECT 70.980 112.035 71.260 112.985 ;
        RECT 71.430 112.125 71.600 113.230 ;
        RECT 71.770 112.445 72.010 113.040 ;
        RECT 72.180 112.975 72.710 113.340 ;
        RECT 72.180 112.275 72.350 112.975 ;
        RECT 72.880 112.895 73.050 113.510 ;
        RECT 73.220 113.155 73.390 113.955 ;
        RECT 73.560 113.455 73.810 113.785 ;
        RECT 74.035 113.485 74.920 113.655 ;
        RECT 72.880 112.805 73.390 112.895 ;
        RECT 71.430 111.995 71.655 112.125 ;
        RECT 71.825 112.055 72.350 112.275 ;
        RECT 72.520 112.635 73.390 112.805 ;
        RECT 71.065 111.405 71.315 111.865 ;
        RECT 71.485 111.855 71.655 111.995 ;
        RECT 72.520 111.855 72.690 112.635 ;
        RECT 73.220 112.565 73.390 112.635 ;
        RECT 72.900 112.385 73.100 112.415 ;
        RECT 73.560 112.385 73.730 113.455 ;
        RECT 73.900 112.565 74.090 113.285 ;
        RECT 72.900 112.085 73.730 112.385 ;
        RECT 74.260 112.355 74.580 113.315 ;
        RECT 71.485 111.685 71.820 111.855 ;
        RECT 72.015 111.685 72.690 111.855 ;
        RECT 73.010 111.405 73.380 111.905 ;
        RECT 73.560 111.855 73.730 112.085 ;
        RECT 74.115 112.025 74.580 112.355 ;
        RECT 74.750 112.645 74.920 113.485 ;
        RECT 75.100 113.455 75.415 113.955 ;
        RECT 75.645 113.225 75.985 113.785 ;
        RECT 75.090 112.850 75.985 113.225 ;
        RECT 76.155 112.945 76.325 113.955 ;
        RECT 75.795 112.645 75.985 112.850 ;
        RECT 76.495 112.895 76.825 113.740 ;
        RECT 77.145 113.025 77.315 113.785 ;
        RECT 77.495 113.195 77.825 113.955 ;
        RECT 76.495 112.815 76.885 112.895 ;
        RECT 77.145 112.855 77.810 113.025 ;
        RECT 77.995 112.880 78.265 113.785 ;
        RECT 76.670 112.765 76.885 112.815 ;
        RECT 74.750 112.315 75.625 112.645 ;
        RECT 75.795 112.315 76.545 112.645 ;
        RECT 74.750 111.855 74.920 112.315 ;
        RECT 75.795 112.145 75.995 112.315 ;
        RECT 76.715 112.185 76.885 112.765 ;
        RECT 77.640 112.710 77.810 112.855 ;
        RECT 77.075 112.305 77.405 112.675 ;
        RECT 77.640 112.380 77.925 112.710 ;
        RECT 76.660 112.145 76.885 112.185 ;
        RECT 73.560 111.685 73.965 111.855 ;
        RECT 74.135 111.685 74.920 111.855 ;
        RECT 75.195 111.405 75.405 111.935 ;
        RECT 75.665 111.620 75.995 112.145 ;
        RECT 76.505 112.060 76.885 112.145 ;
        RECT 77.640 112.125 77.810 112.380 ;
        RECT 76.165 111.405 76.335 112.015 ;
        RECT 76.505 111.625 76.835 112.060 ;
        RECT 77.145 111.955 77.810 112.125 ;
        RECT 78.095 112.080 78.265 112.880 ;
        RECT 78.435 113.195 78.950 113.605 ;
        RECT 79.185 113.195 79.355 113.955 ;
        RECT 79.525 113.615 81.555 113.785 ;
        RECT 78.435 112.385 78.775 113.195 ;
        RECT 79.525 112.950 79.695 113.615 ;
        RECT 80.090 113.275 81.215 113.445 ;
        RECT 78.945 112.760 79.695 112.950 ;
        RECT 79.865 112.935 80.875 113.105 ;
        RECT 78.435 112.215 79.665 112.385 ;
        RECT 77.145 111.575 77.315 111.955 ;
        RECT 77.495 111.405 77.825 111.785 ;
        RECT 78.005 111.575 78.265 112.080 ;
        RECT 78.710 111.610 78.955 112.215 ;
        RECT 79.175 111.405 79.685 111.940 ;
        RECT 79.865 111.575 80.055 112.935 ;
        RECT 80.225 112.595 80.500 112.735 ;
        RECT 80.225 112.425 80.505 112.595 ;
        RECT 80.225 111.575 80.500 112.425 ;
        RECT 80.705 112.135 80.875 112.935 ;
        RECT 81.045 112.145 81.215 113.275 ;
        RECT 81.385 112.645 81.555 113.615 ;
        RECT 81.725 112.815 81.895 113.955 ;
        RECT 82.065 112.815 82.400 113.785 ;
        RECT 81.385 112.315 81.580 112.645 ;
        RECT 81.805 112.315 82.060 112.645 ;
        RECT 81.805 112.145 81.975 112.315 ;
        RECT 82.230 112.145 82.400 112.815 ;
        RECT 81.045 111.975 81.975 112.145 ;
        RECT 81.045 111.940 81.220 111.975 ;
        RECT 80.690 111.575 81.220 111.940 ;
        RECT 81.645 111.405 81.975 111.805 ;
        RECT 82.145 111.575 82.400 112.145 ;
        RECT 82.580 112.815 82.915 113.785 ;
        RECT 83.085 112.815 83.255 113.955 ;
        RECT 83.425 113.615 85.455 113.785 ;
        RECT 82.580 112.145 82.750 112.815 ;
        RECT 83.425 112.645 83.595 113.615 ;
        RECT 82.920 112.315 83.175 112.645 ;
        RECT 83.400 112.315 83.595 112.645 ;
        RECT 83.765 113.275 84.890 113.445 ;
        RECT 83.005 112.145 83.175 112.315 ;
        RECT 83.765 112.145 83.935 113.275 ;
        RECT 82.580 111.575 82.835 112.145 ;
        RECT 83.005 111.975 83.935 112.145 ;
        RECT 84.105 112.935 85.115 113.105 ;
        RECT 84.105 112.135 84.275 112.935 ;
        RECT 84.480 112.595 84.755 112.735 ;
        RECT 84.475 112.425 84.755 112.595 ;
        RECT 83.760 111.940 83.935 111.975 ;
        RECT 83.005 111.405 83.335 111.805 ;
        RECT 83.760 111.575 84.290 111.940 ;
        RECT 84.480 111.575 84.755 112.425 ;
        RECT 84.925 111.575 85.115 112.935 ;
        RECT 85.285 112.950 85.455 113.615 ;
        RECT 85.625 113.195 85.795 113.955 ;
        RECT 86.030 113.195 86.545 113.605 ;
        RECT 85.285 112.760 86.035 112.950 ;
        RECT 86.205 112.385 86.545 113.195 ;
        RECT 87.175 112.790 87.465 113.955 ;
        RECT 88.645 113.285 88.815 113.785 ;
        RECT 88.985 113.455 89.315 113.955 ;
        RECT 88.645 113.115 89.310 113.285 ;
        RECT 85.315 112.215 86.545 112.385 ;
        RECT 88.560 112.295 88.910 112.945 ;
        RECT 85.295 111.405 85.805 111.940 ;
        RECT 86.025 111.610 86.270 112.215 ;
        RECT 87.175 111.405 87.465 112.130 ;
        RECT 89.080 112.125 89.310 113.115 ;
        RECT 88.645 111.955 89.310 112.125 ;
        RECT 88.645 111.665 88.815 111.955 ;
        RECT 88.985 111.405 89.315 111.785 ;
        RECT 89.485 111.665 89.670 113.785 ;
        RECT 89.910 113.495 90.175 113.955 ;
        RECT 90.345 113.360 90.595 113.785 ;
        RECT 90.805 113.510 91.910 113.680 ;
        RECT 90.290 113.230 90.595 113.360 ;
        RECT 89.840 112.035 90.120 112.985 ;
        RECT 90.290 112.125 90.460 113.230 ;
        RECT 90.630 112.445 90.870 113.040 ;
        RECT 91.040 112.975 91.570 113.340 ;
        RECT 91.040 112.275 91.210 112.975 ;
        RECT 91.740 112.895 91.910 113.510 ;
        RECT 92.080 113.155 92.250 113.955 ;
        RECT 92.420 113.455 92.670 113.785 ;
        RECT 92.895 113.485 93.780 113.655 ;
        RECT 91.740 112.805 92.250 112.895 ;
        RECT 90.290 111.995 90.515 112.125 ;
        RECT 90.685 112.055 91.210 112.275 ;
        RECT 91.380 112.635 92.250 112.805 ;
        RECT 89.925 111.405 90.175 111.865 ;
        RECT 90.345 111.855 90.515 111.995 ;
        RECT 91.380 111.855 91.550 112.635 ;
        RECT 92.080 112.565 92.250 112.635 ;
        RECT 91.760 112.385 91.960 112.415 ;
        RECT 92.420 112.385 92.590 113.455 ;
        RECT 92.760 112.565 92.950 113.285 ;
        RECT 91.760 112.085 92.590 112.385 ;
        RECT 93.120 112.355 93.440 113.315 ;
        RECT 90.345 111.685 90.680 111.855 ;
        RECT 90.875 111.685 91.550 111.855 ;
        RECT 91.870 111.405 92.240 111.905 ;
        RECT 92.420 111.855 92.590 112.085 ;
        RECT 92.975 112.025 93.440 112.355 ;
        RECT 93.610 112.645 93.780 113.485 ;
        RECT 93.960 113.455 94.275 113.955 ;
        RECT 94.505 113.225 94.845 113.785 ;
        RECT 93.950 112.850 94.845 113.225 ;
        RECT 95.015 112.945 95.185 113.955 ;
        RECT 94.655 112.645 94.845 112.850 ;
        RECT 95.355 112.895 95.685 113.740 ;
        RECT 95.355 112.815 95.745 112.895 ;
        RECT 95.530 112.765 95.745 112.815 ;
        RECT 93.610 112.315 94.485 112.645 ;
        RECT 94.655 112.315 95.405 112.645 ;
        RECT 93.610 111.855 93.780 112.315 ;
        RECT 94.655 112.145 94.855 112.315 ;
        RECT 95.575 112.185 95.745 112.765 ;
        RECT 95.520 112.145 95.745 112.185 ;
        RECT 92.420 111.685 92.825 111.855 ;
        RECT 92.995 111.685 93.780 111.855 ;
        RECT 94.055 111.405 94.265 111.935 ;
        RECT 94.525 111.620 94.855 112.145 ;
        RECT 95.365 112.060 95.745 112.145 ;
        RECT 95.920 112.815 96.255 113.785 ;
        RECT 96.425 112.815 96.595 113.955 ;
        RECT 96.765 113.615 98.795 113.785 ;
        RECT 95.920 112.145 96.090 112.815 ;
        RECT 96.765 112.645 96.935 113.615 ;
        RECT 96.260 112.315 96.515 112.645 ;
        RECT 96.740 112.315 96.935 112.645 ;
        RECT 97.105 113.275 98.230 113.445 ;
        RECT 96.345 112.145 96.515 112.315 ;
        RECT 97.105 112.145 97.275 113.275 ;
        RECT 95.025 111.405 95.195 112.015 ;
        RECT 95.365 111.625 95.695 112.060 ;
        RECT 95.920 111.575 96.175 112.145 ;
        RECT 96.345 111.975 97.275 112.145 ;
        RECT 97.445 112.935 98.455 113.105 ;
        RECT 97.445 112.135 97.615 112.935 ;
        RECT 97.820 112.255 98.095 112.735 ;
        RECT 97.815 112.085 98.095 112.255 ;
        RECT 97.100 111.940 97.275 111.975 ;
        RECT 96.345 111.405 96.675 111.805 ;
        RECT 97.100 111.575 97.630 111.940 ;
        RECT 97.820 111.575 98.095 112.085 ;
        RECT 98.265 111.575 98.455 112.935 ;
        RECT 98.625 112.950 98.795 113.615 ;
        RECT 98.965 113.195 99.135 113.955 ;
        RECT 99.370 113.195 99.885 113.605 ;
        RECT 98.625 112.760 99.375 112.950 ;
        RECT 99.545 112.385 99.885 113.195 ;
        RECT 100.055 112.865 103.565 113.955 ;
        RECT 103.735 112.865 104.945 113.955 ;
        RECT 98.655 112.215 99.885 112.385 ;
        RECT 98.635 111.405 99.145 111.940 ;
        RECT 99.365 111.610 99.610 112.215 ;
        RECT 100.055 112.175 101.705 112.695 ;
        RECT 101.875 112.345 103.565 112.865 ;
        RECT 100.055 111.405 103.565 112.175 ;
        RECT 103.735 112.155 104.255 112.695 ;
        RECT 104.425 112.325 104.945 112.865 ;
        RECT 105.120 112.815 105.455 113.785 ;
        RECT 105.625 112.815 105.795 113.955 ;
        RECT 105.965 113.615 107.995 113.785 ;
        RECT 103.735 111.405 104.945 112.155 ;
        RECT 105.120 112.145 105.290 112.815 ;
        RECT 105.965 112.645 106.135 113.615 ;
        RECT 105.460 112.315 105.715 112.645 ;
        RECT 105.940 112.315 106.135 112.645 ;
        RECT 106.305 113.275 107.430 113.445 ;
        RECT 105.545 112.145 105.715 112.315 ;
        RECT 106.305 112.145 106.475 113.275 ;
        RECT 105.120 111.575 105.375 112.145 ;
        RECT 105.545 111.975 106.475 112.145 ;
        RECT 106.645 112.935 107.655 113.105 ;
        RECT 106.645 112.135 106.815 112.935 ;
        RECT 106.300 111.940 106.475 111.975 ;
        RECT 105.545 111.405 105.875 111.805 ;
        RECT 106.300 111.575 106.830 111.940 ;
        RECT 107.020 111.915 107.295 112.735 ;
        RECT 107.015 111.745 107.295 111.915 ;
        RECT 107.020 111.575 107.295 111.745 ;
        RECT 107.465 111.575 107.655 112.935 ;
        RECT 107.825 112.950 107.995 113.615 ;
        RECT 108.165 113.195 108.335 113.955 ;
        RECT 108.570 113.195 109.085 113.605 ;
        RECT 107.825 112.760 108.575 112.950 ;
        RECT 108.745 112.385 109.085 113.195 ;
        RECT 107.855 112.215 109.085 112.385 ;
        RECT 109.715 112.880 109.985 113.785 ;
        RECT 110.155 113.195 110.485 113.955 ;
        RECT 110.665 113.025 110.835 113.785 ;
        RECT 107.835 111.405 108.345 111.940 ;
        RECT 108.565 111.610 108.810 112.215 ;
        RECT 109.715 112.080 109.885 112.880 ;
        RECT 110.170 112.855 110.835 113.025 ;
        RECT 111.095 112.865 112.765 113.955 ;
        RECT 110.170 112.710 110.340 112.855 ;
        RECT 110.055 112.380 110.340 112.710 ;
        RECT 110.170 112.125 110.340 112.380 ;
        RECT 110.575 112.305 110.905 112.675 ;
        RECT 111.095 112.175 111.845 112.695 ;
        RECT 112.015 112.345 112.765 112.865 ;
        RECT 112.935 112.790 113.225 113.955 ;
        RECT 113.595 113.285 113.875 113.955 ;
        RECT 114.045 113.065 114.345 113.615 ;
        RECT 114.545 113.235 114.875 113.955 ;
        RECT 115.065 113.235 115.525 113.785 ;
        RECT 113.410 112.645 113.675 113.005 ;
        RECT 114.045 112.895 114.985 113.065 ;
        RECT 114.815 112.645 114.985 112.895 ;
        RECT 113.410 112.395 114.085 112.645 ;
        RECT 114.305 112.395 114.645 112.645 ;
        RECT 114.815 112.315 115.105 112.645 ;
        RECT 114.815 112.225 114.985 112.315 ;
        RECT 109.715 111.575 109.975 112.080 ;
        RECT 110.170 111.955 110.835 112.125 ;
        RECT 110.155 111.405 110.485 111.785 ;
        RECT 110.665 111.575 110.835 111.955 ;
        RECT 111.095 111.405 112.765 112.175 ;
        RECT 112.935 111.405 113.225 112.130 ;
        RECT 113.595 112.035 114.985 112.225 ;
        RECT 113.595 111.675 113.925 112.035 ;
        RECT 115.275 111.865 115.525 113.235 ;
        RECT 115.875 113.040 116.045 113.955 ;
        RECT 116.215 112.895 116.545 113.740 ;
        RECT 116.715 112.945 116.885 113.955 ;
        RECT 117.055 113.225 117.395 113.785 ;
        RECT 117.625 113.455 117.940 113.955 ;
        RECT 118.120 113.485 119.005 113.655 ;
        RECT 116.155 112.815 116.545 112.895 ;
        RECT 117.055 112.850 117.950 113.225 ;
        RECT 116.155 112.765 116.370 112.815 ;
        RECT 116.155 112.185 116.325 112.765 ;
        RECT 117.055 112.645 117.245 112.850 ;
        RECT 118.120 112.645 118.290 113.485 ;
        RECT 119.230 113.455 119.480 113.785 ;
        RECT 116.495 112.315 117.245 112.645 ;
        RECT 117.415 112.315 118.290 112.645 ;
        RECT 116.155 112.145 116.380 112.185 ;
        RECT 117.045 112.145 117.245 112.315 ;
        RECT 116.155 112.060 116.535 112.145 ;
        RECT 114.545 111.405 114.795 111.865 ;
        RECT 114.965 111.575 115.525 111.865 ;
        RECT 115.865 111.405 116.035 111.920 ;
        RECT 116.205 111.625 116.535 112.060 ;
        RECT 116.705 111.405 116.875 112.015 ;
        RECT 117.045 111.620 117.375 112.145 ;
        RECT 117.635 111.405 117.845 111.935 ;
        RECT 118.120 111.855 118.290 112.315 ;
        RECT 118.460 112.355 118.780 113.315 ;
        RECT 118.950 112.565 119.140 113.285 ;
        RECT 119.310 112.385 119.480 113.455 ;
        RECT 119.650 113.155 119.820 113.955 ;
        RECT 119.990 113.510 121.095 113.680 ;
        RECT 119.990 112.895 120.160 113.510 ;
        RECT 121.305 113.360 121.555 113.785 ;
        RECT 121.725 113.495 121.990 113.955 ;
        RECT 120.330 112.975 120.860 113.340 ;
        RECT 121.305 113.230 121.610 113.360 ;
        RECT 119.650 112.805 120.160 112.895 ;
        RECT 119.650 112.635 120.520 112.805 ;
        RECT 119.650 112.565 119.820 112.635 ;
        RECT 119.940 112.385 120.140 112.415 ;
        RECT 118.460 112.025 118.925 112.355 ;
        RECT 119.310 112.085 120.140 112.385 ;
        RECT 119.310 111.855 119.480 112.085 ;
        RECT 118.120 111.685 118.905 111.855 ;
        RECT 119.075 111.685 119.480 111.855 ;
        RECT 119.660 111.405 120.030 111.905 ;
        RECT 120.350 111.855 120.520 112.635 ;
        RECT 120.690 112.275 120.860 112.975 ;
        RECT 121.030 112.445 121.270 113.040 ;
        RECT 120.690 112.055 121.215 112.275 ;
        RECT 121.440 112.125 121.610 113.230 ;
        RECT 121.385 111.995 121.610 112.125 ;
        RECT 121.780 112.035 122.060 112.985 ;
        RECT 121.385 111.855 121.555 111.995 ;
        RECT 120.350 111.685 121.025 111.855 ;
        RECT 121.220 111.685 121.555 111.855 ;
        RECT 121.725 111.405 121.975 111.865 ;
        RECT 122.230 111.665 122.415 113.785 ;
        RECT 122.585 113.455 122.915 113.955 ;
        RECT 123.085 113.285 123.255 113.785 ;
        RECT 122.590 113.115 123.255 113.285 ;
        RECT 122.590 112.125 122.820 113.115 ;
        RECT 122.990 112.295 123.340 112.945 ;
        RECT 123.515 112.865 125.185 113.955 ;
        RECT 125.445 113.285 125.615 113.785 ;
        RECT 125.785 113.455 126.115 113.955 ;
        RECT 125.445 113.115 126.110 113.285 ;
        RECT 123.515 112.175 124.265 112.695 ;
        RECT 124.435 112.345 125.185 112.865 ;
        RECT 125.360 112.295 125.710 112.945 ;
        RECT 122.590 111.955 123.255 112.125 ;
        RECT 122.585 111.405 122.915 111.785 ;
        RECT 123.085 111.665 123.255 111.955 ;
        RECT 123.515 111.405 125.185 112.175 ;
        RECT 125.880 112.125 126.110 113.115 ;
        RECT 125.445 111.955 126.110 112.125 ;
        RECT 125.445 111.665 125.615 111.955 ;
        RECT 125.785 111.405 126.115 111.785 ;
        RECT 126.285 111.665 126.470 113.785 ;
        RECT 126.710 113.495 126.975 113.955 ;
        RECT 127.145 113.360 127.395 113.785 ;
        RECT 127.605 113.510 128.710 113.680 ;
        RECT 127.090 113.230 127.395 113.360 ;
        RECT 126.640 112.035 126.920 112.985 ;
        RECT 127.090 112.125 127.260 113.230 ;
        RECT 127.430 112.445 127.670 113.040 ;
        RECT 127.840 112.975 128.370 113.340 ;
        RECT 127.840 112.275 128.010 112.975 ;
        RECT 128.540 112.895 128.710 113.510 ;
        RECT 128.880 113.155 129.050 113.955 ;
        RECT 129.220 113.455 129.470 113.785 ;
        RECT 129.695 113.485 130.580 113.655 ;
        RECT 128.540 112.805 129.050 112.895 ;
        RECT 127.090 111.995 127.315 112.125 ;
        RECT 127.485 112.055 128.010 112.275 ;
        RECT 128.180 112.635 129.050 112.805 ;
        RECT 126.725 111.405 126.975 111.865 ;
        RECT 127.145 111.855 127.315 111.995 ;
        RECT 128.180 111.855 128.350 112.635 ;
        RECT 128.880 112.565 129.050 112.635 ;
        RECT 128.560 112.385 128.760 112.415 ;
        RECT 129.220 112.385 129.390 113.455 ;
        RECT 129.560 112.565 129.750 113.285 ;
        RECT 128.560 112.085 129.390 112.385 ;
        RECT 129.920 112.355 130.240 113.315 ;
        RECT 127.145 111.685 127.480 111.855 ;
        RECT 127.675 111.685 128.350 111.855 ;
        RECT 128.670 111.405 129.040 111.905 ;
        RECT 129.220 111.855 129.390 112.085 ;
        RECT 129.775 112.025 130.240 112.355 ;
        RECT 130.410 112.645 130.580 113.485 ;
        RECT 130.760 113.455 131.075 113.955 ;
        RECT 131.305 113.225 131.645 113.785 ;
        RECT 130.750 112.850 131.645 113.225 ;
        RECT 131.815 112.945 131.985 113.955 ;
        RECT 131.455 112.645 131.645 112.850 ;
        RECT 132.155 112.895 132.485 113.740 ;
        RECT 132.155 112.815 132.545 112.895 ;
        RECT 132.330 112.765 132.545 112.815 ;
        RECT 130.410 112.315 131.285 112.645 ;
        RECT 131.455 112.315 132.205 112.645 ;
        RECT 130.410 111.855 130.580 112.315 ;
        RECT 131.455 112.145 131.655 112.315 ;
        RECT 132.375 112.185 132.545 112.765 ;
        RECT 132.320 112.145 132.545 112.185 ;
        RECT 129.220 111.685 129.625 111.855 ;
        RECT 129.795 111.685 130.580 111.855 ;
        RECT 130.855 111.405 131.065 111.935 ;
        RECT 131.325 111.620 131.655 112.145 ;
        RECT 132.165 112.060 132.545 112.145 ;
        RECT 131.825 111.405 131.995 112.015 ;
        RECT 132.165 111.625 132.495 112.060 ;
        RECT 133.175 111.685 133.455 113.785 ;
        RECT 133.645 113.195 134.430 113.955 ;
        RECT 134.825 113.125 135.210 113.785 ;
        RECT 134.825 113.025 135.235 113.125 ;
        RECT 133.625 112.815 135.235 113.025 ;
        RECT 135.535 112.935 135.735 113.725 ;
        RECT 133.625 112.215 133.900 112.815 ;
        RECT 135.405 112.765 135.735 112.935 ;
        RECT 135.905 112.775 136.225 113.955 ;
        RECT 136.395 113.235 136.855 113.785 ;
        RECT 137.045 113.235 137.375 113.955 ;
        RECT 135.405 112.645 135.585 112.765 ;
        RECT 134.070 112.395 134.425 112.645 ;
        RECT 134.620 112.595 135.085 112.645 ;
        RECT 134.615 112.425 135.085 112.595 ;
        RECT 134.620 112.395 135.085 112.425 ;
        RECT 135.255 112.395 135.585 112.645 ;
        RECT 135.760 112.395 136.225 112.595 ;
        RECT 133.625 112.035 134.875 112.215 ;
        RECT 134.510 111.965 134.875 112.035 ;
        RECT 135.045 112.015 136.225 112.185 ;
        RECT 133.685 111.405 133.855 111.865 ;
        RECT 135.045 111.795 135.375 112.015 ;
        RECT 134.125 111.615 135.375 111.795 ;
        RECT 135.545 111.405 135.715 111.845 ;
        RECT 135.885 111.600 136.225 112.015 ;
        RECT 136.395 111.865 136.645 113.235 ;
        RECT 137.575 113.065 137.875 113.615 ;
        RECT 138.045 113.285 138.325 113.955 ;
        RECT 136.935 112.895 137.875 113.065 ;
        RECT 136.935 112.645 137.105 112.895 ;
        RECT 138.245 112.645 138.510 113.005 ;
        RECT 138.695 112.790 138.985 113.955 ;
        RECT 139.155 112.815 139.435 113.955 ;
        RECT 139.605 112.805 139.935 113.785 ;
        RECT 140.105 112.815 140.365 113.955 ;
        RECT 140.740 112.985 141.070 113.785 ;
        RECT 141.240 113.155 141.570 113.955 ;
        RECT 141.870 112.985 142.200 113.785 ;
        RECT 142.845 113.155 143.095 113.955 ;
        RECT 140.740 112.815 143.175 112.985 ;
        RECT 143.365 112.815 143.535 113.955 ;
        RECT 143.705 112.815 144.045 113.785 ;
        RECT 136.815 112.315 137.105 112.645 ;
        RECT 137.275 112.395 137.615 112.645 ;
        RECT 137.835 112.395 138.510 112.645 ;
        RECT 139.165 112.375 139.500 112.645 ;
        RECT 136.935 112.225 137.105 112.315 ;
        RECT 136.935 112.035 138.325 112.225 ;
        RECT 139.670 112.205 139.840 112.805 ;
        RECT 140.010 112.395 140.345 112.645 ;
        RECT 140.535 112.395 140.885 112.645 ;
        RECT 136.395 111.575 136.955 111.865 ;
        RECT 137.125 111.405 137.375 111.865 ;
        RECT 137.995 111.675 138.325 112.035 ;
        RECT 138.695 111.405 138.985 112.130 ;
        RECT 139.155 111.405 139.465 112.205 ;
        RECT 139.670 111.575 140.365 112.205 ;
        RECT 141.070 112.185 141.240 112.815 ;
        RECT 141.410 112.395 141.740 112.595 ;
        RECT 141.910 112.395 142.240 112.595 ;
        RECT 142.410 112.395 142.830 112.595 ;
        RECT 143.005 112.565 143.175 112.815 ;
        RECT 143.005 112.395 143.700 112.565 ;
        RECT 140.740 111.575 141.240 112.185 ;
        RECT 141.870 112.055 143.095 112.225 ;
        RECT 143.870 112.205 144.045 112.815 ;
        RECT 141.870 111.575 142.200 112.055 ;
        RECT 142.370 111.405 142.595 111.865 ;
        RECT 142.765 111.575 143.095 112.055 ;
        RECT 143.285 111.405 143.535 112.205 ;
        RECT 143.705 111.575 144.045 112.205 ;
        RECT 144.250 113.165 144.785 113.785 ;
        RECT 144.250 112.145 144.565 113.165 ;
        RECT 144.955 113.155 145.285 113.955 ;
        RECT 145.770 112.985 146.160 113.160 ;
        RECT 146.525 113.145 146.820 113.955 ;
        RECT 144.735 112.815 146.160 112.985 ;
        RECT 144.735 112.315 144.905 112.815 ;
        RECT 144.250 111.575 144.865 112.145 ;
        RECT 145.155 112.085 145.420 112.645 ;
        RECT 145.590 111.915 145.760 112.815 ;
        RECT 147.000 112.645 147.245 113.785 ;
        RECT 147.420 113.145 147.680 113.955 ;
        RECT 148.280 113.950 154.555 113.955 ;
        RECT 147.860 112.645 148.110 113.780 ;
        RECT 148.280 113.155 148.540 113.950 ;
        RECT 148.710 113.055 148.970 113.780 ;
        RECT 149.140 113.225 149.400 113.950 ;
        RECT 149.570 113.055 149.830 113.780 ;
        RECT 150.000 113.225 150.260 113.950 ;
        RECT 150.430 113.055 150.690 113.780 ;
        RECT 150.860 113.225 151.120 113.950 ;
        RECT 151.290 113.055 151.550 113.780 ;
        RECT 151.720 113.225 151.965 113.950 ;
        RECT 152.135 113.055 152.395 113.780 ;
        RECT 152.580 113.225 152.825 113.950 ;
        RECT 152.995 113.055 153.255 113.780 ;
        RECT 153.440 113.225 153.685 113.950 ;
        RECT 153.855 113.055 154.115 113.780 ;
        RECT 154.300 113.225 154.555 113.950 ;
        RECT 148.710 113.040 154.115 113.055 ;
        RECT 154.725 113.040 155.015 113.780 ;
        RECT 155.185 113.210 155.455 113.955 ;
        RECT 148.710 112.815 155.455 113.040 ;
        RECT 145.930 112.085 146.285 112.645 ;
        RECT 146.515 112.085 146.830 112.645 ;
        RECT 147.000 112.395 154.120 112.645 ;
        RECT 145.035 111.405 145.250 111.915 ;
        RECT 145.480 111.585 145.760 111.915 ;
        RECT 145.940 111.405 146.180 111.915 ;
        RECT 146.515 111.405 146.820 111.915 ;
        RECT 147.000 111.585 147.250 112.395 ;
        RECT 147.420 111.405 147.680 111.930 ;
        RECT 147.860 111.585 148.110 112.395 ;
        RECT 154.290 112.225 155.455 112.815 ;
        RECT 155.715 112.865 156.925 113.955 ;
        RECT 155.715 112.325 156.235 112.865 ;
        RECT 148.710 112.055 155.455 112.225 ;
        RECT 156.405 112.155 156.925 112.695 ;
        RECT 148.280 111.405 148.540 111.965 ;
        RECT 148.710 111.600 148.970 112.055 ;
        RECT 149.140 111.405 149.400 111.885 ;
        RECT 149.570 111.600 149.830 112.055 ;
        RECT 150.000 111.405 150.260 111.885 ;
        RECT 150.430 111.600 150.690 112.055 ;
        RECT 150.860 111.405 151.105 111.885 ;
        RECT 151.275 111.600 151.550 112.055 ;
        RECT 151.720 111.405 151.965 111.885 ;
        RECT 152.135 111.600 152.395 112.055 ;
        RECT 152.575 111.405 152.825 111.885 ;
        RECT 152.995 111.600 153.255 112.055 ;
        RECT 153.435 111.405 153.685 111.885 ;
        RECT 153.855 111.600 154.115 112.055 ;
        RECT 154.295 111.405 154.555 111.885 ;
        RECT 154.725 111.600 154.985 112.055 ;
        RECT 155.155 111.405 155.455 111.885 ;
        RECT 155.715 111.405 156.925 112.155 ;
        RECT 22.690 111.235 157.010 111.405 ;
        RECT 22.775 110.485 23.985 111.235 ;
        RECT 24.245 110.685 24.415 110.975 ;
        RECT 24.585 110.855 24.915 111.235 ;
        RECT 24.245 110.515 24.910 110.685 ;
        RECT 22.775 109.945 23.295 110.485 ;
        RECT 23.465 109.775 23.985 110.315 ;
        RECT 22.775 108.685 23.985 109.775 ;
        RECT 24.160 109.695 24.510 110.345 ;
        RECT 24.680 109.525 24.910 110.515 ;
        RECT 24.245 109.355 24.910 109.525 ;
        RECT 24.245 108.855 24.415 109.355 ;
        RECT 24.585 108.685 24.915 109.185 ;
        RECT 25.085 108.855 25.270 110.975 ;
        RECT 25.525 110.775 25.775 111.235 ;
        RECT 25.945 110.785 26.280 110.955 ;
        RECT 26.475 110.785 27.150 110.955 ;
        RECT 25.945 110.645 26.115 110.785 ;
        RECT 25.440 109.655 25.720 110.605 ;
        RECT 25.890 110.515 26.115 110.645 ;
        RECT 25.890 109.410 26.060 110.515 ;
        RECT 26.285 110.365 26.810 110.585 ;
        RECT 26.230 109.600 26.470 110.195 ;
        RECT 26.640 109.665 26.810 110.365 ;
        RECT 26.980 110.005 27.150 110.785 ;
        RECT 27.470 110.735 27.840 111.235 ;
        RECT 28.020 110.785 28.425 110.955 ;
        RECT 28.595 110.785 29.380 110.955 ;
        RECT 28.020 110.555 28.190 110.785 ;
        RECT 27.360 110.255 28.190 110.555 ;
        RECT 28.575 110.285 29.040 110.615 ;
        RECT 27.360 110.225 27.560 110.255 ;
        RECT 27.680 110.005 27.850 110.075 ;
        RECT 26.980 109.835 27.850 110.005 ;
        RECT 27.340 109.745 27.850 109.835 ;
        RECT 25.890 109.280 26.195 109.410 ;
        RECT 26.640 109.300 27.170 109.665 ;
        RECT 25.510 108.685 25.775 109.145 ;
        RECT 25.945 108.855 26.195 109.280 ;
        RECT 27.340 109.130 27.510 109.745 ;
        RECT 26.405 108.960 27.510 109.130 ;
        RECT 27.680 108.685 27.850 109.485 ;
        RECT 28.020 109.185 28.190 110.255 ;
        RECT 28.360 109.355 28.550 110.075 ;
        RECT 28.720 109.325 29.040 110.285 ;
        RECT 29.210 110.325 29.380 110.785 ;
        RECT 29.655 110.705 29.865 111.235 ;
        RECT 30.125 110.495 30.455 111.020 ;
        RECT 30.625 110.625 30.795 111.235 ;
        RECT 30.965 110.580 31.295 111.015 ;
        RECT 30.965 110.495 31.345 110.580 ;
        RECT 30.255 110.325 30.455 110.495 ;
        RECT 31.120 110.455 31.345 110.495 ;
        RECT 29.210 109.995 30.085 110.325 ;
        RECT 30.255 109.995 31.005 110.325 ;
        RECT 28.020 108.855 28.270 109.185 ;
        RECT 29.210 109.155 29.380 109.995 ;
        RECT 30.255 109.790 30.445 109.995 ;
        RECT 31.175 109.875 31.345 110.455 ;
        RECT 31.520 110.395 31.780 111.235 ;
        RECT 31.955 110.490 32.210 111.065 ;
        RECT 32.380 110.855 32.710 111.235 ;
        RECT 32.925 110.685 33.095 111.065 ;
        RECT 32.380 110.515 33.095 110.685 ;
        RECT 33.445 110.685 33.615 110.975 ;
        RECT 33.785 110.855 34.115 111.235 ;
        RECT 33.445 110.515 34.110 110.685 ;
        RECT 31.130 109.825 31.345 109.875 ;
        RECT 29.550 109.415 30.445 109.790 ;
        RECT 30.955 109.745 31.345 109.825 ;
        RECT 28.495 108.985 29.380 109.155 ;
        RECT 29.560 108.685 29.875 109.185 ;
        RECT 30.105 108.855 30.445 109.415 ;
        RECT 30.615 108.685 30.785 109.695 ;
        RECT 30.955 108.900 31.285 109.745 ;
        RECT 31.520 108.685 31.780 109.835 ;
        RECT 31.955 109.760 32.125 110.490 ;
        RECT 32.380 110.325 32.550 110.515 ;
        RECT 32.295 109.995 32.550 110.325 ;
        RECT 32.380 109.785 32.550 109.995 ;
        RECT 32.830 109.965 33.185 110.335 ;
        RECT 31.955 108.855 32.210 109.760 ;
        RECT 32.380 109.615 33.095 109.785 ;
        RECT 33.360 109.695 33.710 110.345 ;
        RECT 32.380 108.685 32.710 109.445 ;
        RECT 32.925 108.855 33.095 109.615 ;
        RECT 33.880 109.525 34.110 110.515 ;
        RECT 33.445 109.355 34.110 109.525 ;
        RECT 33.445 108.855 33.615 109.355 ;
        RECT 33.785 108.685 34.115 109.185 ;
        RECT 34.285 108.855 34.470 110.975 ;
        RECT 34.725 110.775 34.975 111.235 ;
        RECT 35.145 110.785 35.480 110.955 ;
        RECT 35.675 110.785 36.350 110.955 ;
        RECT 35.145 110.645 35.315 110.785 ;
        RECT 34.640 109.655 34.920 110.605 ;
        RECT 35.090 110.515 35.315 110.645 ;
        RECT 35.090 109.410 35.260 110.515 ;
        RECT 35.485 110.365 36.010 110.585 ;
        RECT 35.430 109.600 35.670 110.195 ;
        RECT 35.840 109.665 36.010 110.365 ;
        RECT 36.180 110.005 36.350 110.785 ;
        RECT 36.670 110.735 37.040 111.235 ;
        RECT 37.220 110.785 37.625 110.955 ;
        RECT 37.795 110.785 38.580 110.955 ;
        RECT 37.220 110.555 37.390 110.785 ;
        RECT 36.560 110.255 37.390 110.555 ;
        RECT 37.775 110.285 38.240 110.615 ;
        RECT 36.560 110.225 36.760 110.255 ;
        RECT 36.880 110.005 37.050 110.075 ;
        RECT 36.180 109.835 37.050 110.005 ;
        RECT 36.540 109.745 37.050 109.835 ;
        RECT 35.090 109.280 35.395 109.410 ;
        RECT 35.840 109.300 36.370 109.665 ;
        RECT 34.710 108.685 34.975 109.145 ;
        RECT 35.145 108.855 35.395 109.280 ;
        RECT 36.540 109.130 36.710 109.745 ;
        RECT 35.605 108.960 36.710 109.130 ;
        RECT 36.880 108.685 37.050 109.485 ;
        RECT 37.220 109.185 37.390 110.255 ;
        RECT 37.560 109.355 37.750 110.075 ;
        RECT 37.920 109.325 38.240 110.285 ;
        RECT 38.410 110.325 38.580 110.785 ;
        RECT 38.855 110.705 39.065 111.235 ;
        RECT 39.325 110.495 39.655 111.020 ;
        RECT 39.825 110.625 39.995 111.235 ;
        RECT 40.165 110.580 40.495 111.015 ;
        RECT 40.880 110.725 41.120 111.235 ;
        RECT 41.300 110.725 41.580 111.055 ;
        RECT 41.810 110.725 42.025 111.235 ;
        RECT 40.165 110.495 40.545 110.580 ;
        RECT 39.455 110.325 39.655 110.495 ;
        RECT 40.320 110.455 40.545 110.495 ;
        RECT 38.410 109.995 39.285 110.325 ;
        RECT 39.455 109.995 40.205 110.325 ;
        RECT 37.220 108.855 37.470 109.185 ;
        RECT 38.410 109.155 38.580 109.995 ;
        RECT 39.455 109.790 39.645 109.995 ;
        RECT 40.375 109.875 40.545 110.455 ;
        RECT 40.775 109.995 41.130 110.555 ;
        RECT 40.330 109.825 40.545 109.875 ;
        RECT 41.300 109.825 41.470 110.725 ;
        RECT 41.640 109.995 41.905 110.555 ;
        RECT 42.195 110.495 42.810 111.065 ;
        RECT 42.155 109.825 42.325 110.325 ;
        RECT 38.750 109.415 39.645 109.790 ;
        RECT 40.155 109.745 40.545 109.825 ;
        RECT 37.695 108.985 38.580 109.155 ;
        RECT 38.760 108.685 39.075 109.185 ;
        RECT 39.305 108.855 39.645 109.415 ;
        RECT 39.815 108.685 39.985 109.695 ;
        RECT 40.155 108.900 40.485 109.745 ;
        RECT 40.900 109.655 42.325 109.825 ;
        RECT 40.900 109.480 41.290 109.655 ;
        RECT 41.775 108.685 42.105 109.485 ;
        RECT 42.495 109.475 42.810 110.495 ;
        RECT 42.275 108.855 42.810 109.475 ;
        RECT 43.015 110.435 43.355 111.065 ;
        RECT 43.525 110.435 43.775 111.235 ;
        RECT 43.965 110.585 44.295 111.065 ;
        RECT 44.465 110.775 44.690 111.235 ;
        RECT 44.860 110.585 45.190 111.065 ;
        RECT 43.015 109.825 43.190 110.435 ;
        RECT 43.965 110.415 45.190 110.585 ;
        RECT 45.820 110.455 46.320 111.065 ;
        RECT 46.695 110.465 48.365 111.235 ;
        RECT 48.535 110.510 48.825 111.235 ;
        RECT 49.455 110.495 49.840 111.065 ;
        RECT 50.010 110.775 50.335 111.235 ;
        RECT 50.855 110.605 51.135 111.065 ;
        RECT 43.360 110.075 44.055 110.245 ;
        RECT 43.885 109.825 44.055 110.075 ;
        RECT 44.230 110.045 44.650 110.245 ;
        RECT 44.820 110.045 45.150 110.245 ;
        RECT 45.320 110.045 45.650 110.245 ;
        RECT 45.820 109.825 45.990 110.455 ;
        RECT 46.175 109.995 46.525 110.245 ;
        RECT 46.695 109.945 47.445 110.465 ;
        RECT 43.015 108.855 43.355 109.825 ;
        RECT 43.525 108.685 43.695 109.825 ;
        RECT 43.885 109.655 46.320 109.825 ;
        RECT 47.615 109.775 48.365 110.295 ;
        RECT 43.965 108.685 44.215 109.485 ;
        RECT 44.860 108.855 45.190 109.655 ;
        RECT 45.490 108.685 45.820 109.485 ;
        RECT 45.990 108.855 46.320 109.655 ;
        RECT 46.695 108.685 48.365 109.775 ;
        RECT 48.535 108.685 48.825 109.850 ;
        RECT 49.455 109.825 49.735 110.495 ;
        RECT 50.010 110.435 51.135 110.605 ;
        RECT 50.010 110.325 50.460 110.435 ;
        RECT 49.905 109.995 50.460 110.325 ;
        RECT 51.325 110.265 51.725 111.065 ;
        RECT 52.125 110.775 52.395 111.235 ;
        RECT 52.565 110.605 52.850 111.065 ;
        RECT 53.145 110.735 53.475 111.235 ;
        RECT 49.455 108.855 49.840 109.825 ;
        RECT 50.010 109.535 50.460 109.995 ;
        RECT 50.630 109.705 51.725 110.265 ;
        RECT 50.010 109.315 51.135 109.535 ;
        RECT 50.010 108.685 50.335 109.145 ;
        RECT 50.855 108.855 51.135 109.315 ;
        RECT 51.325 108.855 51.725 109.705 ;
        RECT 51.895 110.435 52.850 110.605 ;
        RECT 53.675 110.665 53.845 111.015 ;
        RECT 54.045 110.835 54.375 111.235 ;
        RECT 54.545 110.665 54.715 111.015 ;
        RECT 54.885 110.835 55.265 111.235 ;
        RECT 51.895 109.535 52.105 110.435 ;
        RECT 52.275 109.705 52.965 110.265 ;
        RECT 53.140 109.995 53.490 110.565 ;
        RECT 53.675 110.495 55.285 110.665 ;
        RECT 55.455 110.560 55.725 110.905 ;
        RECT 55.115 110.325 55.285 110.495 ;
        RECT 53.140 109.535 53.460 109.825 ;
        RECT 53.660 109.705 54.370 110.325 ;
        RECT 54.540 109.995 54.945 110.325 ;
        RECT 55.115 109.995 55.385 110.325 ;
        RECT 55.115 109.825 55.285 109.995 ;
        RECT 55.555 109.825 55.725 110.560 ;
        RECT 54.560 109.655 55.285 109.825 ;
        RECT 54.560 109.535 54.730 109.655 ;
        RECT 51.895 109.315 52.850 109.535 ;
        RECT 53.140 109.365 54.730 109.535 ;
        RECT 52.125 108.685 52.395 109.145 ;
        RECT 52.565 108.855 52.850 109.315 ;
        RECT 53.140 108.905 54.795 109.195 ;
        RECT 54.965 108.685 55.245 109.485 ;
        RECT 55.455 108.855 55.725 109.825 ;
        RECT 55.930 110.495 56.545 111.065 ;
        RECT 56.715 110.725 56.930 111.235 ;
        RECT 57.160 110.725 57.440 111.055 ;
        RECT 57.620 110.725 57.860 111.235 ;
        RECT 55.930 109.475 56.245 110.495 ;
        RECT 56.415 109.825 56.585 110.325 ;
        RECT 56.835 109.995 57.100 110.555 ;
        RECT 57.270 109.825 57.440 110.725 ;
        RECT 57.610 109.995 57.965 110.555 ;
        RECT 58.655 110.495 59.040 111.065 ;
        RECT 59.210 110.775 59.535 111.235 ;
        RECT 60.055 110.605 60.335 111.065 ;
        RECT 58.655 109.825 58.935 110.495 ;
        RECT 59.210 110.435 60.335 110.605 ;
        RECT 59.210 110.325 59.660 110.435 ;
        RECT 59.105 109.995 59.660 110.325 ;
        RECT 60.525 110.265 60.925 111.065 ;
        RECT 61.325 110.775 61.595 111.235 ;
        RECT 61.765 110.605 62.050 111.065 ;
        RECT 56.415 109.655 57.840 109.825 ;
        RECT 55.930 108.855 56.465 109.475 ;
        RECT 56.635 108.685 56.965 109.485 ;
        RECT 57.450 109.480 57.840 109.655 ;
        RECT 58.655 108.855 59.040 109.825 ;
        RECT 59.210 109.535 59.660 109.995 ;
        RECT 59.830 109.705 60.925 110.265 ;
        RECT 59.210 109.315 60.335 109.535 ;
        RECT 59.210 108.685 59.535 109.145 ;
        RECT 60.055 108.855 60.335 109.315 ;
        RECT 60.525 108.855 60.925 109.705 ;
        RECT 61.095 110.435 62.050 110.605 ;
        RECT 62.360 110.585 62.670 111.055 ;
        RECT 62.840 110.755 63.575 111.235 ;
        RECT 63.745 110.665 63.915 111.015 ;
        RECT 64.085 110.835 64.465 111.235 ;
        RECT 61.095 109.535 61.305 110.435 ;
        RECT 62.360 110.415 63.095 110.585 ;
        RECT 63.745 110.495 64.485 110.665 ;
        RECT 64.655 110.560 64.925 110.905 ;
        RECT 62.845 110.325 63.095 110.415 ;
        RECT 64.315 110.325 64.485 110.495 ;
        RECT 61.475 109.705 62.165 110.265 ;
        RECT 62.340 109.995 62.675 110.245 ;
        RECT 62.845 109.995 63.585 110.325 ;
        RECT 64.315 109.995 64.545 110.325 ;
        RECT 61.095 109.315 62.050 109.535 ;
        RECT 61.325 108.685 61.595 109.145 ;
        RECT 61.765 108.855 62.050 109.315 ;
        RECT 62.340 108.685 62.595 109.825 ;
        RECT 62.845 109.435 63.015 109.995 ;
        RECT 64.315 109.825 64.485 109.995 ;
        RECT 64.755 109.825 64.925 110.560 ;
        RECT 65.135 110.415 65.365 111.235 ;
        RECT 65.535 110.435 65.865 111.065 ;
        RECT 65.115 109.995 65.445 110.245 ;
        RECT 65.615 109.835 65.865 110.435 ;
        RECT 66.035 110.415 66.245 111.235 ;
        RECT 66.475 110.495 66.940 111.040 ;
        RECT 63.240 109.655 64.485 109.825 ;
        RECT 63.240 109.405 63.660 109.655 ;
        RECT 62.790 108.905 63.985 109.235 ;
        RECT 64.165 108.685 64.445 109.485 ;
        RECT 64.655 108.855 64.925 109.825 ;
        RECT 65.135 108.685 65.365 109.825 ;
        RECT 65.535 108.855 65.865 109.835 ;
        RECT 66.035 108.685 66.245 109.825 ;
        RECT 66.475 109.535 66.645 110.495 ;
        RECT 67.445 110.415 67.615 111.235 ;
        RECT 67.785 110.585 68.115 111.065 ;
        RECT 68.285 110.845 68.635 111.235 ;
        RECT 68.805 110.665 69.035 111.065 ;
        RECT 68.525 110.585 69.035 110.665 ;
        RECT 67.785 110.495 69.035 110.585 ;
        RECT 69.205 110.495 69.525 110.975 ;
        RECT 69.705 110.505 70.005 111.235 ;
        RECT 67.785 110.415 68.695 110.495 ;
        RECT 66.815 109.875 67.060 110.325 ;
        RECT 67.320 110.045 68.015 110.245 ;
        RECT 68.185 110.075 68.785 110.245 ;
        RECT 68.185 109.875 68.355 110.075 ;
        RECT 69.015 109.905 69.185 110.325 ;
        RECT 66.815 109.705 68.355 109.875 ;
        RECT 68.525 109.735 69.185 109.905 ;
        RECT 68.525 109.535 68.695 109.735 ;
        RECT 69.355 109.565 69.525 110.495 ;
        RECT 70.185 110.325 70.415 110.945 ;
        RECT 70.615 110.675 70.840 111.055 ;
        RECT 71.010 110.845 71.340 111.235 ;
        RECT 70.615 110.495 70.945 110.675 ;
        RECT 69.710 109.995 70.005 110.325 ;
        RECT 70.185 109.995 70.600 110.325 ;
        RECT 70.770 109.825 70.945 110.495 ;
        RECT 71.115 109.995 71.355 110.645 ;
        RECT 71.535 110.465 74.125 111.235 ;
        RECT 74.295 110.510 74.585 111.235 ;
        RECT 75.765 110.585 75.935 111.065 ;
        RECT 76.115 110.755 76.355 111.235 ;
        RECT 76.605 110.585 76.775 111.065 ;
        RECT 76.945 110.755 77.275 111.235 ;
        RECT 77.445 110.585 77.615 111.065 ;
        RECT 71.535 109.945 72.745 110.465 ;
        RECT 75.765 110.415 76.400 110.585 ;
        RECT 76.605 110.415 77.615 110.585 ;
        RECT 77.785 110.435 78.115 111.235 ;
        RECT 79.445 110.685 79.615 110.975 ;
        RECT 79.785 110.855 80.115 111.235 ;
        RECT 79.445 110.515 80.110 110.685 ;
        RECT 66.475 109.365 68.695 109.535 ;
        RECT 68.865 109.365 69.525 109.565 ;
        RECT 69.705 109.465 70.600 109.795 ;
        RECT 70.770 109.635 71.355 109.825 ;
        RECT 72.915 109.775 74.125 110.295 ;
        RECT 76.230 110.245 76.400 110.415 ;
        RECT 75.680 110.005 76.060 110.245 ;
        RECT 76.230 110.075 76.730 110.245 ;
        RECT 66.475 108.685 66.775 109.195 ;
        RECT 66.945 108.855 67.275 109.365 ;
        RECT 68.865 109.195 69.035 109.365 ;
        RECT 69.705 109.295 70.910 109.465 ;
        RECT 67.445 108.685 68.075 109.195 ;
        RECT 68.655 109.025 69.035 109.195 ;
        RECT 69.205 108.685 69.505 109.195 ;
        RECT 69.705 108.865 70.035 109.295 ;
        RECT 70.215 108.685 70.410 109.125 ;
        RECT 70.580 108.865 70.910 109.295 ;
        RECT 71.080 108.865 71.355 109.635 ;
        RECT 71.535 108.685 74.125 109.775 ;
        RECT 74.295 108.685 74.585 109.850 ;
        RECT 76.230 109.835 76.400 110.075 ;
        RECT 77.120 109.875 77.615 110.415 ;
        RECT 75.685 109.665 76.400 109.835 ;
        RECT 76.605 109.705 77.615 109.875 ;
        RECT 75.685 108.855 76.015 109.665 ;
        RECT 76.185 108.685 76.425 109.485 ;
        RECT 76.605 108.855 76.775 109.705 ;
        RECT 76.945 108.685 77.275 109.485 ;
        RECT 77.445 108.855 77.615 109.705 ;
        RECT 77.785 108.685 78.115 109.835 ;
        RECT 79.360 109.695 79.710 110.345 ;
        RECT 79.880 109.525 80.110 110.515 ;
        RECT 79.445 109.355 80.110 109.525 ;
        RECT 79.445 108.855 79.615 109.355 ;
        RECT 79.785 108.685 80.115 109.185 ;
        RECT 80.285 108.855 80.470 110.975 ;
        RECT 80.725 110.775 80.975 111.235 ;
        RECT 81.145 110.785 81.480 110.955 ;
        RECT 81.675 110.785 82.350 110.955 ;
        RECT 81.145 110.645 81.315 110.785 ;
        RECT 80.640 109.655 80.920 110.605 ;
        RECT 81.090 110.515 81.315 110.645 ;
        RECT 81.090 109.410 81.260 110.515 ;
        RECT 81.485 110.365 82.010 110.585 ;
        RECT 81.430 109.600 81.670 110.195 ;
        RECT 81.840 109.665 82.010 110.365 ;
        RECT 82.180 110.005 82.350 110.785 ;
        RECT 82.670 110.735 83.040 111.235 ;
        RECT 83.220 110.785 83.625 110.955 ;
        RECT 83.795 110.785 84.580 110.955 ;
        RECT 83.220 110.555 83.390 110.785 ;
        RECT 82.560 110.255 83.390 110.555 ;
        RECT 83.775 110.285 84.240 110.615 ;
        RECT 82.560 110.225 82.760 110.255 ;
        RECT 82.880 110.005 83.050 110.075 ;
        RECT 82.180 109.835 83.050 110.005 ;
        RECT 82.540 109.745 83.050 109.835 ;
        RECT 81.090 109.280 81.395 109.410 ;
        RECT 81.840 109.300 82.370 109.665 ;
        RECT 80.710 108.685 80.975 109.145 ;
        RECT 81.145 108.855 81.395 109.280 ;
        RECT 82.540 109.130 82.710 109.745 ;
        RECT 81.605 108.960 82.710 109.130 ;
        RECT 82.880 108.685 83.050 109.485 ;
        RECT 83.220 109.185 83.390 110.255 ;
        RECT 83.560 109.355 83.750 110.075 ;
        RECT 83.920 109.325 84.240 110.285 ;
        RECT 84.410 110.325 84.580 110.785 ;
        RECT 84.855 110.705 85.065 111.235 ;
        RECT 85.325 110.495 85.655 111.020 ;
        RECT 85.825 110.625 85.995 111.235 ;
        RECT 86.165 110.580 86.495 111.015 ;
        RECT 86.665 110.720 86.835 111.235 ;
        RECT 87.175 110.775 87.735 111.065 ;
        RECT 87.905 110.775 88.155 111.235 ;
        RECT 86.165 110.495 86.545 110.580 ;
        RECT 85.455 110.325 85.655 110.495 ;
        RECT 86.320 110.455 86.545 110.495 ;
        RECT 84.410 109.995 85.285 110.325 ;
        RECT 85.455 109.995 86.205 110.325 ;
        RECT 83.220 108.855 83.470 109.185 ;
        RECT 84.410 109.155 84.580 109.995 ;
        RECT 85.455 109.790 85.645 109.995 ;
        RECT 86.375 109.875 86.545 110.455 ;
        RECT 86.330 109.825 86.545 109.875 ;
        RECT 84.750 109.415 85.645 109.790 ;
        RECT 86.155 109.745 86.545 109.825 ;
        RECT 83.695 108.985 84.580 109.155 ;
        RECT 84.760 108.685 85.075 109.185 ;
        RECT 85.305 108.855 85.645 109.415 ;
        RECT 85.815 108.685 85.985 109.695 ;
        RECT 86.155 108.900 86.485 109.745 ;
        RECT 86.655 108.685 86.825 109.600 ;
        RECT 87.175 109.405 87.425 110.775 ;
        RECT 88.775 110.605 89.105 110.965 ;
        RECT 87.715 110.415 89.105 110.605 ;
        RECT 90.395 110.560 90.655 111.065 ;
        RECT 90.835 110.855 91.165 111.235 ;
        RECT 91.345 110.685 91.515 111.065 ;
        RECT 87.715 110.325 87.885 110.415 ;
        RECT 87.595 109.995 87.885 110.325 ;
        RECT 88.055 109.995 88.395 110.245 ;
        RECT 88.615 109.995 89.290 110.245 ;
        RECT 87.715 109.745 87.885 109.995 ;
        RECT 87.715 109.575 88.655 109.745 ;
        RECT 89.025 109.635 89.290 109.995 ;
        RECT 90.395 109.760 90.565 110.560 ;
        RECT 90.850 110.515 91.515 110.685 ;
        RECT 90.850 110.260 91.020 110.515 ;
        RECT 91.785 110.425 92.055 111.235 ;
        RECT 92.225 110.425 92.555 111.065 ;
        RECT 92.725 110.425 92.965 111.235 ;
        RECT 93.355 110.605 93.685 110.965 ;
        RECT 94.305 110.775 94.555 111.235 ;
        RECT 94.725 110.775 95.285 111.065 ;
        RECT 90.735 109.930 91.020 110.260 ;
        RECT 91.255 109.965 91.585 110.335 ;
        RECT 91.775 109.995 92.125 110.245 ;
        RECT 90.850 109.785 91.020 109.930 ;
        RECT 92.295 109.825 92.465 110.425 ;
        RECT 93.355 110.415 94.745 110.605 ;
        RECT 94.575 110.325 94.745 110.415 ;
        RECT 92.635 109.995 92.985 110.245 ;
        RECT 93.170 109.995 93.845 110.245 ;
        RECT 94.065 109.995 94.405 110.245 ;
        RECT 94.575 109.995 94.865 110.325 ;
        RECT 87.175 108.855 87.635 109.405 ;
        RECT 87.825 108.685 88.155 109.405 ;
        RECT 88.355 109.025 88.655 109.575 ;
        RECT 88.825 108.685 89.105 109.355 ;
        RECT 90.395 108.855 90.665 109.760 ;
        RECT 90.850 109.615 91.515 109.785 ;
        RECT 90.835 108.685 91.165 109.445 ;
        RECT 91.345 108.855 91.515 109.615 ;
        RECT 91.785 108.685 92.115 109.825 ;
        RECT 92.295 109.655 92.975 109.825 ;
        RECT 92.645 108.870 92.975 109.655 ;
        RECT 93.170 109.635 93.435 109.995 ;
        RECT 94.575 109.745 94.745 109.995 ;
        RECT 93.805 109.575 94.745 109.745 ;
        RECT 93.355 108.685 93.635 109.355 ;
        RECT 93.805 109.025 94.105 109.575 ;
        RECT 95.035 109.405 95.285 110.775 ;
        RECT 95.455 110.465 98.965 111.235 ;
        RECT 100.055 110.510 100.345 111.235 ;
        RECT 100.515 110.465 102.185 111.235 ;
        RECT 102.445 110.685 102.615 111.065 ;
        RECT 102.795 110.855 103.125 111.235 ;
        RECT 102.445 110.515 103.110 110.685 ;
        RECT 103.305 110.560 103.565 111.065 ;
        RECT 95.455 109.945 97.105 110.465 ;
        RECT 97.275 109.775 98.965 110.295 ;
        RECT 100.515 109.945 101.265 110.465 ;
        RECT 94.305 108.685 94.635 109.405 ;
        RECT 94.825 108.855 95.285 109.405 ;
        RECT 95.455 108.685 98.965 109.775 ;
        RECT 100.055 108.685 100.345 109.850 ;
        RECT 101.435 109.775 102.185 110.295 ;
        RECT 102.375 109.965 102.705 110.335 ;
        RECT 102.940 110.260 103.110 110.515 ;
        RECT 102.940 109.930 103.225 110.260 ;
        RECT 102.940 109.785 103.110 109.930 ;
        RECT 100.515 108.685 102.185 109.775 ;
        RECT 102.445 109.615 103.110 109.785 ;
        RECT 103.395 109.760 103.565 110.560 ;
        RECT 103.825 110.685 103.995 110.975 ;
        RECT 104.165 110.855 104.495 111.235 ;
        RECT 103.825 110.515 104.490 110.685 ;
        RECT 102.445 108.855 102.615 109.615 ;
        RECT 102.795 108.685 103.125 109.445 ;
        RECT 103.295 108.855 103.565 109.760 ;
        RECT 103.740 109.695 104.090 110.345 ;
        RECT 104.260 109.525 104.490 110.515 ;
        RECT 103.825 109.355 104.490 109.525 ;
        RECT 103.825 108.855 103.995 109.355 ;
        RECT 104.165 108.685 104.495 109.185 ;
        RECT 104.665 108.855 104.850 110.975 ;
        RECT 105.105 110.775 105.355 111.235 ;
        RECT 105.525 110.785 105.860 110.955 ;
        RECT 106.055 110.785 106.730 110.955 ;
        RECT 105.525 110.645 105.695 110.785 ;
        RECT 105.020 109.655 105.300 110.605 ;
        RECT 105.470 110.515 105.695 110.645 ;
        RECT 105.470 109.410 105.640 110.515 ;
        RECT 105.865 110.365 106.390 110.585 ;
        RECT 105.810 109.600 106.050 110.195 ;
        RECT 106.220 109.665 106.390 110.365 ;
        RECT 106.560 110.005 106.730 110.785 ;
        RECT 107.050 110.735 107.420 111.235 ;
        RECT 107.600 110.785 108.005 110.955 ;
        RECT 108.175 110.785 108.960 110.955 ;
        RECT 107.600 110.555 107.770 110.785 ;
        RECT 106.940 110.255 107.770 110.555 ;
        RECT 108.155 110.285 108.620 110.615 ;
        RECT 106.940 110.225 107.140 110.255 ;
        RECT 107.260 110.005 107.430 110.075 ;
        RECT 106.560 109.835 107.430 110.005 ;
        RECT 106.920 109.745 107.430 109.835 ;
        RECT 105.470 109.280 105.775 109.410 ;
        RECT 106.220 109.300 106.750 109.665 ;
        RECT 105.090 108.685 105.355 109.145 ;
        RECT 105.525 108.855 105.775 109.280 ;
        RECT 106.920 109.130 107.090 109.745 ;
        RECT 105.985 108.960 107.090 109.130 ;
        RECT 107.260 108.685 107.430 109.485 ;
        RECT 107.600 109.185 107.770 110.255 ;
        RECT 107.940 109.355 108.130 110.075 ;
        RECT 108.300 109.325 108.620 110.285 ;
        RECT 108.790 110.325 108.960 110.785 ;
        RECT 109.235 110.705 109.445 111.235 ;
        RECT 109.705 110.495 110.035 111.020 ;
        RECT 110.205 110.625 110.375 111.235 ;
        RECT 110.545 110.580 110.875 111.015 ;
        RECT 111.095 110.775 111.655 111.065 ;
        RECT 111.825 110.775 112.075 111.235 ;
        RECT 110.545 110.495 110.925 110.580 ;
        RECT 109.835 110.325 110.035 110.495 ;
        RECT 110.700 110.455 110.925 110.495 ;
        RECT 108.790 109.995 109.665 110.325 ;
        RECT 109.835 109.995 110.585 110.325 ;
        RECT 107.600 108.855 107.850 109.185 ;
        RECT 108.790 109.155 108.960 109.995 ;
        RECT 109.835 109.790 110.025 109.995 ;
        RECT 110.755 109.875 110.925 110.455 ;
        RECT 110.710 109.825 110.925 109.875 ;
        RECT 109.130 109.415 110.025 109.790 ;
        RECT 110.535 109.745 110.925 109.825 ;
        RECT 108.075 108.985 108.960 109.155 ;
        RECT 109.140 108.685 109.455 109.185 ;
        RECT 109.685 108.855 110.025 109.415 ;
        RECT 110.195 108.685 110.365 109.695 ;
        RECT 110.535 108.900 110.865 109.745 ;
        RECT 111.095 109.405 111.345 110.775 ;
        RECT 112.695 110.605 113.025 110.965 ;
        RECT 111.635 110.415 113.025 110.605 ;
        RECT 113.395 110.465 116.905 111.235 ;
        RECT 117.275 110.605 117.605 110.965 ;
        RECT 118.225 110.775 118.475 111.235 ;
        RECT 118.645 110.775 119.205 111.065 ;
        RECT 111.635 110.325 111.805 110.415 ;
        RECT 111.515 109.995 111.805 110.325 ;
        RECT 111.975 109.995 112.315 110.245 ;
        RECT 112.535 109.995 113.210 110.245 ;
        RECT 111.635 109.745 111.805 109.995 ;
        RECT 111.635 109.575 112.575 109.745 ;
        RECT 112.945 109.635 113.210 109.995 ;
        RECT 113.395 109.945 115.045 110.465 ;
        RECT 117.275 110.415 118.665 110.605 ;
        RECT 118.495 110.325 118.665 110.415 ;
        RECT 115.215 109.775 116.905 110.295 ;
        RECT 111.095 108.855 111.555 109.405 ;
        RECT 111.745 108.685 112.075 109.405 ;
        RECT 112.275 109.025 112.575 109.575 ;
        RECT 112.745 108.685 113.025 109.355 ;
        RECT 113.395 108.685 116.905 109.775 ;
        RECT 117.090 109.995 117.765 110.245 ;
        RECT 117.985 109.995 118.325 110.245 ;
        RECT 118.495 109.995 118.785 110.325 ;
        RECT 117.090 109.635 117.355 109.995 ;
        RECT 118.495 109.745 118.665 109.995 ;
        RECT 117.725 109.575 118.665 109.745 ;
        RECT 117.275 108.685 117.555 109.355 ;
        RECT 117.725 109.025 118.025 109.575 ;
        RECT 118.955 109.405 119.205 110.775 ;
        RECT 119.375 110.690 124.720 111.235 ;
        RECT 120.960 109.860 121.300 110.690 ;
        RECT 125.815 110.510 126.105 111.235 ;
        RECT 126.275 110.690 131.620 111.235 ;
        RECT 118.225 108.685 118.555 109.405 ;
        RECT 118.745 108.855 119.205 109.405 ;
        RECT 122.780 109.120 123.130 110.370 ;
        RECT 127.860 109.860 128.200 110.690 ;
        RECT 131.795 110.485 133.005 111.235 ;
        RECT 133.185 110.505 133.485 111.235 ;
        RECT 119.375 108.685 124.720 109.120 ;
        RECT 125.815 108.685 126.105 109.850 ;
        RECT 129.680 109.120 130.030 110.370 ;
        RECT 131.795 109.945 132.315 110.485 ;
        RECT 133.665 110.325 133.895 110.945 ;
        RECT 134.095 110.675 134.320 111.055 ;
        RECT 134.490 110.845 134.820 111.235 ;
        RECT 134.095 110.495 134.425 110.675 ;
        RECT 132.485 109.775 133.005 110.315 ;
        RECT 133.190 109.995 133.485 110.325 ;
        RECT 133.665 109.995 134.080 110.325 ;
        RECT 134.250 109.825 134.425 110.495 ;
        RECT 134.595 109.995 134.835 110.645 ;
        RECT 135.015 110.465 136.685 111.235 ;
        RECT 135.015 109.945 135.765 110.465 ;
        RECT 136.915 110.415 137.125 111.235 ;
        RECT 137.295 110.435 137.625 111.065 ;
        RECT 126.275 108.685 131.620 109.120 ;
        RECT 131.795 108.685 133.005 109.775 ;
        RECT 133.185 109.465 134.080 109.795 ;
        RECT 134.250 109.635 134.835 109.825 ;
        RECT 135.935 109.775 136.685 110.295 ;
        RECT 137.295 109.835 137.545 110.435 ;
        RECT 137.795 110.415 138.025 111.235 ;
        RECT 138.325 110.685 138.495 110.975 ;
        RECT 138.665 110.855 138.995 111.235 ;
        RECT 138.325 110.515 138.990 110.685 ;
        RECT 137.715 109.995 138.045 110.245 ;
        RECT 133.185 109.295 134.390 109.465 ;
        RECT 133.185 108.865 133.515 109.295 ;
        RECT 133.695 108.685 133.890 109.125 ;
        RECT 134.060 108.865 134.390 109.295 ;
        RECT 134.560 108.865 134.835 109.635 ;
        RECT 135.015 108.685 136.685 109.775 ;
        RECT 136.915 108.685 137.125 109.825 ;
        RECT 137.295 108.855 137.625 109.835 ;
        RECT 137.795 108.685 138.025 109.825 ;
        RECT 138.240 109.695 138.590 110.345 ;
        RECT 138.760 109.525 138.990 110.515 ;
        RECT 138.325 109.355 138.990 109.525 ;
        RECT 138.325 108.855 138.495 109.355 ;
        RECT 138.665 108.685 138.995 109.185 ;
        RECT 139.165 108.855 139.350 110.975 ;
        RECT 139.605 110.775 139.855 111.235 ;
        RECT 140.025 110.785 140.360 110.955 ;
        RECT 140.555 110.785 141.230 110.955 ;
        RECT 140.025 110.645 140.195 110.785 ;
        RECT 139.520 109.655 139.800 110.605 ;
        RECT 139.970 110.515 140.195 110.645 ;
        RECT 139.970 109.410 140.140 110.515 ;
        RECT 140.365 110.365 140.890 110.585 ;
        RECT 140.310 109.600 140.550 110.195 ;
        RECT 140.720 109.665 140.890 110.365 ;
        RECT 141.060 110.005 141.230 110.785 ;
        RECT 141.550 110.735 141.920 111.235 ;
        RECT 142.100 110.785 142.505 110.955 ;
        RECT 142.675 110.785 143.460 110.955 ;
        RECT 142.100 110.555 142.270 110.785 ;
        RECT 141.440 110.255 142.270 110.555 ;
        RECT 142.655 110.285 143.120 110.615 ;
        RECT 141.440 110.225 141.640 110.255 ;
        RECT 141.760 110.005 141.930 110.075 ;
        RECT 141.060 109.835 141.930 110.005 ;
        RECT 141.420 109.745 141.930 109.835 ;
        RECT 139.970 109.280 140.275 109.410 ;
        RECT 140.720 109.300 141.250 109.665 ;
        RECT 139.590 108.685 139.855 109.145 ;
        RECT 140.025 108.855 140.275 109.280 ;
        RECT 141.420 109.130 141.590 109.745 ;
        RECT 140.485 108.960 141.590 109.130 ;
        RECT 141.760 108.685 141.930 109.485 ;
        RECT 142.100 109.185 142.270 110.255 ;
        RECT 142.440 109.355 142.630 110.075 ;
        RECT 142.800 109.325 143.120 110.285 ;
        RECT 143.290 110.325 143.460 110.785 ;
        RECT 143.735 110.705 143.945 111.235 ;
        RECT 144.205 110.495 144.535 111.020 ;
        RECT 144.705 110.625 144.875 111.235 ;
        RECT 145.045 110.580 145.375 111.015 ;
        RECT 145.710 110.605 145.995 111.065 ;
        RECT 146.165 110.775 146.435 111.235 ;
        RECT 145.045 110.495 145.425 110.580 ;
        RECT 144.335 110.325 144.535 110.495 ;
        RECT 145.200 110.455 145.425 110.495 ;
        RECT 143.290 109.995 144.165 110.325 ;
        RECT 144.335 109.995 145.085 110.325 ;
        RECT 142.100 108.855 142.350 109.185 ;
        RECT 143.290 109.155 143.460 109.995 ;
        RECT 144.335 109.790 144.525 109.995 ;
        RECT 145.255 109.875 145.425 110.455 ;
        RECT 145.710 110.435 146.665 110.605 ;
        RECT 145.210 109.825 145.425 109.875 ;
        RECT 143.630 109.415 144.525 109.790 ;
        RECT 145.035 109.745 145.425 109.825 ;
        RECT 142.575 108.985 143.460 109.155 ;
        RECT 143.640 108.685 143.955 109.185 ;
        RECT 144.185 108.855 144.525 109.415 ;
        RECT 144.695 108.685 144.865 109.695 ;
        RECT 145.035 108.900 145.365 109.745 ;
        RECT 145.595 109.705 146.285 110.265 ;
        RECT 146.455 109.535 146.665 110.435 ;
        RECT 145.710 109.315 146.665 109.535 ;
        RECT 146.835 110.265 147.235 111.065 ;
        RECT 147.425 110.605 147.705 111.065 ;
        RECT 148.225 110.775 148.550 111.235 ;
        RECT 147.425 110.435 148.550 110.605 ;
        RECT 148.720 110.495 149.105 111.065 ;
        RECT 148.100 110.325 148.550 110.435 ;
        RECT 146.835 109.705 147.930 110.265 ;
        RECT 148.100 109.995 148.655 110.325 ;
        RECT 145.710 108.855 145.995 109.315 ;
        RECT 146.165 108.685 146.435 109.145 ;
        RECT 146.835 108.855 147.235 109.705 ;
        RECT 148.100 109.535 148.550 109.995 ;
        RECT 148.825 109.825 149.105 110.495 ;
        RECT 149.315 110.415 149.545 111.235 ;
        RECT 149.715 110.435 150.045 111.065 ;
        RECT 149.295 109.995 149.625 110.245 ;
        RECT 149.795 109.835 150.045 110.435 ;
        RECT 150.215 110.415 150.425 111.235 ;
        RECT 151.575 110.510 151.865 111.235 ;
        RECT 152.035 110.465 155.545 111.235 ;
        RECT 155.715 110.485 156.925 111.235 ;
        RECT 152.035 109.945 153.685 110.465 ;
        RECT 147.425 109.315 148.550 109.535 ;
        RECT 147.425 108.855 147.705 109.315 ;
        RECT 148.225 108.685 148.550 109.145 ;
        RECT 148.720 108.855 149.105 109.825 ;
        RECT 149.315 108.685 149.545 109.825 ;
        RECT 149.715 108.855 150.045 109.835 ;
        RECT 150.215 108.685 150.425 109.825 ;
        RECT 151.575 108.685 151.865 109.850 ;
        RECT 153.855 109.775 155.545 110.295 ;
        RECT 152.035 108.685 155.545 109.775 ;
        RECT 155.715 109.775 156.235 110.315 ;
        RECT 156.405 109.945 156.925 110.485 ;
        RECT 155.715 108.685 156.925 109.775 ;
        RECT 22.690 108.515 157.010 108.685 ;
        RECT 22.775 107.425 23.985 108.515 ;
        RECT 22.775 106.715 23.295 107.255 ;
        RECT 23.465 106.885 23.985 107.425 ;
        RECT 25.260 107.545 25.650 107.720 ;
        RECT 26.135 107.715 26.465 108.515 ;
        RECT 26.635 107.725 27.170 108.345 ;
        RECT 25.260 107.375 26.685 107.545 ;
        RECT 22.775 105.965 23.985 106.715 ;
        RECT 25.135 106.645 25.490 107.205 ;
        RECT 25.660 106.475 25.830 107.375 ;
        RECT 26.000 106.645 26.265 107.205 ;
        RECT 26.515 106.875 26.685 107.375 ;
        RECT 26.855 106.705 27.170 107.725 ;
        RECT 25.240 105.965 25.480 106.475 ;
        RECT 25.660 106.145 25.940 106.475 ;
        RECT 26.170 105.965 26.385 106.475 ;
        RECT 26.555 106.135 27.170 106.705 ;
        RECT 27.375 107.375 27.760 108.345 ;
        RECT 27.930 108.055 28.255 108.515 ;
        RECT 28.775 107.885 29.055 108.345 ;
        RECT 27.930 107.665 29.055 107.885 ;
        RECT 27.375 106.705 27.655 107.375 ;
        RECT 27.930 107.205 28.380 107.665 ;
        RECT 29.245 107.495 29.645 108.345 ;
        RECT 30.045 108.055 30.315 108.515 ;
        RECT 30.485 107.885 30.770 108.345 ;
        RECT 27.825 106.875 28.380 107.205 ;
        RECT 28.550 106.935 29.645 107.495 ;
        RECT 27.930 106.765 28.380 106.875 ;
        RECT 27.375 106.135 27.760 106.705 ;
        RECT 27.930 106.595 29.055 106.765 ;
        RECT 27.930 105.965 28.255 106.425 ;
        RECT 28.775 106.135 29.055 106.595 ;
        RECT 29.245 106.135 29.645 106.935 ;
        RECT 29.815 107.665 30.770 107.885 ;
        RECT 29.815 106.765 30.025 107.665 ;
        RECT 30.195 106.935 30.885 107.495 ;
        RECT 31.975 107.375 32.360 108.345 ;
        RECT 32.530 108.055 32.855 108.515 ;
        RECT 33.375 107.885 33.655 108.345 ;
        RECT 32.530 107.665 33.655 107.885 ;
        RECT 29.815 106.595 30.770 106.765 ;
        RECT 30.045 105.965 30.315 106.425 ;
        RECT 30.485 106.135 30.770 106.595 ;
        RECT 31.975 106.705 32.255 107.375 ;
        RECT 32.530 107.205 32.980 107.665 ;
        RECT 33.845 107.495 34.245 108.345 ;
        RECT 34.645 108.055 34.915 108.515 ;
        RECT 35.085 107.885 35.370 108.345 ;
        RECT 32.425 106.875 32.980 107.205 ;
        RECT 33.150 106.935 34.245 107.495 ;
        RECT 32.530 106.765 32.980 106.875 ;
        RECT 31.975 106.135 32.360 106.705 ;
        RECT 32.530 106.595 33.655 106.765 ;
        RECT 32.530 105.965 32.855 106.425 ;
        RECT 33.375 106.135 33.655 106.595 ;
        RECT 33.845 106.135 34.245 106.935 ;
        RECT 34.415 107.665 35.370 107.885 ;
        RECT 34.415 106.765 34.625 107.665 ;
        RECT 34.795 106.935 35.485 107.495 ;
        RECT 35.655 107.350 35.945 108.515 ;
        RECT 37.240 107.545 37.570 108.345 ;
        RECT 37.740 107.715 38.070 108.515 ;
        RECT 38.370 107.545 38.700 108.345 ;
        RECT 39.345 107.715 39.595 108.515 ;
        RECT 37.240 107.375 39.675 107.545 ;
        RECT 39.865 107.375 40.035 108.515 ;
        RECT 40.205 107.375 40.545 108.345 ;
        RECT 40.830 107.885 41.115 108.345 ;
        RECT 41.285 108.055 41.555 108.515 ;
        RECT 40.830 107.665 41.785 107.885 ;
        RECT 37.035 106.955 37.385 107.205 ;
        RECT 34.415 106.595 35.370 106.765 ;
        RECT 37.570 106.745 37.740 107.375 ;
        RECT 37.910 106.955 38.240 107.155 ;
        RECT 38.410 106.955 38.740 107.155 ;
        RECT 38.910 106.955 39.330 107.155 ;
        RECT 39.505 107.125 39.675 107.375 ;
        RECT 39.505 106.955 40.200 107.125 ;
        RECT 34.645 105.965 34.915 106.425 ;
        RECT 35.085 106.135 35.370 106.595 ;
        RECT 35.655 105.965 35.945 106.690 ;
        RECT 37.240 106.135 37.740 106.745 ;
        RECT 38.370 106.615 39.595 106.785 ;
        RECT 40.370 106.765 40.545 107.375 ;
        RECT 40.715 106.935 41.405 107.495 ;
        RECT 41.575 106.765 41.785 107.665 ;
        RECT 38.370 106.135 38.700 106.615 ;
        RECT 38.870 105.965 39.095 106.425 ;
        RECT 39.265 106.135 39.595 106.615 ;
        RECT 39.785 105.965 40.035 106.765 ;
        RECT 40.205 106.135 40.545 106.765 ;
        RECT 40.830 106.595 41.785 106.765 ;
        RECT 41.955 107.495 42.355 108.345 ;
        RECT 42.545 107.885 42.825 108.345 ;
        RECT 43.345 108.055 43.670 108.515 ;
        RECT 42.545 107.665 43.670 107.885 ;
        RECT 41.955 106.935 43.050 107.495 ;
        RECT 43.220 107.205 43.670 107.665 ;
        RECT 43.840 107.375 44.225 108.345 ;
        RECT 40.830 106.135 41.115 106.595 ;
        RECT 41.285 105.965 41.555 106.425 ;
        RECT 41.955 106.135 42.355 106.935 ;
        RECT 43.220 106.875 43.775 107.205 ;
        RECT 43.220 106.765 43.670 106.875 ;
        RECT 42.545 106.595 43.670 106.765 ;
        RECT 43.945 106.705 44.225 107.375 ;
        RECT 42.545 106.135 42.825 106.595 ;
        RECT 43.345 105.965 43.670 106.425 ;
        RECT 43.840 106.135 44.225 106.705 ;
        RECT 44.395 107.375 44.735 108.345 ;
        RECT 44.905 107.375 45.075 108.515 ;
        RECT 45.345 107.715 45.595 108.515 ;
        RECT 46.240 107.545 46.570 108.345 ;
        RECT 46.870 107.715 47.200 108.515 ;
        RECT 47.370 107.545 47.700 108.345 ;
        RECT 48.190 107.885 48.475 108.345 ;
        RECT 48.645 108.055 48.915 108.515 ;
        RECT 48.190 107.665 49.145 107.885 ;
        RECT 45.265 107.375 47.700 107.545 ;
        RECT 44.395 107.325 44.625 107.375 ;
        RECT 44.395 106.765 44.570 107.325 ;
        RECT 45.265 107.125 45.435 107.375 ;
        RECT 44.740 106.955 45.435 107.125 ;
        RECT 45.610 106.955 46.030 107.155 ;
        RECT 46.200 106.955 46.530 107.155 ;
        RECT 46.700 106.955 47.030 107.155 ;
        RECT 44.395 106.135 44.735 106.765 ;
        RECT 44.905 105.965 45.155 106.765 ;
        RECT 45.345 106.615 46.570 106.785 ;
        RECT 45.345 106.135 45.675 106.615 ;
        RECT 45.845 105.965 46.070 106.425 ;
        RECT 46.240 106.135 46.570 106.615 ;
        RECT 47.200 106.745 47.370 107.375 ;
        RECT 47.555 106.955 47.905 107.205 ;
        RECT 48.075 106.935 48.765 107.495 ;
        RECT 48.935 106.765 49.145 107.665 ;
        RECT 47.200 106.135 47.700 106.745 ;
        RECT 48.190 106.595 49.145 106.765 ;
        RECT 49.315 107.495 49.715 108.345 ;
        RECT 49.905 107.885 50.185 108.345 ;
        RECT 50.705 108.055 51.030 108.515 ;
        RECT 49.905 107.665 51.030 107.885 ;
        RECT 49.315 106.935 50.410 107.495 ;
        RECT 50.580 107.205 51.030 107.665 ;
        RECT 51.200 107.375 51.585 108.345 ;
        RECT 48.190 106.135 48.475 106.595 ;
        RECT 48.645 105.965 48.915 106.425 ;
        RECT 49.315 106.135 49.715 106.935 ;
        RECT 50.580 106.875 51.135 107.205 ;
        RECT 50.580 106.765 51.030 106.875 ;
        RECT 49.905 106.595 51.030 106.765 ;
        RECT 51.305 106.705 51.585 107.375 ;
        RECT 49.905 106.135 50.185 106.595 ;
        RECT 50.705 105.965 51.030 106.425 ;
        RECT 51.200 106.135 51.585 106.705 ;
        RECT 51.755 107.375 52.095 108.345 ;
        RECT 52.265 107.375 52.435 108.515 ;
        RECT 52.705 107.715 52.955 108.515 ;
        RECT 53.600 107.545 53.930 108.345 ;
        RECT 54.230 107.715 54.560 108.515 ;
        RECT 54.730 107.545 55.060 108.345 ;
        RECT 52.625 107.375 55.060 107.545 ;
        RECT 55.470 107.725 56.005 108.345 ;
        RECT 51.755 106.765 51.930 107.375 ;
        RECT 52.625 107.125 52.795 107.375 ;
        RECT 52.100 106.955 52.795 107.125 ;
        RECT 52.970 106.955 53.390 107.155 ;
        RECT 53.560 106.955 53.890 107.155 ;
        RECT 54.060 106.955 54.390 107.155 ;
        RECT 51.755 106.135 52.095 106.765 ;
        RECT 52.265 105.965 52.515 106.765 ;
        RECT 52.705 106.615 53.930 106.785 ;
        RECT 52.705 106.135 53.035 106.615 ;
        RECT 53.205 105.965 53.430 106.425 ;
        RECT 53.600 106.135 53.930 106.615 ;
        RECT 54.560 106.745 54.730 107.375 ;
        RECT 54.915 106.955 55.265 107.205 ;
        RECT 54.560 106.135 55.060 106.745 ;
        RECT 55.470 106.705 55.785 107.725 ;
        RECT 56.175 107.715 56.505 108.515 ;
        RECT 56.990 107.545 57.380 107.720 ;
        RECT 55.955 107.375 57.380 107.545 ;
        RECT 57.920 107.545 58.310 107.720 ;
        RECT 58.795 107.715 59.125 108.515 ;
        RECT 59.295 107.725 59.830 108.345 ;
        RECT 57.920 107.375 59.345 107.545 ;
        RECT 55.955 106.875 56.125 107.375 ;
        RECT 55.470 106.135 56.085 106.705 ;
        RECT 56.375 106.645 56.640 107.205 ;
        RECT 56.810 106.475 56.980 107.375 ;
        RECT 57.150 106.645 57.505 107.205 ;
        RECT 57.795 106.645 58.150 107.205 ;
        RECT 58.320 106.475 58.490 107.375 ;
        RECT 58.660 106.645 58.925 107.205 ;
        RECT 59.175 106.875 59.345 107.375 ;
        RECT 59.515 106.705 59.830 107.725 ;
        RECT 56.255 105.965 56.470 106.475 ;
        RECT 56.700 106.145 56.980 106.475 ;
        RECT 57.160 105.965 57.400 106.475 ;
        RECT 57.900 105.965 58.140 106.475 ;
        RECT 58.320 106.145 58.600 106.475 ;
        RECT 58.830 105.965 59.045 106.475 ;
        RECT 59.215 106.135 59.830 106.705 ;
        RECT 60.035 107.440 60.305 108.345 ;
        RECT 60.475 107.755 60.805 108.515 ;
        RECT 60.985 107.585 61.155 108.345 ;
        RECT 60.035 106.640 60.205 107.440 ;
        RECT 60.490 107.415 61.155 107.585 ;
        RECT 60.490 107.270 60.660 107.415 ;
        RECT 61.415 107.350 61.705 108.515 ;
        RECT 61.875 107.425 65.385 108.515 ;
        RECT 66.020 107.715 66.275 108.515 ;
        RECT 66.475 107.665 66.805 108.345 ;
        RECT 60.375 106.940 60.660 107.270 ;
        RECT 60.490 106.685 60.660 106.940 ;
        RECT 60.895 106.865 61.225 107.235 ;
        RECT 61.875 106.735 63.525 107.255 ;
        RECT 63.695 106.905 65.385 107.425 ;
        RECT 66.020 107.175 66.265 107.535 ;
        RECT 66.455 107.385 66.805 107.665 ;
        RECT 66.455 107.005 66.625 107.385 ;
        RECT 66.985 107.205 67.180 108.255 ;
        RECT 67.360 107.375 67.680 108.515 ;
        RECT 67.855 107.375 68.240 108.345 ;
        RECT 68.410 108.055 68.735 108.515 ;
        RECT 69.255 107.885 69.535 108.345 ;
        RECT 68.410 107.665 69.535 107.885 ;
        RECT 66.105 106.835 66.625 107.005 ;
        RECT 66.795 106.875 67.180 107.205 ;
        RECT 67.360 107.155 67.620 107.205 ;
        RECT 67.360 106.985 67.625 107.155 ;
        RECT 67.360 106.875 67.620 106.985 ;
        RECT 66.105 106.815 66.275 106.835 ;
        RECT 60.035 106.135 60.295 106.640 ;
        RECT 60.490 106.515 61.155 106.685 ;
        RECT 60.475 105.965 60.805 106.345 ;
        RECT 60.985 106.135 61.155 106.515 ;
        RECT 61.415 105.965 61.705 106.690 ;
        RECT 61.875 105.965 65.385 106.735 ;
        RECT 66.075 106.645 66.275 106.815 ;
        RECT 67.855 106.705 68.135 107.375 ;
        RECT 68.410 107.205 68.860 107.665 ;
        RECT 69.725 107.495 70.125 108.345 ;
        RECT 70.525 108.055 70.795 108.515 ;
        RECT 70.965 107.885 71.250 108.345 ;
        RECT 68.305 106.875 68.860 107.205 ;
        RECT 69.030 106.935 70.125 107.495 ;
        RECT 68.410 106.765 68.860 106.875 ;
        RECT 66.105 106.270 66.275 106.645 ;
        RECT 66.465 106.495 67.680 106.665 ;
        RECT 66.465 106.190 66.695 106.495 ;
        RECT 66.865 105.965 67.195 106.325 ;
        RECT 67.390 106.145 67.680 106.495 ;
        RECT 67.855 106.135 68.240 106.705 ;
        RECT 68.410 106.595 69.535 106.765 ;
        RECT 68.410 105.965 68.735 106.425 ;
        RECT 69.255 106.135 69.535 106.595 ;
        RECT 69.725 106.135 70.125 106.935 ;
        RECT 70.295 107.665 71.250 107.885 ;
        RECT 71.650 107.885 71.935 108.345 ;
        RECT 72.105 108.055 72.375 108.515 ;
        RECT 71.650 107.665 72.605 107.885 ;
        RECT 70.295 106.765 70.505 107.665 ;
        RECT 70.675 106.935 71.365 107.495 ;
        RECT 71.535 106.935 72.225 107.495 ;
        RECT 72.395 106.765 72.605 107.665 ;
        RECT 70.295 106.595 71.250 106.765 ;
        RECT 70.525 105.965 70.795 106.425 ;
        RECT 70.965 106.135 71.250 106.595 ;
        RECT 71.650 106.595 72.605 106.765 ;
        RECT 72.775 107.495 73.175 108.345 ;
        RECT 73.365 107.885 73.645 108.345 ;
        RECT 74.165 108.055 74.490 108.515 ;
        RECT 73.365 107.665 74.490 107.885 ;
        RECT 72.775 106.935 73.870 107.495 ;
        RECT 74.040 107.205 74.490 107.665 ;
        RECT 74.660 107.375 75.045 108.345 ;
        RECT 75.215 107.425 78.725 108.515 ;
        RECT 71.650 106.135 71.935 106.595 ;
        RECT 72.105 105.965 72.375 106.425 ;
        RECT 72.775 106.135 73.175 106.935 ;
        RECT 74.040 106.875 74.595 107.205 ;
        RECT 74.040 106.765 74.490 106.875 ;
        RECT 73.365 106.595 74.490 106.765 ;
        RECT 74.765 106.705 75.045 107.375 ;
        RECT 73.365 106.135 73.645 106.595 ;
        RECT 74.165 105.965 74.490 106.425 ;
        RECT 74.660 106.135 75.045 106.705 ;
        RECT 75.215 106.735 76.865 107.255 ;
        RECT 77.035 106.905 78.725 107.425 ;
        RECT 79.360 107.370 79.655 108.515 ;
        RECT 75.215 105.965 78.725 106.735 ;
        RECT 79.360 105.965 79.655 106.785 ;
        RECT 79.825 106.515 80.055 108.215 ;
        RECT 80.270 107.710 80.525 108.515 ;
        RECT 80.725 107.900 81.055 108.345 ;
        RECT 81.225 108.070 81.500 108.515 ;
        RECT 81.735 107.900 82.065 108.345 ;
        RECT 80.725 107.720 82.065 107.900 ;
        RECT 82.525 107.540 82.855 108.205 ;
        RECT 80.270 107.370 82.855 107.540 ;
        RECT 83.035 107.425 85.625 108.515 ;
        RECT 80.270 106.755 80.580 107.370 ;
        RECT 80.750 106.925 81.080 107.155 ;
        RECT 81.250 106.925 81.720 107.155 ;
        RECT 81.890 106.985 82.345 107.155 ;
        RECT 81.890 106.925 82.340 106.985 ;
        RECT 82.530 106.925 82.865 107.155 ;
        RECT 80.270 106.575 82.855 106.755 ;
        RECT 79.825 106.135 80.045 106.515 ;
        RECT 80.215 105.965 81.065 106.325 ;
        RECT 81.545 106.155 81.875 106.575 ;
        RECT 82.080 105.965 82.355 106.405 ;
        RECT 82.525 106.155 82.855 106.575 ;
        RECT 83.035 106.735 84.245 107.255 ;
        RECT 84.415 106.905 85.625 107.425 ;
        RECT 85.805 107.375 86.135 108.515 ;
        RECT 86.665 107.545 86.995 108.330 ;
        RECT 86.315 107.375 86.995 107.545 ;
        RECT 85.795 106.955 86.145 107.205 ;
        RECT 86.315 106.775 86.485 107.375 ;
        RECT 87.175 107.350 87.465 108.515 ;
        RECT 87.635 108.080 92.980 108.515 ;
        RECT 86.655 106.955 87.005 107.205 ;
        RECT 83.035 105.965 85.625 106.735 ;
        RECT 85.805 105.965 86.075 106.775 ;
        RECT 86.245 106.135 86.575 106.775 ;
        RECT 86.745 105.965 86.985 106.775 ;
        RECT 87.175 105.965 87.465 106.690 ;
        RECT 89.220 106.510 89.560 107.340 ;
        RECT 91.040 106.830 91.390 108.080 ;
        RECT 93.615 107.440 93.885 108.345 ;
        RECT 94.055 107.755 94.385 108.515 ;
        RECT 94.565 107.585 94.735 108.345 ;
        RECT 93.615 106.640 93.785 107.440 ;
        RECT 94.070 107.415 94.735 107.585 ;
        RECT 95.915 107.795 96.375 108.345 ;
        RECT 96.565 107.795 96.895 108.515 ;
        RECT 94.070 107.270 94.240 107.415 ;
        RECT 93.955 106.940 94.240 107.270 ;
        RECT 94.070 106.685 94.240 106.940 ;
        RECT 94.475 106.865 94.805 107.235 ;
        RECT 87.635 105.965 92.980 106.510 ;
        RECT 93.615 106.135 93.875 106.640 ;
        RECT 94.070 106.515 94.735 106.685 ;
        RECT 94.055 105.965 94.385 106.345 ;
        RECT 94.565 106.135 94.735 106.515 ;
        RECT 95.915 106.425 96.165 107.795 ;
        RECT 97.095 107.625 97.395 108.175 ;
        RECT 97.565 107.845 97.845 108.515 ;
        RECT 96.455 107.455 97.395 107.625 ;
        RECT 96.455 107.205 96.625 107.455 ;
        RECT 97.765 107.205 98.030 107.565 ;
        RECT 98.215 107.425 99.885 108.515 ;
        RECT 96.335 106.875 96.625 107.205 ;
        RECT 96.795 106.955 97.135 107.205 ;
        RECT 97.355 106.955 98.030 107.205 ;
        RECT 96.455 106.785 96.625 106.875 ;
        RECT 96.455 106.595 97.845 106.785 ;
        RECT 95.915 106.135 96.475 106.425 ;
        RECT 96.645 105.965 96.895 106.425 ;
        RECT 97.515 106.235 97.845 106.595 ;
        RECT 98.215 106.735 98.965 107.255 ;
        RECT 99.135 106.905 99.885 107.425 ;
        RECT 100.145 107.585 100.315 108.345 ;
        RECT 100.495 107.755 100.825 108.515 ;
        RECT 100.145 107.415 100.810 107.585 ;
        RECT 100.995 107.440 101.265 108.345 ;
        RECT 101.435 108.080 106.780 108.515 ;
        RECT 106.955 108.080 112.300 108.515 ;
        RECT 100.640 107.270 100.810 107.415 ;
        RECT 100.075 106.865 100.405 107.235 ;
        RECT 100.640 106.940 100.925 107.270 ;
        RECT 98.215 105.965 99.885 106.735 ;
        RECT 100.640 106.685 100.810 106.940 ;
        RECT 100.145 106.515 100.810 106.685 ;
        RECT 101.095 106.640 101.265 107.440 ;
        RECT 100.145 106.135 100.315 106.515 ;
        RECT 100.495 105.965 100.825 106.345 ;
        RECT 101.005 106.135 101.265 106.640 ;
        RECT 103.020 106.510 103.360 107.340 ;
        RECT 104.840 106.830 105.190 108.080 ;
        RECT 108.540 106.510 108.880 107.340 ;
        RECT 110.360 106.830 110.710 108.080 ;
        RECT 112.935 107.350 113.225 108.515 ;
        RECT 113.405 107.545 113.735 108.330 ;
        RECT 113.405 107.375 114.085 107.545 ;
        RECT 114.265 107.375 114.595 108.515 ;
        RECT 114.785 107.375 115.115 108.515 ;
        RECT 115.645 107.545 115.975 108.330 ;
        RECT 115.295 107.375 115.975 107.545 ;
        RECT 116.155 107.425 117.365 108.515 ;
        RECT 117.735 107.845 118.015 108.515 ;
        RECT 118.185 107.625 118.485 108.175 ;
        RECT 118.685 107.795 119.015 108.515 ;
        RECT 119.205 107.795 119.665 108.345 ;
        RECT 113.395 106.955 113.745 107.205 ;
        RECT 113.915 106.775 114.085 107.375 ;
        RECT 114.255 106.955 114.605 107.205 ;
        RECT 114.775 106.955 115.125 107.205 ;
        RECT 115.295 106.775 115.465 107.375 ;
        RECT 115.635 106.955 115.985 107.205 ;
        RECT 101.435 105.965 106.780 106.510 ;
        RECT 106.955 105.965 112.300 106.510 ;
        RECT 112.935 105.965 113.225 106.690 ;
        RECT 113.415 105.965 113.655 106.775 ;
        RECT 113.825 106.135 114.155 106.775 ;
        RECT 114.325 105.965 114.595 106.775 ;
        RECT 114.785 105.965 115.055 106.775 ;
        RECT 115.225 106.135 115.555 106.775 ;
        RECT 115.725 105.965 115.965 106.775 ;
        RECT 116.155 106.715 116.675 107.255 ;
        RECT 116.845 106.885 117.365 107.425 ;
        RECT 117.550 107.205 117.815 107.565 ;
        RECT 118.185 107.455 119.125 107.625 ;
        RECT 118.955 107.205 119.125 107.455 ;
        RECT 117.550 106.955 118.225 107.205 ;
        RECT 118.445 106.955 118.785 107.205 ;
        RECT 118.955 106.875 119.245 107.205 ;
        RECT 118.955 106.785 119.125 106.875 ;
        RECT 116.155 105.965 117.365 106.715 ;
        RECT 117.735 106.595 119.125 106.785 ;
        RECT 117.735 106.235 118.065 106.595 ;
        RECT 119.415 106.425 119.665 107.795 ;
        RECT 119.835 107.425 121.505 108.515 ;
        RECT 118.685 105.965 118.935 106.425 ;
        RECT 119.105 106.135 119.665 106.425 ;
        RECT 119.835 106.735 120.585 107.255 ;
        RECT 120.755 106.905 121.505 107.425 ;
        RECT 121.675 107.375 122.015 108.345 ;
        RECT 122.185 107.375 122.355 108.515 ;
        RECT 122.625 107.715 122.875 108.515 ;
        RECT 123.520 107.545 123.850 108.345 ;
        RECT 124.150 107.715 124.480 108.515 ;
        RECT 124.650 107.545 124.980 108.345 ;
        RECT 122.545 107.375 124.980 107.545 ;
        RECT 125.355 107.375 125.740 108.345 ;
        RECT 125.910 108.055 126.235 108.515 ;
        RECT 126.755 107.885 127.035 108.345 ;
        RECT 125.910 107.665 127.035 107.885 ;
        RECT 121.675 106.815 121.850 107.375 ;
        RECT 122.545 107.125 122.715 107.375 ;
        RECT 122.020 106.955 122.715 107.125 ;
        RECT 122.890 106.955 123.310 107.155 ;
        RECT 123.480 106.955 123.810 107.155 ;
        RECT 123.980 106.955 124.310 107.155 ;
        RECT 121.675 106.765 121.905 106.815 ;
        RECT 119.835 105.965 121.505 106.735 ;
        RECT 121.675 106.135 122.015 106.765 ;
        RECT 122.185 105.965 122.435 106.765 ;
        RECT 122.625 106.615 123.850 106.785 ;
        RECT 122.625 106.135 122.955 106.615 ;
        RECT 123.125 105.965 123.350 106.425 ;
        RECT 123.520 106.135 123.850 106.615 ;
        RECT 124.480 106.745 124.650 107.375 ;
        RECT 124.835 106.955 125.185 107.205 ;
        RECT 124.480 106.135 124.980 106.745 ;
        RECT 125.355 106.705 125.635 107.375 ;
        RECT 125.910 107.205 126.360 107.665 ;
        RECT 127.225 107.495 127.625 108.345 ;
        RECT 128.025 108.055 128.295 108.515 ;
        RECT 128.465 107.885 128.750 108.345 ;
        RECT 125.805 106.875 126.360 107.205 ;
        RECT 126.530 106.935 127.625 107.495 ;
        RECT 125.910 106.765 126.360 106.875 ;
        RECT 125.355 106.135 125.740 106.705 ;
        RECT 125.910 106.595 127.035 106.765 ;
        RECT 125.910 105.965 126.235 106.425 ;
        RECT 126.755 106.135 127.035 106.595 ;
        RECT 127.225 106.135 127.625 106.935 ;
        RECT 127.795 107.665 128.750 107.885 ;
        RECT 127.795 106.765 128.005 107.665 ;
        RECT 129.125 107.605 129.295 108.335 ;
        RECT 129.475 107.785 129.805 108.515 ;
        RECT 129.975 107.605 130.165 108.335 ;
        RECT 128.175 106.935 128.865 107.495 ;
        RECT 129.125 107.405 130.165 107.605 ;
        RECT 130.335 107.225 130.665 108.335 ;
        RECT 130.855 108.105 131.185 108.515 ;
        RECT 131.355 107.925 131.615 108.315 ;
        RECT 131.795 108.080 137.140 108.515 ;
        RECT 129.070 106.875 129.360 107.225 ;
        RECT 129.555 106.875 129.950 107.225 ;
        RECT 130.130 106.925 130.665 107.225 ;
        RECT 130.855 107.725 131.615 107.925 ;
        RECT 130.855 107.045 131.195 107.725 ;
        RECT 127.795 106.595 128.750 106.765 ;
        RECT 128.025 105.965 128.295 106.425 ;
        RECT 128.465 106.135 128.750 106.595 ;
        RECT 129.055 105.965 129.385 106.695 ;
        RECT 129.555 106.255 129.765 106.875 ;
        RECT 130.130 106.675 130.375 106.925 ;
        RECT 129.945 106.145 130.375 106.675 ;
        RECT 130.555 105.965 130.785 106.745 ;
        RECT 130.965 106.595 131.195 107.045 ;
        RECT 131.375 106.855 131.605 107.545 ;
        RECT 130.965 106.145 131.345 106.595 ;
        RECT 133.380 106.510 133.720 107.340 ;
        RECT 135.200 106.830 135.550 108.080 ;
        RECT 137.315 107.425 138.525 108.515 ;
        RECT 137.315 106.715 137.835 107.255 ;
        RECT 138.005 106.885 138.525 107.425 ;
        RECT 138.695 107.350 138.985 108.515 ;
        RECT 139.155 107.425 142.665 108.515 ;
        RECT 142.835 107.425 144.045 108.515 ;
        RECT 139.155 106.735 140.805 107.255 ;
        RECT 140.975 106.905 142.665 107.425 ;
        RECT 131.795 105.965 137.140 106.510 ;
        RECT 137.315 105.965 138.525 106.715 ;
        RECT 138.695 105.965 138.985 106.690 ;
        RECT 139.155 105.965 142.665 106.735 ;
        RECT 142.835 106.715 143.355 107.255 ;
        RECT 143.525 106.885 144.045 107.425 ;
        RECT 144.215 107.375 144.475 108.515 ;
        RECT 144.645 107.365 144.975 108.345 ;
        RECT 145.145 107.375 145.425 108.515 ;
        RECT 145.595 108.080 150.940 108.515 ;
        RECT 144.235 106.955 144.570 107.205 ;
        RECT 144.740 106.765 144.910 107.365 ;
        RECT 145.080 106.935 145.415 107.205 ;
        RECT 142.835 105.965 144.045 106.715 ;
        RECT 144.215 106.135 144.910 106.765 ;
        RECT 145.115 105.965 145.425 106.765 ;
        RECT 147.180 106.510 147.520 107.340 ;
        RECT 149.000 106.830 149.350 108.080 ;
        RECT 151.115 107.425 154.625 108.515 ;
        RECT 151.115 106.735 152.765 107.255 ;
        RECT 152.935 106.905 154.625 107.425 ;
        RECT 155.715 107.425 156.925 108.515 ;
        RECT 155.715 106.885 156.235 107.425 ;
        RECT 145.595 105.965 150.940 106.510 ;
        RECT 151.115 105.965 154.625 106.735 ;
        RECT 156.405 106.715 156.925 107.255 ;
        RECT 155.715 105.965 156.925 106.715 ;
        RECT 22.690 105.795 157.010 105.965 ;
        RECT 22.775 105.045 23.985 105.795 ;
        RECT 22.775 104.505 23.295 105.045 ;
        RECT 24.155 105.025 25.825 105.795 ;
        RECT 23.465 104.335 23.985 104.875 ;
        RECT 24.155 104.505 24.905 105.025 ;
        RECT 26.200 105.015 26.700 105.625 ;
        RECT 25.075 104.335 25.825 104.855 ;
        RECT 25.995 104.555 26.345 104.805 ;
        RECT 26.530 104.385 26.700 105.015 ;
        RECT 27.330 105.145 27.660 105.625 ;
        RECT 27.830 105.335 28.055 105.795 ;
        RECT 28.225 105.145 28.555 105.625 ;
        RECT 27.330 104.975 28.555 105.145 ;
        RECT 28.745 104.995 28.995 105.795 ;
        RECT 29.165 104.995 29.505 105.625 ;
        RECT 30.685 105.245 30.855 105.535 ;
        RECT 31.025 105.415 31.355 105.795 ;
        RECT 30.685 105.075 31.350 105.245 ;
        RECT 26.870 104.605 27.200 104.805 ;
        RECT 27.370 104.605 27.700 104.805 ;
        RECT 27.870 104.605 28.290 104.805 ;
        RECT 28.465 104.635 29.160 104.805 ;
        RECT 28.465 104.385 28.635 104.635 ;
        RECT 29.330 104.385 29.505 104.995 ;
        RECT 22.775 103.245 23.985 104.335 ;
        RECT 24.155 103.245 25.825 104.335 ;
        RECT 26.200 104.215 28.635 104.385 ;
        RECT 26.200 103.415 26.530 104.215 ;
        RECT 26.700 103.245 27.030 104.045 ;
        RECT 27.330 103.415 27.660 104.215 ;
        RECT 28.305 103.245 28.555 104.045 ;
        RECT 28.825 103.245 28.995 104.385 ;
        RECT 29.165 103.415 29.505 104.385 ;
        RECT 30.600 104.255 30.950 104.905 ;
        RECT 31.120 104.085 31.350 105.075 ;
        RECT 30.685 103.915 31.350 104.085 ;
        RECT 30.685 103.415 30.855 103.915 ;
        RECT 31.025 103.245 31.355 103.745 ;
        RECT 31.525 103.415 31.710 105.535 ;
        RECT 31.965 105.335 32.215 105.795 ;
        RECT 32.385 105.345 32.720 105.515 ;
        RECT 32.915 105.345 33.590 105.515 ;
        RECT 32.385 105.205 32.555 105.345 ;
        RECT 31.880 104.215 32.160 105.165 ;
        RECT 32.330 105.075 32.555 105.205 ;
        RECT 32.330 103.970 32.500 105.075 ;
        RECT 32.725 104.925 33.250 105.145 ;
        RECT 32.670 104.160 32.910 104.755 ;
        RECT 33.080 104.225 33.250 104.925 ;
        RECT 33.420 104.565 33.590 105.345 ;
        RECT 33.910 105.295 34.280 105.795 ;
        RECT 34.460 105.345 34.865 105.515 ;
        RECT 35.035 105.345 35.820 105.515 ;
        RECT 34.460 105.115 34.630 105.345 ;
        RECT 33.800 104.815 34.630 105.115 ;
        RECT 35.015 104.845 35.480 105.175 ;
        RECT 33.800 104.785 34.000 104.815 ;
        RECT 34.120 104.565 34.290 104.635 ;
        RECT 33.420 104.395 34.290 104.565 ;
        RECT 33.780 104.305 34.290 104.395 ;
        RECT 32.330 103.840 32.635 103.970 ;
        RECT 33.080 103.860 33.610 104.225 ;
        RECT 31.950 103.245 32.215 103.705 ;
        RECT 32.385 103.415 32.635 103.840 ;
        RECT 33.780 103.690 33.950 104.305 ;
        RECT 32.845 103.520 33.950 103.690 ;
        RECT 34.120 103.245 34.290 104.045 ;
        RECT 34.460 103.745 34.630 104.815 ;
        RECT 34.800 103.915 34.990 104.635 ;
        RECT 35.160 103.885 35.480 104.845 ;
        RECT 35.650 104.885 35.820 105.345 ;
        RECT 36.095 105.265 36.305 105.795 ;
        RECT 36.565 105.055 36.895 105.580 ;
        RECT 37.065 105.185 37.235 105.795 ;
        RECT 37.405 105.140 37.735 105.575 ;
        RECT 37.955 105.285 38.260 105.795 ;
        RECT 37.405 105.055 37.785 105.140 ;
        RECT 36.695 104.885 36.895 105.055 ;
        RECT 37.560 105.015 37.785 105.055 ;
        RECT 35.650 104.555 36.525 104.885 ;
        RECT 36.695 104.555 37.445 104.885 ;
        RECT 34.460 103.415 34.710 103.745 ;
        RECT 35.650 103.715 35.820 104.555 ;
        RECT 36.695 104.350 36.885 104.555 ;
        RECT 37.615 104.435 37.785 105.015 ;
        RECT 37.955 104.555 38.270 105.115 ;
        RECT 38.440 104.805 38.690 105.615 ;
        RECT 38.860 105.270 39.120 105.795 ;
        RECT 39.300 104.805 39.550 105.615 ;
        RECT 39.720 105.235 39.980 105.795 ;
        RECT 40.150 105.145 40.410 105.600 ;
        RECT 40.580 105.315 40.840 105.795 ;
        RECT 41.010 105.145 41.270 105.600 ;
        RECT 41.440 105.315 41.700 105.795 ;
        RECT 41.870 105.145 42.130 105.600 ;
        RECT 42.300 105.315 42.545 105.795 ;
        RECT 42.715 105.145 42.990 105.600 ;
        RECT 43.160 105.315 43.405 105.795 ;
        RECT 43.575 105.145 43.835 105.600 ;
        RECT 44.015 105.315 44.265 105.795 ;
        RECT 44.435 105.145 44.695 105.600 ;
        RECT 44.875 105.315 45.125 105.795 ;
        RECT 45.295 105.145 45.555 105.600 ;
        RECT 45.735 105.315 45.995 105.795 ;
        RECT 46.165 105.145 46.425 105.600 ;
        RECT 46.595 105.315 46.895 105.795 ;
        RECT 40.150 104.975 46.895 105.145 ;
        RECT 38.440 104.555 45.560 104.805 ;
        RECT 37.570 104.385 37.785 104.435 ;
        RECT 35.990 103.975 36.885 104.350 ;
        RECT 37.395 104.305 37.785 104.385 ;
        RECT 34.935 103.545 35.820 103.715 ;
        RECT 36.000 103.245 36.315 103.745 ;
        RECT 36.545 103.415 36.885 103.975 ;
        RECT 37.055 103.245 37.225 104.255 ;
        RECT 37.395 103.460 37.725 104.305 ;
        RECT 37.965 103.245 38.260 104.055 ;
        RECT 38.440 103.415 38.685 104.555 ;
        RECT 38.860 103.245 39.120 104.055 ;
        RECT 39.300 103.420 39.550 104.555 ;
        RECT 45.730 104.385 46.895 104.975 ;
        RECT 47.155 105.045 48.365 105.795 ;
        RECT 48.535 105.070 48.825 105.795 ;
        RECT 49.005 105.295 49.335 105.795 ;
        RECT 49.535 105.225 49.705 105.575 ;
        RECT 49.905 105.395 50.235 105.795 ;
        RECT 50.405 105.225 50.575 105.575 ;
        RECT 50.745 105.395 51.125 105.795 ;
        RECT 47.155 104.505 47.675 105.045 ;
        RECT 40.150 104.160 46.895 104.385 ;
        RECT 47.845 104.335 48.365 104.875 ;
        RECT 49.000 104.555 49.350 105.125 ;
        RECT 49.535 105.055 51.145 105.225 ;
        RECT 51.315 105.120 51.585 105.465 ;
        RECT 50.975 104.885 51.145 105.055 ;
        RECT 40.150 104.145 45.555 104.160 ;
        RECT 39.720 103.250 39.980 104.045 ;
        RECT 40.150 103.420 40.410 104.145 ;
        RECT 40.580 103.250 40.840 103.975 ;
        RECT 41.010 103.420 41.270 104.145 ;
        RECT 41.440 103.250 41.700 103.975 ;
        RECT 41.870 103.420 42.130 104.145 ;
        RECT 42.300 103.250 42.560 103.975 ;
        RECT 42.730 103.420 42.990 104.145 ;
        RECT 43.160 103.250 43.405 103.975 ;
        RECT 43.575 103.420 43.835 104.145 ;
        RECT 44.020 103.250 44.265 103.975 ;
        RECT 44.435 103.420 44.695 104.145 ;
        RECT 44.880 103.250 45.125 103.975 ;
        RECT 45.295 103.420 45.555 104.145 ;
        RECT 45.740 103.250 45.995 103.975 ;
        RECT 46.165 103.420 46.455 104.160 ;
        RECT 39.720 103.245 45.995 103.250 ;
        RECT 46.625 103.245 46.895 103.990 ;
        RECT 47.155 103.245 48.365 104.335 ;
        RECT 48.535 103.245 48.825 104.410 ;
        RECT 49.000 104.095 49.320 104.385 ;
        RECT 49.520 104.265 50.230 104.885 ;
        RECT 50.400 104.555 50.805 104.885 ;
        RECT 50.975 104.555 51.245 104.885 ;
        RECT 50.975 104.385 51.145 104.555 ;
        RECT 51.415 104.385 51.585 105.120 ;
        RECT 50.420 104.215 51.145 104.385 ;
        RECT 50.420 104.095 50.590 104.215 ;
        RECT 49.000 103.925 50.590 104.095 ;
        RECT 49.000 103.465 50.655 103.755 ;
        RECT 50.825 103.245 51.105 104.045 ;
        RECT 51.315 103.415 51.585 104.385 ;
        RECT 52.215 105.055 52.600 105.625 ;
        RECT 52.770 105.335 53.095 105.795 ;
        RECT 53.615 105.165 53.895 105.625 ;
        RECT 52.215 104.385 52.495 105.055 ;
        RECT 52.770 104.995 53.895 105.165 ;
        RECT 52.770 104.885 53.220 104.995 ;
        RECT 52.665 104.555 53.220 104.885 ;
        RECT 54.085 104.825 54.485 105.625 ;
        RECT 54.885 105.335 55.155 105.795 ;
        RECT 55.325 105.165 55.610 105.625 ;
        RECT 52.215 103.415 52.600 104.385 ;
        RECT 52.770 104.095 53.220 104.555 ;
        RECT 53.390 104.265 54.485 104.825 ;
        RECT 52.770 103.875 53.895 104.095 ;
        RECT 52.770 103.245 53.095 103.705 ;
        RECT 53.615 103.415 53.895 103.875 ;
        RECT 54.085 103.415 54.485 104.265 ;
        RECT 54.655 104.995 55.610 105.165 ;
        RECT 55.985 105.245 56.155 105.535 ;
        RECT 56.325 105.415 56.655 105.795 ;
        RECT 55.985 105.075 56.650 105.245 ;
        RECT 54.655 104.095 54.865 104.995 ;
        RECT 55.035 104.265 55.725 104.825 ;
        RECT 55.900 104.255 56.250 104.905 ;
        RECT 54.655 103.875 55.610 104.095 ;
        RECT 56.420 104.085 56.650 105.075 ;
        RECT 54.885 103.245 55.155 103.705 ;
        RECT 55.325 103.415 55.610 103.875 ;
        RECT 55.985 103.915 56.650 104.085 ;
        RECT 55.985 103.415 56.155 103.915 ;
        RECT 56.325 103.245 56.655 103.745 ;
        RECT 56.825 103.415 57.010 105.535 ;
        RECT 57.265 105.335 57.515 105.795 ;
        RECT 57.685 105.345 58.020 105.515 ;
        RECT 58.215 105.345 58.890 105.515 ;
        RECT 57.685 105.205 57.855 105.345 ;
        RECT 57.180 104.215 57.460 105.165 ;
        RECT 57.630 105.075 57.855 105.205 ;
        RECT 57.630 103.970 57.800 105.075 ;
        RECT 58.025 104.925 58.550 105.145 ;
        RECT 57.970 104.160 58.210 104.755 ;
        RECT 58.380 104.225 58.550 104.925 ;
        RECT 58.720 104.565 58.890 105.345 ;
        RECT 59.210 105.295 59.580 105.795 ;
        RECT 59.760 105.345 60.165 105.515 ;
        RECT 60.335 105.345 61.120 105.515 ;
        RECT 59.760 105.115 59.930 105.345 ;
        RECT 59.100 104.815 59.930 105.115 ;
        RECT 60.315 104.845 60.780 105.175 ;
        RECT 59.100 104.785 59.300 104.815 ;
        RECT 59.420 104.565 59.590 104.635 ;
        RECT 58.720 104.395 59.590 104.565 ;
        RECT 59.080 104.305 59.590 104.395 ;
        RECT 57.630 103.840 57.935 103.970 ;
        RECT 58.380 103.860 58.910 104.225 ;
        RECT 57.250 103.245 57.515 103.705 ;
        RECT 57.685 103.415 57.935 103.840 ;
        RECT 59.080 103.690 59.250 104.305 ;
        RECT 58.145 103.520 59.250 103.690 ;
        RECT 59.420 103.245 59.590 104.045 ;
        RECT 59.760 103.745 59.930 104.815 ;
        RECT 60.100 103.915 60.290 104.635 ;
        RECT 60.460 103.885 60.780 104.845 ;
        RECT 60.950 104.885 61.120 105.345 ;
        RECT 61.395 105.265 61.605 105.795 ;
        RECT 61.865 105.055 62.195 105.580 ;
        RECT 62.365 105.185 62.535 105.795 ;
        RECT 62.705 105.140 63.035 105.575 ;
        RECT 63.205 105.280 63.375 105.795 ;
        RECT 62.705 105.055 63.085 105.140 ;
        RECT 61.995 104.885 62.195 105.055 ;
        RECT 62.860 105.015 63.085 105.055 ;
        RECT 60.950 104.555 61.825 104.885 ;
        RECT 61.995 104.555 62.745 104.885 ;
        RECT 59.760 103.415 60.010 103.745 ;
        RECT 60.950 103.715 61.120 104.555 ;
        RECT 61.995 104.350 62.185 104.555 ;
        RECT 62.915 104.435 63.085 105.015 ;
        RECT 62.870 104.385 63.085 104.435 ;
        RECT 61.290 103.975 62.185 104.350 ;
        RECT 62.695 104.305 63.085 104.385 ;
        RECT 63.750 105.055 64.365 105.625 ;
        RECT 64.535 105.285 64.750 105.795 ;
        RECT 64.980 105.285 65.260 105.615 ;
        RECT 65.440 105.285 65.680 105.795 ;
        RECT 60.235 103.545 61.120 103.715 ;
        RECT 61.300 103.245 61.615 103.745 ;
        RECT 61.845 103.415 62.185 103.975 ;
        RECT 62.355 103.245 62.525 104.255 ;
        RECT 62.695 103.460 63.025 104.305 ;
        RECT 63.195 103.245 63.365 104.160 ;
        RECT 63.750 104.035 64.065 105.055 ;
        RECT 64.235 104.385 64.405 104.885 ;
        RECT 64.655 104.555 64.920 105.115 ;
        RECT 65.090 104.385 65.260 105.285 ;
        RECT 66.985 105.140 67.315 105.575 ;
        RECT 67.485 105.185 67.655 105.795 ;
        RECT 65.430 104.555 65.785 105.115 ;
        RECT 66.935 105.055 67.315 105.140 ;
        RECT 67.825 105.055 68.155 105.580 ;
        RECT 68.415 105.265 68.625 105.795 ;
        RECT 68.900 105.345 69.685 105.515 ;
        RECT 69.855 105.345 70.260 105.515 ;
        RECT 66.935 105.015 67.160 105.055 ;
        RECT 66.935 104.435 67.105 105.015 ;
        RECT 67.825 104.885 68.025 105.055 ;
        RECT 68.900 104.885 69.070 105.345 ;
        RECT 67.275 104.555 68.025 104.885 ;
        RECT 68.195 104.555 69.070 104.885 ;
        RECT 66.935 104.385 67.150 104.435 ;
        RECT 64.235 104.215 65.660 104.385 ;
        RECT 66.935 104.305 67.325 104.385 ;
        RECT 63.750 103.415 64.285 104.035 ;
        RECT 64.455 103.245 64.785 104.045 ;
        RECT 65.270 104.040 65.660 104.215 ;
        RECT 66.995 103.460 67.325 104.305 ;
        RECT 67.835 104.350 68.025 104.555 ;
        RECT 67.495 103.245 67.665 104.255 ;
        RECT 67.835 103.975 68.730 104.350 ;
        RECT 67.835 103.415 68.175 103.975 ;
        RECT 68.405 103.245 68.720 103.745 ;
        RECT 68.900 103.715 69.070 104.555 ;
        RECT 69.240 104.845 69.705 105.175 ;
        RECT 70.090 105.115 70.260 105.345 ;
        RECT 70.440 105.295 70.810 105.795 ;
        RECT 71.130 105.345 71.805 105.515 ;
        RECT 72.000 105.345 72.335 105.515 ;
        RECT 69.240 103.885 69.560 104.845 ;
        RECT 70.090 104.815 70.920 105.115 ;
        RECT 69.730 103.915 69.920 104.635 ;
        RECT 70.090 103.745 70.260 104.815 ;
        RECT 70.720 104.785 70.920 104.815 ;
        RECT 70.430 104.565 70.600 104.635 ;
        RECT 71.130 104.565 71.300 105.345 ;
        RECT 72.165 105.205 72.335 105.345 ;
        RECT 72.505 105.335 72.755 105.795 ;
        RECT 70.430 104.395 71.300 104.565 ;
        RECT 71.470 104.925 71.995 105.145 ;
        RECT 72.165 105.075 72.390 105.205 ;
        RECT 70.430 104.305 70.940 104.395 ;
        RECT 68.900 103.545 69.785 103.715 ;
        RECT 70.010 103.415 70.260 103.745 ;
        RECT 70.430 103.245 70.600 104.045 ;
        RECT 70.770 103.690 70.940 104.305 ;
        RECT 71.470 104.225 71.640 104.925 ;
        RECT 71.110 103.860 71.640 104.225 ;
        RECT 71.810 104.160 72.050 104.755 ;
        RECT 72.220 103.970 72.390 105.075 ;
        RECT 72.560 104.215 72.840 105.165 ;
        RECT 72.085 103.840 72.390 103.970 ;
        RECT 70.770 103.520 71.875 103.690 ;
        RECT 72.085 103.415 72.335 103.840 ;
        RECT 72.505 103.245 72.770 103.705 ;
        RECT 73.010 103.415 73.195 105.535 ;
        RECT 73.365 105.415 73.695 105.795 ;
        RECT 73.865 105.245 74.035 105.535 ;
        RECT 73.370 105.075 74.035 105.245 ;
        RECT 73.370 104.085 73.600 105.075 ;
        RECT 74.295 105.070 74.585 105.795 ;
        RECT 74.775 105.405 75.950 105.625 ;
        RECT 74.755 104.985 75.530 105.235 ;
        RECT 75.700 105.155 75.950 105.405 ;
        RECT 76.120 105.325 76.290 105.795 ;
        RECT 76.460 105.155 76.790 105.625 ;
        RECT 73.770 104.255 74.120 104.905 ;
        RECT 73.370 103.915 74.035 104.085 ;
        RECT 73.365 103.245 73.695 103.745 ;
        RECT 73.865 103.415 74.035 103.915 ;
        RECT 74.295 103.245 74.585 104.410 ;
        RECT 74.755 104.095 74.985 104.985 ;
        RECT 75.700 104.975 76.790 105.155 ;
        RECT 77.100 104.975 77.270 105.795 ;
        RECT 77.440 105.155 77.770 105.625 ;
        RECT 77.940 105.325 78.110 105.795 ;
        RECT 78.280 105.155 78.645 105.625 ;
        RECT 78.815 105.325 78.985 105.795 ;
        RECT 79.255 105.405 80.565 105.575 ;
        RECT 79.675 105.155 80.005 105.235 ;
        RECT 77.440 104.975 80.005 105.155 ;
        RECT 75.155 104.595 75.630 104.805 ;
        RECT 75.925 104.605 77.375 104.805 ;
        RECT 75.460 104.435 75.630 104.595 ;
        RECT 77.600 104.595 78.625 104.805 ;
        RECT 79.305 104.635 79.965 104.805 ;
        RECT 77.600 104.435 77.770 104.595 ;
        RECT 75.460 104.265 77.770 104.435 ;
        RECT 79.305 104.425 79.475 104.635 ;
        RECT 80.175 104.465 80.565 105.405 ;
        RECT 80.735 105.025 82.405 105.795 ;
        RECT 80.735 104.505 81.485 105.025 ;
        RECT 83.040 104.975 83.335 105.795 ;
        RECT 83.505 105.245 83.725 105.625 ;
        RECT 83.895 105.435 84.745 105.795 ;
        RECT 77.980 104.255 79.475 104.425 ;
        RECT 79.715 104.255 80.565 104.465 ;
        RECT 81.655 104.335 82.405 104.855 ;
        RECT 77.980 104.095 78.150 104.255 ;
        RECT 74.755 103.925 78.150 104.095 ;
        RECT 79.715 104.085 79.965 104.255 ;
        RECT 74.755 103.915 76.750 103.925 ;
        RECT 74.755 103.415 75.070 103.915 ;
        RECT 75.240 103.245 75.490 103.745 ;
        RECT 75.660 103.415 75.910 103.915 ;
        RECT 76.080 103.245 76.330 103.745 ;
        RECT 76.500 103.415 76.750 103.915 ;
        RECT 78.395 103.915 79.965 104.085 ;
        RECT 78.395 103.755 78.605 103.915 ;
        RECT 79.715 103.755 79.965 103.915 ;
        RECT 77.060 103.415 77.310 103.755 ;
        RECT 77.480 103.245 77.730 103.745 ;
        RECT 77.900 103.585 78.225 103.755 ;
        RECT 78.775 103.585 79.025 103.745 ;
        RECT 77.900 103.415 79.025 103.585 ;
        RECT 79.295 103.245 79.545 103.745 ;
        RECT 80.135 103.245 80.565 104.085 ;
        RECT 80.735 103.245 82.405 104.335 ;
        RECT 83.040 103.245 83.335 104.390 ;
        RECT 83.505 103.545 83.735 105.245 ;
        RECT 85.225 105.185 85.555 105.605 ;
        RECT 85.760 105.355 86.035 105.795 ;
        RECT 86.205 105.185 86.535 105.605 ;
        RECT 83.950 105.005 86.535 105.185 ;
        RECT 83.950 104.390 84.260 105.005 ;
        RECT 86.725 104.985 86.995 105.795 ;
        RECT 87.165 104.985 87.495 105.625 ;
        RECT 87.665 104.985 87.905 105.795 ;
        RECT 84.430 104.605 84.760 104.835 ;
        RECT 84.930 104.605 85.400 104.835 ;
        RECT 85.570 104.775 86.020 104.835 ;
        RECT 85.570 104.605 86.025 104.775 ;
        RECT 86.210 104.605 86.545 104.835 ;
        RECT 86.715 104.555 87.065 104.805 ;
        RECT 83.950 104.220 86.535 104.390 ;
        RECT 87.235 104.385 87.405 104.985 ;
        RECT 88.560 104.975 88.855 105.795 ;
        RECT 89.025 105.245 89.245 105.625 ;
        RECT 89.415 105.435 90.265 105.795 ;
        RECT 87.575 104.555 87.925 104.805 ;
        RECT 83.950 103.245 84.205 104.050 ;
        RECT 84.405 103.860 85.745 104.040 ;
        RECT 84.405 103.415 84.735 103.860 ;
        RECT 84.905 103.245 85.180 103.690 ;
        RECT 85.415 103.415 85.745 103.860 ;
        RECT 86.205 103.555 86.535 104.220 ;
        RECT 86.725 103.245 87.055 104.385 ;
        RECT 87.235 104.215 87.915 104.385 ;
        RECT 87.585 103.430 87.915 104.215 ;
        RECT 88.560 103.245 88.855 104.390 ;
        RECT 89.025 103.545 89.255 105.245 ;
        RECT 90.745 105.185 91.075 105.605 ;
        RECT 91.280 105.355 91.555 105.795 ;
        RECT 91.725 105.185 92.055 105.605 ;
        RECT 89.470 105.005 92.055 105.185 ;
        RECT 92.325 105.245 92.495 105.535 ;
        RECT 92.665 105.415 92.995 105.795 ;
        RECT 92.325 105.075 92.990 105.245 ;
        RECT 89.470 104.390 89.780 105.005 ;
        RECT 89.950 104.605 90.280 104.835 ;
        RECT 90.450 104.605 90.920 104.835 ;
        RECT 91.090 104.775 91.540 104.835 ;
        RECT 91.090 104.605 91.545 104.775 ;
        RECT 91.730 104.605 92.065 104.835 ;
        RECT 89.470 104.220 92.055 104.390 ;
        RECT 92.240 104.255 92.590 104.905 ;
        RECT 89.470 103.245 89.725 104.050 ;
        RECT 89.925 103.860 91.265 104.040 ;
        RECT 89.925 103.415 90.255 103.860 ;
        RECT 90.425 103.245 90.700 103.690 ;
        RECT 90.935 103.415 91.265 103.860 ;
        RECT 91.725 103.555 92.055 104.220 ;
        RECT 92.760 104.085 92.990 105.075 ;
        RECT 92.325 103.915 92.990 104.085 ;
        RECT 92.325 103.415 92.495 103.915 ;
        RECT 92.665 103.245 92.995 103.745 ;
        RECT 93.165 103.415 93.350 105.535 ;
        RECT 93.605 105.335 93.855 105.795 ;
        RECT 94.025 105.345 94.360 105.515 ;
        RECT 94.555 105.345 95.230 105.515 ;
        RECT 94.025 105.205 94.195 105.345 ;
        RECT 93.520 104.215 93.800 105.165 ;
        RECT 93.970 105.075 94.195 105.205 ;
        RECT 93.970 103.970 94.140 105.075 ;
        RECT 94.365 104.925 94.890 105.145 ;
        RECT 94.310 104.160 94.550 104.755 ;
        RECT 94.720 104.225 94.890 104.925 ;
        RECT 95.060 104.565 95.230 105.345 ;
        RECT 95.550 105.295 95.920 105.795 ;
        RECT 96.100 105.345 96.505 105.515 ;
        RECT 96.675 105.345 97.460 105.515 ;
        RECT 96.100 105.115 96.270 105.345 ;
        RECT 95.440 104.815 96.270 105.115 ;
        RECT 96.655 104.845 97.120 105.175 ;
        RECT 95.440 104.785 95.640 104.815 ;
        RECT 95.760 104.565 95.930 104.635 ;
        RECT 95.060 104.395 95.930 104.565 ;
        RECT 95.420 104.305 95.930 104.395 ;
        RECT 93.970 103.840 94.275 103.970 ;
        RECT 94.720 103.860 95.250 104.225 ;
        RECT 93.590 103.245 93.855 103.705 ;
        RECT 94.025 103.415 94.275 103.840 ;
        RECT 95.420 103.690 95.590 104.305 ;
        RECT 94.485 103.520 95.590 103.690 ;
        RECT 95.760 103.245 95.930 104.045 ;
        RECT 96.100 103.745 96.270 104.815 ;
        RECT 96.440 103.915 96.630 104.635 ;
        RECT 96.800 103.885 97.120 104.845 ;
        RECT 97.290 104.885 97.460 105.345 ;
        RECT 97.735 105.265 97.945 105.795 ;
        RECT 98.205 105.055 98.535 105.580 ;
        RECT 98.705 105.185 98.875 105.795 ;
        RECT 99.045 105.140 99.375 105.575 ;
        RECT 99.045 105.055 99.425 105.140 ;
        RECT 100.055 105.070 100.345 105.795 ;
        RECT 98.335 104.885 98.535 105.055 ;
        RECT 99.200 105.015 99.425 105.055 ;
        RECT 97.290 104.555 98.165 104.885 ;
        RECT 98.335 104.555 99.085 104.885 ;
        RECT 96.100 103.415 96.350 103.745 ;
        RECT 97.290 103.715 97.460 104.555 ;
        RECT 98.335 104.350 98.525 104.555 ;
        RECT 99.255 104.435 99.425 105.015 ;
        RECT 99.210 104.385 99.425 104.435 ;
        RECT 100.520 105.055 100.775 105.625 ;
        RECT 100.945 105.395 101.275 105.795 ;
        RECT 101.700 105.260 102.230 105.625 ;
        RECT 101.700 105.225 101.875 105.260 ;
        RECT 100.945 105.055 101.875 105.225 ;
        RECT 102.420 105.115 102.695 105.625 ;
        RECT 97.630 103.975 98.525 104.350 ;
        RECT 99.035 104.305 99.425 104.385 ;
        RECT 96.575 103.545 97.460 103.715 ;
        RECT 97.640 103.245 97.955 103.745 ;
        RECT 98.185 103.415 98.525 103.975 ;
        RECT 98.695 103.245 98.865 104.255 ;
        RECT 99.035 103.460 99.365 104.305 ;
        RECT 100.055 103.245 100.345 104.410 ;
        RECT 100.520 104.385 100.690 105.055 ;
        RECT 100.945 104.885 101.115 105.055 ;
        RECT 100.860 104.555 101.115 104.885 ;
        RECT 101.340 104.555 101.535 104.885 ;
        RECT 100.520 103.415 100.855 104.385 ;
        RECT 101.025 103.245 101.195 104.385 ;
        RECT 101.365 103.585 101.535 104.555 ;
        RECT 101.705 103.925 101.875 105.055 ;
        RECT 102.045 104.265 102.215 105.065 ;
        RECT 102.415 104.945 102.695 105.115 ;
        RECT 102.420 104.465 102.695 104.945 ;
        RECT 102.865 104.265 103.055 105.625 ;
        RECT 103.235 105.260 103.745 105.795 ;
        RECT 103.965 104.985 104.210 105.590 ;
        RECT 104.655 105.025 106.325 105.795 ;
        RECT 106.960 105.055 107.215 105.625 ;
        RECT 107.385 105.395 107.715 105.795 ;
        RECT 108.140 105.260 108.670 105.625 ;
        RECT 108.140 105.225 108.315 105.260 ;
        RECT 107.385 105.055 108.315 105.225 ;
        RECT 103.255 104.815 104.485 104.985 ;
        RECT 102.045 104.095 103.055 104.265 ;
        RECT 103.225 104.250 103.975 104.440 ;
        RECT 101.705 103.755 102.830 103.925 ;
        RECT 103.225 103.585 103.395 104.250 ;
        RECT 104.145 104.005 104.485 104.815 ;
        RECT 104.655 104.505 105.405 105.025 ;
        RECT 105.575 104.335 106.325 104.855 ;
        RECT 101.365 103.415 103.395 103.585 ;
        RECT 103.565 103.245 103.735 104.005 ;
        RECT 103.970 103.595 104.485 104.005 ;
        RECT 104.655 103.245 106.325 104.335 ;
        RECT 106.960 104.385 107.130 105.055 ;
        RECT 107.385 104.885 107.555 105.055 ;
        RECT 107.300 104.555 107.555 104.885 ;
        RECT 107.780 104.555 107.975 104.885 ;
        RECT 106.960 103.415 107.295 104.385 ;
        RECT 107.465 103.245 107.635 104.385 ;
        RECT 107.805 103.585 107.975 104.555 ;
        RECT 108.145 103.925 108.315 105.055 ;
        RECT 108.485 104.265 108.655 105.065 ;
        RECT 108.860 104.775 109.135 105.625 ;
        RECT 108.855 104.605 109.135 104.775 ;
        RECT 108.860 104.465 109.135 104.605 ;
        RECT 109.305 104.265 109.495 105.625 ;
        RECT 109.675 105.260 110.185 105.795 ;
        RECT 110.405 104.985 110.650 105.590 ;
        RECT 109.695 104.815 110.925 104.985 ;
        RECT 111.100 104.975 111.395 105.795 ;
        RECT 111.565 105.245 111.785 105.625 ;
        RECT 111.955 105.435 112.805 105.795 ;
        RECT 108.485 104.095 109.495 104.265 ;
        RECT 109.665 104.250 110.415 104.440 ;
        RECT 108.145 103.755 109.270 103.925 ;
        RECT 109.665 103.585 109.835 104.250 ;
        RECT 110.585 104.005 110.925 104.815 ;
        RECT 107.805 103.415 109.835 103.585 ;
        RECT 110.005 103.245 110.175 104.005 ;
        RECT 110.410 103.595 110.925 104.005 ;
        RECT 111.100 103.245 111.395 104.390 ;
        RECT 111.565 103.545 111.795 105.245 ;
        RECT 113.285 105.185 113.615 105.605 ;
        RECT 113.820 105.355 114.095 105.795 ;
        RECT 114.265 105.185 114.595 105.605 ;
        RECT 112.010 105.005 114.595 105.185 ;
        RECT 115.235 105.120 115.495 105.625 ;
        RECT 115.675 105.415 116.005 105.795 ;
        RECT 116.185 105.245 116.355 105.625 ;
        RECT 112.010 104.390 112.320 105.005 ;
        RECT 112.490 104.605 112.820 104.835 ;
        RECT 112.990 104.605 113.460 104.835 ;
        RECT 113.630 104.775 114.080 104.835 ;
        RECT 113.630 104.605 114.085 104.775 ;
        RECT 114.270 104.605 114.605 104.835 ;
        RECT 112.010 104.220 114.595 104.390 ;
        RECT 112.010 103.245 112.265 104.050 ;
        RECT 112.465 103.860 113.805 104.040 ;
        RECT 112.465 103.415 112.795 103.860 ;
        RECT 112.965 103.245 113.240 103.690 ;
        RECT 113.475 103.415 113.805 103.860 ;
        RECT 114.265 103.555 114.595 104.220 ;
        RECT 115.235 104.320 115.405 105.120 ;
        RECT 115.690 105.075 116.355 105.245 ;
        RECT 115.690 104.820 115.860 105.075 ;
        RECT 116.620 105.055 116.875 105.625 ;
        RECT 117.045 105.395 117.375 105.795 ;
        RECT 117.800 105.260 118.330 105.625 ;
        RECT 118.520 105.455 118.795 105.625 ;
        RECT 118.515 105.285 118.795 105.455 ;
        RECT 117.800 105.225 117.975 105.260 ;
        RECT 117.045 105.055 117.975 105.225 ;
        RECT 115.575 104.490 115.860 104.820 ;
        RECT 116.095 104.525 116.425 104.895 ;
        RECT 115.690 104.345 115.860 104.490 ;
        RECT 116.620 104.385 116.790 105.055 ;
        RECT 117.045 104.885 117.215 105.055 ;
        RECT 116.960 104.555 117.215 104.885 ;
        RECT 117.440 104.555 117.635 104.885 ;
        RECT 115.235 103.415 115.505 104.320 ;
        RECT 115.690 104.175 116.355 104.345 ;
        RECT 115.675 103.245 116.005 104.005 ;
        RECT 116.185 103.415 116.355 104.175 ;
        RECT 116.620 103.415 116.955 104.385 ;
        RECT 117.125 103.245 117.295 104.385 ;
        RECT 117.465 103.585 117.635 104.555 ;
        RECT 117.805 103.925 117.975 105.055 ;
        RECT 118.145 104.265 118.315 105.065 ;
        RECT 118.520 104.465 118.795 105.285 ;
        RECT 118.965 104.265 119.155 105.625 ;
        RECT 119.335 105.260 119.845 105.795 ;
        RECT 120.065 104.985 120.310 105.590 ;
        RECT 120.755 105.025 122.425 105.795 ;
        RECT 122.645 105.405 122.975 105.795 ;
        RECT 123.145 105.225 123.315 105.545 ;
        RECT 123.485 105.405 123.815 105.795 ;
        RECT 124.230 105.395 125.185 105.565 ;
        RECT 122.595 105.055 124.845 105.225 ;
        RECT 119.355 104.815 120.585 104.985 ;
        RECT 118.145 104.095 119.155 104.265 ;
        RECT 119.325 104.250 120.075 104.440 ;
        RECT 117.805 103.755 118.930 103.925 ;
        RECT 119.325 103.585 119.495 104.250 ;
        RECT 120.245 104.005 120.585 104.815 ;
        RECT 120.755 104.505 121.505 105.025 ;
        RECT 121.675 104.335 122.425 104.855 ;
        RECT 117.465 103.415 119.495 103.585 ;
        RECT 119.665 103.245 119.835 104.005 ;
        RECT 120.070 103.595 120.585 104.005 ;
        RECT 120.755 103.245 122.425 104.335 ;
        RECT 122.595 104.095 122.765 105.055 ;
        RECT 122.935 104.435 123.180 104.885 ;
        RECT 123.350 104.605 123.900 104.805 ;
        RECT 124.070 104.635 124.445 104.805 ;
        RECT 124.070 104.435 124.240 104.635 ;
        RECT 124.615 104.555 124.845 105.055 ;
        RECT 122.935 104.265 124.240 104.435 ;
        RECT 125.015 104.515 125.185 105.395 ;
        RECT 125.355 104.960 125.645 105.795 ;
        RECT 125.815 105.070 126.105 105.795 ;
        RECT 126.325 105.140 126.655 105.575 ;
        RECT 126.825 105.185 126.995 105.795 ;
        RECT 126.275 105.055 126.655 105.140 ;
        RECT 127.165 105.055 127.495 105.580 ;
        RECT 127.755 105.265 127.965 105.795 ;
        RECT 128.240 105.345 129.025 105.515 ;
        RECT 129.195 105.345 129.600 105.515 ;
        RECT 126.275 105.015 126.500 105.055 ;
        RECT 125.015 104.345 125.645 104.515 ;
        RECT 126.275 104.435 126.445 105.015 ;
        RECT 127.165 104.885 127.365 105.055 ;
        RECT 128.240 104.885 128.410 105.345 ;
        RECT 126.615 104.555 127.365 104.885 ;
        RECT 127.535 104.555 128.410 104.885 ;
        RECT 122.595 103.415 122.975 104.095 ;
        RECT 123.565 103.245 123.735 104.095 ;
        RECT 123.905 103.925 125.145 104.095 ;
        RECT 123.905 103.415 124.235 103.925 ;
        RECT 124.405 103.245 124.575 103.755 ;
        RECT 124.745 103.415 125.145 103.925 ;
        RECT 125.325 103.415 125.645 104.345 ;
        RECT 125.815 103.245 126.105 104.410 ;
        RECT 126.275 104.385 126.490 104.435 ;
        RECT 126.275 104.305 126.665 104.385 ;
        RECT 126.335 103.460 126.665 104.305 ;
        RECT 127.175 104.350 127.365 104.555 ;
        RECT 126.835 103.245 127.005 104.255 ;
        RECT 127.175 103.975 128.070 104.350 ;
        RECT 127.175 103.415 127.515 103.975 ;
        RECT 127.745 103.245 128.060 103.745 ;
        RECT 128.240 103.715 128.410 104.555 ;
        RECT 128.580 104.845 129.045 105.175 ;
        RECT 129.430 105.115 129.600 105.345 ;
        RECT 129.780 105.295 130.150 105.795 ;
        RECT 130.470 105.345 131.145 105.515 ;
        RECT 131.340 105.345 131.675 105.515 ;
        RECT 128.580 103.885 128.900 104.845 ;
        RECT 129.430 104.815 130.260 105.115 ;
        RECT 129.070 103.915 129.260 104.635 ;
        RECT 129.430 103.745 129.600 104.815 ;
        RECT 130.060 104.785 130.260 104.815 ;
        RECT 129.770 104.565 129.940 104.635 ;
        RECT 130.470 104.565 130.640 105.345 ;
        RECT 131.505 105.205 131.675 105.345 ;
        RECT 131.845 105.335 132.095 105.795 ;
        RECT 129.770 104.395 130.640 104.565 ;
        RECT 130.810 104.925 131.335 105.145 ;
        RECT 131.505 105.075 131.730 105.205 ;
        RECT 129.770 104.305 130.280 104.395 ;
        RECT 128.240 103.545 129.125 103.715 ;
        RECT 129.350 103.415 129.600 103.745 ;
        RECT 129.770 103.245 129.940 104.045 ;
        RECT 130.110 103.690 130.280 104.305 ;
        RECT 130.810 104.225 130.980 104.925 ;
        RECT 130.450 103.860 130.980 104.225 ;
        RECT 131.150 104.160 131.390 104.755 ;
        RECT 131.560 103.970 131.730 105.075 ;
        RECT 131.900 104.215 132.180 105.165 ;
        RECT 131.425 103.840 131.730 103.970 ;
        RECT 130.110 103.520 131.215 103.690 ;
        RECT 131.425 103.415 131.675 103.840 ;
        RECT 131.845 103.245 132.110 103.705 ;
        RECT 132.350 103.415 132.535 105.535 ;
        RECT 132.705 105.415 133.035 105.795 ;
        RECT 133.205 105.245 133.375 105.535 ;
        RECT 133.635 105.250 138.980 105.795 ;
        RECT 132.710 105.075 133.375 105.245 ;
        RECT 132.710 104.085 132.940 105.075 ;
        RECT 133.110 104.255 133.460 104.905 ;
        RECT 135.220 104.420 135.560 105.250 ;
        RECT 139.155 105.025 142.665 105.795 ;
        RECT 143.385 105.245 143.555 105.625 ;
        RECT 143.735 105.415 144.065 105.795 ;
        RECT 143.385 105.075 144.050 105.245 ;
        RECT 144.245 105.120 144.505 105.625 ;
        RECT 144.675 105.250 150.020 105.795 ;
        RECT 132.710 103.915 133.375 104.085 ;
        RECT 132.705 103.245 133.035 103.745 ;
        RECT 133.205 103.415 133.375 103.915 ;
        RECT 137.040 103.680 137.390 104.930 ;
        RECT 139.155 104.505 140.805 105.025 ;
        RECT 140.975 104.335 142.665 104.855 ;
        RECT 143.315 104.525 143.645 104.895 ;
        RECT 143.880 104.820 144.050 105.075 ;
        RECT 143.880 104.490 144.165 104.820 ;
        RECT 143.880 104.345 144.050 104.490 ;
        RECT 133.635 103.245 138.980 103.680 ;
        RECT 139.155 103.245 142.665 104.335 ;
        RECT 143.385 104.175 144.050 104.345 ;
        RECT 144.335 104.320 144.505 105.120 ;
        RECT 146.260 104.420 146.600 105.250 ;
        RECT 150.195 105.045 151.405 105.795 ;
        RECT 151.575 105.070 151.865 105.795 ;
        RECT 143.385 103.415 143.555 104.175 ;
        RECT 143.735 103.245 144.065 104.005 ;
        RECT 144.235 103.415 144.505 104.320 ;
        RECT 148.080 103.680 148.430 104.930 ;
        RECT 150.195 104.505 150.715 105.045 ;
        RECT 152.035 105.025 155.545 105.795 ;
        RECT 155.715 105.045 156.925 105.795 ;
        RECT 150.885 104.335 151.405 104.875 ;
        RECT 152.035 104.505 153.685 105.025 ;
        RECT 144.675 103.245 150.020 103.680 ;
        RECT 150.195 103.245 151.405 104.335 ;
        RECT 151.575 103.245 151.865 104.410 ;
        RECT 153.855 104.335 155.545 104.855 ;
        RECT 152.035 103.245 155.545 104.335 ;
        RECT 155.715 104.335 156.235 104.875 ;
        RECT 156.405 104.505 156.925 105.045 ;
        RECT 155.715 103.245 156.925 104.335 ;
        RECT 22.690 103.075 157.010 103.245 ;
        RECT 22.775 101.985 23.985 103.075 ;
        RECT 24.215 102.015 24.545 102.860 ;
        RECT 24.715 102.065 24.885 103.075 ;
        RECT 25.055 102.345 25.395 102.905 ;
        RECT 25.625 102.575 25.940 103.075 ;
        RECT 26.120 102.605 27.005 102.775 ;
        RECT 22.775 101.275 23.295 101.815 ;
        RECT 23.465 101.445 23.985 101.985 ;
        RECT 24.155 101.935 24.545 102.015 ;
        RECT 25.055 101.970 25.950 102.345 ;
        RECT 24.155 101.885 24.370 101.935 ;
        RECT 24.155 101.305 24.325 101.885 ;
        RECT 25.055 101.765 25.245 101.970 ;
        RECT 26.120 101.765 26.290 102.605 ;
        RECT 27.230 102.575 27.480 102.905 ;
        RECT 24.495 101.435 25.245 101.765 ;
        RECT 25.415 101.435 26.290 101.765 ;
        RECT 22.775 100.525 23.985 101.275 ;
        RECT 24.155 101.265 24.380 101.305 ;
        RECT 25.045 101.265 25.245 101.435 ;
        RECT 24.155 101.180 24.535 101.265 ;
        RECT 24.205 100.745 24.535 101.180 ;
        RECT 24.705 100.525 24.875 101.135 ;
        RECT 25.045 100.740 25.375 101.265 ;
        RECT 25.635 100.525 25.845 101.055 ;
        RECT 26.120 100.975 26.290 101.435 ;
        RECT 26.460 101.475 26.780 102.435 ;
        RECT 26.950 101.685 27.140 102.405 ;
        RECT 27.310 101.505 27.480 102.575 ;
        RECT 27.650 102.275 27.820 103.075 ;
        RECT 27.990 102.630 29.095 102.800 ;
        RECT 27.990 102.015 28.160 102.630 ;
        RECT 29.305 102.480 29.555 102.905 ;
        RECT 29.725 102.615 29.990 103.075 ;
        RECT 28.330 102.095 28.860 102.460 ;
        RECT 29.305 102.350 29.610 102.480 ;
        RECT 27.650 101.925 28.160 102.015 ;
        RECT 27.650 101.755 28.520 101.925 ;
        RECT 27.650 101.685 27.820 101.755 ;
        RECT 27.940 101.505 28.140 101.535 ;
        RECT 26.460 101.145 26.925 101.475 ;
        RECT 27.310 101.205 28.140 101.505 ;
        RECT 27.310 100.975 27.480 101.205 ;
        RECT 26.120 100.805 26.905 100.975 ;
        RECT 27.075 100.805 27.480 100.975 ;
        RECT 27.660 100.525 28.030 101.025 ;
        RECT 28.350 100.975 28.520 101.755 ;
        RECT 28.690 101.395 28.860 102.095 ;
        RECT 29.030 101.565 29.270 102.160 ;
        RECT 28.690 101.175 29.215 101.395 ;
        RECT 29.440 101.245 29.610 102.350 ;
        RECT 29.385 101.115 29.610 101.245 ;
        RECT 29.780 101.155 30.060 102.105 ;
        RECT 29.385 100.975 29.555 101.115 ;
        RECT 28.350 100.805 29.025 100.975 ;
        RECT 29.220 100.805 29.555 100.975 ;
        RECT 29.725 100.525 29.975 100.985 ;
        RECT 30.230 100.785 30.415 102.905 ;
        RECT 30.585 102.575 30.915 103.075 ;
        RECT 31.085 102.405 31.255 102.905 ;
        RECT 30.590 102.235 31.255 102.405 ;
        RECT 30.590 101.245 30.820 102.235 ;
        RECT 32.180 102.105 32.510 102.905 ;
        RECT 32.680 102.275 33.010 103.075 ;
        RECT 33.310 102.105 33.640 102.905 ;
        RECT 34.285 102.275 34.535 103.075 ;
        RECT 30.990 101.415 31.340 102.065 ;
        RECT 32.180 101.935 34.615 102.105 ;
        RECT 34.805 101.935 34.975 103.075 ;
        RECT 35.145 101.935 35.485 102.905 ;
        RECT 31.975 101.515 32.325 101.765 ;
        RECT 32.510 101.305 32.680 101.935 ;
        RECT 32.850 101.515 33.180 101.715 ;
        RECT 33.350 101.515 33.680 101.715 ;
        RECT 33.850 101.515 34.270 101.715 ;
        RECT 34.445 101.685 34.615 101.935 ;
        RECT 34.445 101.515 35.140 101.685 ;
        RECT 30.590 101.075 31.255 101.245 ;
        RECT 30.585 100.525 30.915 100.905 ;
        RECT 31.085 100.785 31.255 101.075 ;
        RECT 32.180 100.695 32.680 101.305 ;
        RECT 33.310 101.175 34.535 101.345 ;
        RECT 35.310 101.325 35.485 101.935 ;
        RECT 35.655 101.910 35.945 103.075 ;
        RECT 36.760 102.105 37.150 102.280 ;
        RECT 37.635 102.275 37.965 103.075 ;
        RECT 38.135 102.285 38.670 102.905 ;
        RECT 36.760 101.935 38.185 102.105 ;
        RECT 33.310 100.695 33.640 101.175 ;
        RECT 33.810 100.525 34.035 100.985 ;
        RECT 34.205 100.695 34.535 101.175 ;
        RECT 34.725 100.525 34.975 101.325 ;
        RECT 35.145 100.695 35.485 101.325 ;
        RECT 35.655 100.525 35.945 101.250 ;
        RECT 36.635 101.205 36.990 101.765 ;
        RECT 37.160 101.035 37.330 101.935 ;
        RECT 37.500 101.205 37.765 101.765 ;
        RECT 38.015 101.435 38.185 101.935 ;
        RECT 38.355 101.265 38.670 102.285 ;
        RECT 36.740 100.525 36.980 101.035 ;
        RECT 37.160 100.705 37.440 101.035 ;
        RECT 37.670 100.525 37.885 101.035 ;
        RECT 38.055 100.695 38.670 101.265 ;
        RECT 38.875 101.935 39.260 102.905 ;
        RECT 39.430 102.615 39.755 103.075 ;
        RECT 40.275 102.445 40.555 102.905 ;
        RECT 39.430 102.225 40.555 102.445 ;
        RECT 38.875 101.265 39.155 101.935 ;
        RECT 39.430 101.765 39.880 102.225 ;
        RECT 40.745 102.055 41.145 102.905 ;
        RECT 41.545 102.615 41.815 103.075 ;
        RECT 41.985 102.445 42.270 102.905 ;
        RECT 39.325 101.435 39.880 101.765 ;
        RECT 40.050 101.495 41.145 102.055 ;
        RECT 39.430 101.325 39.880 101.435 ;
        RECT 38.875 100.695 39.260 101.265 ;
        RECT 39.430 101.155 40.555 101.325 ;
        RECT 39.430 100.525 39.755 100.985 ;
        RECT 40.275 100.695 40.555 101.155 ;
        RECT 40.745 100.695 41.145 101.495 ;
        RECT 41.315 102.225 42.270 102.445 ;
        RECT 42.645 102.405 42.815 102.905 ;
        RECT 42.985 102.575 43.315 103.075 ;
        RECT 42.645 102.235 43.310 102.405 ;
        RECT 41.315 101.325 41.525 102.225 ;
        RECT 41.695 101.495 42.385 102.055 ;
        RECT 42.560 101.415 42.910 102.065 ;
        RECT 41.315 101.155 42.270 101.325 ;
        RECT 43.080 101.245 43.310 102.235 ;
        RECT 41.545 100.525 41.815 100.985 ;
        RECT 41.985 100.695 42.270 101.155 ;
        RECT 42.645 101.075 43.310 101.245 ;
        RECT 42.645 100.785 42.815 101.075 ;
        RECT 42.985 100.525 43.315 100.905 ;
        RECT 43.485 100.785 43.670 102.905 ;
        RECT 43.910 102.615 44.175 103.075 ;
        RECT 44.345 102.480 44.595 102.905 ;
        RECT 44.805 102.630 45.910 102.800 ;
        RECT 44.290 102.350 44.595 102.480 ;
        RECT 43.840 101.155 44.120 102.105 ;
        RECT 44.290 101.245 44.460 102.350 ;
        RECT 44.630 101.565 44.870 102.160 ;
        RECT 45.040 102.095 45.570 102.460 ;
        RECT 45.040 101.395 45.210 102.095 ;
        RECT 45.740 102.015 45.910 102.630 ;
        RECT 46.080 102.275 46.250 103.075 ;
        RECT 46.420 102.575 46.670 102.905 ;
        RECT 46.895 102.605 47.780 102.775 ;
        RECT 45.740 101.925 46.250 102.015 ;
        RECT 44.290 101.115 44.515 101.245 ;
        RECT 44.685 101.175 45.210 101.395 ;
        RECT 45.380 101.755 46.250 101.925 ;
        RECT 43.925 100.525 44.175 100.985 ;
        RECT 44.345 100.975 44.515 101.115 ;
        RECT 45.380 100.975 45.550 101.755 ;
        RECT 46.080 101.685 46.250 101.755 ;
        RECT 45.760 101.505 45.960 101.535 ;
        RECT 46.420 101.505 46.590 102.575 ;
        RECT 46.760 101.685 46.950 102.405 ;
        RECT 45.760 101.205 46.590 101.505 ;
        RECT 47.120 101.475 47.440 102.435 ;
        RECT 44.345 100.805 44.680 100.975 ;
        RECT 44.875 100.805 45.550 100.975 ;
        RECT 45.870 100.525 46.240 101.025 ;
        RECT 46.420 100.975 46.590 101.205 ;
        RECT 46.975 101.145 47.440 101.475 ;
        RECT 47.610 101.765 47.780 102.605 ;
        RECT 47.960 102.575 48.275 103.075 ;
        RECT 48.505 102.345 48.845 102.905 ;
        RECT 47.950 101.970 48.845 102.345 ;
        RECT 49.015 102.065 49.185 103.075 ;
        RECT 48.655 101.765 48.845 101.970 ;
        RECT 49.355 102.015 49.685 102.860 ;
        RECT 50.005 102.405 50.175 102.905 ;
        RECT 50.345 102.575 50.675 103.075 ;
        RECT 50.005 102.235 50.670 102.405 ;
        RECT 49.355 101.935 49.745 102.015 ;
        RECT 49.530 101.885 49.745 101.935 ;
        RECT 47.610 101.435 48.485 101.765 ;
        RECT 48.655 101.435 49.405 101.765 ;
        RECT 47.610 100.975 47.780 101.435 ;
        RECT 48.655 101.265 48.855 101.435 ;
        RECT 49.575 101.305 49.745 101.885 ;
        RECT 49.920 101.415 50.270 102.065 ;
        RECT 49.520 101.265 49.745 101.305 ;
        RECT 46.420 100.805 46.825 100.975 ;
        RECT 46.995 100.805 47.780 100.975 ;
        RECT 48.055 100.525 48.265 101.055 ;
        RECT 48.525 100.740 48.855 101.265 ;
        RECT 49.365 101.180 49.745 101.265 ;
        RECT 50.440 101.245 50.670 102.235 ;
        RECT 49.025 100.525 49.195 101.135 ;
        RECT 49.365 100.745 49.695 101.180 ;
        RECT 50.005 101.075 50.670 101.245 ;
        RECT 50.005 100.785 50.175 101.075 ;
        RECT 50.345 100.525 50.675 100.905 ;
        RECT 50.845 100.785 51.030 102.905 ;
        RECT 51.270 102.615 51.535 103.075 ;
        RECT 51.705 102.480 51.955 102.905 ;
        RECT 52.165 102.630 53.270 102.800 ;
        RECT 51.650 102.350 51.955 102.480 ;
        RECT 51.200 101.155 51.480 102.105 ;
        RECT 51.650 101.245 51.820 102.350 ;
        RECT 51.990 101.565 52.230 102.160 ;
        RECT 52.400 102.095 52.930 102.460 ;
        RECT 52.400 101.395 52.570 102.095 ;
        RECT 53.100 102.015 53.270 102.630 ;
        RECT 53.440 102.275 53.610 103.075 ;
        RECT 53.780 102.575 54.030 102.905 ;
        RECT 54.255 102.605 55.140 102.775 ;
        RECT 53.100 101.925 53.610 102.015 ;
        RECT 51.650 101.115 51.875 101.245 ;
        RECT 52.045 101.175 52.570 101.395 ;
        RECT 52.740 101.755 53.610 101.925 ;
        RECT 51.285 100.525 51.535 100.985 ;
        RECT 51.705 100.975 51.875 101.115 ;
        RECT 52.740 100.975 52.910 101.755 ;
        RECT 53.440 101.685 53.610 101.755 ;
        RECT 53.120 101.505 53.320 101.535 ;
        RECT 53.780 101.505 53.950 102.575 ;
        RECT 54.120 101.685 54.310 102.405 ;
        RECT 53.120 101.205 53.950 101.505 ;
        RECT 54.480 101.475 54.800 102.435 ;
        RECT 51.705 100.805 52.040 100.975 ;
        RECT 52.235 100.805 52.910 100.975 ;
        RECT 53.230 100.525 53.600 101.025 ;
        RECT 53.780 100.975 53.950 101.205 ;
        RECT 54.335 101.145 54.800 101.475 ;
        RECT 54.970 101.765 55.140 102.605 ;
        RECT 55.320 102.575 55.635 103.075 ;
        RECT 55.865 102.345 56.205 102.905 ;
        RECT 55.310 101.970 56.205 102.345 ;
        RECT 56.375 102.065 56.545 103.075 ;
        RECT 56.015 101.765 56.205 101.970 ;
        RECT 56.715 102.015 57.045 102.860 ;
        RECT 58.195 102.565 58.455 103.075 ;
        RECT 56.715 101.935 57.105 102.015 ;
        RECT 56.890 101.885 57.105 101.935 ;
        RECT 54.970 101.435 55.845 101.765 ;
        RECT 56.015 101.435 56.765 101.765 ;
        RECT 54.970 100.975 55.140 101.435 ;
        RECT 56.015 101.265 56.215 101.435 ;
        RECT 56.935 101.305 57.105 101.885 ;
        RECT 58.195 101.515 58.535 102.395 ;
        RECT 58.705 101.685 58.875 102.905 ;
        RECT 59.115 102.570 59.730 103.075 ;
        RECT 59.115 102.035 59.365 102.400 ;
        RECT 59.535 102.395 59.730 102.570 ;
        RECT 59.900 102.565 60.375 102.905 ;
        RECT 60.545 102.530 60.760 103.075 ;
        RECT 59.535 102.205 59.865 102.395 ;
        RECT 60.085 102.035 60.800 102.330 ;
        RECT 60.970 102.205 61.245 102.905 ;
        RECT 59.115 101.865 60.905 102.035 ;
        RECT 58.705 101.435 59.500 101.685 ;
        RECT 58.705 101.345 58.955 101.435 ;
        RECT 56.880 101.265 57.105 101.305 ;
        RECT 53.780 100.805 54.185 100.975 ;
        RECT 54.355 100.805 55.140 100.975 ;
        RECT 55.415 100.525 55.625 101.055 ;
        RECT 55.885 100.740 56.215 101.265 ;
        RECT 56.725 101.180 57.105 101.265 ;
        RECT 56.385 100.525 56.555 101.135 ;
        RECT 56.725 100.745 57.055 101.180 ;
        RECT 58.195 100.525 58.455 101.345 ;
        RECT 58.625 100.925 58.955 101.345 ;
        RECT 59.670 101.010 59.925 101.865 ;
        RECT 59.135 100.745 59.925 101.010 ;
        RECT 60.095 101.165 60.505 101.685 ;
        RECT 60.675 101.435 60.905 101.865 ;
        RECT 61.075 101.175 61.245 102.205 ;
        RECT 61.415 101.910 61.705 103.075 ;
        RECT 61.875 101.985 63.085 103.075 ;
        RECT 63.555 102.435 63.885 102.865 ;
        RECT 61.875 101.275 62.395 101.815 ;
        RECT 62.565 101.445 63.085 101.985 ;
        RECT 63.430 102.265 63.885 102.435 ;
        RECT 64.065 102.435 64.315 102.855 ;
        RECT 64.545 102.605 64.875 103.075 ;
        RECT 65.105 102.435 65.355 102.855 ;
        RECT 64.065 102.265 65.355 102.435 ;
        RECT 60.095 100.745 60.295 101.165 ;
        RECT 60.485 100.525 60.815 100.985 ;
        RECT 60.985 100.695 61.245 101.175 ;
        RECT 61.415 100.525 61.705 101.250 ;
        RECT 61.875 100.525 63.085 101.275 ;
        RECT 63.430 101.265 63.600 102.265 ;
        RECT 63.770 101.435 64.015 102.095 ;
        RECT 64.230 101.435 64.495 102.095 ;
        RECT 64.690 101.435 64.975 102.095 ;
        RECT 65.150 101.765 65.365 102.095 ;
        RECT 65.545 101.935 65.795 103.075 ;
        RECT 65.965 102.015 66.295 102.865 ;
        RECT 65.150 101.435 65.455 101.765 ;
        RECT 65.625 101.435 65.935 101.765 ;
        RECT 65.625 101.265 65.795 101.435 ;
        RECT 63.430 101.095 65.795 101.265 ;
        RECT 66.105 101.250 66.295 102.015 ;
        RECT 63.585 100.525 63.915 100.925 ;
        RECT 64.085 100.755 64.415 101.095 ;
        RECT 65.465 100.525 65.795 100.925 ;
        RECT 65.965 100.740 66.295 101.250 ;
        RECT 66.475 102.645 66.815 102.905 ;
        RECT 66.475 101.245 66.735 102.645 ;
        RECT 66.985 102.275 67.315 103.075 ;
        RECT 67.780 102.105 68.030 102.905 ;
        RECT 68.215 102.355 68.545 103.075 ;
        RECT 68.765 102.105 69.015 102.905 ;
        RECT 69.185 102.695 69.520 103.075 ;
        RECT 66.925 101.935 69.115 102.105 ;
        RECT 66.925 101.765 67.240 101.935 ;
        RECT 66.910 101.515 67.240 101.765 ;
        RECT 66.475 100.735 66.815 101.245 ;
        RECT 66.985 100.525 67.255 101.325 ;
        RECT 67.435 100.795 67.715 101.765 ;
        RECT 67.895 100.795 68.195 101.765 ;
        RECT 68.375 100.800 68.725 101.765 ;
        RECT 68.945 101.025 69.115 101.935 ;
        RECT 69.285 101.205 69.525 102.515 ;
        RECT 69.695 102.205 69.970 102.905 ;
        RECT 70.140 102.530 70.395 103.075 ;
        RECT 70.565 102.565 71.045 102.905 ;
        RECT 71.220 102.520 71.825 103.075 ;
        RECT 71.210 102.420 71.825 102.520 ;
        RECT 71.210 102.395 71.395 102.420 ;
        RECT 69.695 101.175 69.865 102.205 ;
        RECT 70.140 102.075 70.895 102.325 ;
        RECT 71.065 102.150 71.395 102.395 ;
        RECT 70.140 102.040 70.910 102.075 ;
        RECT 70.140 102.030 70.925 102.040 ;
        RECT 70.035 102.015 70.930 102.030 ;
        RECT 70.035 102.000 70.950 102.015 ;
        RECT 70.035 101.990 70.970 102.000 ;
        RECT 70.035 101.980 70.995 101.990 ;
        RECT 70.035 101.950 71.065 101.980 ;
        RECT 70.035 101.920 71.085 101.950 ;
        RECT 70.035 101.890 71.105 101.920 ;
        RECT 70.035 101.865 71.135 101.890 ;
        RECT 70.035 101.830 71.170 101.865 ;
        RECT 70.035 101.825 71.200 101.830 ;
        RECT 70.035 101.430 70.265 101.825 ;
        RECT 70.810 101.820 71.200 101.825 ;
        RECT 70.835 101.810 71.200 101.820 ;
        RECT 70.850 101.805 71.200 101.810 ;
        RECT 70.865 101.800 71.200 101.805 ;
        RECT 71.565 101.800 71.825 102.250 ;
        RECT 71.995 101.985 73.665 103.075 ;
        RECT 70.865 101.795 71.825 101.800 ;
        RECT 70.875 101.785 71.825 101.795 ;
        RECT 70.885 101.780 71.825 101.785 ;
        RECT 70.895 101.770 71.825 101.780 ;
        RECT 70.900 101.760 71.825 101.770 ;
        RECT 70.905 101.755 71.825 101.760 ;
        RECT 70.915 101.740 71.825 101.755 ;
        RECT 70.920 101.725 71.825 101.740 ;
        RECT 70.930 101.700 71.825 101.725 ;
        RECT 70.435 101.230 70.765 101.655 ;
        RECT 68.945 100.695 69.440 101.025 ;
        RECT 69.695 100.695 69.955 101.175 ;
        RECT 70.125 100.525 70.375 101.065 ;
        RECT 70.545 100.745 70.765 101.230 ;
        RECT 70.935 101.630 71.825 101.700 ;
        RECT 70.935 100.905 71.105 101.630 ;
        RECT 71.275 101.075 71.825 101.460 ;
        RECT 71.995 101.295 72.745 101.815 ;
        RECT 72.915 101.465 73.665 101.985 ;
        RECT 73.835 102.405 74.150 102.905 ;
        RECT 74.320 102.575 74.570 103.075 ;
        RECT 74.740 102.405 74.990 102.905 ;
        RECT 75.160 102.575 75.410 103.075 ;
        RECT 75.580 102.405 75.830 102.905 ;
        RECT 76.140 102.565 76.390 102.905 ;
        RECT 76.560 102.575 76.810 103.075 ;
        RECT 76.980 102.735 78.105 102.905 ;
        RECT 76.980 102.565 77.305 102.735 ;
        RECT 77.855 102.575 78.105 102.735 ;
        RECT 78.375 102.575 78.625 103.075 ;
        RECT 73.835 102.395 75.830 102.405 ;
        RECT 77.475 102.405 77.685 102.565 ;
        RECT 78.795 102.405 79.045 102.565 ;
        RECT 73.835 102.225 77.230 102.395 ;
        RECT 77.475 102.235 79.045 102.405 ;
        RECT 79.215 102.235 79.645 103.075 ;
        RECT 73.835 101.335 74.065 102.225 ;
        RECT 77.060 102.065 77.230 102.225 ;
        RECT 78.795 102.065 79.045 102.235 ;
        RECT 74.540 101.885 76.850 102.055 ;
        RECT 77.060 101.895 78.555 102.065 ;
        RECT 74.540 101.725 74.710 101.885 ;
        RECT 74.235 101.515 74.710 101.725 ;
        RECT 76.680 101.725 76.850 101.885 ;
        RECT 75.005 101.515 76.455 101.715 ;
        RECT 76.680 101.515 77.705 101.725 ;
        RECT 78.385 101.685 78.555 101.895 ;
        RECT 78.795 101.855 79.645 102.065 ;
        RECT 79.815 101.985 81.485 103.075 ;
        RECT 78.385 101.515 79.045 101.685 ;
        RECT 70.935 100.735 71.825 100.905 ;
        RECT 71.995 100.525 73.665 101.295 ;
        RECT 73.835 101.085 74.610 101.335 ;
        RECT 74.780 101.165 75.870 101.345 ;
        RECT 74.780 100.915 75.030 101.165 ;
        RECT 73.855 100.695 75.030 100.915 ;
        RECT 75.200 100.525 75.370 100.995 ;
        RECT 75.540 100.695 75.870 101.165 ;
        RECT 76.180 100.525 76.350 101.345 ;
        RECT 76.520 101.165 79.085 101.345 ;
        RECT 76.520 100.695 76.850 101.165 ;
        RECT 77.020 100.525 77.190 100.995 ;
        RECT 77.360 100.695 77.725 101.165 ;
        RECT 78.755 101.085 79.085 101.165 ;
        RECT 77.895 100.525 78.065 100.995 ;
        RECT 79.255 100.915 79.645 101.855 ;
        RECT 78.335 100.745 79.645 100.915 ;
        RECT 79.815 101.295 80.565 101.815 ;
        RECT 80.735 101.465 81.485 101.985 ;
        RECT 82.125 101.935 82.455 103.075 ;
        RECT 82.985 102.105 83.315 102.890 ;
        RECT 82.635 101.935 83.315 102.105 ;
        RECT 83.495 101.985 85.165 103.075 ;
        RECT 82.115 101.515 82.465 101.765 ;
        RECT 82.635 101.335 82.805 101.935 ;
        RECT 82.975 101.515 83.325 101.765 ;
        RECT 79.815 100.525 81.485 101.295 ;
        RECT 82.125 100.525 82.395 101.335 ;
        RECT 82.565 100.695 82.895 101.335 ;
        RECT 83.065 100.525 83.305 101.335 ;
        RECT 83.495 101.295 84.245 101.815 ;
        RECT 84.415 101.465 85.165 101.985 ;
        RECT 85.805 102.105 86.135 102.890 ;
        RECT 85.805 101.935 86.485 102.105 ;
        RECT 86.665 101.935 86.995 103.075 ;
        RECT 85.795 101.515 86.145 101.765 ;
        RECT 86.315 101.335 86.485 101.935 ;
        RECT 87.175 101.910 87.465 103.075 ;
        RECT 87.635 101.985 88.845 103.075 ;
        RECT 86.655 101.515 87.005 101.765 ;
        RECT 83.495 100.525 85.165 101.295 ;
        RECT 85.815 100.525 86.055 101.335 ;
        RECT 86.225 100.695 86.555 101.335 ;
        RECT 86.725 100.525 86.995 101.335 ;
        RECT 87.635 101.275 88.155 101.815 ;
        RECT 88.325 101.445 88.845 101.985 ;
        RECT 89.020 101.930 89.315 103.075 ;
        RECT 87.175 100.525 87.465 101.250 ;
        RECT 87.635 100.525 88.845 101.275 ;
        RECT 89.020 100.525 89.315 101.345 ;
        RECT 89.485 101.075 89.715 102.775 ;
        RECT 89.930 102.270 90.185 103.075 ;
        RECT 90.385 102.460 90.715 102.905 ;
        RECT 90.885 102.630 91.160 103.075 ;
        RECT 91.395 102.460 91.725 102.905 ;
        RECT 90.385 102.280 91.725 102.460 ;
        RECT 92.185 102.100 92.515 102.765 ;
        RECT 89.930 101.930 92.515 102.100 ;
        RECT 92.695 101.985 94.365 103.075 ;
        RECT 89.930 101.315 90.240 101.930 ;
        RECT 90.410 101.485 90.740 101.715 ;
        RECT 90.910 101.485 91.380 101.715 ;
        RECT 91.550 101.545 92.005 101.715 ;
        RECT 91.550 101.485 92.000 101.545 ;
        RECT 92.190 101.485 92.525 101.715 ;
        RECT 89.930 101.135 92.515 101.315 ;
        RECT 89.485 100.695 89.705 101.075 ;
        RECT 89.875 100.525 90.725 100.885 ;
        RECT 91.205 100.715 91.535 101.135 ;
        RECT 91.740 100.525 92.015 100.965 ;
        RECT 92.185 100.715 92.515 101.135 ;
        RECT 92.695 101.295 93.445 101.815 ;
        RECT 93.615 101.465 94.365 101.985 ;
        RECT 94.540 101.935 94.875 102.905 ;
        RECT 95.045 101.935 95.215 103.075 ;
        RECT 95.385 102.735 97.415 102.905 ;
        RECT 92.695 100.525 94.365 101.295 ;
        RECT 94.540 101.265 94.710 101.935 ;
        RECT 95.385 101.765 95.555 102.735 ;
        RECT 94.880 101.435 95.135 101.765 ;
        RECT 95.360 101.435 95.555 101.765 ;
        RECT 95.725 102.395 96.850 102.565 ;
        RECT 94.965 101.265 95.135 101.435 ;
        RECT 95.725 101.265 95.895 102.395 ;
        RECT 94.540 100.695 94.795 101.265 ;
        RECT 94.965 101.095 95.895 101.265 ;
        RECT 96.065 102.055 97.075 102.225 ;
        RECT 96.065 101.255 96.235 102.055 ;
        RECT 96.440 101.715 96.715 101.855 ;
        RECT 96.435 101.545 96.715 101.715 ;
        RECT 95.720 101.060 95.895 101.095 ;
        RECT 94.965 100.525 95.295 100.925 ;
        RECT 95.720 100.695 96.250 101.060 ;
        RECT 96.440 100.695 96.715 101.545 ;
        RECT 96.885 100.695 97.075 102.055 ;
        RECT 97.245 102.070 97.415 102.735 ;
        RECT 97.585 102.315 97.755 103.075 ;
        RECT 97.990 102.315 98.505 102.725 ;
        RECT 97.245 101.880 97.995 102.070 ;
        RECT 98.165 101.505 98.505 102.315 ;
        RECT 99.195 102.015 99.525 102.860 ;
        RECT 99.695 102.065 99.865 103.075 ;
        RECT 100.035 102.345 100.375 102.905 ;
        RECT 100.605 102.575 100.920 103.075 ;
        RECT 101.100 102.605 101.985 102.775 ;
        RECT 97.275 101.335 98.505 101.505 ;
        RECT 99.135 101.935 99.525 102.015 ;
        RECT 100.035 101.970 100.930 102.345 ;
        RECT 99.135 101.885 99.350 101.935 ;
        RECT 97.255 100.525 97.765 101.060 ;
        RECT 97.985 100.730 98.230 101.335 ;
        RECT 99.135 101.305 99.305 101.885 ;
        RECT 100.035 101.765 100.225 101.970 ;
        RECT 101.100 101.765 101.270 102.605 ;
        RECT 102.210 102.575 102.460 102.905 ;
        RECT 99.475 101.435 100.225 101.765 ;
        RECT 100.395 101.435 101.270 101.765 ;
        RECT 99.135 101.265 99.360 101.305 ;
        RECT 100.025 101.265 100.225 101.435 ;
        RECT 99.135 101.180 99.515 101.265 ;
        RECT 99.185 100.745 99.515 101.180 ;
        RECT 99.685 100.525 99.855 101.135 ;
        RECT 100.025 100.740 100.355 101.265 ;
        RECT 100.615 100.525 100.825 101.055 ;
        RECT 101.100 100.975 101.270 101.435 ;
        RECT 101.440 101.475 101.760 102.435 ;
        RECT 101.930 101.685 102.120 102.405 ;
        RECT 102.290 101.505 102.460 102.575 ;
        RECT 102.630 102.275 102.800 103.075 ;
        RECT 102.970 102.630 104.075 102.800 ;
        RECT 102.970 102.015 103.140 102.630 ;
        RECT 104.285 102.480 104.535 102.905 ;
        RECT 104.705 102.615 104.970 103.075 ;
        RECT 103.310 102.095 103.840 102.460 ;
        RECT 104.285 102.350 104.590 102.480 ;
        RECT 102.630 101.925 103.140 102.015 ;
        RECT 102.630 101.755 103.500 101.925 ;
        RECT 102.630 101.685 102.800 101.755 ;
        RECT 102.920 101.505 103.120 101.535 ;
        RECT 101.440 101.145 101.905 101.475 ;
        RECT 102.290 101.205 103.120 101.505 ;
        RECT 102.290 100.975 102.460 101.205 ;
        RECT 101.100 100.805 101.885 100.975 ;
        RECT 102.055 100.805 102.460 100.975 ;
        RECT 102.640 100.525 103.010 101.025 ;
        RECT 103.330 100.975 103.500 101.755 ;
        RECT 103.670 101.395 103.840 102.095 ;
        RECT 104.010 101.565 104.250 102.160 ;
        RECT 103.670 101.175 104.195 101.395 ;
        RECT 104.420 101.245 104.590 102.350 ;
        RECT 104.365 101.115 104.590 101.245 ;
        RECT 104.760 101.155 105.040 102.105 ;
        RECT 104.365 100.975 104.535 101.115 ;
        RECT 103.330 100.805 104.005 100.975 ;
        RECT 104.200 100.805 104.535 100.975 ;
        RECT 104.705 100.525 104.955 100.985 ;
        RECT 105.210 100.785 105.395 102.905 ;
        RECT 105.565 102.575 105.895 103.075 ;
        RECT 106.065 102.405 106.235 102.905 ;
        RECT 105.570 102.235 106.235 102.405 ;
        RECT 105.570 101.245 105.800 102.235 ;
        RECT 105.970 101.415 106.320 102.065 ;
        RECT 106.955 102.000 107.225 102.905 ;
        RECT 107.395 102.315 107.725 103.075 ;
        RECT 107.905 102.145 108.075 102.905 ;
        RECT 105.570 101.075 106.235 101.245 ;
        RECT 105.565 100.525 105.895 100.905 ;
        RECT 106.065 100.785 106.235 101.075 ;
        RECT 106.955 101.200 107.125 102.000 ;
        RECT 107.410 101.975 108.075 102.145 ;
        RECT 109.255 102.355 109.715 102.905 ;
        RECT 109.905 102.355 110.235 103.075 ;
        RECT 107.410 101.830 107.580 101.975 ;
        RECT 107.295 101.500 107.580 101.830 ;
        RECT 107.410 101.245 107.580 101.500 ;
        RECT 107.815 101.425 108.145 101.795 ;
        RECT 106.955 100.695 107.215 101.200 ;
        RECT 107.410 101.075 108.075 101.245 ;
        RECT 107.395 100.525 107.725 100.905 ;
        RECT 107.905 100.695 108.075 101.075 ;
        RECT 109.255 100.985 109.505 102.355 ;
        RECT 110.435 102.185 110.735 102.735 ;
        RECT 110.905 102.405 111.185 103.075 ;
        RECT 109.795 102.015 110.735 102.185 ;
        RECT 109.795 101.765 109.965 102.015 ;
        RECT 111.105 101.765 111.370 102.125 ;
        RECT 111.555 101.985 112.765 103.075 ;
        RECT 109.675 101.435 109.965 101.765 ;
        RECT 110.135 101.515 110.475 101.765 ;
        RECT 110.695 101.515 111.370 101.765 ;
        RECT 109.795 101.345 109.965 101.435 ;
        RECT 109.795 101.155 111.185 101.345 ;
        RECT 109.255 100.695 109.815 100.985 ;
        RECT 109.985 100.525 110.235 100.985 ;
        RECT 110.855 100.795 111.185 101.155 ;
        RECT 111.555 101.275 112.075 101.815 ;
        RECT 112.245 101.445 112.765 101.985 ;
        RECT 112.935 101.910 113.225 103.075 ;
        RECT 113.395 101.985 114.605 103.075 ;
        RECT 114.865 102.405 115.035 102.905 ;
        RECT 115.205 102.575 115.535 103.075 ;
        RECT 114.865 102.235 115.530 102.405 ;
        RECT 113.395 101.275 113.915 101.815 ;
        RECT 114.085 101.445 114.605 101.985 ;
        RECT 114.780 101.415 115.130 102.065 ;
        RECT 111.555 100.525 112.765 101.275 ;
        RECT 112.935 100.525 113.225 101.250 ;
        RECT 113.395 100.525 114.605 101.275 ;
        RECT 115.300 101.245 115.530 102.235 ;
        RECT 114.865 101.075 115.530 101.245 ;
        RECT 114.865 100.785 115.035 101.075 ;
        RECT 115.205 100.525 115.535 100.905 ;
        RECT 115.705 100.785 115.890 102.905 ;
        RECT 116.130 102.615 116.395 103.075 ;
        RECT 116.565 102.480 116.815 102.905 ;
        RECT 117.025 102.630 118.130 102.800 ;
        RECT 116.510 102.350 116.815 102.480 ;
        RECT 116.060 101.155 116.340 102.105 ;
        RECT 116.510 101.245 116.680 102.350 ;
        RECT 116.850 101.565 117.090 102.160 ;
        RECT 117.260 102.095 117.790 102.460 ;
        RECT 117.260 101.395 117.430 102.095 ;
        RECT 117.960 102.015 118.130 102.630 ;
        RECT 118.300 102.275 118.470 103.075 ;
        RECT 118.640 102.575 118.890 102.905 ;
        RECT 119.115 102.605 120.000 102.775 ;
        RECT 117.960 101.925 118.470 102.015 ;
        RECT 116.510 101.115 116.735 101.245 ;
        RECT 116.905 101.175 117.430 101.395 ;
        RECT 117.600 101.755 118.470 101.925 ;
        RECT 116.145 100.525 116.395 100.985 ;
        RECT 116.565 100.975 116.735 101.115 ;
        RECT 117.600 100.975 117.770 101.755 ;
        RECT 118.300 101.685 118.470 101.755 ;
        RECT 117.980 101.505 118.180 101.535 ;
        RECT 118.640 101.505 118.810 102.575 ;
        RECT 118.980 101.685 119.170 102.405 ;
        RECT 117.980 101.205 118.810 101.505 ;
        RECT 119.340 101.475 119.660 102.435 ;
        RECT 116.565 100.805 116.900 100.975 ;
        RECT 117.095 100.805 117.770 100.975 ;
        RECT 118.090 100.525 118.460 101.025 ;
        RECT 118.640 100.975 118.810 101.205 ;
        RECT 119.195 101.145 119.660 101.475 ;
        RECT 119.830 101.765 120.000 102.605 ;
        RECT 120.180 102.575 120.495 103.075 ;
        RECT 120.725 102.345 121.065 102.905 ;
        RECT 120.170 101.970 121.065 102.345 ;
        RECT 121.235 102.065 121.405 103.075 ;
        RECT 120.875 101.765 121.065 101.970 ;
        RECT 121.575 102.015 121.905 102.860 ;
        RECT 121.575 101.935 121.965 102.015 ;
        RECT 121.750 101.885 121.965 101.935 ;
        RECT 119.830 101.435 120.705 101.765 ;
        RECT 120.875 101.435 121.625 101.765 ;
        RECT 119.830 100.975 120.000 101.435 ;
        RECT 120.875 101.265 121.075 101.435 ;
        RECT 121.795 101.305 121.965 101.885 ;
        RECT 121.740 101.265 121.965 101.305 ;
        RECT 118.640 100.805 119.045 100.975 ;
        RECT 119.215 100.805 120.000 100.975 ;
        RECT 120.275 100.525 120.485 101.055 ;
        RECT 120.745 100.740 121.075 101.265 ;
        RECT 121.585 101.180 121.965 101.265 ;
        RECT 121.245 100.525 121.415 101.135 ;
        RECT 121.585 100.745 121.915 101.180 ;
        RECT 123.065 100.705 123.325 102.895 ;
        RECT 123.495 102.345 123.835 103.075 ;
        RECT 124.015 102.165 124.285 102.895 ;
        RECT 123.515 101.945 124.285 102.165 ;
        RECT 124.465 102.185 124.695 102.895 ;
        RECT 124.865 102.365 125.195 103.075 ;
        RECT 125.365 102.185 125.625 102.895 ;
        RECT 126.285 102.355 126.615 103.075 ;
        RECT 124.465 101.945 125.625 102.185 ;
        RECT 123.515 101.275 123.805 101.945 ;
        RECT 123.985 101.455 124.450 101.765 ;
        RECT 124.630 101.455 125.155 101.765 ;
        RECT 123.515 101.075 124.745 101.275 ;
        RECT 123.585 100.525 124.255 100.895 ;
        RECT 124.435 100.705 124.745 101.075 ;
        RECT 124.925 100.815 125.155 101.455 ;
        RECT 125.335 101.435 125.635 101.765 ;
        RECT 126.275 101.715 126.505 102.055 ;
        RECT 126.795 101.715 127.010 102.830 ;
        RECT 127.205 102.130 127.535 102.905 ;
        RECT 127.705 102.300 128.415 103.075 ;
        RECT 127.205 101.915 128.355 102.130 ;
        RECT 126.275 101.515 126.605 101.715 ;
        RECT 126.795 101.535 127.245 101.715 ;
        RECT 126.915 101.515 127.245 101.535 ;
        RECT 127.415 101.515 127.885 101.745 ;
        RECT 128.070 101.345 128.355 101.915 ;
        RECT 128.585 101.470 128.865 102.905 ;
        RECT 129.035 101.985 132.545 103.075 ;
        RECT 132.715 102.565 133.015 103.075 ;
        RECT 133.185 102.395 133.515 102.905 ;
        RECT 133.685 102.565 134.315 103.075 ;
        RECT 134.895 102.565 135.275 102.735 ;
        RECT 135.445 102.565 135.745 103.075 ;
        RECT 135.105 102.395 135.275 102.565 ;
        RECT 125.335 100.525 125.625 101.255 ;
        RECT 126.275 101.155 127.455 101.345 ;
        RECT 126.275 100.695 126.615 101.155 ;
        RECT 127.125 101.075 127.455 101.155 ;
        RECT 127.645 101.155 128.355 101.345 ;
        RECT 127.645 101.015 127.945 101.155 ;
        RECT 127.630 101.005 127.945 101.015 ;
        RECT 127.620 100.995 127.945 101.005 ;
        RECT 127.610 100.990 127.945 100.995 ;
        RECT 126.785 100.525 126.955 100.985 ;
        RECT 127.605 100.980 127.945 100.990 ;
        RECT 127.600 100.975 127.945 100.980 ;
        RECT 127.595 100.965 127.945 100.975 ;
        RECT 127.590 100.960 127.945 100.965 ;
        RECT 127.585 100.695 127.945 100.960 ;
        RECT 128.185 100.525 128.355 100.985 ;
        RECT 128.525 100.695 128.865 101.470 ;
        RECT 129.035 101.295 130.685 101.815 ;
        RECT 130.855 101.465 132.545 101.985 ;
        RECT 132.715 102.225 134.935 102.395 ;
        RECT 129.035 100.525 132.545 101.295 ;
        RECT 132.715 101.265 132.885 102.225 ;
        RECT 133.055 101.885 134.595 102.055 ;
        RECT 133.055 101.435 133.300 101.885 ;
        RECT 133.560 101.515 134.255 101.715 ;
        RECT 134.425 101.685 134.595 101.885 ;
        RECT 134.765 102.025 134.935 102.225 ;
        RECT 135.105 102.195 135.765 102.395 ;
        RECT 134.765 101.855 135.425 102.025 ;
        RECT 134.425 101.515 135.025 101.685 ;
        RECT 135.255 101.435 135.425 101.855 ;
        RECT 132.715 100.720 133.180 101.265 ;
        RECT 133.685 100.525 133.855 101.345 ;
        RECT 134.025 101.265 134.935 101.345 ;
        RECT 135.595 101.265 135.765 102.195 ;
        RECT 135.935 101.985 138.525 103.075 ;
        RECT 134.025 101.175 135.275 101.265 ;
        RECT 134.025 100.695 134.355 101.175 ;
        RECT 134.765 101.095 135.275 101.175 ;
        RECT 134.525 100.525 134.875 100.915 ;
        RECT 135.045 100.695 135.275 101.095 ;
        RECT 135.445 100.785 135.765 101.265 ;
        RECT 135.935 101.295 137.145 101.815 ;
        RECT 137.315 101.465 138.525 101.985 ;
        RECT 138.695 101.910 138.985 103.075 ;
        RECT 139.155 102.565 139.455 103.075 ;
        RECT 139.625 102.395 139.955 102.905 ;
        RECT 140.125 102.565 140.755 103.075 ;
        RECT 141.335 102.565 141.715 102.735 ;
        RECT 141.885 102.565 142.185 103.075 ;
        RECT 141.545 102.395 141.715 102.565 ;
        RECT 139.155 102.225 141.375 102.395 ;
        RECT 135.935 100.525 138.525 101.295 ;
        RECT 139.155 101.265 139.325 102.225 ;
        RECT 139.495 101.885 141.035 102.055 ;
        RECT 139.495 101.435 139.740 101.885 ;
        RECT 140.000 101.515 140.695 101.715 ;
        RECT 140.865 101.685 141.035 101.885 ;
        RECT 141.205 102.025 141.375 102.225 ;
        RECT 141.545 102.195 142.205 102.395 ;
        RECT 141.205 101.855 141.865 102.025 ;
        RECT 140.865 101.515 141.465 101.685 ;
        RECT 141.695 101.435 141.865 101.855 ;
        RECT 138.695 100.525 138.985 101.250 ;
        RECT 139.155 100.720 139.620 101.265 ;
        RECT 140.125 100.525 140.295 101.345 ;
        RECT 140.465 101.265 141.375 101.345 ;
        RECT 142.035 101.265 142.205 102.195 ;
        RECT 142.895 102.015 143.225 102.860 ;
        RECT 143.395 102.065 143.565 103.075 ;
        RECT 143.735 102.345 144.075 102.905 ;
        RECT 144.305 102.575 144.620 103.075 ;
        RECT 144.800 102.605 145.685 102.775 ;
        RECT 140.465 101.175 141.715 101.265 ;
        RECT 140.465 100.695 140.795 101.175 ;
        RECT 141.205 101.095 141.715 101.175 ;
        RECT 140.965 100.525 141.315 100.915 ;
        RECT 141.485 100.695 141.715 101.095 ;
        RECT 141.885 100.785 142.205 101.265 ;
        RECT 142.835 101.935 143.225 102.015 ;
        RECT 143.735 101.970 144.630 102.345 ;
        RECT 142.835 101.885 143.050 101.935 ;
        RECT 142.835 101.305 143.005 101.885 ;
        RECT 143.735 101.765 143.925 101.970 ;
        RECT 144.800 101.765 144.970 102.605 ;
        RECT 145.910 102.575 146.160 102.905 ;
        RECT 143.175 101.435 143.925 101.765 ;
        RECT 144.095 101.435 144.970 101.765 ;
        RECT 142.835 101.265 143.060 101.305 ;
        RECT 143.725 101.265 143.925 101.435 ;
        RECT 142.835 101.180 143.215 101.265 ;
        RECT 142.885 100.745 143.215 101.180 ;
        RECT 143.385 100.525 143.555 101.135 ;
        RECT 143.725 100.740 144.055 101.265 ;
        RECT 144.315 100.525 144.525 101.055 ;
        RECT 144.800 100.975 144.970 101.435 ;
        RECT 145.140 101.475 145.460 102.435 ;
        RECT 145.630 101.685 145.820 102.405 ;
        RECT 145.990 101.505 146.160 102.575 ;
        RECT 146.330 102.275 146.500 103.075 ;
        RECT 146.670 102.630 147.775 102.800 ;
        RECT 146.670 102.015 146.840 102.630 ;
        RECT 147.985 102.480 148.235 102.905 ;
        RECT 148.405 102.615 148.670 103.075 ;
        RECT 147.010 102.095 147.540 102.460 ;
        RECT 147.985 102.350 148.290 102.480 ;
        RECT 146.330 101.925 146.840 102.015 ;
        RECT 146.330 101.755 147.200 101.925 ;
        RECT 146.330 101.685 146.500 101.755 ;
        RECT 146.620 101.505 146.820 101.535 ;
        RECT 145.140 101.145 145.605 101.475 ;
        RECT 145.990 101.205 146.820 101.505 ;
        RECT 145.990 100.975 146.160 101.205 ;
        RECT 144.800 100.805 145.585 100.975 ;
        RECT 145.755 100.805 146.160 100.975 ;
        RECT 146.340 100.525 146.710 101.025 ;
        RECT 147.030 100.975 147.200 101.755 ;
        RECT 147.370 101.395 147.540 102.095 ;
        RECT 147.710 101.565 147.950 102.160 ;
        RECT 147.370 101.175 147.895 101.395 ;
        RECT 148.120 101.245 148.290 102.350 ;
        RECT 148.065 101.115 148.290 101.245 ;
        RECT 148.460 101.155 148.740 102.105 ;
        RECT 148.065 100.975 148.235 101.115 ;
        RECT 147.030 100.805 147.705 100.975 ;
        RECT 147.900 100.805 148.235 100.975 ;
        RECT 148.405 100.525 148.655 100.985 ;
        RECT 148.910 100.785 149.095 102.905 ;
        RECT 149.265 102.575 149.595 103.075 ;
        RECT 149.765 102.405 149.935 102.905 ;
        RECT 150.195 102.640 155.540 103.075 ;
        RECT 149.270 102.235 149.935 102.405 ;
        RECT 149.270 101.245 149.500 102.235 ;
        RECT 149.670 101.415 150.020 102.065 ;
        RECT 149.270 101.075 149.935 101.245 ;
        RECT 149.265 100.525 149.595 100.905 ;
        RECT 149.765 100.785 149.935 101.075 ;
        RECT 151.780 101.070 152.120 101.900 ;
        RECT 153.600 101.390 153.950 102.640 ;
        RECT 155.715 101.985 156.925 103.075 ;
        RECT 155.715 101.445 156.235 101.985 ;
        RECT 156.405 101.275 156.925 101.815 ;
        RECT 150.195 100.525 155.540 101.070 ;
        RECT 155.715 100.525 156.925 101.275 ;
        RECT 22.690 100.355 157.010 100.525 ;
        RECT 22.775 99.605 23.985 100.355 ;
        RECT 22.775 99.065 23.295 99.605 ;
        RECT 24.155 99.585 25.825 100.355 ;
        RECT 25.995 99.615 26.380 100.185 ;
        RECT 26.550 99.895 26.875 100.355 ;
        RECT 27.395 99.725 27.675 100.185 ;
        RECT 23.465 98.895 23.985 99.435 ;
        RECT 24.155 99.065 24.905 99.585 ;
        RECT 25.075 98.895 25.825 99.415 ;
        RECT 22.775 97.805 23.985 98.895 ;
        RECT 24.155 97.805 25.825 98.895 ;
        RECT 25.995 98.945 26.275 99.615 ;
        RECT 26.550 99.555 27.675 99.725 ;
        RECT 26.550 99.445 27.000 99.555 ;
        RECT 26.445 99.115 27.000 99.445 ;
        RECT 27.865 99.385 28.265 100.185 ;
        RECT 28.665 99.895 28.935 100.355 ;
        RECT 29.105 99.725 29.390 100.185 ;
        RECT 25.995 97.975 26.380 98.945 ;
        RECT 26.550 98.655 27.000 99.115 ;
        RECT 27.170 98.825 28.265 99.385 ;
        RECT 26.550 98.435 27.675 98.655 ;
        RECT 26.550 97.805 26.875 98.265 ;
        RECT 27.395 97.975 27.675 98.435 ;
        RECT 27.865 97.975 28.265 98.825 ;
        RECT 28.435 99.555 29.390 99.725 ;
        RECT 29.880 99.575 30.380 100.185 ;
        RECT 28.435 98.655 28.645 99.555 ;
        RECT 28.815 98.825 29.505 99.385 ;
        RECT 29.675 99.115 30.025 99.365 ;
        RECT 30.210 98.945 30.380 99.575 ;
        RECT 31.010 99.705 31.340 100.185 ;
        RECT 31.510 99.895 31.735 100.355 ;
        RECT 31.905 99.705 32.235 100.185 ;
        RECT 31.010 99.535 32.235 99.705 ;
        RECT 32.425 99.555 32.675 100.355 ;
        RECT 32.845 99.555 33.185 100.185 ;
        RECT 33.375 99.625 33.665 100.355 ;
        RECT 30.550 99.165 30.880 99.365 ;
        RECT 31.050 99.165 31.380 99.365 ;
        RECT 31.550 99.165 31.970 99.365 ;
        RECT 32.145 99.195 32.840 99.365 ;
        RECT 32.145 98.945 32.315 99.195 ;
        RECT 33.010 98.995 33.185 99.555 ;
        RECT 33.365 99.115 33.665 99.445 ;
        RECT 33.845 99.425 34.075 100.065 ;
        RECT 34.255 99.805 34.565 100.175 ;
        RECT 34.745 99.985 35.415 100.355 ;
        RECT 34.255 99.605 35.485 99.805 ;
        RECT 33.845 99.115 34.370 99.425 ;
        RECT 34.550 99.115 35.015 99.425 ;
        RECT 32.955 98.945 33.185 98.995 ;
        RECT 29.880 98.775 32.315 98.945 ;
        RECT 28.435 98.435 29.390 98.655 ;
        RECT 28.665 97.805 28.935 98.265 ;
        RECT 29.105 97.975 29.390 98.435 ;
        RECT 29.880 97.975 30.210 98.775 ;
        RECT 30.380 97.805 30.710 98.605 ;
        RECT 31.010 97.975 31.340 98.775 ;
        RECT 31.985 97.805 32.235 98.605 ;
        RECT 32.505 97.805 32.675 98.945 ;
        RECT 32.845 97.975 33.185 98.945 ;
        RECT 35.195 98.935 35.485 99.605 ;
        RECT 33.375 98.695 34.535 98.935 ;
        RECT 33.375 97.985 33.635 98.695 ;
        RECT 33.805 97.805 34.135 98.515 ;
        RECT 34.305 97.985 34.535 98.695 ;
        RECT 34.715 98.715 35.485 98.935 ;
        RECT 34.715 97.985 34.985 98.715 ;
        RECT 35.165 97.805 35.505 98.535 ;
        RECT 35.675 97.985 35.935 100.175 ;
        RECT 37.070 99.615 37.685 100.185 ;
        RECT 37.855 99.845 38.070 100.355 ;
        RECT 38.300 99.845 38.580 100.175 ;
        RECT 38.760 99.845 39.000 100.355 ;
        RECT 37.070 98.595 37.385 99.615 ;
        RECT 37.555 98.945 37.725 99.445 ;
        RECT 37.975 99.115 38.240 99.675 ;
        RECT 38.410 98.945 38.580 99.845 ;
        RECT 39.425 99.805 39.595 100.095 ;
        RECT 39.765 99.975 40.095 100.355 ;
        RECT 38.750 99.115 39.105 99.675 ;
        RECT 39.425 99.635 40.090 99.805 ;
        RECT 37.555 98.775 38.980 98.945 ;
        RECT 39.340 98.815 39.690 99.465 ;
        RECT 37.070 97.975 37.605 98.595 ;
        RECT 37.775 97.805 38.105 98.605 ;
        RECT 38.590 98.600 38.980 98.775 ;
        RECT 39.860 98.645 40.090 99.635 ;
        RECT 39.425 98.475 40.090 98.645 ;
        RECT 39.425 97.975 39.595 98.475 ;
        RECT 39.765 97.805 40.095 98.305 ;
        RECT 40.265 97.975 40.450 100.095 ;
        RECT 40.705 99.895 40.955 100.355 ;
        RECT 41.125 99.905 41.460 100.075 ;
        RECT 41.655 99.905 42.330 100.075 ;
        RECT 41.125 99.765 41.295 99.905 ;
        RECT 40.620 98.775 40.900 99.725 ;
        RECT 41.070 99.635 41.295 99.765 ;
        RECT 41.070 98.530 41.240 99.635 ;
        RECT 41.465 99.485 41.990 99.705 ;
        RECT 41.410 98.720 41.650 99.315 ;
        RECT 41.820 98.785 41.990 99.485 ;
        RECT 42.160 99.125 42.330 99.905 ;
        RECT 42.650 99.855 43.020 100.355 ;
        RECT 43.200 99.905 43.605 100.075 ;
        RECT 43.775 99.905 44.560 100.075 ;
        RECT 43.200 99.675 43.370 99.905 ;
        RECT 42.540 99.375 43.370 99.675 ;
        RECT 43.755 99.405 44.220 99.735 ;
        RECT 42.540 99.345 42.740 99.375 ;
        RECT 42.860 99.125 43.030 99.195 ;
        RECT 42.160 98.955 43.030 99.125 ;
        RECT 42.520 98.865 43.030 98.955 ;
        RECT 41.070 98.400 41.375 98.530 ;
        RECT 41.820 98.420 42.350 98.785 ;
        RECT 40.690 97.805 40.955 98.265 ;
        RECT 41.125 97.975 41.375 98.400 ;
        RECT 42.520 98.250 42.690 98.865 ;
        RECT 41.585 98.080 42.690 98.250 ;
        RECT 42.860 97.805 43.030 98.605 ;
        RECT 43.200 98.305 43.370 99.375 ;
        RECT 43.540 98.475 43.730 99.195 ;
        RECT 43.900 98.445 44.220 99.405 ;
        RECT 44.390 99.445 44.560 99.905 ;
        RECT 44.835 99.825 45.045 100.355 ;
        RECT 45.305 99.615 45.635 100.140 ;
        RECT 45.805 99.745 45.975 100.355 ;
        RECT 46.145 99.700 46.475 100.135 ;
        RECT 46.145 99.615 46.525 99.700 ;
        RECT 45.435 99.445 45.635 99.615 ;
        RECT 46.300 99.575 46.525 99.615 ;
        RECT 44.390 99.115 45.265 99.445 ;
        RECT 45.435 99.115 46.185 99.445 ;
        RECT 43.200 97.975 43.450 98.305 ;
        RECT 44.390 98.275 44.560 99.115 ;
        RECT 45.435 98.910 45.625 99.115 ;
        RECT 46.355 98.995 46.525 99.575 ;
        RECT 46.695 99.585 48.365 100.355 ;
        RECT 48.535 99.630 48.825 100.355 ;
        RECT 48.995 99.810 54.340 100.355 ;
        RECT 46.695 99.065 47.445 99.585 ;
        RECT 46.310 98.945 46.525 98.995 ;
        RECT 44.730 98.535 45.625 98.910 ;
        RECT 46.135 98.865 46.525 98.945 ;
        RECT 47.615 98.895 48.365 99.415 ;
        RECT 50.580 98.980 50.920 99.810 ;
        RECT 54.515 99.585 57.105 100.355 ;
        RECT 57.555 99.725 57.935 100.175 ;
        RECT 43.675 98.105 44.560 98.275 ;
        RECT 44.740 97.805 45.055 98.305 ;
        RECT 45.285 97.975 45.625 98.535 ;
        RECT 45.795 97.805 45.965 98.815 ;
        RECT 46.135 98.020 46.465 98.865 ;
        RECT 46.695 97.805 48.365 98.895 ;
        RECT 48.535 97.805 48.825 98.970 ;
        RECT 52.400 98.240 52.750 99.490 ;
        RECT 54.515 99.065 55.725 99.585 ;
        RECT 55.895 98.895 57.105 99.415 ;
        RECT 48.995 97.805 54.340 98.240 ;
        RECT 54.515 97.805 57.105 98.895 ;
        RECT 57.295 98.775 57.525 99.465 ;
        RECT 57.705 99.275 57.935 99.725 ;
        RECT 58.115 99.575 58.345 100.355 ;
        RECT 58.525 99.645 58.955 100.175 ;
        RECT 58.525 99.395 58.770 99.645 ;
        RECT 59.135 99.445 59.345 100.065 ;
        RECT 59.515 99.625 59.845 100.355 ;
        RECT 57.705 98.595 58.045 99.275 ;
        RECT 57.285 98.395 58.045 98.595 ;
        RECT 58.235 99.095 58.770 99.395 ;
        RECT 58.950 99.095 59.345 99.445 ;
        RECT 59.540 99.095 59.830 99.445 ;
        RECT 60.035 99.410 60.375 100.185 ;
        RECT 60.545 99.895 60.715 100.355 ;
        RECT 60.955 99.920 61.315 100.185 ;
        RECT 60.955 99.915 61.310 99.920 ;
        RECT 60.955 99.905 61.305 99.915 ;
        RECT 60.955 99.900 61.300 99.905 ;
        RECT 60.955 99.890 61.295 99.900 ;
        RECT 61.945 99.895 62.115 100.355 ;
        RECT 60.955 99.885 61.290 99.890 ;
        RECT 60.955 99.875 61.280 99.885 ;
        RECT 60.955 99.865 61.270 99.875 ;
        RECT 60.955 99.725 61.255 99.865 ;
        RECT 60.545 99.535 61.255 99.725 ;
        RECT 61.445 99.725 61.775 99.805 ;
        RECT 62.285 99.725 62.625 100.185 ;
        RECT 61.445 99.535 62.625 99.725 ;
        RECT 62.795 99.895 63.355 100.185 ;
        RECT 63.525 99.895 63.775 100.355 ;
        RECT 57.285 98.005 57.545 98.395 ;
        RECT 57.715 97.805 58.045 98.215 ;
        RECT 58.235 97.985 58.565 99.095 ;
        RECT 58.735 98.715 59.775 98.915 ;
        RECT 58.735 97.985 58.925 98.715 ;
        RECT 59.095 97.805 59.425 98.535 ;
        RECT 59.605 97.985 59.775 98.715 ;
        RECT 60.035 97.975 60.315 99.410 ;
        RECT 60.545 98.965 60.830 99.535 ;
        RECT 61.015 99.135 61.485 99.365 ;
        RECT 61.655 99.345 61.985 99.365 ;
        RECT 61.655 99.165 62.105 99.345 ;
        RECT 62.295 99.165 62.625 99.365 ;
        RECT 60.545 98.750 61.695 98.965 ;
        RECT 60.485 97.805 61.195 98.580 ;
        RECT 61.365 97.975 61.695 98.750 ;
        RECT 61.890 98.050 62.105 99.165 ;
        RECT 62.395 98.825 62.625 99.165 ;
        RECT 62.795 98.525 63.045 99.895 ;
        RECT 64.395 99.725 64.725 100.085 ;
        RECT 63.335 99.535 64.725 99.725 ;
        RECT 65.095 99.535 65.355 100.355 ;
        RECT 65.525 99.535 65.855 99.955 ;
        RECT 66.035 99.870 66.825 100.135 ;
        RECT 63.335 99.445 63.505 99.535 ;
        RECT 63.215 99.115 63.505 99.445 ;
        RECT 65.605 99.445 65.855 99.535 ;
        RECT 63.675 99.115 64.015 99.365 ;
        RECT 64.235 99.115 64.910 99.365 ;
        RECT 63.335 98.865 63.505 99.115 ;
        RECT 63.335 98.695 64.275 98.865 ;
        RECT 64.645 98.755 64.910 99.115 ;
        RECT 62.285 97.805 62.615 98.525 ;
        RECT 62.795 97.975 63.255 98.525 ;
        RECT 63.445 97.805 63.775 98.525 ;
        RECT 63.975 98.145 64.275 98.695 ;
        RECT 65.095 98.485 65.435 99.365 ;
        RECT 65.605 99.195 66.400 99.445 ;
        RECT 64.445 97.805 64.725 98.475 ;
        RECT 65.095 97.805 65.355 98.315 ;
        RECT 65.605 97.975 65.775 99.195 ;
        RECT 66.570 99.015 66.825 99.870 ;
        RECT 66.995 99.715 67.195 100.135 ;
        RECT 67.385 99.895 67.715 100.355 ;
        RECT 66.995 99.195 67.405 99.715 ;
        RECT 67.885 99.705 68.145 100.185 ;
        RECT 68.315 99.810 73.660 100.355 ;
        RECT 67.575 99.015 67.805 99.445 ;
        RECT 66.015 98.845 67.805 99.015 ;
        RECT 66.015 98.480 66.265 98.845 ;
        RECT 66.435 98.485 66.765 98.675 ;
        RECT 66.985 98.550 67.700 98.845 ;
        RECT 67.975 98.675 68.145 99.705 ;
        RECT 69.900 98.980 70.240 99.810 ;
        RECT 74.295 99.630 74.585 100.355 ;
        RECT 74.840 99.965 76.850 100.185 ;
        RECT 74.755 99.535 76.430 99.795 ;
        RECT 76.600 99.715 76.850 99.965 ;
        RECT 77.020 99.885 77.190 100.355 ;
        RECT 77.360 99.715 77.690 100.185 ;
        RECT 77.860 99.885 78.030 100.355 ;
        RECT 78.200 99.715 78.530 100.185 ;
        RECT 76.600 99.535 78.530 99.715 ;
        RECT 78.705 99.535 78.980 100.355 ;
        RECT 79.150 99.715 79.480 100.185 ;
        RECT 79.650 99.885 79.820 100.355 ;
        RECT 79.990 99.715 80.320 100.185 ;
        RECT 80.490 99.885 80.660 100.355 ;
        RECT 80.830 99.715 81.160 100.185 ;
        RECT 81.330 99.885 81.500 100.355 ;
        RECT 81.670 99.715 82.000 100.185 ;
        RECT 82.170 99.885 82.440 100.355 ;
        RECT 82.630 99.965 84.640 100.135 ;
        RECT 79.150 99.705 82.100 99.715 ;
        RECT 82.630 99.705 82.880 99.965 ;
        RECT 79.150 99.535 82.880 99.705 ;
        RECT 83.050 99.535 84.705 99.795 ;
        RECT 84.885 99.745 85.215 100.165 ;
        RECT 85.385 99.915 85.660 100.355 ;
        RECT 85.865 99.745 86.195 100.165 ;
        RECT 86.675 99.995 87.525 100.355 ;
        RECT 87.695 99.805 87.915 100.185 ;
        RECT 84.885 99.565 87.470 99.745 ;
        RECT 66.435 98.310 66.630 98.485 ;
        RECT 66.015 97.805 66.630 98.310 ;
        RECT 66.800 97.975 67.275 98.315 ;
        RECT 67.445 97.805 67.660 98.350 ;
        RECT 67.870 97.975 68.145 98.675 ;
        RECT 71.720 98.240 72.070 99.490 ;
        RECT 74.755 98.995 74.990 99.535 ;
        RECT 75.160 99.165 76.525 99.365 ;
        RECT 76.845 99.165 80.060 99.365 ;
        RECT 80.230 99.165 82.100 99.365 ;
        RECT 82.270 99.165 84.315 99.365 ;
        RECT 76.355 98.995 76.525 99.165 ;
        RECT 80.230 98.995 80.400 99.165 ;
        RECT 82.270 98.995 82.440 99.165 ;
        RECT 84.485 98.995 84.705 99.535 ;
        RECT 84.875 99.165 85.210 99.395 ;
        RECT 85.400 99.335 85.850 99.395 ;
        RECT 85.395 99.165 85.850 99.335 ;
        RECT 86.020 99.165 86.490 99.395 ;
        RECT 86.660 99.165 86.990 99.395 ;
        RECT 68.315 97.805 73.660 98.240 ;
        RECT 74.295 97.805 74.585 98.970 ;
        RECT 74.755 98.825 75.970 98.995 ;
        RECT 76.355 98.825 80.400 98.995 ;
        RECT 80.570 98.825 82.440 98.995 ;
        RECT 74.755 97.975 75.130 98.825 ;
        RECT 75.720 98.655 75.970 98.825 ;
        RECT 82.630 98.775 84.705 98.995 ;
        RECT 87.160 98.950 87.470 99.565 ;
        RECT 82.630 98.655 82.920 98.775 ;
        RECT 75.300 97.805 75.550 98.605 ;
        RECT 75.720 98.435 78.490 98.655 ;
        RECT 75.720 97.975 75.970 98.435 ;
        RECT 76.140 97.805 76.390 98.265 ;
        RECT 76.560 97.975 76.810 98.435 ;
        RECT 76.980 97.805 77.230 98.265 ;
        RECT 77.400 97.975 77.650 98.435 ;
        RECT 77.820 97.805 78.070 98.265 ;
        RECT 78.240 97.975 78.490 98.435 ;
        RECT 78.705 98.435 80.660 98.655 ;
        RECT 78.705 97.975 79.020 98.435 ;
        RECT 79.190 97.805 79.440 98.265 ;
        RECT 79.610 97.975 79.860 98.435 ;
        RECT 80.030 97.805 80.280 98.265 ;
        RECT 80.450 98.225 80.660 98.435 ;
        RECT 80.830 98.395 82.920 98.655 ;
        RECT 80.450 97.975 82.420 98.225 ;
        RECT 82.630 97.975 82.920 98.395 ;
        RECT 83.090 97.805 83.340 98.605 ;
        RECT 83.510 97.975 83.760 98.775 ;
        RECT 83.930 97.805 84.180 98.605 ;
        RECT 84.350 97.975 84.705 98.775 ;
        RECT 84.885 98.780 87.470 98.950 ;
        RECT 84.885 98.115 85.215 98.780 ;
        RECT 85.675 98.420 87.015 98.600 ;
        RECT 85.675 97.975 86.005 98.420 ;
        RECT 86.240 97.805 86.515 98.250 ;
        RECT 86.685 97.975 87.015 98.420 ;
        RECT 87.215 97.805 87.470 98.610 ;
        RECT 87.685 98.105 87.915 99.805 ;
        RECT 88.085 99.535 88.380 100.355 ;
        RECT 88.560 99.535 88.855 100.355 ;
        RECT 89.025 99.805 89.245 100.185 ;
        RECT 89.415 99.995 90.265 100.355 ;
        RECT 88.085 97.805 88.380 98.950 ;
        RECT 88.560 97.805 88.855 98.950 ;
        RECT 89.025 98.105 89.255 99.805 ;
        RECT 90.745 99.745 91.075 100.165 ;
        RECT 91.280 99.915 91.555 100.355 ;
        RECT 91.725 99.745 92.055 100.165 ;
        RECT 89.470 99.565 92.055 99.745 ;
        RECT 89.470 98.950 89.780 99.565 ;
        RECT 93.165 99.545 93.435 100.355 ;
        RECT 93.605 99.545 93.935 100.185 ;
        RECT 94.105 99.545 94.345 100.355 ;
        RECT 94.545 99.545 94.815 100.355 ;
        RECT 94.985 99.545 95.315 100.185 ;
        RECT 95.485 99.545 95.725 100.355 ;
        RECT 95.915 99.585 99.425 100.355 ;
        RECT 100.055 99.630 100.345 100.355 ;
        RECT 101.175 99.725 101.505 100.085 ;
        RECT 102.125 99.895 102.375 100.355 ;
        RECT 102.545 99.895 103.105 100.185 ;
        RECT 89.950 99.165 90.280 99.395 ;
        RECT 90.450 99.165 90.920 99.395 ;
        RECT 91.090 99.335 91.540 99.395 ;
        RECT 91.090 99.165 91.545 99.335 ;
        RECT 91.730 99.165 92.065 99.395 ;
        RECT 93.155 99.115 93.505 99.365 ;
        RECT 89.470 98.780 92.055 98.950 ;
        RECT 93.675 98.945 93.845 99.545 ;
        RECT 94.015 99.115 94.365 99.365 ;
        RECT 94.535 99.115 94.885 99.365 ;
        RECT 95.055 98.945 95.225 99.545 ;
        RECT 95.395 99.115 95.745 99.365 ;
        RECT 95.915 99.065 97.565 99.585 ;
        RECT 101.175 99.535 102.565 99.725 ;
        RECT 102.395 99.445 102.565 99.535 ;
        RECT 89.470 97.805 89.725 98.610 ;
        RECT 89.925 98.420 91.265 98.600 ;
        RECT 89.925 97.975 90.255 98.420 ;
        RECT 90.425 97.805 90.700 98.250 ;
        RECT 90.935 97.975 91.265 98.420 ;
        RECT 91.725 98.115 92.055 98.780 ;
        RECT 93.165 97.805 93.495 98.945 ;
        RECT 93.675 98.775 94.355 98.945 ;
        RECT 94.025 97.990 94.355 98.775 ;
        RECT 94.545 97.805 94.875 98.945 ;
        RECT 95.055 98.775 95.735 98.945 ;
        RECT 97.735 98.895 99.425 99.415 ;
        RECT 100.990 99.115 101.665 99.365 ;
        RECT 101.885 99.115 102.225 99.365 ;
        RECT 102.395 99.115 102.685 99.445 ;
        RECT 95.405 97.990 95.735 98.775 ;
        RECT 95.915 97.805 99.425 98.895 ;
        RECT 100.055 97.805 100.345 98.970 ;
        RECT 100.990 98.755 101.255 99.115 ;
        RECT 102.395 98.865 102.565 99.115 ;
        RECT 101.625 98.695 102.565 98.865 ;
        RECT 101.175 97.805 101.455 98.475 ;
        RECT 101.625 98.145 101.925 98.695 ;
        RECT 102.855 98.525 103.105 99.895 ;
        RECT 103.275 99.585 104.945 100.355 ;
        RECT 105.665 99.805 105.835 100.095 ;
        RECT 106.005 99.975 106.335 100.355 ;
        RECT 105.665 99.635 106.330 99.805 ;
        RECT 103.275 99.065 104.025 99.585 ;
        RECT 104.195 98.895 104.945 99.415 ;
        RECT 102.125 97.805 102.455 98.525 ;
        RECT 102.645 97.975 103.105 98.525 ;
        RECT 103.275 97.805 104.945 98.895 ;
        RECT 105.580 98.815 105.930 99.465 ;
        RECT 106.100 98.645 106.330 99.635 ;
        RECT 105.665 98.475 106.330 98.645 ;
        RECT 105.665 97.975 105.835 98.475 ;
        RECT 106.005 97.805 106.335 98.305 ;
        RECT 106.505 97.975 106.690 100.095 ;
        RECT 106.945 99.895 107.195 100.355 ;
        RECT 107.365 99.905 107.700 100.075 ;
        RECT 107.895 99.905 108.570 100.075 ;
        RECT 107.365 99.765 107.535 99.905 ;
        RECT 106.860 98.775 107.140 99.725 ;
        RECT 107.310 99.635 107.535 99.765 ;
        RECT 107.310 98.530 107.480 99.635 ;
        RECT 107.705 99.485 108.230 99.705 ;
        RECT 107.650 98.720 107.890 99.315 ;
        RECT 108.060 98.785 108.230 99.485 ;
        RECT 108.400 99.125 108.570 99.905 ;
        RECT 108.890 99.855 109.260 100.355 ;
        RECT 109.440 99.905 109.845 100.075 ;
        RECT 110.015 99.905 110.800 100.075 ;
        RECT 109.440 99.675 109.610 99.905 ;
        RECT 108.780 99.375 109.610 99.675 ;
        RECT 109.995 99.405 110.460 99.735 ;
        RECT 108.780 99.345 108.980 99.375 ;
        RECT 109.100 99.125 109.270 99.195 ;
        RECT 108.400 98.955 109.270 99.125 ;
        RECT 108.760 98.865 109.270 98.955 ;
        RECT 107.310 98.400 107.615 98.530 ;
        RECT 108.060 98.420 108.590 98.785 ;
        RECT 106.930 97.805 107.195 98.265 ;
        RECT 107.365 97.975 107.615 98.400 ;
        RECT 108.760 98.250 108.930 98.865 ;
        RECT 107.825 98.080 108.930 98.250 ;
        RECT 109.100 97.805 109.270 98.605 ;
        RECT 109.440 98.305 109.610 99.375 ;
        RECT 109.780 98.475 109.970 99.195 ;
        RECT 110.140 98.445 110.460 99.405 ;
        RECT 110.630 99.445 110.800 99.905 ;
        RECT 111.075 99.825 111.285 100.355 ;
        RECT 111.545 99.615 111.875 100.140 ;
        RECT 112.045 99.745 112.215 100.355 ;
        RECT 112.385 99.700 112.715 100.135 ;
        RECT 112.945 99.745 113.275 100.165 ;
        RECT 113.445 99.915 113.720 100.355 ;
        RECT 113.925 99.745 114.255 100.165 ;
        RECT 114.735 99.995 115.585 100.355 ;
        RECT 115.755 99.805 115.975 100.185 ;
        RECT 112.385 99.615 112.765 99.700 ;
        RECT 111.675 99.445 111.875 99.615 ;
        RECT 112.540 99.575 112.765 99.615 ;
        RECT 110.630 99.115 111.505 99.445 ;
        RECT 111.675 99.115 112.425 99.445 ;
        RECT 109.440 97.975 109.690 98.305 ;
        RECT 110.630 98.275 110.800 99.115 ;
        RECT 111.675 98.910 111.865 99.115 ;
        RECT 112.595 98.995 112.765 99.575 ;
        RECT 112.945 99.565 115.530 99.745 ;
        RECT 112.935 99.165 113.270 99.395 ;
        RECT 113.460 99.335 113.910 99.395 ;
        RECT 113.455 99.165 113.910 99.335 ;
        RECT 114.080 99.165 114.550 99.395 ;
        RECT 114.720 99.165 115.050 99.395 ;
        RECT 112.550 98.945 112.765 98.995 ;
        RECT 115.220 98.950 115.530 99.565 ;
        RECT 110.970 98.535 111.865 98.910 ;
        RECT 112.375 98.865 112.765 98.945 ;
        RECT 109.915 98.105 110.800 98.275 ;
        RECT 110.980 97.805 111.295 98.305 ;
        RECT 111.525 97.975 111.865 98.535 ;
        RECT 112.035 97.805 112.205 98.815 ;
        RECT 112.375 98.020 112.705 98.865 ;
        RECT 112.945 98.780 115.530 98.950 ;
        RECT 112.945 98.115 113.275 98.780 ;
        RECT 113.735 98.420 115.075 98.600 ;
        RECT 113.735 97.975 114.065 98.420 ;
        RECT 114.300 97.805 114.575 98.250 ;
        RECT 114.745 97.975 115.075 98.420 ;
        RECT 115.275 97.805 115.530 98.610 ;
        RECT 115.745 98.105 115.975 99.805 ;
        RECT 116.145 99.535 116.440 100.355 ;
        RECT 116.620 99.535 116.915 100.355 ;
        RECT 117.085 99.805 117.305 100.185 ;
        RECT 117.475 99.995 118.325 100.355 ;
        RECT 116.145 97.805 116.440 98.950 ;
        RECT 116.620 97.805 116.915 98.950 ;
        RECT 117.085 98.105 117.315 99.805 ;
        RECT 118.805 99.745 119.135 100.165 ;
        RECT 119.340 99.915 119.615 100.355 ;
        RECT 119.785 99.745 120.115 100.165 ;
        RECT 117.530 99.565 120.115 99.745 ;
        RECT 117.530 98.950 117.840 99.565 ;
        RECT 120.305 99.545 120.575 100.355 ;
        RECT 120.745 99.545 121.075 100.185 ;
        RECT 121.245 99.545 121.485 100.355 ;
        RECT 121.675 99.585 125.185 100.355 ;
        RECT 125.815 99.630 126.105 100.355 ;
        RECT 126.275 99.810 131.620 100.355 ;
        RECT 118.010 99.165 118.340 99.395 ;
        RECT 118.510 99.165 118.980 99.395 ;
        RECT 119.150 99.335 119.600 99.395 ;
        RECT 119.150 99.165 119.605 99.335 ;
        RECT 119.790 99.165 120.125 99.395 ;
        RECT 120.295 99.115 120.645 99.365 ;
        RECT 117.530 98.780 120.115 98.950 ;
        RECT 120.815 98.945 120.985 99.545 ;
        RECT 121.155 99.115 121.505 99.365 ;
        RECT 121.675 99.065 123.325 99.585 ;
        RECT 117.530 97.805 117.785 98.610 ;
        RECT 117.985 98.420 119.325 98.600 ;
        RECT 117.985 97.975 118.315 98.420 ;
        RECT 118.485 97.805 118.760 98.250 ;
        RECT 118.995 97.975 119.325 98.420 ;
        RECT 119.785 98.115 120.115 98.780 ;
        RECT 120.305 97.805 120.635 98.945 ;
        RECT 120.815 98.775 121.495 98.945 ;
        RECT 123.495 98.895 125.185 99.415 ;
        RECT 127.860 98.980 128.200 99.810 ;
        RECT 132.255 99.615 132.695 100.175 ;
        RECT 132.865 99.615 133.315 100.355 ;
        RECT 133.485 99.785 133.655 100.185 ;
        RECT 133.825 99.955 134.245 100.355 ;
        RECT 134.415 99.785 134.645 100.185 ;
        RECT 133.485 99.615 134.645 99.785 ;
        RECT 134.815 99.615 135.305 100.185 ;
        RECT 121.165 97.990 121.495 98.775 ;
        RECT 121.675 97.805 125.185 98.895 ;
        RECT 125.815 97.805 126.105 98.970 ;
        RECT 129.680 98.240 130.030 99.490 ;
        RECT 132.255 98.605 132.565 99.615 ;
        RECT 132.735 98.995 132.905 99.445 ;
        RECT 133.075 99.165 133.465 99.445 ;
        RECT 133.650 99.115 133.895 99.445 ;
        RECT 132.735 98.825 133.525 98.995 ;
        RECT 126.275 97.805 131.620 98.240 ;
        RECT 132.255 97.975 132.695 98.605 ;
        RECT 132.870 97.805 133.185 98.655 ;
        RECT 133.355 98.145 133.525 98.825 ;
        RECT 133.695 98.315 133.895 99.115 ;
        RECT 134.095 98.315 134.345 99.445 ;
        RECT 134.560 99.115 134.965 99.445 ;
        RECT 135.135 98.945 135.305 99.615 ;
        RECT 134.535 98.775 135.305 98.945 ;
        RECT 135.475 99.555 135.815 100.185 ;
        RECT 135.985 99.555 136.235 100.355 ;
        RECT 136.425 99.705 136.755 100.185 ;
        RECT 136.925 99.895 137.150 100.355 ;
        RECT 137.320 99.705 137.650 100.185 ;
        RECT 135.475 98.945 135.650 99.555 ;
        RECT 136.425 99.535 137.650 99.705 ;
        RECT 138.280 99.575 138.780 100.185 ;
        RECT 139.155 99.585 141.745 100.355 ;
        RECT 142.115 99.725 142.445 100.085 ;
        RECT 143.065 99.895 143.315 100.355 ;
        RECT 143.485 99.895 144.045 100.185 ;
        RECT 135.820 99.195 136.515 99.365 ;
        RECT 136.345 98.945 136.515 99.195 ;
        RECT 136.690 99.165 137.110 99.365 ;
        RECT 137.280 99.165 137.610 99.365 ;
        RECT 137.780 99.165 138.110 99.365 ;
        RECT 138.280 98.945 138.450 99.575 ;
        RECT 138.635 99.115 138.985 99.365 ;
        RECT 139.155 99.065 140.365 99.585 ;
        RECT 142.115 99.535 143.505 99.725 ;
        RECT 143.335 99.445 143.505 99.535 ;
        RECT 134.535 98.145 134.785 98.775 ;
        RECT 133.355 97.975 134.785 98.145 ;
        RECT 134.965 97.805 135.295 98.605 ;
        RECT 135.475 97.975 135.815 98.945 ;
        RECT 135.985 97.805 136.155 98.945 ;
        RECT 136.345 98.775 138.780 98.945 ;
        RECT 140.535 98.895 141.745 99.415 ;
        RECT 136.425 97.805 136.675 98.605 ;
        RECT 137.320 97.975 137.650 98.775 ;
        RECT 137.950 97.805 138.280 98.605 ;
        RECT 138.450 97.975 138.780 98.775 ;
        RECT 139.155 97.805 141.745 98.895 ;
        RECT 141.930 99.115 142.605 99.365 ;
        RECT 142.825 99.115 143.165 99.365 ;
        RECT 143.335 99.115 143.625 99.445 ;
        RECT 141.930 98.755 142.195 99.115 ;
        RECT 143.335 98.865 143.505 99.115 ;
        RECT 142.565 98.695 143.505 98.865 ;
        RECT 142.115 97.805 142.395 98.475 ;
        RECT 142.565 98.145 142.865 98.695 ;
        RECT 143.795 98.525 144.045 99.895 ;
        RECT 144.215 99.810 149.560 100.355 ;
        RECT 145.800 98.980 146.140 99.810 ;
        RECT 149.735 99.585 151.405 100.355 ;
        RECT 151.575 99.630 151.865 100.355 ;
        RECT 152.035 99.585 155.545 100.355 ;
        RECT 155.715 99.605 156.925 100.355 ;
        RECT 143.065 97.805 143.395 98.525 ;
        RECT 143.585 97.975 144.045 98.525 ;
        RECT 147.620 98.240 147.970 99.490 ;
        RECT 149.735 99.065 150.485 99.585 ;
        RECT 150.655 98.895 151.405 99.415 ;
        RECT 152.035 99.065 153.685 99.585 ;
        RECT 144.215 97.805 149.560 98.240 ;
        RECT 149.735 97.805 151.405 98.895 ;
        RECT 151.575 97.805 151.865 98.970 ;
        RECT 153.855 98.895 155.545 99.415 ;
        RECT 152.035 97.805 155.545 98.895 ;
        RECT 155.715 98.895 156.235 99.435 ;
        RECT 156.405 99.065 156.925 99.605 ;
        RECT 155.715 97.805 156.925 98.895 ;
        RECT 22.690 97.635 157.010 97.805 ;
        RECT 22.775 96.545 23.985 97.635 ;
        RECT 24.165 97.045 24.425 97.435 ;
        RECT 24.595 97.225 24.925 97.635 ;
        RECT 24.165 96.845 24.925 97.045 ;
        RECT 22.775 95.835 23.295 96.375 ;
        RECT 23.465 96.005 23.985 96.545 ;
        RECT 24.175 95.975 24.405 96.665 ;
        RECT 24.585 96.165 24.925 96.845 ;
        RECT 25.115 96.345 25.445 97.455 ;
        RECT 25.615 96.725 25.805 97.455 ;
        RECT 25.975 96.905 26.305 97.635 ;
        RECT 26.485 96.725 26.655 97.455 ;
        RECT 25.615 96.525 26.655 96.725 ;
        RECT 26.915 96.535 27.235 97.465 ;
        RECT 27.415 96.955 27.815 97.465 ;
        RECT 27.985 97.125 28.155 97.635 ;
        RECT 28.325 96.955 28.655 97.465 ;
        RECT 27.415 96.785 28.655 96.955 ;
        RECT 28.825 96.785 28.995 97.635 ;
        RECT 29.585 96.785 29.965 97.465 ;
        RECT 26.915 96.365 27.545 96.535 ;
        RECT 22.775 95.085 23.985 95.835 ;
        RECT 24.585 95.715 24.815 96.165 ;
        RECT 25.115 96.045 25.650 96.345 ;
        RECT 24.435 95.265 24.815 95.715 ;
        RECT 24.995 95.085 25.225 95.865 ;
        RECT 25.405 95.795 25.650 96.045 ;
        RECT 25.830 95.995 26.225 96.345 ;
        RECT 26.420 95.995 26.710 96.345 ;
        RECT 25.405 95.265 25.835 95.795 ;
        RECT 26.015 95.375 26.225 95.995 ;
        RECT 26.395 95.085 26.725 95.815 ;
        RECT 26.915 95.085 27.205 95.920 ;
        RECT 27.375 95.485 27.545 96.365 ;
        RECT 28.320 96.445 29.625 96.615 ;
        RECT 27.715 95.825 27.945 96.325 ;
        RECT 28.320 96.245 28.490 96.445 ;
        RECT 28.115 96.075 28.490 96.245 ;
        RECT 28.660 96.075 29.210 96.275 ;
        RECT 29.380 95.995 29.625 96.445 ;
        RECT 29.795 95.825 29.965 96.785 ;
        RECT 27.715 95.655 29.965 95.825 ;
        RECT 30.135 96.030 30.415 97.465 ;
        RECT 30.585 96.860 31.295 97.635 ;
        RECT 31.465 96.690 31.795 97.465 ;
        RECT 30.645 96.475 31.795 96.690 ;
        RECT 27.375 95.315 28.330 95.485 ;
        RECT 28.745 95.085 29.075 95.475 ;
        RECT 29.245 95.335 29.415 95.655 ;
        RECT 29.585 95.085 29.915 95.475 ;
        RECT 30.135 95.255 30.475 96.030 ;
        RECT 30.645 95.905 30.930 96.475 ;
        RECT 31.115 96.075 31.585 96.305 ;
        RECT 31.990 96.275 32.205 97.390 ;
        RECT 32.385 96.915 32.715 97.635 ;
        RECT 32.930 96.845 33.465 97.465 ;
        RECT 32.495 96.275 32.725 96.615 ;
        RECT 31.755 96.095 32.205 96.275 ;
        RECT 31.755 96.075 32.085 96.095 ;
        RECT 32.395 96.075 32.725 96.275 ;
        RECT 30.645 95.715 31.355 95.905 ;
        RECT 31.055 95.575 31.355 95.715 ;
        RECT 31.545 95.715 32.725 95.905 ;
        RECT 31.545 95.635 31.875 95.715 ;
        RECT 31.055 95.565 31.370 95.575 ;
        RECT 31.055 95.555 31.380 95.565 ;
        RECT 31.055 95.550 31.390 95.555 ;
        RECT 30.645 95.085 30.815 95.545 ;
        RECT 31.055 95.540 31.395 95.550 ;
        RECT 31.055 95.535 31.400 95.540 ;
        RECT 31.055 95.525 31.405 95.535 ;
        RECT 31.055 95.520 31.410 95.525 ;
        RECT 31.055 95.255 31.415 95.520 ;
        RECT 32.045 95.085 32.215 95.545 ;
        RECT 32.385 95.255 32.725 95.715 ;
        RECT 32.930 95.825 33.245 96.845 ;
        RECT 33.635 96.835 33.965 97.635 ;
        RECT 34.450 96.665 34.840 96.840 ;
        RECT 33.415 96.495 34.840 96.665 ;
        RECT 33.415 95.995 33.585 96.495 ;
        RECT 32.930 95.255 33.545 95.825 ;
        RECT 33.835 95.765 34.100 96.325 ;
        RECT 34.270 95.595 34.440 96.495 ;
        RECT 35.655 96.470 35.945 97.635 ;
        RECT 36.205 96.965 36.375 97.465 ;
        RECT 36.545 97.135 36.875 97.635 ;
        RECT 36.205 96.795 36.870 96.965 ;
        RECT 34.610 95.765 34.965 96.325 ;
        RECT 36.120 95.975 36.470 96.625 ;
        RECT 33.715 95.085 33.930 95.595 ;
        RECT 34.160 95.265 34.440 95.595 ;
        RECT 34.620 95.085 34.860 95.595 ;
        RECT 35.655 95.085 35.945 95.810 ;
        RECT 36.640 95.805 36.870 96.795 ;
        RECT 36.205 95.635 36.870 95.805 ;
        RECT 36.205 95.345 36.375 95.635 ;
        RECT 36.545 95.085 36.875 95.465 ;
        RECT 37.045 95.345 37.230 97.465 ;
        RECT 37.470 97.175 37.735 97.635 ;
        RECT 37.905 97.040 38.155 97.465 ;
        RECT 38.365 97.190 39.470 97.360 ;
        RECT 37.850 96.910 38.155 97.040 ;
        RECT 37.400 95.715 37.680 96.665 ;
        RECT 37.850 95.805 38.020 96.910 ;
        RECT 38.190 96.125 38.430 96.720 ;
        RECT 38.600 96.655 39.130 97.020 ;
        RECT 38.600 95.955 38.770 96.655 ;
        RECT 39.300 96.575 39.470 97.190 ;
        RECT 39.640 96.835 39.810 97.635 ;
        RECT 39.980 97.135 40.230 97.465 ;
        RECT 40.455 97.165 41.340 97.335 ;
        RECT 39.300 96.485 39.810 96.575 ;
        RECT 37.850 95.675 38.075 95.805 ;
        RECT 38.245 95.735 38.770 95.955 ;
        RECT 38.940 96.315 39.810 96.485 ;
        RECT 37.485 95.085 37.735 95.545 ;
        RECT 37.905 95.535 38.075 95.675 ;
        RECT 38.940 95.535 39.110 96.315 ;
        RECT 39.640 96.245 39.810 96.315 ;
        RECT 39.320 96.065 39.520 96.095 ;
        RECT 39.980 96.065 40.150 97.135 ;
        RECT 40.320 96.245 40.510 96.965 ;
        RECT 39.320 95.765 40.150 96.065 ;
        RECT 40.680 96.035 41.000 96.995 ;
        RECT 37.905 95.365 38.240 95.535 ;
        RECT 38.435 95.365 39.110 95.535 ;
        RECT 39.430 95.085 39.800 95.585 ;
        RECT 39.980 95.535 40.150 95.765 ;
        RECT 40.535 95.705 41.000 96.035 ;
        RECT 41.170 96.325 41.340 97.165 ;
        RECT 41.520 97.135 41.835 97.635 ;
        RECT 42.065 96.905 42.405 97.465 ;
        RECT 41.510 96.530 42.405 96.905 ;
        RECT 42.575 96.625 42.745 97.635 ;
        RECT 42.215 96.325 42.405 96.530 ;
        RECT 42.915 96.575 43.245 97.420 ;
        RECT 42.915 96.495 43.305 96.575 ;
        RECT 43.475 96.545 46.065 97.635 ;
        RECT 46.325 96.965 46.495 97.465 ;
        RECT 46.665 97.135 46.995 97.635 ;
        RECT 46.325 96.795 46.990 96.965 ;
        RECT 43.090 96.445 43.305 96.495 ;
        RECT 41.170 95.995 42.045 96.325 ;
        RECT 42.215 95.995 42.965 96.325 ;
        RECT 41.170 95.535 41.340 95.995 ;
        RECT 42.215 95.825 42.415 95.995 ;
        RECT 43.135 95.865 43.305 96.445 ;
        RECT 43.080 95.825 43.305 95.865 ;
        RECT 39.980 95.365 40.385 95.535 ;
        RECT 40.555 95.365 41.340 95.535 ;
        RECT 41.615 95.085 41.825 95.615 ;
        RECT 42.085 95.300 42.415 95.825 ;
        RECT 42.925 95.740 43.305 95.825 ;
        RECT 43.475 95.855 44.685 96.375 ;
        RECT 44.855 96.025 46.065 96.545 ;
        RECT 46.240 95.975 46.590 96.625 ;
        RECT 42.585 95.085 42.755 95.695 ;
        RECT 42.925 95.305 43.255 95.740 ;
        RECT 43.475 95.085 46.065 95.855 ;
        RECT 46.760 95.805 46.990 96.795 ;
        RECT 46.325 95.635 46.990 95.805 ;
        RECT 46.325 95.345 46.495 95.635 ;
        RECT 46.665 95.085 46.995 95.465 ;
        RECT 47.165 95.345 47.350 97.465 ;
        RECT 47.590 97.175 47.855 97.635 ;
        RECT 48.025 97.040 48.275 97.465 ;
        RECT 48.485 97.190 49.590 97.360 ;
        RECT 47.970 96.910 48.275 97.040 ;
        RECT 47.520 95.715 47.800 96.665 ;
        RECT 47.970 95.805 48.140 96.910 ;
        RECT 48.310 96.125 48.550 96.720 ;
        RECT 48.720 96.655 49.250 97.020 ;
        RECT 48.720 95.955 48.890 96.655 ;
        RECT 49.420 96.575 49.590 97.190 ;
        RECT 49.760 96.835 49.930 97.635 ;
        RECT 50.100 97.135 50.350 97.465 ;
        RECT 50.575 97.165 51.460 97.335 ;
        RECT 49.420 96.485 49.930 96.575 ;
        RECT 47.970 95.675 48.195 95.805 ;
        RECT 48.365 95.735 48.890 95.955 ;
        RECT 49.060 96.315 49.930 96.485 ;
        RECT 47.605 95.085 47.855 95.545 ;
        RECT 48.025 95.535 48.195 95.675 ;
        RECT 49.060 95.535 49.230 96.315 ;
        RECT 49.760 96.245 49.930 96.315 ;
        RECT 49.440 96.065 49.640 96.095 ;
        RECT 50.100 96.065 50.270 97.135 ;
        RECT 50.440 96.245 50.630 96.965 ;
        RECT 49.440 95.765 50.270 96.065 ;
        RECT 50.800 96.035 51.120 96.995 ;
        RECT 48.025 95.365 48.360 95.535 ;
        RECT 48.555 95.365 49.230 95.535 ;
        RECT 49.550 95.085 49.920 95.585 ;
        RECT 50.100 95.535 50.270 95.765 ;
        RECT 50.655 95.705 51.120 96.035 ;
        RECT 51.290 96.325 51.460 97.165 ;
        RECT 51.640 97.135 51.955 97.635 ;
        RECT 52.185 96.905 52.525 97.465 ;
        RECT 51.630 96.530 52.525 96.905 ;
        RECT 52.695 96.625 52.865 97.635 ;
        RECT 52.335 96.325 52.525 96.530 ;
        RECT 53.035 96.575 53.365 97.420 ;
        RECT 53.685 96.965 53.855 97.465 ;
        RECT 54.025 97.135 54.355 97.635 ;
        RECT 53.685 96.795 54.350 96.965 ;
        RECT 53.035 96.495 53.425 96.575 ;
        RECT 53.210 96.445 53.425 96.495 ;
        RECT 51.290 95.995 52.165 96.325 ;
        RECT 52.335 95.995 53.085 96.325 ;
        RECT 51.290 95.535 51.460 95.995 ;
        RECT 52.335 95.825 52.535 95.995 ;
        RECT 53.255 95.865 53.425 96.445 ;
        RECT 53.600 95.975 53.950 96.625 ;
        RECT 53.200 95.825 53.425 95.865 ;
        RECT 50.100 95.365 50.505 95.535 ;
        RECT 50.675 95.365 51.460 95.535 ;
        RECT 51.735 95.085 51.945 95.615 ;
        RECT 52.205 95.300 52.535 95.825 ;
        RECT 53.045 95.740 53.425 95.825 ;
        RECT 54.120 95.805 54.350 96.795 ;
        RECT 52.705 95.085 52.875 95.695 ;
        RECT 53.045 95.305 53.375 95.740 ;
        RECT 53.685 95.635 54.350 95.805 ;
        RECT 53.685 95.345 53.855 95.635 ;
        RECT 54.025 95.085 54.355 95.465 ;
        RECT 54.525 95.345 54.710 97.465 ;
        RECT 54.950 97.175 55.215 97.635 ;
        RECT 55.385 97.040 55.635 97.465 ;
        RECT 55.845 97.190 56.950 97.360 ;
        RECT 55.330 96.910 55.635 97.040 ;
        RECT 54.880 95.715 55.160 96.665 ;
        RECT 55.330 95.805 55.500 96.910 ;
        RECT 55.670 96.125 55.910 96.720 ;
        RECT 56.080 96.655 56.610 97.020 ;
        RECT 56.080 95.955 56.250 96.655 ;
        RECT 56.780 96.575 56.950 97.190 ;
        RECT 57.120 96.835 57.290 97.635 ;
        RECT 57.460 97.135 57.710 97.465 ;
        RECT 57.935 97.165 58.820 97.335 ;
        RECT 56.780 96.485 57.290 96.575 ;
        RECT 55.330 95.675 55.555 95.805 ;
        RECT 55.725 95.735 56.250 95.955 ;
        RECT 56.420 96.315 57.290 96.485 ;
        RECT 54.965 95.085 55.215 95.545 ;
        RECT 55.385 95.535 55.555 95.675 ;
        RECT 56.420 95.535 56.590 96.315 ;
        RECT 57.120 96.245 57.290 96.315 ;
        RECT 56.800 96.065 57.000 96.095 ;
        RECT 57.460 96.065 57.630 97.135 ;
        RECT 57.800 96.245 57.990 96.965 ;
        RECT 56.800 95.765 57.630 96.065 ;
        RECT 58.160 96.035 58.480 96.995 ;
        RECT 55.385 95.365 55.720 95.535 ;
        RECT 55.915 95.365 56.590 95.535 ;
        RECT 56.910 95.085 57.280 95.585 ;
        RECT 57.460 95.535 57.630 95.765 ;
        RECT 58.015 95.705 58.480 96.035 ;
        RECT 58.650 96.325 58.820 97.165 ;
        RECT 59.000 97.135 59.315 97.635 ;
        RECT 59.545 96.905 59.885 97.465 ;
        RECT 58.990 96.530 59.885 96.905 ;
        RECT 60.055 96.625 60.225 97.635 ;
        RECT 59.695 96.325 59.885 96.530 ;
        RECT 60.395 96.575 60.725 97.420 ;
        RECT 60.895 96.720 61.065 97.635 ;
        RECT 60.395 96.495 60.785 96.575 ;
        RECT 60.570 96.445 60.785 96.495 ;
        RECT 61.415 96.470 61.705 97.635 ;
        RECT 61.875 96.545 65.385 97.635 ;
        RECT 66.105 96.965 66.275 97.465 ;
        RECT 66.445 97.135 66.775 97.635 ;
        RECT 66.105 96.795 66.770 96.965 ;
        RECT 58.650 95.995 59.525 96.325 ;
        RECT 59.695 95.995 60.445 96.325 ;
        RECT 58.650 95.535 58.820 95.995 ;
        RECT 59.695 95.825 59.895 95.995 ;
        RECT 60.615 95.865 60.785 96.445 ;
        RECT 60.560 95.825 60.785 95.865 ;
        RECT 57.460 95.365 57.865 95.535 ;
        RECT 58.035 95.365 58.820 95.535 ;
        RECT 59.095 95.085 59.305 95.615 ;
        RECT 59.565 95.300 59.895 95.825 ;
        RECT 60.405 95.740 60.785 95.825 ;
        RECT 61.875 95.855 63.525 96.375 ;
        RECT 63.695 96.025 65.385 96.545 ;
        RECT 66.020 95.975 66.370 96.625 ;
        RECT 60.065 95.085 60.235 95.695 ;
        RECT 60.405 95.305 60.735 95.740 ;
        RECT 60.905 95.085 61.075 95.600 ;
        RECT 61.415 95.085 61.705 95.810 ;
        RECT 61.875 95.085 65.385 95.855 ;
        RECT 66.540 95.805 66.770 96.795 ;
        RECT 66.105 95.635 66.770 95.805 ;
        RECT 66.105 95.345 66.275 95.635 ;
        RECT 66.445 95.085 66.775 95.465 ;
        RECT 66.945 95.345 67.130 97.465 ;
        RECT 67.370 97.175 67.635 97.635 ;
        RECT 67.805 97.040 68.055 97.465 ;
        RECT 68.265 97.190 69.370 97.360 ;
        RECT 67.750 96.910 68.055 97.040 ;
        RECT 67.300 95.715 67.580 96.665 ;
        RECT 67.750 95.805 67.920 96.910 ;
        RECT 68.090 96.125 68.330 96.720 ;
        RECT 68.500 96.655 69.030 97.020 ;
        RECT 68.500 95.955 68.670 96.655 ;
        RECT 69.200 96.575 69.370 97.190 ;
        RECT 69.540 96.835 69.710 97.635 ;
        RECT 69.880 97.135 70.130 97.465 ;
        RECT 70.355 97.165 71.240 97.335 ;
        RECT 69.200 96.485 69.710 96.575 ;
        RECT 67.750 95.675 67.975 95.805 ;
        RECT 68.145 95.735 68.670 95.955 ;
        RECT 68.840 96.315 69.710 96.485 ;
        RECT 67.385 95.085 67.635 95.545 ;
        RECT 67.805 95.535 67.975 95.675 ;
        RECT 68.840 95.535 69.010 96.315 ;
        RECT 69.540 96.245 69.710 96.315 ;
        RECT 69.220 96.065 69.420 96.095 ;
        RECT 69.880 96.065 70.050 97.135 ;
        RECT 70.220 96.245 70.410 96.965 ;
        RECT 69.220 95.765 70.050 96.065 ;
        RECT 70.580 96.035 70.900 96.995 ;
        RECT 67.805 95.365 68.140 95.535 ;
        RECT 68.335 95.365 69.010 95.535 ;
        RECT 69.330 95.085 69.700 95.585 ;
        RECT 69.880 95.535 70.050 95.765 ;
        RECT 70.435 95.705 70.900 96.035 ;
        RECT 71.070 96.325 71.240 97.165 ;
        RECT 71.420 97.135 71.735 97.635 ;
        RECT 71.965 96.905 72.305 97.465 ;
        RECT 71.410 96.530 72.305 96.905 ;
        RECT 72.475 96.625 72.645 97.635 ;
        RECT 72.115 96.325 72.305 96.530 ;
        RECT 72.815 96.575 73.145 97.420 ;
        RECT 73.375 96.965 73.690 97.465 ;
        RECT 73.860 97.135 74.110 97.635 ;
        RECT 74.280 96.965 74.530 97.465 ;
        RECT 74.700 97.135 74.950 97.635 ;
        RECT 75.120 96.965 75.370 97.465 ;
        RECT 75.680 97.125 75.930 97.465 ;
        RECT 76.100 97.135 76.350 97.635 ;
        RECT 76.520 97.295 77.645 97.465 ;
        RECT 76.520 97.125 76.845 97.295 ;
        RECT 77.395 97.135 77.645 97.295 ;
        RECT 77.915 97.135 78.165 97.635 ;
        RECT 73.375 96.955 75.370 96.965 ;
        RECT 77.015 96.965 77.225 97.125 ;
        RECT 78.335 96.965 78.585 97.125 ;
        RECT 73.375 96.785 76.770 96.955 ;
        RECT 77.015 96.795 78.585 96.965 ;
        RECT 78.755 96.795 79.185 97.635 ;
        RECT 72.815 96.495 73.205 96.575 ;
        RECT 72.990 96.445 73.205 96.495 ;
        RECT 71.070 95.995 71.945 96.325 ;
        RECT 72.115 95.995 72.865 96.325 ;
        RECT 71.070 95.535 71.240 95.995 ;
        RECT 72.115 95.825 72.315 95.995 ;
        RECT 73.035 95.865 73.205 96.445 ;
        RECT 72.980 95.825 73.205 95.865 ;
        RECT 69.880 95.365 70.285 95.535 ;
        RECT 70.455 95.365 71.240 95.535 ;
        RECT 71.515 95.085 71.725 95.615 ;
        RECT 71.985 95.300 72.315 95.825 ;
        RECT 72.825 95.740 73.205 95.825 ;
        RECT 73.375 95.895 73.605 96.785 ;
        RECT 76.600 96.625 76.770 96.785 ;
        RECT 78.335 96.625 78.585 96.795 ;
        RECT 74.080 96.445 76.390 96.615 ;
        RECT 76.600 96.455 78.095 96.625 ;
        RECT 74.080 96.285 74.250 96.445 ;
        RECT 73.775 96.075 74.250 96.285 ;
        RECT 76.220 96.285 76.390 96.445 ;
        RECT 74.545 96.075 75.995 96.275 ;
        RECT 76.220 96.075 77.245 96.285 ;
        RECT 77.925 96.245 78.095 96.455 ;
        RECT 78.335 96.415 79.185 96.625 ;
        RECT 79.355 96.545 81.945 97.635 ;
        RECT 82.175 97.285 84.245 97.455 ;
        RECT 82.175 96.785 82.435 97.285 ;
        RECT 83.105 97.255 84.245 97.285 ;
        RECT 82.605 96.785 82.935 97.105 ;
        RECT 83.105 96.785 83.295 97.255 ;
        RECT 77.925 96.075 78.585 96.245 ;
        RECT 72.485 95.085 72.655 95.695 ;
        RECT 72.825 95.305 73.155 95.740 ;
        RECT 73.375 95.645 74.150 95.895 ;
        RECT 74.320 95.725 75.410 95.905 ;
        RECT 74.320 95.475 74.570 95.725 ;
        RECT 73.395 95.255 74.570 95.475 ;
        RECT 74.740 95.085 74.910 95.555 ;
        RECT 75.080 95.255 75.410 95.725 ;
        RECT 75.720 95.085 75.890 95.905 ;
        RECT 76.060 95.725 78.625 95.905 ;
        RECT 76.060 95.255 76.390 95.725 ;
        RECT 76.560 95.085 76.730 95.555 ;
        RECT 76.900 95.255 77.265 95.725 ;
        RECT 78.295 95.645 78.625 95.725 ;
        RECT 77.435 95.085 77.605 95.555 ;
        RECT 78.795 95.475 79.185 96.415 ;
        RECT 77.875 95.305 79.185 95.475 ;
        RECT 79.355 95.855 80.565 96.375 ;
        RECT 80.735 96.025 81.945 96.545 ;
        RECT 82.130 95.995 82.435 96.615 ;
        RECT 82.605 95.855 82.885 96.785 ;
        RECT 83.465 96.655 83.795 97.075 ;
        RECT 83.965 96.835 84.245 97.255 ;
        RECT 84.465 96.835 84.695 97.635 ;
        RECT 84.875 96.655 85.145 97.465 ;
        RECT 85.325 96.835 85.555 97.635 ;
        RECT 85.735 96.655 86.005 97.465 ;
        RECT 86.185 96.835 86.415 97.635 ;
        RECT 83.065 96.285 83.285 96.615 ;
        RECT 83.465 96.455 86.005 96.655 ;
        RECT 86.205 96.285 86.530 96.655 ;
        RECT 87.175 96.470 87.465 97.635 ;
        RECT 87.635 96.545 90.225 97.635 ;
        RECT 90.400 97.255 94.135 97.465 ;
        RECT 94.305 97.275 94.635 97.635 ;
        RECT 93.965 97.105 94.135 97.255 ;
        RECT 94.805 97.105 94.975 97.465 ;
        RECT 95.145 97.275 95.475 97.635 ;
        RECT 95.645 97.105 95.815 97.465 ;
        RECT 95.985 97.275 96.315 97.635 ;
        RECT 96.485 97.105 96.655 97.465 ;
        RECT 96.825 97.255 97.155 97.635 ;
        RECT 93.965 97.085 96.655 97.105 ;
        RECT 97.325 97.085 97.575 97.465 ;
        RECT 83.065 96.035 83.815 96.285 ;
        RECT 84.400 96.035 85.110 96.285 ;
        RECT 85.770 96.035 86.530 96.285 ;
        RECT 84.015 95.855 84.185 95.935 ;
        RECT 87.635 95.855 88.845 96.375 ;
        RECT 89.015 96.025 90.225 96.545 ;
        RECT 90.395 96.865 92.500 97.085 ;
        RECT 90.395 96.495 90.740 96.865 ;
        RECT 92.760 96.785 93.795 97.085 ;
        RECT 93.965 96.795 97.575 97.085 ;
        RECT 92.760 96.695 93.040 96.785 ;
        RECT 79.355 95.085 81.945 95.855 ;
        RECT 82.175 95.085 82.425 95.815 ;
        RECT 82.605 95.655 85.175 95.855 ;
        RECT 82.605 95.255 82.865 95.655 ;
        RECT 83.035 95.085 83.365 95.475 ;
        RECT 83.535 95.285 83.725 95.655 ;
        RECT 85.355 95.635 86.465 95.855 ;
        RECT 85.355 95.475 85.525 95.635 ;
        RECT 83.895 95.085 84.225 95.475 ;
        RECT 84.415 95.265 85.525 95.475 ;
        RECT 85.705 95.085 86.035 95.455 ;
        RECT 86.215 95.265 86.465 95.635 ;
        RECT 87.175 95.085 87.465 95.810 ;
        RECT 87.635 95.085 90.225 95.855 ;
        RECT 90.395 95.825 90.565 96.495 ;
        RECT 90.910 96.325 91.080 96.615 ;
        RECT 90.735 95.995 91.080 96.325 ;
        RECT 91.320 96.275 91.540 96.695 ;
        RECT 91.710 96.445 93.040 96.695 ;
        RECT 93.210 96.275 93.925 96.615 ;
        RECT 91.320 96.035 92.670 96.275 ;
        RECT 92.915 96.035 93.925 96.275 ;
        RECT 94.095 96.445 97.570 96.625 ;
        RECT 97.755 96.545 100.345 97.635 ;
        RECT 94.095 96.035 94.425 96.445 ;
        RECT 94.595 96.245 96.010 96.275 ;
        RECT 94.595 96.105 96.015 96.245 ;
        RECT 94.665 96.075 96.015 96.105 ;
        RECT 94.665 96.035 96.010 96.075 ;
        RECT 96.285 96.035 97.570 96.445 ;
        RECT 91.315 95.825 95.895 95.865 ;
        RECT 90.395 95.695 95.895 95.825 ;
        RECT 90.395 95.625 93.795 95.695 ;
        RECT 94.340 95.675 95.895 95.695 ;
        RECT 96.065 95.695 97.105 95.865 ;
        RECT 90.395 95.615 91.955 95.625 ;
        RECT 90.400 95.085 90.755 95.445 ;
        RECT 91.285 95.085 91.615 95.445 ;
        RECT 91.785 95.255 91.955 95.615 ;
        RECT 92.625 95.615 93.795 95.625 ;
        RECT 92.125 95.085 92.455 95.445 ;
        RECT 92.625 95.255 92.795 95.615 ;
        RECT 92.975 95.085 93.305 95.445 ;
        RECT 93.475 95.255 93.795 95.615 ;
        RECT 93.965 95.085 94.135 95.525 ;
        RECT 96.065 95.505 96.315 95.695 ;
        RECT 96.895 95.530 97.105 95.695 ;
        RECT 97.755 95.855 98.965 96.375 ;
        RECT 99.135 96.025 100.345 96.545 ;
        RECT 101.065 96.705 101.235 97.465 ;
        RECT 101.415 96.875 101.745 97.635 ;
        RECT 101.065 96.535 101.730 96.705 ;
        RECT 101.915 96.560 102.185 97.465 ;
        RECT 101.560 96.390 101.730 96.535 ;
        RECT 100.995 95.985 101.325 96.355 ;
        RECT 101.560 96.060 101.845 96.390 ;
        RECT 94.305 95.255 96.315 95.505 ;
        RECT 96.485 95.085 96.720 95.525 ;
        RECT 97.275 95.085 97.575 95.585 ;
        RECT 97.755 95.085 100.345 95.855 ;
        RECT 101.560 95.805 101.730 96.060 ;
        RECT 101.065 95.635 101.730 95.805 ;
        RECT 102.015 95.760 102.185 96.560 ;
        RECT 102.355 96.545 105.865 97.635 ;
        RECT 101.065 95.255 101.235 95.635 ;
        RECT 101.415 95.085 101.745 95.465 ;
        RECT 101.925 95.255 102.185 95.760 ;
        RECT 102.355 95.855 104.005 96.375 ;
        RECT 104.175 96.025 105.865 96.545 ;
        RECT 107.045 96.705 107.215 97.465 ;
        RECT 107.395 96.875 107.725 97.635 ;
        RECT 107.045 96.535 107.710 96.705 ;
        RECT 107.895 96.560 108.165 97.465 ;
        RECT 107.540 96.390 107.710 96.535 ;
        RECT 106.975 95.985 107.305 96.355 ;
        RECT 107.540 96.060 107.825 96.390 ;
        RECT 102.355 95.085 105.865 95.855 ;
        RECT 107.540 95.805 107.710 96.060 ;
        RECT 107.045 95.635 107.710 95.805 ;
        RECT 107.995 95.760 108.165 96.560 ;
        RECT 108.335 96.545 110.925 97.635 ;
        RECT 107.045 95.255 107.215 95.635 ;
        RECT 107.395 95.085 107.725 95.465 ;
        RECT 107.905 95.255 108.165 95.760 ;
        RECT 108.335 95.855 109.545 96.375 ;
        RECT 109.715 96.025 110.925 96.545 ;
        RECT 111.565 96.665 111.895 97.450 ;
        RECT 111.565 96.495 112.245 96.665 ;
        RECT 112.425 96.495 112.755 97.635 ;
        RECT 111.555 96.075 111.905 96.325 ;
        RECT 112.075 95.895 112.245 96.495 ;
        RECT 112.935 96.470 113.225 97.635 ;
        RECT 113.485 96.890 113.755 97.635 ;
        RECT 114.385 97.630 120.660 97.635 ;
        RECT 113.925 96.720 114.215 97.460 ;
        RECT 114.385 96.905 114.640 97.630 ;
        RECT 114.825 96.735 115.085 97.460 ;
        RECT 115.255 96.905 115.500 97.630 ;
        RECT 115.685 96.735 115.945 97.460 ;
        RECT 116.115 96.905 116.360 97.630 ;
        RECT 116.545 96.735 116.805 97.460 ;
        RECT 116.975 96.905 117.220 97.630 ;
        RECT 117.390 96.735 117.650 97.460 ;
        RECT 117.820 96.905 118.080 97.630 ;
        RECT 118.250 96.735 118.510 97.460 ;
        RECT 118.680 96.905 118.940 97.630 ;
        RECT 119.110 96.735 119.370 97.460 ;
        RECT 119.540 96.905 119.800 97.630 ;
        RECT 119.970 96.735 120.230 97.460 ;
        RECT 120.400 96.835 120.660 97.630 ;
        RECT 114.825 96.720 120.230 96.735 ;
        RECT 113.485 96.495 120.230 96.720 ;
        RECT 112.415 96.075 112.765 96.325 ;
        RECT 113.485 95.905 114.650 96.495 ;
        RECT 120.830 96.325 121.080 97.460 ;
        RECT 121.260 96.825 121.520 97.635 ;
        RECT 121.695 96.325 121.940 97.465 ;
        RECT 122.120 96.825 122.415 97.635 ;
        RECT 123.065 97.045 123.325 97.435 ;
        RECT 123.495 97.225 123.825 97.635 ;
        RECT 123.065 96.845 123.825 97.045 ;
        RECT 114.820 96.075 121.940 96.325 ;
        RECT 108.335 95.085 110.925 95.855 ;
        RECT 111.575 95.085 111.815 95.895 ;
        RECT 111.985 95.255 112.315 95.895 ;
        RECT 112.485 95.085 112.755 95.895 ;
        RECT 112.935 95.085 113.225 95.810 ;
        RECT 113.485 95.735 120.230 95.905 ;
        RECT 113.485 95.085 113.785 95.565 ;
        RECT 113.955 95.280 114.215 95.735 ;
        RECT 114.385 95.085 114.645 95.565 ;
        RECT 114.825 95.280 115.085 95.735 ;
        RECT 115.255 95.085 115.505 95.565 ;
        RECT 115.685 95.280 115.945 95.735 ;
        RECT 116.115 95.085 116.365 95.565 ;
        RECT 116.545 95.280 116.805 95.735 ;
        RECT 116.975 95.085 117.220 95.565 ;
        RECT 117.390 95.280 117.665 95.735 ;
        RECT 117.835 95.085 118.080 95.565 ;
        RECT 118.250 95.280 118.510 95.735 ;
        RECT 118.680 95.085 118.940 95.565 ;
        RECT 119.110 95.280 119.370 95.735 ;
        RECT 119.540 95.085 119.800 95.565 ;
        RECT 119.970 95.280 120.230 95.735 ;
        RECT 120.400 95.085 120.660 95.645 ;
        RECT 120.830 95.265 121.080 96.075 ;
        RECT 121.260 95.085 121.520 95.610 ;
        RECT 121.690 95.265 121.940 96.075 ;
        RECT 122.110 95.765 122.425 96.325 ;
        RECT 123.075 95.975 123.305 96.665 ;
        RECT 123.485 96.165 123.825 96.845 ;
        RECT 124.015 96.345 124.345 97.455 ;
        RECT 124.515 96.725 124.705 97.455 ;
        RECT 124.875 96.905 125.205 97.635 ;
        RECT 125.385 96.725 125.555 97.455 ;
        RECT 124.515 96.525 125.555 96.725 ;
        RECT 126.735 96.495 127.005 97.465 ;
        RECT 127.215 96.835 127.495 97.635 ;
        RECT 127.675 97.085 128.870 97.415 ;
        RECT 128.000 96.665 128.420 96.915 ;
        RECT 127.175 96.495 128.420 96.665 ;
        RECT 123.485 95.715 123.715 96.165 ;
        RECT 124.015 96.045 124.550 96.345 ;
        RECT 122.120 95.085 122.425 95.595 ;
        RECT 123.335 95.265 123.715 95.715 ;
        RECT 123.895 95.085 124.125 95.865 ;
        RECT 124.305 95.795 124.550 96.045 ;
        RECT 124.730 95.995 125.125 96.345 ;
        RECT 125.320 95.995 125.610 96.345 ;
        RECT 124.305 95.265 124.735 95.795 ;
        RECT 124.915 95.375 125.125 95.995 ;
        RECT 125.295 95.085 125.625 95.815 ;
        RECT 126.735 95.760 126.905 96.495 ;
        RECT 127.175 96.325 127.345 96.495 ;
        RECT 128.645 96.325 128.815 96.885 ;
        RECT 129.065 96.495 129.320 97.635 ;
        RECT 129.500 96.835 129.755 97.635 ;
        RECT 129.955 96.785 130.285 97.465 ;
        RECT 127.115 95.995 127.345 96.325 ;
        RECT 128.075 95.995 128.815 96.325 ;
        RECT 128.985 96.075 129.320 96.325 ;
        RECT 129.500 96.295 129.745 96.655 ;
        RECT 129.935 96.505 130.285 96.785 ;
        RECT 129.935 96.125 130.105 96.505 ;
        RECT 130.465 96.325 130.660 97.375 ;
        RECT 130.840 96.495 131.160 97.635 ;
        RECT 131.335 96.545 133.925 97.635 ;
        RECT 127.175 95.825 127.345 95.995 ;
        RECT 128.565 95.905 128.815 95.995 ;
        RECT 129.585 95.955 130.105 96.125 ;
        RECT 130.275 95.995 130.660 96.325 ;
        RECT 130.840 96.275 131.100 96.325 ;
        RECT 130.840 96.105 131.105 96.275 ;
        RECT 130.840 95.995 131.100 96.105 ;
        RECT 126.735 95.415 127.005 95.760 ;
        RECT 127.175 95.655 127.915 95.825 ;
        RECT 128.565 95.735 129.300 95.905 ;
        RECT 127.195 95.085 127.575 95.485 ;
        RECT 127.745 95.305 127.915 95.655 ;
        RECT 128.085 95.085 128.820 95.565 ;
        RECT 128.990 95.265 129.300 95.735 ;
        RECT 129.585 95.595 129.755 95.955 ;
        RECT 131.335 95.855 132.545 96.375 ;
        RECT 132.715 96.025 133.925 96.545 ;
        RECT 134.565 96.685 134.840 97.455 ;
        RECT 135.010 97.025 135.340 97.455 ;
        RECT 135.510 97.195 135.705 97.635 ;
        RECT 135.885 97.025 136.215 97.455 ;
        RECT 135.010 96.855 136.215 97.025 ;
        RECT 134.565 96.495 135.150 96.685 ;
        RECT 135.320 96.525 136.215 96.855 ;
        RECT 137.315 96.495 137.595 97.635 ;
        RECT 129.555 95.425 129.755 95.595 ;
        RECT 129.585 95.390 129.755 95.425 ;
        RECT 129.945 95.615 131.160 95.785 ;
        RECT 129.945 95.310 130.175 95.615 ;
        RECT 130.345 95.085 130.675 95.445 ;
        RECT 130.870 95.265 131.160 95.615 ;
        RECT 131.335 95.085 133.925 95.855 ;
        RECT 134.565 95.675 134.805 96.325 ;
        RECT 134.975 95.825 135.150 96.495 ;
        RECT 137.765 96.485 138.095 97.465 ;
        RECT 138.265 96.495 138.525 97.635 ;
        RECT 135.320 95.995 135.735 96.325 ;
        RECT 135.915 95.995 136.210 96.325 ;
        RECT 137.325 96.055 137.660 96.325 ;
        RECT 134.975 95.645 135.305 95.825 ;
        RECT 134.580 95.085 134.910 95.475 ;
        RECT 135.080 95.265 135.305 95.645 ;
        RECT 135.505 95.375 135.735 95.995 ;
        RECT 137.830 95.885 138.000 96.485 ;
        RECT 138.695 96.470 138.985 97.635 ;
        RECT 139.160 96.495 139.480 97.635 ;
        RECT 139.660 96.325 139.855 97.375 ;
        RECT 140.035 96.785 140.365 97.465 ;
        RECT 140.565 96.835 140.820 97.635 ;
        RECT 140.035 96.505 140.385 96.785 ;
        RECT 138.170 96.075 138.505 96.325 ;
        RECT 139.220 96.275 139.480 96.325 ;
        RECT 139.215 96.105 139.480 96.275 ;
        RECT 139.220 95.995 139.480 96.105 ;
        RECT 139.660 95.995 140.045 96.325 ;
        RECT 140.215 96.125 140.385 96.505 ;
        RECT 140.575 96.295 140.820 96.655 ;
        RECT 140.995 96.495 141.255 97.635 ;
        RECT 141.425 96.485 141.755 97.465 ;
        RECT 141.925 96.495 142.205 97.635 ;
        RECT 142.375 96.545 143.585 97.635 ;
        RECT 143.845 97.015 144.015 97.445 ;
        RECT 144.185 97.185 144.515 97.635 ;
        RECT 143.845 96.785 144.520 97.015 ;
        RECT 140.215 95.955 140.735 96.125 ;
        RECT 141.015 96.075 141.350 96.325 ;
        RECT 135.915 95.085 136.215 95.815 ;
        RECT 137.315 95.085 137.625 95.885 ;
        RECT 137.830 95.255 138.525 95.885 ;
        RECT 138.695 95.085 138.985 95.810 ;
        RECT 139.160 95.615 140.375 95.785 ;
        RECT 139.160 95.265 139.450 95.615 ;
        RECT 139.645 95.085 139.975 95.445 ;
        RECT 140.145 95.310 140.375 95.615 ;
        RECT 140.565 95.390 140.735 95.955 ;
        RECT 141.520 95.885 141.690 96.485 ;
        RECT 141.860 96.055 142.195 96.325 ;
        RECT 140.995 95.255 141.690 95.885 ;
        RECT 141.895 95.085 142.205 95.885 ;
        RECT 142.375 95.835 142.895 96.375 ;
        RECT 143.065 96.005 143.585 96.545 ;
        RECT 142.375 95.085 143.585 95.835 ;
        RECT 143.815 95.765 144.115 96.615 ;
        RECT 144.285 96.135 144.520 96.785 ;
        RECT 144.690 96.475 144.975 97.420 ;
        RECT 145.155 97.165 145.840 97.635 ;
        RECT 145.150 96.645 145.845 96.955 ;
        RECT 146.020 96.580 146.325 97.365 ;
        RECT 147.175 96.965 147.455 97.635 ;
        RECT 147.625 96.745 147.925 97.295 ;
        RECT 148.125 96.915 148.455 97.635 ;
        RECT 148.645 96.915 149.105 97.465 ;
        RECT 149.275 97.200 154.620 97.635 ;
        RECT 144.690 96.325 145.550 96.475 ;
        RECT 144.690 96.305 145.975 96.325 ;
        RECT 144.285 95.805 144.820 96.135 ;
        RECT 144.990 95.945 145.975 96.305 ;
        RECT 144.285 95.655 144.505 95.805 ;
        RECT 143.760 95.085 144.095 95.590 ;
        RECT 144.265 95.280 144.505 95.655 ;
        RECT 144.990 95.610 145.160 95.945 ;
        RECT 146.150 95.775 146.325 96.580 ;
        RECT 146.990 96.325 147.255 96.685 ;
        RECT 147.625 96.575 148.565 96.745 ;
        RECT 148.395 96.325 148.565 96.575 ;
        RECT 146.990 96.075 147.665 96.325 ;
        RECT 147.885 96.075 148.225 96.325 ;
        RECT 148.395 95.995 148.685 96.325 ;
        RECT 148.395 95.905 148.565 95.995 ;
        RECT 144.785 95.415 145.160 95.610 ;
        RECT 144.785 95.270 144.955 95.415 ;
        RECT 145.520 95.085 145.915 95.580 ;
        RECT 146.085 95.255 146.325 95.775 ;
        RECT 147.175 95.715 148.565 95.905 ;
        RECT 147.175 95.355 147.505 95.715 ;
        RECT 148.855 95.545 149.105 96.915 ;
        RECT 150.860 95.630 151.200 96.460 ;
        RECT 152.680 95.950 153.030 97.200 ;
        RECT 155.715 96.545 156.925 97.635 ;
        RECT 155.715 96.005 156.235 96.545 ;
        RECT 156.405 95.835 156.925 96.375 ;
        RECT 148.125 95.085 148.375 95.545 ;
        RECT 148.545 95.255 149.105 95.545 ;
        RECT 149.275 95.085 154.620 95.630 ;
        RECT 155.715 95.085 156.925 95.835 ;
        RECT 22.690 94.915 157.010 95.085 ;
        RECT 22.775 94.165 23.985 94.915 ;
        RECT 24.155 94.370 29.500 94.915 ;
        RECT 22.775 93.625 23.295 94.165 ;
        RECT 23.465 93.455 23.985 93.995 ;
        RECT 25.740 93.540 26.080 94.370 ;
        RECT 29.675 94.145 32.265 94.915 ;
        RECT 32.525 94.235 32.695 94.610 ;
        RECT 22.775 92.365 23.985 93.455 ;
        RECT 27.560 92.800 27.910 94.050 ;
        RECT 29.675 93.625 30.885 94.145 ;
        RECT 32.495 94.065 32.695 94.235 ;
        RECT 32.885 94.385 33.115 94.690 ;
        RECT 33.285 94.555 33.615 94.915 ;
        RECT 33.810 94.385 34.100 94.735 ;
        RECT 34.300 94.525 34.630 94.915 ;
        RECT 32.885 94.215 34.100 94.385 ;
        RECT 34.800 94.355 35.025 94.735 ;
        RECT 32.525 94.045 32.695 94.065 ;
        RECT 31.055 93.455 32.265 93.975 ;
        RECT 32.525 93.875 33.045 94.045 ;
        RECT 24.155 92.365 29.500 92.800 ;
        RECT 29.675 92.365 32.265 93.455 ;
        RECT 32.440 93.345 32.685 93.705 ;
        RECT 32.875 93.495 33.045 93.875 ;
        RECT 33.215 93.675 33.600 94.005 ;
        RECT 33.780 93.895 34.040 94.005 ;
        RECT 33.780 93.725 34.045 93.895 ;
        RECT 33.780 93.675 34.040 93.725 ;
        RECT 34.285 93.675 34.525 94.325 ;
        RECT 34.695 94.175 35.025 94.355 ;
        RECT 32.875 93.215 33.225 93.495 ;
        RECT 32.440 92.365 32.695 93.165 ;
        RECT 32.895 92.535 33.225 93.215 ;
        RECT 33.405 92.625 33.600 93.675 ;
        RECT 34.695 93.505 34.870 94.175 ;
        RECT 35.225 94.005 35.455 94.625 ;
        RECT 35.635 94.185 35.935 94.915 ;
        RECT 36.150 94.175 36.765 94.745 ;
        RECT 36.935 94.405 37.150 94.915 ;
        RECT 37.380 94.405 37.660 94.735 ;
        RECT 37.840 94.405 38.080 94.915 ;
        RECT 35.040 93.675 35.455 94.005 ;
        RECT 35.635 93.675 35.930 94.005 ;
        RECT 33.780 92.365 34.100 93.505 ;
        RECT 34.285 93.315 34.870 93.505 ;
        RECT 34.285 92.545 34.560 93.315 ;
        RECT 35.040 93.145 35.935 93.475 ;
        RECT 34.730 92.975 35.935 93.145 ;
        RECT 34.730 92.545 35.060 92.975 ;
        RECT 35.230 92.365 35.425 92.805 ;
        RECT 35.605 92.545 35.935 92.975 ;
        RECT 36.150 93.155 36.465 94.175 ;
        RECT 36.635 93.505 36.805 94.005 ;
        RECT 37.055 93.675 37.320 94.235 ;
        RECT 37.490 93.505 37.660 94.405 ;
        RECT 37.830 93.675 38.185 94.235 ;
        RECT 38.910 94.175 39.525 94.745 ;
        RECT 39.695 94.405 39.910 94.915 ;
        RECT 40.140 94.405 40.420 94.735 ;
        RECT 40.600 94.405 40.840 94.915 ;
        RECT 36.635 93.335 38.060 93.505 ;
        RECT 36.150 92.535 36.685 93.155 ;
        RECT 36.855 92.365 37.185 93.165 ;
        RECT 37.670 93.160 38.060 93.335 ;
        RECT 38.910 93.155 39.225 94.175 ;
        RECT 39.395 93.505 39.565 94.005 ;
        RECT 39.815 93.675 40.080 94.235 ;
        RECT 40.250 93.505 40.420 94.405 ;
        RECT 40.590 93.675 40.945 94.235 ;
        RECT 41.175 94.175 41.640 94.720 ;
        RECT 39.395 93.335 40.820 93.505 ;
        RECT 38.910 92.535 39.445 93.155 ;
        RECT 39.615 92.365 39.945 93.165 ;
        RECT 40.430 93.160 40.820 93.335 ;
        RECT 41.175 93.215 41.345 94.175 ;
        RECT 42.145 94.095 42.315 94.915 ;
        RECT 42.485 94.265 42.815 94.745 ;
        RECT 42.985 94.525 43.335 94.915 ;
        RECT 43.505 94.345 43.735 94.745 ;
        RECT 43.225 94.265 43.735 94.345 ;
        RECT 42.485 94.175 43.735 94.265 ;
        RECT 43.905 94.175 44.225 94.655 ;
        RECT 42.485 94.095 43.395 94.175 ;
        RECT 41.515 93.555 41.760 94.005 ;
        RECT 42.020 93.725 42.715 93.925 ;
        RECT 42.885 93.755 43.485 93.925 ;
        RECT 42.885 93.555 43.055 93.755 ;
        RECT 43.715 93.585 43.885 94.005 ;
        RECT 41.515 93.385 43.055 93.555 ;
        RECT 43.225 93.415 43.885 93.585 ;
        RECT 43.225 93.215 43.395 93.415 ;
        RECT 44.055 93.245 44.225 94.175 ;
        RECT 44.395 94.115 45.090 94.745 ;
        RECT 45.295 94.115 45.605 94.915 ;
        RECT 45.775 94.455 46.335 94.745 ;
        RECT 46.505 94.455 46.755 94.915 ;
        RECT 44.415 93.675 44.750 93.925 ;
        RECT 44.920 93.515 45.090 94.115 ;
        RECT 45.260 93.675 45.595 93.945 ;
        RECT 41.175 93.045 43.395 93.215 ;
        RECT 43.565 93.045 44.225 93.245 ;
        RECT 41.175 92.365 41.475 92.875 ;
        RECT 41.645 92.535 41.975 93.045 ;
        RECT 43.565 92.875 43.735 93.045 ;
        RECT 42.145 92.365 42.775 92.875 ;
        RECT 43.355 92.705 43.735 92.875 ;
        RECT 43.905 92.365 44.205 92.875 ;
        RECT 44.395 92.365 44.655 93.505 ;
        RECT 44.825 92.535 45.155 93.515 ;
        RECT 45.325 92.365 45.605 93.505 ;
        RECT 45.775 93.085 46.025 94.455 ;
        RECT 47.375 94.285 47.705 94.645 ;
        RECT 46.315 94.095 47.705 94.285 ;
        RECT 48.535 94.190 48.825 94.915 ;
        RECT 48.995 94.145 51.585 94.915 ;
        RECT 51.755 94.240 52.015 94.745 ;
        RECT 52.195 94.535 52.525 94.915 ;
        RECT 52.705 94.365 52.875 94.745 ;
        RECT 46.315 94.005 46.485 94.095 ;
        RECT 46.195 93.675 46.485 94.005 ;
        RECT 46.655 93.675 46.995 93.925 ;
        RECT 47.215 93.675 47.890 93.925 ;
        RECT 46.315 93.425 46.485 93.675 ;
        RECT 46.315 93.255 47.255 93.425 ;
        RECT 47.625 93.315 47.890 93.675 ;
        RECT 48.995 93.625 50.205 94.145 ;
        RECT 45.775 92.535 46.235 93.085 ;
        RECT 46.425 92.365 46.755 93.085 ;
        RECT 46.955 92.705 47.255 93.255 ;
        RECT 47.425 92.365 47.705 93.035 ;
        RECT 48.535 92.365 48.825 93.530 ;
        RECT 50.375 93.455 51.585 93.975 ;
        RECT 48.995 92.365 51.585 93.455 ;
        RECT 51.755 93.440 51.925 94.240 ;
        RECT 52.210 94.195 52.875 94.365 ;
        RECT 53.135 94.455 53.695 94.745 ;
        RECT 53.865 94.455 54.115 94.915 ;
        RECT 52.210 93.940 52.380 94.195 ;
        RECT 52.095 93.610 52.380 93.940 ;
        RECT 52.615 93.645 52.945 94.015 ;
        RECT 52.210 93.465 52.380 93.610 ;
        RECT 51.755 92.535 52.025 93.440 ;
        RECT 52.210 93.295 52.875 93.465 ;
        RECT 52.195 92.365 52.525 93.125 ;
        RECT 52.705 92.535 52.875 93.295 ;
        RECT 53.135 93.085 53.385 94.455 ;
        RECT 54.735 94.285 55.065 94.645 ;
        RECT 55.435 94.370 60.780 94.915 ;
        RECT 60.955 94.370 66.300 94.915 ;
        RECT 53.675 94.095 55.065 94.285 ;
        RECT 53.675 94.005 53.845 94.095 ;
        RECT 53.555 93.675 53.845 94.005 ;
        RECT 54.015 93.675 54.355 93.925 ;
        RECT 54.575 93.675 55.250 93.925 ;
        RECT 53.675 93.425 53.845 93.675 ;
        RECT 53.675 93.255 54.615 93.425 ;
        RECT 54.985 93.315 55.250 93.675 ;
        RECT 57.020 93.540 57.360 94.370 ;
        RECT 53.135 92.535 53.595 93.085 ;
        RECT 53.785 92.365 54.115 93.085 ;
        RECT 54.315 92.705 54.615 93.255 ;
        RECT 54.785 92.365 55.065 93.035 ;
        RECT 58.840 92.800 59.190 94.050 ;
        RECT 62.540 93.540 62.880 94.370 ;
        RECT 67.395 94.240 67.655 94.745 ;
        RECT 67.835 94.535 68.165 94.915 ;
        RECT 68.345 94.365 68.515 94.745 ;
        RECT 68.775 94.370 74.120 94.915 ;
        RECT 64.360 92.800 64.710 94.050 ;
        RECT 67.395 93.440 67.565 94.240 ;
        RECT 67.850 94.195 68.515 94.365 ;
        RECT 67.850 93.940 68.020 94.195 ;
        RECT 67.735 93.610 68.020 93.940 ;
        RECT 68.255 93.645 68.585 94.015 ;
        RECT 67.850 93.465 68.020 93.610 ;
        RECT 70.360 93.540 70.700 94.370 ;
        RECT 74.295 94.190 74.585 94.915 ;
        RECT 74.755 94.145 77.345 94.915 ;
        RECT 77.795 94.285 78.175 94.735 ;
        RECT 55.435 92.365 60.780 92.800 ;
        RECT 60.955 92.365 66.300 92.800 ;
        RECT 67.395 92.535 67.665 93.440 ;
        RECT 67.850 93.295 68.515 93.465 ;
        RECT 67.835 92.365 68.165 93.125 ;
        RECT 68.345 92.535 68.515 93.295 ;
        RECT 72.180 92.800 72.530 94.050 ;
        RECT 74.755 93.625 75.965 94.145 ;
        RECT 68.775 92.365 74.120 92.800 ;
        RECT 74.295 92.365 74.585 93.530 ;
        RECT 76.135 93.455 77.345 93.975 ;
        RECT 74.755 92.365 77.345 93.455 ;
        RECT 77.535 93.335 77.765 94.025 ;
        RECT 77.945 93.835 78.175 94.285 ;
        RECT 78.355 94.135 78.585 94.915 ;
        RECT 78.765 94.205 79.195 94.735 ;
        RECT 78.765 93.955 79.010 94.205 ;
        RECT 79.375 94.005 79.585 94.625 ;
        RECT 79.755 94.185 80.085 94.915 ;
        RECT 77.945 93.155 78.285 93.835 ;
        RECT 77.525 92.955 78.285 93.155 ;
        RECT 78.475 93.655 79.010 93.955 ;
        RECT 79.190 93.655 79.585 94.005 ;
        RECT 79.780 93.655 80.070 94.005 ;
        RECT 77.525 92.565 77.785 92.955 ;
        RECT 77.955 92.365 78.285 92.775 ;
        RECT 78.475 92.545 78.805 93.655 ;
        RECT 78.975 93.275 80.015 93.475 ;
        RECT 78.975 92.545 79.165 93.275 ;
        RECT 79.335 92.365 79.665 93.095 ;
        RECT 79.845 92.545 80.015 93.275 ;
        RECT 80.280 93.315 80.615 94.735 ;
        RECT 80.795 94.545 81.540 94.915 ;
        RECT 82.105 94.375 82.360 94.735 ;
        RECT 82.540 94.545 82.870 94.915 ;
        RECT 83.050 94.375 83.275 94.735 ;
        RECT 80.790 94.185 83.275 94.375 ;
        RECT 83.495 94.370 88.840 94.915 ;
        RECT 80.790 93.495 81.015 94.185 ;
        RECT 81.215 93.675 81.495 94.005 ;
        RECT 81.675 93.675 82.250 94.005 ;
        RECT 82.430 93.675 82.865 94.005 ;
        RECT 83.045 93.675 83.315 94.005 ;
        RECT 85.080 93.540 85.420 94.370 ;
        RECT 89.480 94.095 89.775 94.915 ;
        RECT 89.945 94.365 90.165 94.745 ;
        RECT 90.335 94.555 91.185 94.915 ;
        RECT 80.790 93.315 83.285 93.495 ;
        RECT 80.280 92.545 80.545 93.315 ;
        RECT 80.715 92.365 81.045 93.085 ;
        RECT 81.235 92.905 82.425 93.135 ;
        RECT 81.235 92.545 81.495 92.905 ;
        RECT 81.665 92.365 81.995 92.735 ;
        RECT 82.165 92.545 82.425 92.905 ;
        RECT 82.995 92.545 83.285 93.315 ;
        RECT 86.900 92.800 87.250 94.050 ;
        RECT 83.495 92.365 88.840 92.800 ;
        RECT 89.480 92.365 89.775 93.510 ;
        RECT 89.945 92.665 90.175 94.365 ;
        RECT 91.665 94.305 91.995 94.725 ;
        RECT 92.200 94.475 92.475 94.915 ;
        RECT 92.645 94.305 92.975 94.725 ;
        RECT 90.390 94.125 92.975 94.305 ;
        RECT 93.155 94.175 93.620 94.720 ;
        RECT 90.390 93.510 90.700 94.125 ;
        RECT 90.870 93.725 91.200 93.955 ;
        RECT 91.370 93.725 91.840 93.955 ;
        RECT 92.010 93.895 92.460 93.955 ;
        RECT 92.010 93.725 92.465 93.895 ;
        RECT 92.650 93.725 92.985 93.955 ;
        RECT 90.390 93.340 92.975 93.510 ;
        RECT 90.390 92.365 90.645 93.170 ;
        RECT 90.845 92.980 92.185 93.160 ;
        RECT 90.845 92.535 91.175 92.980 ;
        RECT 91.345 92.365 91.620 92.810 ;
        RECT 91.855 92.535 92.185 92.980 ;
        RECT 92.645 92.675 92.975 93.340 ;
        RECT 93.155 93.215 93.325 94.175 ;
        RECT 94.125 94.095 94.295 94.915 ;
        RECT 94.465 94.265 94.795 94.745 ;
        RECT 94.965 94.525 95.315 94.915 ;
        RECT 95.485 94.345 95.715 94.745 ;
        RECT 95.205 94.265 95.715 94.345 ;
        RECT 94.465 94.175 95.715 94.265 ;
        RECT 95.885 94.175 96.205 94.655 ;
        RECT 94.465 94.095 95.375 94.175 ;
        RECT 93.495 93.555 93.740 94.005 ;
        RECT 94.000 93.725 94.695 93.925 ;
        RECT 94.865 93.755 95.465 93.925 ;
        RECT 94.865 93.555 95.035 93.755 ;
        RECT 95.695 93.585 95.865 94.005 ;
        RECT 93.495 93.385 95.035 93.555 ;
        RECT 95.205 93.415 95.865 93.585 ;
        RECT 95.205 93.215 95.375 93.415 ;
        RECT 96.035 93.245 96.205 94.175 ;
        RECT 93.155 93.045 95.375 93.215 ;
        RECT 95.545 93.045 96.205 93.245 ;
        RECT 96.375 94.175 96.840 94.720 ;
        RECT 96.375 93.215 96.545 94.175 ;
        RECT 97.345 94.095 97.515 94.915 ;
        RECT 97.685 94.265 98.015 94.745 ;
        RECT 98.185 94.525 98.535 94.915 ;
        RECT 98.705 94.345 98.935 94.745 ;
        RECT 98.425 94.265 98.935 94.345 ;
        RECT 97.685 94.175 98.935 94.265 ;
        RECT 99.105 94.175 99.425 94.655 ;
        RECT 100.055 94.190 100.345 94.915 ;
        RECT 100.565 94.260 100.895 94.695 ;
        RECT 101.065 94.305 101.235 94.915 ;
        RECT 97.685 94.095 98.595 94.175 ;
        RECT 96.715 93.555 96.960 94.005 ;
        RECT 97.220 93.725 97.915 93.925 ;
        RECT 98.085 93.755 98.685 93.925 ;
        RECT 98.085 93.555 98.255 93.755 ;
        RECT 98.915 93.585 99.085 94.005 ;
        RECT 96.715 93.385 98.255 93.555 ;
        RECT 98.425 93.415 99.085 93.585 ;
        RECT 98.425 93.215 98.595 93.415 ;
        RECT 99.255 93.245 99.425 94.175 ;
        RECT 100.515 94.175 100.895 94.260 ;
        RECT 101.405 94.175 101.735 94.700 ;
        RECT 101.995 94.385 102.205 94.915 ;
        RECT 102.480 94.465 103.265 94.635 ;
        RECT 103.435 94.465 103.840 94.635 ;
        RECT 100.515 94.135 100.740 94.175 ;
        RECT 100.515 93.555 100.685 94.135 ;
        RECT 101.405 94.005 101.605 94.175 ;
        RECT 102.480 94.005 102.650 94.465 ;
        RECT 100.855 93.675 101.605 94.005 ;
        RECT 101.775 93.675 102.650 94.005 ;
        RECT 96.375 93.045 98.595 93.215 ;
        RECT 98.765 93.045 99.425 93.245 ;
        RECT 93.155 92.365 93.455 92.875 ;
        RECT 93.625 92.535 93.955 93.045 ;
        RECT 95.545 92.875 95.715 93.045 ;
        RECT 94.125 92.365 94.755 92.875 ;
        RECT 95.335 92.705 95.715 92.875 ;
        RECT 95.885 92.365 96.185 92.875 ;
        RECT 96.375 92.365 96.675 92.875 ;
        RECT 96.845 92.535 97.175 93.045 ;
        RECT 98.765 92.875 98.935 93.045 ;
        RECT 97.345 92.365 97.975 92.875 ;
        RECT 98.555 92.705 98.935 92.875 ;
        RECT 99.105 92.365 99.405 92.875 ;
        RECT 100.055 92.365 100.345 93.530 ;
        RECT 100.515 93.505 100.730 93.555 ;
        RECT 100.515 93.425 100.905 93.505 ;
        RECT 100.575 92.580 100.905 93.425 ;
        RECT 101.415 93.470 101.605 93.675 ;
        RECT 101.075 92.365 101.245 93.375 ;
        RECT 101.415 93.095 102.310 93.470 ;
        RECT 101.415 92.535 101.755 93.095 ;
        RECT 101.985 92.365 102.300 92.865 ;
        RECT 102.480 92.835 102.650 93.675 ;
        RECT 102.820 93.965 103.285 94.295 ;
        RECT 103.670 94.235 103.840 94.465 ;
        RECT 104.020 94.415 104.390 94.915 ;
        RECT 104.710 94.465 105.385 94.635 ;
        RECT 105.580 94.465 105.915 94.635 ;
        RECT 102.820 93.005 103.140 93.965 ;
        RECT 103.670 93.935 104.500 94.235 ;
        RECT 103.310 93.035 103.500 93.755 ;
        RECT 103.670 92.865 103.840 93.935 ;
        RECT 104.300 93.905 104.500 93.935 ;
        RECT 104.010 93.685 104.180 93.755 ;
        RECT 104.710 93.685 104.880 94.465 ;
        RECT 105.745 94.325 105.915 94.465 ;
        RECT 106.085 94.455 106.335 94.915 ;
        RECT 104.010 93.515 104.880 93.685 ;
        RECT 105.050 94.045 105.575 94.265 ;
        RECT 105.745 94.195 105.970 94.325 ;
        RECT 104.010 93.425 104.520 93.515 ;
        RECT 102.480 92.665 103.365 92.835 ;
        RECT 103.590 92.535 103.840 92.865 ;
        RECT 104.010 92.365 104.180 93.165 ;
        RECT 104.350 92.810 104.520 93.425 ;
        RECT 105.050 93.345 105.220 94.045 ;
        RECT 104.690 92.980 105.220 93.345 ;
        RECT 105.390 93.280 105.630 93.875 ;
        RECT 105.800 93.090 105.970 94.195 ;
        RECT 106.140 93.335 106.420 94.285 ;
        RECT 105.665 92.960 105.970 93.090 ;
        RECT 104.350 92.640 105.455 92.810 ;
        RECT 105.665 92.535 105.915 92.960 ;
        RECT 106.085 92.365 106.350 92.825 ;
        RECT 106.590 92.535 106.775 94.655 ;
        RECT 106.945 94.535 107.275 94.915 ;
        RECT 107.445 94.365 107.615 94.655 ;
        RECT 106.950 94.195 107.615 94.365 ;
        RECT 107.925 94.260 108.255 94.695 ;
        RECT 108.425 94.305 108.595 94.915 ;
        RECT 106.950 93.205 107.180 94.195 ;
        RECT 107.875 94.175 108.255 94.260 ;
        RECT 108.765 94.175 109.095 94.700 ;
        RECT 109.355 94.385 109.565 94.915 ;
        RECT 109.840 94.465 110.625 94.635 ;
        RECT 110.795 94.465 111.200 94.635 ;
        RECT 107.875 94.135 108.100 94.175 ;
        RECT 107.350 93.375 107.700 94.025 ;
        RECT 107.875 93.555 108.045 94.135 ;
        RECT 108.765 94.005 108.965 94.175 ;
        RECT 109.840 94.005 110.010 94.465 ;
        RECT 108.215 93.675 108.965 94.005 ;
        RECT 109.135 93.675 110.010 94.005 ;
        RECT 107.875 93.505 108.090 93.555 ;
        RECT 107.875 93.425 108.265 93.505 ;
        RECT 106.950 93.035 107.615 93.205 ;
        RECT 106.945 92.365 107.275 92.865 ;
        RECT 107.445 92.535 107.615 93.035 ;
        RECT 107.935 92.580 108.265 93.425 ;
        RECT 108.775 93.470 108.965 93.675 ;
        RECT 108.435 92.365 108.605 93.375 ;
        RECT 108.775 93.095 109.670 93.470 ;
        RECT 108.775 92.535 109.115 93.095 ;
        RECT 109.345 92.365 109.660 92.865 ;
        RECT 109.840 92.835 110.010 93.675 ;
        RECT 110.180 93.965 110.645 94.295 ;
        RECT 111.030 94.235 111.200 94.465 ;
        RECT 111.380 94.415 111.750 94.915 ;
        RECT 112.070 94.465 112.745 94.635 ;
        RECT 112.940 94.465 113.275 94.635 ;
        RECT 110.180 93.005 110.500 93.965 ;
        RECT 111.030 93.935 111.860 94.235 ;
        RECT 110.670 93.035 110.860 93.755 ;
        RECT 111.030 92.865 111.200 93.935 ;
        RECT 111.660 93.905 111.860 93.935 ;
        RECT 111.370 93.685 111.540 93.755 ;
        RECT 112.070 93.685 112.240 94.465 ;
        RECT 113.105 94.325 113.275 94.465 ;
        RECT 113.445 94.455 113.695 94.915 ;
        RECT 111.370 93.515 112.240 93.685 ;
        RECT 112.410 94.045 112.935 94.265 ;
        RECT 113.105 94.195 113.330 94.325 ;
        RECT 111.370 93.425 111.880 93.515 ;
        RECT 109.840 92.665 110.725 92.835 ;
        RECT 110.950 92.535 111.200 92.865 ;
        RECT 111.370 92.365 111.540 93.165 ;
        RECT 111.710 92.810 111.880 93.425 ;
        RECT 112.410 93.345 112.580 94.045 ;
        RECT 112.050 92.980 112.580 93.345 ;
        RECT 112.750 93.280 112.990 93.875 ;
        RECT 113.160 93.090 113.330 94.195 ;
        RECT 113.500 93.335 113.780 94.285 ;
        RECT 113.025 92.960 113.330 93.090 ;
        RECT 111.710 92.640 112.815 92.810 ;
        RECT 113.025 92.535 113.275 92.960 ;
        RECT 113.445 92.365 113.710 92.825 ;
        RECT 113.950 92.535 114.135 94.655 ;
        RECT 114.305 94.535 114.635 94.915 ;
        RECT 114.805 94.365 114.975 94.655 ;
        RECT 114.310 94.195 114.975 94.365 ;
        RECT 115.285 94.375 115.510 94.735 ;
        RECT 115.690 94.545 116.020 94.915 ;
        RECT 116.200 94.375 116.455 94.735 ;
        RECT 117.020 94.545 117.765 94.915 ;
        RECT 114.310 93.205 114.540 94.195 ;
        RECT 115.285 94.185 117.770 94.375 ;
        RECT 114.710 93.375 115.060 94.025 ;
        RECT 115.245 93.675 115.515 94.005 ;
        RECT 115.695 93.675 116.130 94.005 ;
        RECT 116.310 93.675 116.885 94.005 ;
        RECT 117.065 93.675 117.345 94.005 ;
        RECT 117.545 93.495 117.770 94.185 ;
        RECT 115.275 93.315 117.770 93.495 ;
        RECT 117.945 93.315 118.280 94.735 ;
        RECT 118.545 94.365 118.715 94.655 ;
        RECT 118.885 94.535 119.215 94.915 ;
        RECT 118.545 94.195 119.210 94.365 ;
        RECT 118.460 93.375 118.810 94.025 ;
        RECT 114.310 93.035 114.975 93.205 ;
        RECT 114.305 92.365 114.635 92.865 ;
        RECT 114.805 92.535 114.975 93.035 ;
        RECT 115.275 92.545 115.565 93.315 ;
        RECT 116.135 92.905 117.325 93.135 ;
        RECT 116.135 92.545 116.395 92.905 ;
        RECT 116.565 92.365 116.895 92.735 ;
        RECT 117.065 92.545 117.325 92.905 ;
        RECT 117.515 92.365 117.845 93.085 ;
        RECT 118.015 92.545 118.280 93.315 ;
        RECT 118.980 93.205 119.210 94.195 ;
        RECT 118.545 93.035 119.210 93.205 ;
        RECT 118.545 92.535 118.715 93.035 ;
        RECT 118.885 92.365 119.215 92.865 ;
        RECT 119.385 92.535 119.570 94.655 ;
        RECT 119.825 94.455 120.075 94.915 ;
        RECT 120.245 94.465 120.580 94.635 ;
        RECT 120.775 94.465 121.450 94.635 ;
        RECT 120.245 94.325 120.415 94.465 ;
        RECT 119.740 93.335 120.020 94.285 ;
        RECT 120.190 94.195 120.415 94.325 ;
        RECT 120.190 93.090 120.360 94.195 ;
        RECT 120.585 94.045 121.110 94.265 ;
        RECT 120.530 93.280 120.770 93.875 ;
        RECT 120.940 93.345 121.110 94.045 ;
        RECT 121.280 93.685 121.450 94.465 ;
        RECT 121.770 94.415 122.140 94.915 ;
        RECT 122.320 94.465 122.725 94.635 ;
        RECT 122.895 94.465 123.680 94.635 ;
        RECT 122.320 94.235 122.490 94.465 ;
        RECT 121.660 93.935 122.490 94.235 ;
        RECT 122.875 93.965 123.340 94.295 ;
        RECT 121.660 93.905 121.860 93.935 ;
        RECT 121.980 93.685 122.150 93.755 ;
        RECT 121.280 93.515 122.150 93.685 ;
        RECT 121.640 93.425 122.150 93.515 ;
        RECT 120.190 92.960 120.495 93.090 ;
        RECT 120.940 92.980 121.470 93.345 ;
        RECT 119.810 92.365 120.075 92.825 ;
        RECT 120.245 92.535 120.495 92.960 ;
        RECT 121.640 92.810 121.810 93.425 ;
        RECT 120.705 92.640 121.810 92.810 ;
        RECT 121.980 92.365 122.150 93.165 ;
        RECT 122.320 92.865 122.490 93.935 ;
        RECT 122.660 93.035 122.850 93.755 ;
        RECT 123.020 93.005 123.340 93.965 ;
        RECT 123.510 94.005 123.680 94.465 ;
        RECT 123.955 94.385 124.165 94.915 ;
        RECT 124.425 94.175 124.755 94.700 ;
        RECT 124.925 94.305 125.095 94.915 ;
        RECT 125.265 94.260 125.595 94.695 ;
        RECT 125.265 94.175 125.645 94.260 ;
        RECT 125.815 94.190 126.105 94.915 ;
        RECT 124.555 94.005 124.755 94.175 ;
        RECT 125.420 94.135 125.645 94.175 ;
        RECT 123.510 93.675 124.385 94.005 ;
        RECT 124.555 93.675 125.305 94.005 ;
        RECT 122.320 92.535 122.570 92.865 ;
        RECT 123.510 92.835 123.680 93.675 ;
        RECT 124.555 93.470 124.745 93.675 ;
        RECT 125.475 93.555 125.645 94.135 ;
        RECT 125.430 93.505 125.645 93.555 ;
        RECT 126.275 93.970 126.615 94.745 ;
        RECT 126.785 94.455 126.955 94.915 ;
        RECT 127.195 94.480 127.555 94.745 ;
        RECT 127.195 94.475 127.550 94.480 ;
        RECT 127.195 94.465 127.545 94.475 ;
        RECT 127.195 94.460 127.540 94.465 ;
        RECT 127.195 94.450 127.535 94.460 ;
        RECT 128.185 94.455 128.355 94.915 ;
        RECT 127.195 94.445 127.530 94.450 ;
        RECT 127.195 94.435 127.520 94.445 ;
        RECT 127.195 94.425 127.510 94.435 ;
        RECT 127.195 94.285 127.495 94.425 ;
        RECT 126.785 94.095 127.495 94.285 ;
        RECT 127.685 94.285 128.015 94.365 ;
        RECT 128.525 94.285 128.865 94.745 ;
        RECT 127.685 94.095 128.865 94.285 ;
        RECT 129.055 94.105 129.295 94.915 ;
        RECT 129.465 94.105 129.795 94.745 ;
        RECT 129.965 94.105 130.235 94.915 ;
        RECT 130.415 94.115 130.725 94.915 ;
        RECT 130.930 94.115 131.625 94.745 ;
        RECT 132.740 94.525 133.070 94.915 ;
        RECT 133.240 94.355 133.465 94.735 ;
        RECT 123.850 93.095 124.745 93.470 ;
        RECT 125.255 93.425 125.645 93.505 ;
        RECT 122.795 92.665 123.680 92.835 ;
        RECT 123.860 92.365 124.175 92.865 ;
        RECT 124.405 92.535 124.745 93.095 ;
        RECT 124.915 92.365 125.085 93.375 ;
        RECT 125.255 92.580 125.585 93.425 ;
        RECT 125.815 92.365 126.105 93.530 ;
        RECT 126.275 92.535 126.555 93.970 ;
        RECT 126.785 93.525 127.070 94.095 ;
        RECT 127.255 93.695 127.725 93.925 ;
        RECT 127.895 93.905 128.225 93.925 ;
        RECT 127.895 93.725 128.345 93.905 ;
        RECT 128.535 93.725 128.865 93.925 ;
        RECT 126.785 93.310 127.935 93.525 ;
        RECT 126.725 92.365 127.435 93.140 ;
        RECT 127.605 92.535 127.935 93.310 ;
        RECT 128.130 92.610 128.345 93.725 ;
        RECT 128.635 93.385 128.865 93.725 ;
        RECT 129.035 93.675 129.385 93.925 ;
        RECT 129.555 93.505 129.725 94.105 ;
        RECT 129.895 93.675 130.245 93.925 ;
        RECT 130.425 93.675 130.760 93.945 ;
        RECT 130.930 93.515 131.100 94.115 ;
        RECT 131.270 93.675 131.605 93.925 ;
        RECT 132.725 93.675 132.965 94.325 ;
        RECT 133.135 94.175 133.465 94.355 ;
        RECT 129.045 93.335 129.725 93.505 ;
        RECT 128.525 92.365 128.855 93.085 ;
        RECT 129.045 92.550 129.375 93.335 ;
        RECT 129.905 92.365 130.235 93.505 ;
        RECT 130.415 92.365 130.695 93.505 ;
        RECT 130.865 92.535 131.195 93.515 ;
        RECT 133.135 93.505 133.310 94.175 ;
        RECT 133.665 94.005 133.895 94.625 ;
        RECT 134.075 94.185 134.375 94.915 ;
        RECT 134.645 94.235 134.815 94.610 ;
        RECT 134.615 94.065 134.815 94.235 ;
        RECT 135.005 94.385 135.235 94.690 ;
        RECT 135.405 94.555 135.735 94.915 ;
        RECT 135.930 94.385 136.220 94.735 ;
        RECT 137.480 94.405 137.720 94.915 ;
        RECT 137.900 94.405 138.180 94.735 ;
        RECT 138.410 94.405 138.625 94.915 ;
        RECT 135.005 94.215 136.220 94.385 ;
        RECT 134.645 94.045 134.815 94.065 ;
        RECT 133.480 93.675 133.895 94.005 ;
        RECT 134.075 93.675 134.370 94.005 ;
        RECT 134.645 93.875 135.165 94.045 ;
        RECT 131.365 92.365 131.625 93.505 ;
        RECT 132.725 93.315 133.310 93.505 ;
        RECT 132.725 92.545 133.000 93.315 ;
        RECT 133.480 93.145 134.375 93.475 ;
        RECT 134.560 93.345 134.805 93.705 ;
        RECT 134.995 93.495 135.165 93.875 ;
        RECT 135.335 93.675 135.720 94.005 ;
        RECT 135.900 93.895 136.160 94.005 ;
        RECT 135.900 93.725 136.165 93.895 ;
        RECT 135.900 93.675 136.160 93.725 ;
        RECT 137.375 93.675 137.730 94.235 ;
        RECT 134.995 93.215 135.345 93.495 ;
        RECT 133.170 92.975 134.375 93.145 ;
        RECT 133.170 92.545 133.500 92.975 ;
        RECT 133.670 92.365 133.865 92.805 ;
        RECT 134.045 92.545 134.375 92.975 ;
        RECT 134.560 92.365 134.815 93.165 ;
        RECT 135.015 92.535 135.345 93.215 ;
        RECT 135.525 92.625 135.720 93.675 ;
        RECT 137.900 93.505 138.070 94.405 ;
        RECT 138.240 93.675 138.505 94.235 ;
        RECT 138.795 94.175 139.410 94.745 ;
        RECT 138.755 93.505 138.925 94.005 ;
        RECT 135.900 92.365 136.220 93.505 ;
        RECT 137.500 93.335 138.925 93.505 ;
        RECT 137.500 93.160 137.890 93.335 ;
        RECT 138.375 92.365 138.705 93.165 ;
        RECT 139.095 93.155 139.410 94.175 ;
        RECT 140.085 94.105 140.355 94.915 ;
        RECT 140.525 94.105 140.855 94.745 ;
        RECT 141.025 94.105 141.265 94.915 ;
        RECT 140.075 93.675 140.425 93.925 ;
        RECT 140.595 93.505 140.765 94.105 ;
        RECT 141.455 93.970 141.795 94.745 ;
        RECT 141.965 94.455 142.135 94.915 ;
        RECT 142.375 94.480 142.735 94.745 ;
        RECT 142.375 94.475 142.730 94.480 ;
        RECT 142.375 94.465 142.725 94.475 ;
        RECT 142.375 94.460 142.720 94.465 ;
        RECT 142.375 94.450 142.715 94.460 ;
        RECT 143.365 94.455 143.535 94.915 ;
        RECT 142.375 94.445 142.710 94.450 ;
        RECT 142.375 94.435 142.700 94.445 ;
        RECT 142.375 94.425 142.690 94.435 ;
        RECT 142.375 94.285 142.675 94.425 ;
        RECT 141.965 94.095 142.675 94.285 ;
        RECT 142.865 94.285 143.195 94.365 ;
        RECT 143.705 94.285 144.045 94.745 ;
        RECT 142.865 94.095 144.045 94.285 ;
        RECT 144.265 94.260 144.595 94.695 ;
        RECT 144.765 94.305 144.935 94.915 ;
        RECT 144.215 94.175 144.595 94.260 ;
        RECT 145.105 94.175 145.435 94.700 ;
        RECT 145.695 94.385 145.905 94.915 ;
        RECT 146.180 94.465 146.965 94.635 ;
        RECT 147.135 94.465 147.540 94.635 ;
        RECT 144.215 94.135 144.440 94.175 ;
        RECT 140.935 93.675 141.285 93.925 ;
        RECT 138.875 92.535 139.410 93.155 ;
        RECT 140.085 92.365 140.415 93.505 ;
        RECT 140.595 93.335 141.275 93.505 ;
        RECT 140.945 92.550 141.275 93.335 ;
        RECT 141.455 92.535 141.735 93.970 ;
        RECT 141.965 93.525 142.250 94.095 ;
        RECT 142.435 93.695 142.905 93.925 ;
        RECT 143.075 93.905 143.405 93.925 ;
        RECT 143.075 93.725 143.525 93.905 ;
        RECT 143.715 93.725 144.045 93.925 ;
        RECT 141.965 93.310 143.115 93.525 ;
        RECT 141.905 92.365 142.615 93.140 ;
        RECT 142.785 92.535 143.115 93.310 ;
        RECT 143.310 92.610 143.525 93.725 ;
        RECT 143.815 93.385 144.045 93.725 ;
        RECT 144.215 93.555 144.385 94.135 ;
        RECT 145.105 94.005 145.305 94.175 ;
        RECT 146.180 94.005 146.350 94.465 ;
        RECT 144.555 93.675 145.305 94.005 ;
        RECT 145.475 93.675 146.350 94.005 ;
        RECT 144.215 93.505 144.430 93.555 ;
        RECT 144.215 93.425 144.605 93.505 ;
        RECT 143.705 92.365 144.035 93.085 ;
        RECT 144.275 92.580 144.605 93.425 ;
        RECT 145.115 93.470 145.305 93.675 ;
        RECT 144.775 92.365 144.945 93.375 ;
        RECT 145.115 93.095 146.010 93.470 ;
        RECT 145.115 92.535 145.455 93.095 ;
        RECT 145.685 92.365 146.000 92.865 ;
        RECT 146.180 92.835 146.350 93.675 ;
        RECT 146.520 93.965 146.985 94.295 ;
        RECT 147.370 94.235 147.540 94.465 ;
        RECT 147.720 94.415 148.090 94.915 ;
        RECT 148.410 94.465 149.085 94.635 ;
        RECT 149.280 94.465 149.615 94.635 ;
        RECT 146.520 93.005 146.840 93.965 ;
        RECT 147.370 93.935 148.200 94.235 ;
        RECT 147.010 93.035 147.200 93.755 ;
        RECT 147.370 92.865 147.540 93.935 ;
        RECT 148.000 93.905 148.200 93.935 ;
        RECT 147.710 93.685 147.880 93.755 ;
        RECT 148.410 93.685 148.580 94.465 ;
        RECT 149.445 94.325 149.615 94.465 ;
        RECT 149.785 94.455 150.035 94.915 ;
        RECT 147.710 93.515 148.580 93.685 ;
        RECT 148.750 94.045 149.275 94.265 ;
        RECT 149.445 94.195 149.670 94.325 ;
        RECT 147.710 93.425 148.220 93.515 ;
        RECT 146.180 92.665 147.065 92.835 ;
        RECT 147.290 92.535 147.540 92.865 ;
        RECT 147.710 92.365 147.880 93.165 ;
        RECT 148.050 92.810 148.220 93.425 ;
        RECT 148.750 93.345 148.920 94.045 ;
        RECT 148.390 92.980 148.920 93.345 ;
        RECT 149.090 93.280 149.330 93.875 ;
        RECT 149.500 93.090 149.670 94.195 ;
        RECT 149.840 93.335 150.120 94.285 ;
        RECT 149.365 92.960 149.670 93.090 ;
        RECT 148.050 92.640 149.155 92.810 ;
        RECT 149.365 92.535 149.615 92.960 ;
        RECT 149.785 92.365 150.050 92.825 ;
        RECT 150.290 92.535 150.475 94.655 ;
        RECT 150.645 94.535 150.975 94.915 ;
        RECT 151.145 94.365 151.315 94.655 ;
        RECT 150.650 94.195 151.315 94.365 ;
        RECT 150.650 93.205 150.880 94.195 ;
        RECT 151.575 94.190 151.865 94.915 ;
        RECT 152.035 94.240 152.295 94.745 ;
        RECT 152.475 94.535 152.805 94.915 ;
        RECT 152.985 94.365 153.155 94.745 ;
        RECT 151.050 93.375 151.400 94.025 ;
        RECT 150.650 93.035 151.315 93.205 ;
        RECT 150.645 92.365 150.975 92.865 ;
        RECT 151.145 92.535 151.315 93.035 ;
        RECT 151.575 92.365 151.865 93.530 ;
        RECT 152.035 93.440 152.205 94.240 ;
        RECT 152.490 94.195 153.155 94.365 ;
        RECT 152.490 93.940 152.660 94.195 ;
        RECT 153.415 94.145 155.085 94.915 ;
        RECT 155.715 94.165 156.925 94.915 ;
        RECT 152.375 93.610 152.660 93.940 ;
        RECT 152.895 93.645 153.225 94.015 ;
        RECT 153.415 93.625 154.165 94.145 ;
        RECT 152.490 93.465 152.660 93.610 ;
        RECT 152.035 92.535 152.305 93.440 ;
        RECT 152.490 93.295 153.155 93.465 ;
        RECT 154.335 93.455 155.085 93.975 ;
        RECT 152.475 92.365 152.805 93.125 ;
        RECT 152.985 92.535 153.155 93.295 ;
        RECT 153.415 92.365 155.085 93.455 ;
        RECT 155.715 93.455 156.235 93.995 ;
        RECT 156.405 93.625 156.925 94.165 ;
        RECT 155.715 92.365 156.925 93.455 ;
        RECT 22.690 92.195 157.010 92.365 ;
        RECT 22.775 91.105 23.985 92.195 ;
        RECT 24.155 91.105 26.745 92.195 ;
        RECT 26.925 91.605 27.185 91.995 ;
        RECT 27.355 91.785 27.685 92.195 ;
        RECT 26.925 91.405 27.685 91.605 ;
        RECT 22.775 90.395 23.295 90.935 ;
        RECT 23.465 90.565 23.985 91.105 ;
        RECT 24.155 90.415 25.365 90.935 ;
        RECT 25.535 90.585 26.745 91.105 ;
        RECT 26.935 90.535 27.165 91.225 ;
        RECT 27.345 90.725 27.685 91.405 ;
        RECT 27.875 90.905 28.205 92.015 ;
        RECT 28.375 91.285 28.565 92.015 ;
        RECT 28.735 91.465 29.065 92.195 ;
        RECT 29.245 91.285 29.415 92.015 ;
        RECT 29.695 91.345 30.025 92.195 ;
        RECT 30.195 91.855 31.305 92.025 ;
        RECT 30.195 91.345 30.415 91.855 ;
        RECT 31.115 91.695 31.305 91.855 ;
        RECT 31.500 91.735 31.830 92.195 ;
        RECT 30.585 91.525 30.885 91.685 ;
        RECT 32.000 91.525 32.235 92.025 ;
        RECT 30.585 91.345 32.235 91.525 ;
        RECT 28.375 91.085 29.415 91.285 ;
        RECT 29.710 91.005 31.685 91.175 ;
        RECT 22.775 89.645 23.985 90.395 ;
        RECT 24.155 89.645 26.745 90.415 ;
        RECT 27.345 90.275 27.575 90.725 ;
        RECT 27.875 90.605 28.410 90.905 ;
        RECT 27.195 89.825 27.575 90.275 ;
        RECT 27.755 89.645 27.985 90.425 ;
        RECT 28.165 90.355 28.410 90.605 ;
        RECT 28.590 90.555 28.985 90.905 ;
        RECT 29.180 90.555 29.470 90.905 ;
        RECT 29.710 90.615 30.040 91.005 ;
        RECT 31.190 90.835 31.685 91.005 ;
        RECT 30.210 90.635 31.010 90.835 ;
        RECT 31.190 90.665 31.745 90.835 ;
        RECT 31.190 90.635 31.685 90.665 ;
        RECT 28.165 89.825 28.595 90.355 ;
        RECT 28.775 89.935 28.985 90.555 ;
        RECT 29.155 89.645 29.485 90.375 ;
        RECT 29.695 90.275 31.855 90.445 ;
        RECT 29.695 89.815 30.025 90.275 ;
        RECT 30.205 89.645 30.375 90.105 ;
        RECT 30.555 89.815 30.885 90.275 ;
        RECT 31.115 89.645 31.285 90.105 ;
        RECT 31.525 89.985 31.855 90.275 ;
        RECT 32.025 90.155 32.235 91.345 ;
        RECT 32.405 91.130 32.715 92.195 ;
        RECT 32.895 91.105 35.485 92.195 ;
        RECT 32.405 90.325 32.720 90.960 ;
        RECT 32.895 90.415 34.105 90.935 ;
        RECT 34.275 90.585 35.485 91.105 ;
        RECT 35.655 91.030 35.945 92.195 ;
        RECT 36.115 91.395 36.555 92.025 ;
        RECT 32.405 89.985 32.715 90.155 ;
        RECT 31.525 89.815 32.715 89.985 ;
        RECT 32.895 89.645 35.485 90.415 ;
        RECT 36.115 90.385 36.425 91.395 ;
        RECT 36.730 91.345 37.045 92.195 ;
        RECT 37.215 91.855 38.645 92.025 ;
        RECT 37.215 91.175 37.385 91.855 ;
        RECT 36.595 91.005 37.385 91.175 ;
        RECT 36.595 90.555 36.765 91.005 ;
        RECT 37.555 90.885 37.755 91.685 ;
        RECT 36.935 90.555 37.325 90.835 ;
        RECT 37.510 90.555 37.755 90.885 ;
        RECT 37.955 90.555 38.205 91.685 ;
        RECT 38.395 91.225 38.645 91.855 ;
        RECT 38.825 91.395 39.155 92.195 ;
        RECT 38.395 91.055 39.165 91.225 ;
        RECT 40.260 91.055 40.580 92.195 ;
        RECT 38.420 90.555 38.825 90.885 ;
        RECT 38.995 90.385 39.165 91.055 ;
        RECT 40.760 90.885 40.955 91.935 ;
        RECT 41.135 91.345 41.465 92.025 ;
        RECT 41.665 91.395 41.920 92.195 ;
        RECT 41.135 91.065 41.485 91.345 ;
        RECT 40.320 90.835 40.580 90.885 ;
        RECT 40.315 90.665 40.580 90.835 ;
        RECT 40.320 90.555 40.580 90.665 ;
        RECT 40.760 90.555 41.145 90.885 ;
        RECT 41.315 90.685 41.485 91.065 ;
        RECT 41.675 90.855 41.920 91.215 ;
        RECT 42.095 91.055 42.355 92.195 ;
        RECT 42.525 91.045 42.855 92.025 ;
        RECT 43.025 91.055 43.305 92.195 ;
        RECT 43.475 91.105 46.065 92.195 ;
        RECT 41.315 90.515 41.835 90.685 ;
        RECT 42.115 90.635 42.450 90.885 ;
        RECT 35.655 89.645 35.945 90.370 ;
        RECT 36.115 89.825 36.555 90.385 ;
        RECT 36.725 89.645 37.175 90.385 ;
        RECT 37.345 90.215 38.505 90.385 ;
        RECT 37.345 89.815 37.515 90.215 ;
        RECT 37.685 89.645 38.105 90.045 ;
        RECT 38.275 89.815 38.505 90.215 ;
        RECT 38.675 89.815 39.165 90.385 ;
        RECT 40.260 90.175 41.475 90.345 ;
        RECT 40.260 89.825 40.550 90.175 ;
        RECT 40.745 89.645 41.075 90.005 ;
        RECT 41.245 89.870 41.475 90.175 ;
        RECT 41.665 89.950 41.835 90.515 ;
        RECT 42.620 90.445 42.790 91.045 ;
        RECT 42.960 90.615 43.295 90.885 ;
        RECT 42.095 89.815 42.790 90.445 ;
        RECT 42.995 89.645 43.305 90.445 ;
        RECT 43.475 90.415 44.685 90.935 ;
        RECT 44.855 90.585 46.065 91.105 ;
        RECT 46.325 91.265 46.495 92.025 ;
        RECT 46.675 91.435 47.005 92.195 ;
        RECT 46.325 91.095 46.990 91.265 ;
        RECT 47.175 91.120 47.445 92.025 ;
        RECT 46.820 90.950 46.990 91.095 ;
        RECT 46.255 90.545 46.585 90.915 ;
        RECT 46.820 90.620 47.105 90.950 ;
        RECT 43.475 89.645 46.065 90.415 ;
        RECT 46.820 90.365 46.990 90.620 ;
        RECT 46.325 90.195 46.990 90.365 ;
        RECT 47.275 90.320 47.445 91.120 ;
        RECT 47.615 91.105 51.125 92.195 ;
        RECT 51.295 91.105 52.505 92.195 ;
        RECT 52.695 91.685 52.995 92.195 ;
        RECT 53.165 91.685 53.545 91.855 ;
        RECT 54.125 91.685 54.755 92.195 ;
        RECT 53.165 91.515 53.335 91.685 ;
        RECT 54.925 91.515 55.255 92.025 ;
        RECT 55.425 91.685 55.725 92.195 ;
        RECT 55.895 91.760 61.240 92.195 ;
        RECT 46.325 89.815 46.495 90.195 ;
        RECT 46.675 89.645 47.005 90.025 ;
        RECT 47.185 89.815 47.445 90.320 ;
        RECT 47.615 90.415 49.265 90.935 ;
        RECT 49.435 90.585 51.125 91.105 ;
        RECT 47.615 89.645 51.125 90.415 ;
        RECT 51.295 90.395 51.815 90.935 ;
        RECT 51.985 90.565 52.505 91.105 ;
        RECT 52.675 91.315 53.335 91.515 ;
        RECT 53.505 91.345 55.725 91.515 ;
        RECT 51.295 89.645 52.505 90.395 ;
        RECT 52.675 90.385 52.845 91.315 ;
        RECT 53.505 91.145 53.675 91.345 ;
        RECT 53.015 90.975 53.675 91.145 ;
        RECT 53.845 91.005 55.385 91.175 ;
        RECT 53.015 90.555 53.185 90.975 ;
        RECT 53.845 90.805 54.015 91.005 ;
        RECT 53.415 90.635 54.015 90.805 ;
        RECT 54.185 90.635 54.880 90.835 ;
        RECT 55.140 90.555 55.385 91.005 ;
        RECT 53.505 90.385 54.415 90.465 ;
        RECT 52.675 89.905 52.995 90.385 ;
        RECT 53.165 90.295 54.415 90.385 ;
        RECT 53.165 90.215 53.675 90.295 ;
        RECT 53.165 89.815 53.395 90.215 ;
        RECT 53.565 89.645 53.915 90.035 ;
        RECT 54.085 89.815 54.415 90.295 ;
        RECT 54.585 89.645 54.755 90.465 ;
        RECT 55.555 90.385 55.725 91.345 ;
        RECT 55.260 89.840 55.725 90.385 ;
        RECT 57.480 90.190 57.820 91.020 ;
        RECT 59.300 90.510 59.650 91.760 ;
        RECT 61.415 91.030 61.705 92.195 ;
        RECT 62.335 91.475 62.795 92.025 ;
        RECT 62.985 91.475 63.315 92.195 ;
        RECT 55.895 89.645 61.240 90.190 ;
        RECT 61.415 89.645 61.705 90.370 ;
        RECT 62.335 90.105 62.585 91.475 ;
        RECT 63.515 91.305 63.815 91.855 ;
        RECT 63.985 91.525 64.265 92.195 ;
        RECT 62.875 91.135 63.815 91.305 ;
        RECT 62.875 90.885 63.045 91.135 ;
        RECT 64.185 90.885 64.450 91.245 ;
        RECT 64.635 91.105 68.145 92.195 ;
        RECT 62.755 90.555 63.045 90.885 ;
        RECT 63.215 90.635 63.555 90.885 ;
        RECT 63.775 90.635 64.450 90.885 ;
        RECT 62.875 90.465 63.045 90.555 ;
        RECT 62.875 90.275 64.265 90.465 ;
        RECT 62.335 89.815 62.895 90.105 ;
        RECT 63.065 89.645 63.315 90.105 ;
        RECT 63.935 89.915 64.265 90.275 ;
        RECT 64.635 90.415 66.285 90.935 ;
        RECT 66.455 90.585 68.145 91.105 ;
        RECT 69.235 91.055 69.575 92.025 ;
        RECT 69.745 91.055 69.915 92.195 ;
        RECT 70.185 91.395 70.435 92.195 ;
        RECT 71.080 91.225 71.410 92.025 ;
        RECT 71.710 91.395 72.040 92.195 ;
        RECT 72.210 91.225 72.540 92.025 ;
        RECT 70.105 91.055 72.540 91.225 ;
        RECT 72.915 91.105 74.585 92.195 ;
        RECT 75.275 91.135 75.605 91.980 ;
        RECT 75.775 91.185 75.945 92.195 ;
        RECT 76.115 91.465 76.455 92.025 ;
        RECT 76.685 91.695 77.000 92.195 ;
        RECT 77.180 91.725 78.065 91.895 ;
        RECT 69.235 90.495 69.410 91.055 ;
        RECT 70.105 90.805 70.275 91.055 ;
        RECT 69.580 90.635 70.275 90.805 ;
        RECT 70.450 90.635 70.870 90.835 ;
        RECT 71.040 90.635 71.370 90.835 ;
        RECT 71.540 90.635 71.870 90.835 ;
        RECT 69.235 90.445 69.465 90.495 ;
        RECT 64.635 89.645 68.145 90.415 ;
        RECT 69.235 89.815 69.575 90.445 ;
        RECT 69.745 89.645 69.995 90.445 ;
        RECT 70.185 90.295 71.410 90.465 ;
        RECT 70.185 89.815 70.515 90.295 ;
        RECT 70.685 89.645 70.910 90.105 ;
        RECT 71.080 89.815 71.410 90.295 ;
        RECT 72.040 90.425 72.210 91.055 ;
        RECT 72.395 90.635 72.745 90.885 ;
        RECT 72.040 89.815 72.540 90.425 ;
        RECT 72.915 90.415 73.665 90.935 ;
        RECT 73.835 90.585 74.585 91.105 ;
        RECT 75.215 91.055 75.605 91.135 ;
        RECT 76.115 91.090 77.010 91.465 ;
        RECT 75.215 91.005 75.430 91.055 ;
        RECT 75.215 90.425 75.385 91.005 ;
        RECT 76.115 90.885 76.305 91.090 ;
        RECT 77.180 90.885 77.350 91.725 ;
        RECT 78.290 91.695 78.540 92.025 ;
        RECT 75.555 90.555 76.305 90.885 ;
        RECT 76.475 90.555 77.350 90.885 ;
        RECT 72.915 89.645 74.585 90.415 ;
        RECT 75.215 90.385 75.440 90.425 ;
        RECT 76.105 90.385 76.305 90.555 ;
        RECT 75.215 90.300 75.595 90.385 ;
        RECT 75.265 89.865 75.595 90.300 ;
        RECT 75.765 89.645 75.935 90.255 ;
        RECT 76.105 89.860 76.435 90.385 ;
        RECT 76.695 89.645 76.905 90.175 ;
        RECT 77.180 90.095 77.350 90.555 ;
        RECT 77.520 90.595 77.840 91.555 ;
        RECT 78.010 90.805 78.200 91.525 ;
        RECT 78.370 90.625 78.540 91.695 ;
        RECT 78.710 91.395 78.880 92.195 ;
        RECT 79.050 91.750 80.155 91.920 ;
        RECT 79.050 91.135 79.220 91.750 ;
        RECT 80.365 91.600 80.615 92.025 ;
        RECT 80.785 91.735 81.050 92.195 ;
        RECT 79.390 91.215 79.920 91.580 ;
        RECT 80.365 91.470 80.670 91.600 ;
        RECT 78.710 91.045 79.220 91.135 ;
        RECT 78.710 90.875 79.580 91.045 ;
        RECT 78.710 90.805 78.880 90.875 ;
        RECT 79.000 90.625 79.200 90.655 ;
        RECT 77.520 90.265 77.985 90.595 ;
        RECT 78.370 90.325 79.200 90.625 ;
        RECT 78.370 90.095 78.540 90.325 ;
        RECT 77.180 89.925 77.965 90.095 ;
        RECT 78.135 89.925 78.540 90.095 ;
        RECT 78.720 89.645 79.090 90.145 ;
        RECT 79.410 90.095 79.580 90.875 ;
        RECT 79.750 90.515 79.920 91.215 ;
        RECT 80.090 90.685 80.330 91.280 ;
        RECT 79.750 90.295 80.275 90.515 ;
        RECT 80.500 90.365 80.670 91.470 ;
        RECT 80.445 90.235 80.670 90.365 ;
        RECT 80.840 90.275 81.120 91.225 ;
        RECT 80.445 90.095 80.615 90.235 ;
        RECT 79.410 89.925 80.085 90.095 ;
        RECT 80.280 89.925 80.615 90.095 ;
        RECT 80.785 89.645 81.035 90.105 ;
        RECT 81.290 89.905 81.475 92.025 ;
        RECT 81.645 91.695 81.975 92.195 ;
        RECT 82.145 91.525 82.315 92.025 ;
        RECT 81.650 91.355 82.315 91.525 ;
        RECT 81.650 90.365 81.880 91.355 ;
        RECT 82.050 90.535 82.400 91.185 ;
        RECT 82.575 90.590 82.855 92.025 ;
        RECT 83.025 91.420 83.735 92.195 ;
        RECT 83.905 91.250 84.235 92.025 ;
        RECT 83.085 91.035 84.235 91.250 ;
        RECT 81.650 90.195 82.315 90.365 ;
        RECT 81.645 89.645 81.975 90.025 ;
        RECT 82.145 89.905 82.315 90.195 ;
        RECT 82.575 89.815 82.915 90.590 ;
        RECT 83.085 90.465 83.370 91.035 ;
        RECT 83.555 90.635 84.025 90.865 ;
        RECT 84.430 90.835 84.645 91.950 ;
        RECT 84.825 91.475 85.155 92.195 ;
        RECT 84.935 90.835 85.165 91.175 ;
        RECT 85.335 91.105 87.005 92.195 ;
        RECT 84.195 90.655 84.645 90.835 ;
        RECT 84.195 90.635 84.525 90.655 ;
        RECT 84.835 90.635 85.165 90.835 ;
        RECT 83.085 90.275 83.795 90.465 ;
        RECT 83.495 90.135 83.795 90.275 ;
        RECT 83.985 90.275 85.165 90.465 ;
        RECT 83.985 90.195 84.315 90.275 ;
        RECT 83.495 90.125 83.810 90.135 ;
        RECT 83.495 90.115 83.820 90.125 ;
        RECT 83.495 90.110 83.830 90.115 ;
        RECT 83.085 89.645 83.255 90.105 ;
        RECT 83.495 90.100 83.835 90.110 ;
        RECT 83.495 90.095 83.840 90.100 ;
        RECT 83.495 90.085 83.845 90.095 ;
        RECT 83.495 90.080 83.850 90.085 ;
        RECT 83.495 89.815 83.855 90.080 ;
        RECT 84.485 89.645 84.655 90.105 ;
        RECT 84.825 89.815 85.165 90.275 ;
        RECT 85.335 90.415 86.085 90.935 ;
        RECT 86.255 90.585 87.005 91.105 ;
        RECT 87.175 91.030 87.465 92.195 ;
        RECT 87.635 91.760 92.980 92.195 ;
        RECT 93.155 91.760 98.500 92.195 ;
        RECT 85.335 89.645 87.005 90.415 ;
        RECT 87.175 89.645 87.465 90.370 ;
        RECT 89.220 90.190 89.560 91.020 ;
        RECT 91.040 90.510 91.390 91.760 ;
        RECT 94.740 90.190 95.080 91.020 ;
        RECT 96.560 90.510 96.910 91.760 ;
        RECT 99.795 91.525 100.075 92.195 ;
        RECT 100.245 91.305 100.545 91.855 ;
        RECT 100.745 91.475 101.075 92.195 ;
        RECT 101.265 91.475 101.725 92.025 ;
        RECT 99.610 90.885 99.875 91.245 ;
        RECT 100.245 91.135 101.185 91.305 ;
        RECT 101.015 90.885 101.185 91.135 ;
        RECT 99.610 90.635 100.285 90.885 ;
        RECT 100.505 90.635 100.845 90.885 ;
        RECT 101.015 90.555 101.305 90.885 ;
        RECT 101.015 90.465 101.185 90.555 ;
        RECT 99.795 90.275 101.185 90.465 ;
        RECT 87.635 89.645 92.980 90.190 ;
        RECT 93.155 89.645 98.500 90.190 ;
        RECT 99.795 89.915 100.125 90.275 ;
        RECT 101.475 90.105 101.725 91.475 ;
        RECT 101.895 91.105 105.405 92.195 ;
        RECT 106.235 91.525 106.515 92.195 ;
        RECT 106.685 91.305 106.985 91.855 ;
        RECT 107.185 91.475 107.515 92.195 ;
        RECT 107.705 91.475 108.165 92.025 ;
        RECT 100.745 89.645 100.995 90.105 ;
        RECT 101.165 89.815 101.725 90.105 ;
        RECT 101.895 90.415 103.545 90.935 ;
        RECT 103.715 90.585 105.405 91.105 ;
        RECT 106.050 90.885 106.315 91.245 ;
        RECT 106.685 91.135 107.625 91.305 ;
        RECT 107.455 90.885 107.625 91.135 ;
        RECT 106.050 90.635 106.725 90.885 ;
        RECT 106.945 90.635 107.285 90.885 ;
        RECT 107.455 90.555 107.745 90.885 ;
        RECT 107.455 90.465 107.625 90.555 ;
        RECT 101.895 89.645 105.405 90.415 ;
        RECT 106.235 90.275 107.625 90.465 ;
        RECT 106.235 89.915 106.565 90.275 ;
        RECT 107.915 90.105 108.165 91.475 ;
        RECT 108.335 91.105 111.845 92.195 ;
        RECT 107.185 89.645 107.435 90.105 ;
        RECT 107.605 89.815 108.165 90.105 ;
        RECT 108.335 90.415 109.985 90.935 ;
        RECT 110.155 90.585 111.845 91.105 ;
        RECT 112.935 91.030 113.225 92.195 ;
        RECT 113.395 91.105 114.605 92.195 ;
        RECT 114.905 91.395 115.135 92.195 ;
        RECT 115.315 91.215 115.585 92.025 ;
        RECT 115.765 91.395 115.995 92.195 ;
        RECT 116.175 91.215 116.445 92.025 ;
        RECT 116.625 91.395 116.855 92.195 ;
        RECT 117.075 91.845 119.145 92.015 ;
        RECT 117.075 91.815 118.215 91.845 ;
        RECT 117.075 91.395 117.355 91.815 ;
        RECT 117.525 91.215 117.855 91.635 ;
        RECT 118.025 91.345 118.215 91.815 ;
        RECT 118.385 91.345 118.715 91.665 ;
        RECT 118.885 91.345 119.145 91.845 ;
        RECT 119.375 91.760 124.720 92.195 ;
        RECT 108.335 89.645 111.845 90.415 ;
        RECT 113.395 90.395 113.915 90.935 ;
        RECT 114.085 90.565 114.605 91.105 ;
        RECT 114.790 90.845 115.115 91.215 ;
        RECT 115.315 91.015 117.855 91.215 ;
        RECT 118.035 90.845 118.255 91.175 ;
        RECT 114.790 90.595 115.550 90.845 ;
        RECT 116.210 90.595 116.920 90.845 ;
        RECT 117.505 90.595 118.255 90.845 ;
        RECT 118.435 90.415 118.715 91.345 ;
        RECT 118.885 90.555 119.190 91.175 ;
        RECT 112.935 89.645 113.225 90.370 ;
        RECT 113.395 89.645 114.605 90.395 ;
        RECT 114.855 90.195 115.965 90.415 ;
        RECT 116.145 90.215 118.715 90.415 ;
        RECT 114.855 89.825 115.105 90.195 ;
        RECT 115.795 90.035 115.965 90.195 ;
        RECT 115.285 89.645 115.615 90.015 ;
        RECT 115.795 89.825 116.905 90.035 ;
        RECT 117.095 89.645 117.425 90.035 ;
        RECT 117.595 89.845 117.785 90.215 ;
        RECT 117.955 89.645 118.285 90.035 ;
        RECT 118.455 89.815 118.715 90.215 ;
        RECT 118.895 89.645 119.145 90.375 ;
        RECT 120.960 90.190 121.300 91.020 ;
        RECT 122.780 90.510 123.130 91.760 ;
        RECT 124.895 91.105 127.485 92.195 ;
        RECT 124.895 90.415 126.105 90.935 ;
        RECT 126.275 90.585 127.485 91.105 ;
        RECT 128.115 90.475 128.635 92.025 ;
        RECT 128.805 91.470 129.135 92.195 ;
        RECT 119.375 89.645 124.720 90.190 ;
        RECT 124.895 89.645 127.485 90.415 ;
        RECT 128.295 89.645 128.635 90.305 ;
        RECT 128.805 89.815 129.325 91.300 ;
        RECT 129.495 91.105 131.165 92.195 ;
        RECT 131.425 91.525 131.595 92.025 ;
        RECT 131.765 91.695 132.095 92.195 ;
        RECT 131.425 91.355 132.090 91.525 ;
        RECT 129.495 90.415 130.245 90.935 ;
        RECT 130.415 90.585 131.165 91.105 ;
        RECT 131.340 90.535 131.690 91.185 ;
        RECT 129.495 89.645 131.165 90.415 ;
        RECT 131.860 90.365 132.090 91.355 ;
        RECT 131.425 90.195 132.090 90.365 ;
        RECT 131.425 89.905 131.595 90.195 ;
        RECT 131.765 89.645 132.095 90.025 ;
        RECT 132.265 89.905 132.450 92.025 ;
        RECT 132.690 91.735 132.955 92.195 ;
        RECT 133.125 91.600 133.375 92.025 ;
        RECT 133.585 91.750 134.690 91.920 ;
        RECT 133.070 91.470 133.375 91.600 ;
        RECT 132.620 90.275 132.900 91.225 ;
        RECT 133.070 90.365 133.240 91.470 ;
        RECT 133.410 90.685 133.650 91.280 ;
        RECT 133.820 91.215 134.350 91.580 ;
        RECT 133.820 90.515 133.990 91.215 ;
        RECT 134.520 91.135 134.690 91.750 ;
        RECT 134.860 91.395 135.030 92.195 ;
        RECT 135.200 91.695 135.450 92.025 ;
        RECT 135.675 91.725 136.560 91.895 ;
        RECT 134.520 91.045 135.030 91.135 ;
        RECT 133.070 90.235 133.295 90.365 ;
        RECT 133.465 90.295 133.990 90.515 ;
        RECT 134.160 90.875 135.030 91.045 ;
        RECT 132.705 89.645 132.955 90.105 ;
        RECT 133.125 90.095 133.295 90.235 ;
        RECT 134.160 90.095 134.330 90.875 ;
        RECT 134.860 90.805 135.030 90.875 ;
        RECT 134.540 90.625 134.740 90.655 ;
        RECT 135.200 90.625 135.370 91.695 ;
        RECT 135.540 90.805 135.730 91.525 ;
        RECT 134.540 90.325 135.370 90.625 ;
        RECT 135.900 90.595 136.220 91.555 ;
        RECT 133.125 89.925 133.460 90.095 ;
        RECT 133.655 89.925 134.330 90.095 ;
        RECT 134.650 89.645 135.020 90.145 ;
        RECT 135.200 90.095 135.370 90.325 ;
        RECT 135.755 90.265 136.220 90.595 ;
        RECT 136.390 90.885 136.560 91.725 ;
        RECT 136.740 91.695 137.055 92.195 ;
        RECT 137.285 91.465 137.625 92.025 ;
        RECT 136.730 91.090 137.625 91.465 ;
        RECT 137.795 91.185 137.965 92.195 ;
        RECT 137.435 90.885 137.625 91.090 ;
        RECT 138.135 91.135 138.465 91.980 ;
        RECT 138.135 91.055 138.525 91.135 ;
        RECT 138.310 91.005 138.525 91.055 ;
        RECT 138.695 91.030 138.985 92.195 ;
        RECT 139.155 91.105 142.665 92.195 ;
        RECT 142.835 91.105 144.045 92.195 ;
        RECT 144.215 91.685 144.515 92.195 ;
        RECT 144.685 91.515 145.015 92.025 ;
        RECT 145.185 91.685 145.815 92.195 ;
        RECT 146.395 91.685 146.775 91.855 ;
        RECT 146.945 91.685 147.245 92.195 ;
        RECT 146.605 91.515 146.775 91.685 ;
        RECT 136.390 90.555 137.265 90.885 ;
        RECT 137.435 90.555 138.185 90.885 ;
        RECT 136.390 90.095 136.560 90.555 ;
        RECT 137.435 90.385 137.635 90.555 ;
        RECT 138.355 90.425 138.525 91.005 ;
        RECT 138.300 90.385 138.525 90.425 ;
        RECT 135.200 89.925 135.605 90.095 ;
        RECT 135.775 89.925 136.560 90.095 ;
        RECT 136.835 89.645 137.045 90.175 ;
        RECT 137.305 89.860 137.635 90.385 ;
        RECT 138.145 90.300 138.525 90.385 ;
        RECT 139.155 90.415 140.805 90.935 ;
        RECT 140.975 90.585 142.665 91.105 ;
        RECT 137.805 89.645 137.975 90.255 ;
        RECT 138.145 89.865 138.475 90.300 ;
        RECT 138.695 89.645 138.985 90.370 ;
        RECT 139.155 89.645 142.665 90.415 ;
        RECT 142.835 90.395 143.355 90.935 ;
        RECT 143.525 90.565 144.045 91.105 ;
        RECT 144.215 91.345 146.435 91.515 ;
        RECT 142.835 89.645 144.045 90.395 ;
        RECT 144.215 90.385 144.385 91.345 ;
        RECT 144.555 91.005 146.095 91.175 ;
        RECT 144.555 90.555 144.800 91.005 ;
        RECT 145.060 90.635 145.755 90.835 ;
        RECT 145.925 90.805 146.095 91.005 ;
        RECT 146.265 91.145 146.435 91.345 ;
        RECT 146.605 91.315 147.265 91.515 ;
        RECT 146.265 90.975 146.925 91.145 ;
        RECT 145.925 90.635 146.525 90.805 ;
        RECT 146.755 90.555 146.925 90.975 ;
        RECT 144.215 89.840 144.680 90.385 ;
        RECT 145.185 89.645 145.355 90.465 ;
        RECT 145.525 90.385 146.435 90.465 ;
        RECT 147.095 90.385 147.265 91.315 ;
        RECT 147.435 91.055 147.695 92.195 ;
        RECT 147.865 91.045 148.195 92.025 ;
        RECT 148.365 91.055 148.645 92.195 ;
        RECT 148.815 91.760 154.160 92.195 ;
        RECT 147.455 90.635 147.790 90.885 ;
        RECT 147.960 90.445 148.130 91.045 ;
        RECT 148.300 90.615 148.635 90.885 ;
        RECT 145.525 90.295 146.775 90.385 ;
        RECT 145.525 89.815 145.855 90.295 ;
        RECT 146.265 90.215 146.775 90.295 ;
        RECT 146.025 89.645 146.375 90.035 ;
        RECT 146.545 89.815 146.775 90.215 ;
        RECT 146.945 89.905 147.265 90.385 ;
        RECT 147.435 89.815 148.130 90.445 ;
        RECT 148.335 89.645 148.645 90.445 ;
        RECT 150.400 90.190 150.740 91.020 ;
        RECT 152.220 90.510 152.570 91.760 ;
        RECT 154.335 91.105 155.545 92.195 ;
        RECT 154.335 90.395 154.855 90.935 ;
        RECT 155.025 90.565 155.545 91.105 ;
        RECT 155.715 91.105 156.925 92.195 ;
        RECT 155.715 90.565 156.235 91.105 ;
        RECT 156.405 90.395 156.925 90.935 ;
        RECT 148.815 89.645 154.160 90.190 ;
        RECT 154.335 89.645 155.545 90.395 ;
        RECT 155.715 89.645 156.925 90.395 ;
        RECT 22.690 89.475 157.010 89.645 ;
        RECT 22.775 88.725 23.985 89.475 ;
        RECT 24.245 88.925 24.415 89.215 ;
        RECT 24.585 89.095 24.915 89.475 ;
        RECT 24.245 88.755 24.910 88.925 ;
        RECT 22.775 88.185 23.295 88.725 ;
        RECT 23.465 88.015 23.985 88.555 ;
        RECT 22.775 86.925 23.985 88.015 ;
        RECT 24.160 87.935 24.510 88.585 ;
        RECT 24.680 87.765 24.910 88.755 ;
        RECT 24.245 87.595 24.910 87.765 ;
        RECT 24.245 87.095 24.415 87.595 ;
        RECT 24.585 86.925 24.915 87.425 ;
        RECT 25.085 87.095 25.270 89.215 ;
        RECT 25.525 89.015 25.775 89.475 ;
        RECT 25.945 89.025 26.280 89.195 ;
        RECT 26.475 89.025 27.150 89.195 ;
        RECT 25.945 88.885 26.115 89.025 ;
        RECT 25.440 87.895 25.720 88.845 ;
        RECT 25.890 88.755 26.115 88.885 ;
        RECT 25.890 87.650 26.060 88.755 ;
        RECT 26.285 88.605 26.810 88.825 ;
        RECT 26.230 87.840 26.470 88.435 ;
        RECT 26.640 87.905 26.810 88.605 ;
        RECT 26.980 88.245 27.150 89.025 ;
        RECT 27.470 88.975 27.840 89.475 ;
        RECT 28.020 89.025 28.425 89.195 ;
        RECT 28.595 89.025 29.380 89.195 ;
        RECT 28.020 88.795 28.190 89.025 ;
        RECT 27.360 88.495 28.190 88.795 ;
        RECT 28.575 88.525 29.040 88.855 ;
        RECT 27.360 88.465 27.560 88.495 ;
        RECT 27.680 88.245 27.850 88.315 ;
        RECT 26.980 88.075 27.850 88.245 ;
        RECT 27.340 87.985 27.850 88.075 ;
        RECT 25.890 87.520 26.195 87.650 ;
        RECT 26.640 87.540 27.170 87.905 ;
        RECT 25.510 86.925 25.775 87.385 ;
        RECT 25.945 87.095 26.195 87.520 ;
        RECT 27.340 87.370 27.510 87.985 ;
        RECT 26.405 87.200 27.510 87.370 ;
        RECT 27.680 86.925 27.850 87.725 ;
        RECT 28.020 87.425 28.190 88.495 ;
        RECT 28.360 87.595 28.550 88.315 ;
        RECT 28.720 87.565 29.040 88.525 ;
        RECT 29.210 88.565 29.380 89.025 ;
        RECT 29.655 88.945 29.865 89.475 ;
        RECT 30.125 88.735 30.455 89.260 ;
        RECT 30.625 88.865 30.795 89.475 ;
        RECT 30.965 88.820 31.295 89.255 ;
        RECT 30.965 88.735 31.345 88.820 ;
        RECT 30.255 88.565 30.455 88.735 ;
        RECT 31.120 88.695 31.345 88.735 ;
        RECT 29.210 88.235 30.085 88.565 ;
        RECT 30.255 88.235 31.005 88.565 ;
        RECT 28.020 87.095 28.270 87.425 ;
        RECT 29.210 87.395 29.380 88.235 ;
        RECT 30.255 88.030 30.445 88.235 ;
        RECT 31.175 88.115 31.345 88.695 ;
        RECT 31.130 88.065 31.345 88.115 ;
        RECT 29.550 87.655 30.445 88.030 ;
        RECT 30.955 87.985 31.345 88.065 ;
        RECT 31.515 88.800 31.785 89.145 ;
        RECT 31.975 89.075 32.355 89.475 ;
        RECT 32.525 88.905 32.695 89.255 ;
        RECT 32.865 88.995 33.600 89.475 ;
        RECT 31.515 88.065 31.685 88.800 ;
        RECT 31.955 88.735 32.695 88.905 ;
        RECT 33.770 88.825 34.080 89.295 ;
        RECT 31.955 88.565 32.125 88.735 ;
        RECT 33.345 88.655 34.080 88.825 ;
        RECT 34.275 88.725 35.485 89.475 ;
        RECT 35.665 88.745 35.965 89.475 ;
        RECT 33.345 88.565 33.595 88.655 ;
        RECT 31.895 88.235 32.125 88.565 ;
        RECT 32.855 88.235 33.595 88.565 ;
        RECT 33.765 88.235 34.100 88.485 ;
        RECT 31.955 88.065 32.125 88.235 ;
        RECT 28.495 87.225 29.380 87.395 ;
        RECT 29.560 86.925 29.875 87.425 ;
        RECT 30.105 87.095 30.445 87.655 ;
        RECT 30.615 86.925 30.785 87.935 ;
        RECT 30.955 87.140 31.285 87.985 ;
        RECT 31.515 87.095 31.785 88.065 ;
        RECT 31.955 87.895 33.200 88.065 ;
        RECT 31.995 86.925 32.275 87.725 ;
        RECT 32.780 87.645 33.200 87.895 ;
        RECT 33.425 87.675 33.595 88.235 ;
        RECT 34.275 88.185 34.795 88.725 ;
        RECT 36.145 88.565 36.375 89.185 ;
        RECT 36.575 88.915 36.800 89.295 ;
        RECT 36.970 89.085 37.300 89.475 ;
        RECT 36.575 88.735 36.905 88.915 ;
        RECT 32.455 87.145 33.650 87.475 ;
        RECT 33.845 86.925 34.100 88.065 ;
        RECT 34.965 88.015 35.485 88.555 ;
        RECT 35.670 88.235 35.965 88.565 ;
        RECT 36.145 88.235 36.560 88.565 ;
        RECT 36.730 88.065 36.905 88.735 ;
        RECT 37.075 88.235 37.315 88.885 ;
        RECT 37.495 88.675 37.835 89.305 ;
        RECT 38.005 88.675 38.255 89.475 ;
        RECT 38.445 88.825 38.775 89.305 ;
        RECT 38.945 89.015 39.170 89.475 ;
        RECT 39.340 88.825 39.670 89.305 ;
        RECT 37.495 88.115 37.670 88.675 ;
        RECT 38.445 88.655 39.670 88.825 ;
        RECT 40.300 88.695 40.800 89.305 ;
        RECT 41.225 88.820 41.555 89.255 ;
        RECT 41.725 88.865 41.895 89.475 ;
        RECT 41.175 88.735 41.555 88.820 ;
        RECT 42.065 88.735 42.395 89.260 ;
        RECT 42.655 88.945 42.865 89.475 ;
        RECT 43.140 89.025 43.925 89.195 ;
        RECT 44.095 89.025 44.500 89.195 ;
        RECT 41.175 88.695 41.400 88.735 ;
        RECT 37.840 88.315 38.535 88.485 ;
        RECT 37.495 88.065 37.725 88.115 ;
        RECT 38.365 88.065 38.535 88.315 ;
        RECT 38.710 88.285 39.130 88.485 ;
        RECT 39.300 88.285 39.630 88.485 ;
        RECT 39.800 88.285 40.130 88.485 ;
        RECT 40.300 88.065 40.470 88.695 ;
        RECT 40.655 88.235 41.005 88.485 ;
        RECT 41.175 88.115 41.345 88.695 ;
        RECT 42.065 88.565 42.265 88.735 ;
        RECT 43.140 88.565 43.310 89.025 ;
        RECT 41.515 88.235 42.265 88.565 ;
        RECT 42.435 88.235 43.310 88.565 ;
        RECT 41.175 88.065 41.390 88.115 ;
        RECT 34.275 86.925 35.485 88.015 ;
        RECT 35.665 87.705 36.560 88.035 ;
        RECT 36.730 87.875 37.315 88.065 ;
        RECT 35.665 87.535 36.870 87.705 ;
        RECT 35.665 87.105 35.995 87.535 ;
        RECT 36.175 86.925 36.370 87.365 ;
        RECT 36.540 87.105 36.870 87.535 ;
        RECT 37.040 87.105 37.315 87.875 ;
        RECT 37.495 87.095 37.835 88.065 ;
        RECT 38.005 86.925 38.175 88.065 ;
        RECT 38.365 87.895 40.800 88.065 ;
        RECT 41.175 87.985 41.565 88.065 ;
        RECT 38.445 86.925 38.695 87.725 ;
        RECT 39.340 87.095 39.670 87.895 ;
        RECT 39.970 86.925 40.300 87.725 ;
        RECT 40.470 87.095 40.800 87.895 ;
        RECT 41.235 87.140 41.565 87.985 ;
        RECT 42.075 88.030 42.265 88.235 ;
        RECT 41.735 86.925 41.905 87.935 ;
        RECT 42.075 87.655 42.970 88.030 ;
        RECT 42.075 87.095 42.415 87.655 ;
        RECT 42.645 86.925 42.960 87.425 ;
        RECT 43.140 87.395 43.310 88.235 ;
        RECT 43.480 88.525 43.945 88.855 ;
        RECT 44.330 88.795 44.500 89.025 ;
        RECT 44.680 88.975 45.050 89.475 ;
        RECT 45.370 89.025 46.045 89.195 ;
        RECT 46.240 89.025 46.575 89.195 ;
        RECT 43.480 87.565 43.800 88.525 ;
        RECT 44.330 88.495 45.160 88.795 ;
        RECT 43.970 87.595 44.160 88.315 ;
        RECT 44.330 87.425 44.500 88.495 ;
        RECT 44.960 88.465 45.160 88.495 ;
        RECT 44.670 88.245 44.840 88.315 ;
        RECT 45.370 88.245 45.540 89.025 ;
        RECT 46.405 88.885 46.575 89.025 ;
        RECT 46.745 89.015 46.995 89.475 ;
        RECT 44.670 88.075 45.540 88.245 ;
        RECT 45.710 88.605 46.235 88.825 ;
        RECT 46.405 88.755 46.630 88.885 ;
        RECT 44.670 87.985 45.180 88.075 ;
        RECT 43.140 87.225 44.025 87.395 ;
        RECT 44.250 87.095 44.500 87.425 ;
        RECT 44.670 86.925 44.840 87.725 ;
        RECT 45.010 87.370 45.180 87.985 ;
        RECT 45.710 87.905 45.880 88.605 ;
        RECT 45.350 87.540 45.880 87.905 ;
        RECT 46.050 87.840 46.290 88.435 ;
        RECT 46.460 87.650 46.630 88.755 ;
        RECT 46.800 87.895 47.080 88.845 ;
        RECT 46.325 87.520 46.630 87.650 ;
        RECT 45.010 87.200 46.115 87.370 ;
        RECT 46.325 87.095 46.575 87.520 ;
        RECT 46.745 86.925 47.010 87.385 ;
        RECT 47.250 87.095 47.435 89.215 ;
        RECT 47.605 89.095 47.935 89.475 ;
        RECT 48.105 88.925 48.275 89.215 ;
        RECT 47.610 88.755 48.275 88.925 ;
        RECT 47.610 87.765 47.840 88.755 ;
        RECT 48.535 88.750 48.825 89.475 ;
        RECT 48.995 88.705 50.665 89.475 ;
        RECT 48.010 87.935 48.360 88.585 ;
        RECT 48.995 88.185 49.745 88.705 ;
        RECT 50.845 88.665 51.115 89.475 ;
        RECT 51.285 88.665 51.615 89.305 ;
        RECT 51.785 88.665 52.025 89.475 ;
        RECT 52.220 88.970 52.555 89.475 ;
        RECT 52.725 88.905 52.965 89.280 ;
        RECT 53.245 89.145 53.415 89.290 ;
        RECT 53.245 88.950 53.620 89.145 ;
        RECT 53.980 88.980 54.375 89.475 ;
        RECT 47.610 87.595 48.275 87.765 ;
        RECT 47.605 86.925 47.935 87.425 ;
        RECT 48.105 87.095 48.275 87.595 ;
        RECT 48.535 86.925 48.825 88.090 ;
        RECT 49.915 88.015 50.665 88.535 ;
        RECT 50.835 88.235 51.185 88.485 ;
        RECT 51.355 88.065 51.525 88.665 ;
        RECT 51.695 88.235 52.045 88.485 ;
        RECT 48.995 86.925 50.665 88.015 ;
        RECT 50.845 86.925 51.175 88.065 ;
        RECT 51.355 87.895 52.035 88.065 ;
        RECT 52.275 87.945 52.575 88.795 ;
        RECT 52.745 88.755 52.965 88.905 ;
        RECT 52.745 88.425 53.280 88.755 ;
        RECT 53.450 88.615 53.620 88.950 ;
        RECT 54.545 88.785 54.785 89.305 ;
        RECT 51.705 87.110 52.035 87.895 ;
        RECT 52.745 87.775 52.980 88.425 ;
        RECT 53.450 88.255 54.435 88.615 ;
        RECT 52.305 87.545 52.980 87.775 ;
        RECT 53.150 88.235 54.435 88.255 ;
        RECT 53.150 88.085 54.010 88.235 ;
        RECT 52.305 87.115 52.475 87.545 ;
        RECT 52.645 86.925 52.975 87.375 ;
        RECT 53.150 87.140 53.435 88.085 ;
        RECT 54.610 87.980 54.785 88.785 ;
        RECT 54.975 88.845 55.315 89.305 ;
        RECT 55.485 89.015 55.655 89.475 ;
        RECT 56.285 89.040 56.645 89.305 ;
        RECT 56.290 89.035 56.645 89.040 ;
        RECT 56.295 89.025 56.645 89.035 ;
        RECT 56.300 89.020 56.645 89.025 ;
        RECT 56.305 89.010 56.645 89.020 ;
        RECT 56.885 89.015 57.055 89.475 ;
        RECT 56.310 89.005 56.645 89.010 ;
        RECT 56.320 88.995 56.645 89.005 ;
        RECT 56.330 88.985 56.645 88.995 ;
        RECT 55.825 88.845 56.155 88.925 ;
        RECT 54.975 88.655 56.155 88.845 ;
        RECT 56.345 88.845 56.645 88.985 ;
        RECT 56.345 88.655 57.055 88.845 ;
        RECT 53.610 87.605 54.305 87.915 ;
        RECT 53.615 86.925 54.300 87.395 ;
        RECT 54.480 87.195 54.785 87.980 ;
        RECT 54.975 88.285 55.305 88.485 ;
        RECT 55.615 88.465 55.945 88.485 ;
        RECT 55.495 88.285 55.945 88.465 ;
        RECT 54.975 87.945 55.205 88.285 ;
        RECT 54.985 86.925 55.315 87.645 ;
        RECT 55.495 87.170 55.710 88.285 ;
        RECT 56.115 88.255 56.585 88.485 ;
        RECT 56.770 88.085 57.055 88.655 ;
        RECT 57.225 88.530 57.565 89.305 ;
        RECT 58.285 88.925 58.455 89.305 ;
        RECT 58.635 89.095 58.965 89.475 ;
        RECT 58.285 88.755 58.950 88.925 ;
        RECT 59.145 88.800 59.405 89.305 ;
        RECT 59.625 88.820 59.955 89.255 ;
        RECT 60.125 88.865 60.295 89.475 ;
        RECT 55.905 87.870 57.055 88.085 ;
        RECT 55.905 87.095 56.235 87.870 ;
        RECT 56.405 86.925 57.115 87.700 ;
        RECT 57.285 87.095 57.565 88.530 ;
        RECT 58.215 88.205 58.545 88.575 ;
        RECT 58.780 88.500 58.950 88.755 ;
        RECT 58.780 88.170 59.065 88.500 ;
        RECT 58.780 88.025 58.950 88.170 ;
        RECT 58.285 87.855 58.950 88.025 ;
        RECT 59.235 88.000 59.405 88.800 ;
        RECT 58.285 87.095 58.455 87.855 ;
        RECT 58.635 86.925 58.965 87.685 ;
        RECT 59.135 87.095 59.405 88.000 ;
        RECT 59.575 88.735 59.955 88.820 ;
        RECT 60.465 88.735 60.795 89.260 ;
        RECT 61.055 88.945 61.265 89.475 ;
        RECT 61.540 89.025 62.325 89.195 ;
        RECT 62.495 89.025 62.900 89.195 ;
        RECT 59.575 88.695 59.800 88.735 ;
        RECT 59.575 88.115 59.745 88.695 ;
        RECT 60.465 88.565 60.665 88.735 ;
        RECT 61.540 88.565 61.710 89.025 ;
        RECT 59.915 88.235 60.665 88.565 ;
        RECT 60.835 88.235 61.710 88.565 ;
        RECT 59.575 88.065 59.790 88.115 ;
        RECT 59.575 87.985 59.965 88.065 ;
        RECT 59.635 87.140 59.965 87.985 ;
        RECT 60.475 88.030 60.665 88.235 ;
        RECT 60.135 86.925 60.305 87.935 ;
        RECT 60.475 87.655 61.370 88.030 ;
        RECT 60.475 87.095 60.815 87.655 ;
        RECT 61.045 86.925 61.360 87.425 ;
        RECT 61.540 87.395 61.710 88.235 ;
        RECT 61.880 88.525 62.345 88.855 ;
        RECT 62.730 88.795 62.900 89.025 ;
        RECT 63.080 88.975 63.450 89.475 ;
        RECT 63.770 89.025 64.445 89.195 ;
        RECT 64.640 89.025 64.975 89.195 ;
        RECT 61.880 87.565 62.200 88.525 ;
        RECT 62.730 88.495 63.560 88.795 ;
        RECT 62.370 87.595 62.560 88.315 ;
        RECT 62.730 87.425 62.900 88.495 ;
        RECT 63.360 88.465 63.560 88.495 ;
        RECT 63.070 88.245 63.240 88.315 ;
        RECT 63.770 88.245 63.940 89.025 ;
        RECT 64.805 88.885 64.975 89.025 ;
        RECT 65.145 89.015 65.395 89.475 ;
        RECT 63.070 88.075 63.940 88.245 ;
        RECT 64.110 88.605 64.635 88.825 ;
        RECT 64.805 88.755 65.030 88.885 ;
        RECT 63.070 87.985 63.580 88.075 ;
        RECT 61.540 87.225 62.425 87.395 ;
        RECT 62.650 87.095 62.900 87.425 ;
        RECT 63.070 86.925 63.240 87.725 ;
        RECT 63.410 87.370 63.580 87.985 ;
        RECT 64.110 87.905 64.280 88.605 ;
        RECT 63.750 87.540 64.280 87.905 ;
        RECT 64.450 87.840 64.690 88.435 ;
        RECT 64.860 87.650 65.030 88.755 ;
        RECT 65.200 87.895 65.480 88.845 ;
        RECT 64.725 87.520 65.030 87.650 ;
        RECT 63.410 87.200 64.515 87.370 ;
        RECT 64.725 87.095 64.975 87.520 ;
        RECT 65.145 86.925 65.410 87.385 ;
        RECT 65.650 87.095 65.835 89.215 ;
        RECT 66.005 89.095 66.335 89.475 ;
        RECT 66.505 88.925 66.675 89.215 ;
        RECT 66.010 88.755 66.675 88.925 ;
        RECT 66.010 87.765 66.240 88.755 ;
        RECT 66.935 88.705 69.525 89.475 ;
        RECT 69.715 88.745 70.005 89.475 ;
        RECT 66.410 87.935 66.760 88.585 ;
        RECT 66.935 88.185 68.145 88.705 ;
        RECT 68.315 88.015 69.525 88.535 ;
        RECT 69.705 88.235 70.005 88.565 ;
        RECT 70.185 88.545 70.415 89.185 ;
        RECT 70.595 88.925 70.905 89.295 ;
        RECT 71.085 89.105 71.755 89.475 ;
        RECT 70.595 88.725 71.825 88.925 ;
        RECT 70.185 88.235 70.710 88.545 ;
        RECT 70.890 88.235 71.355 88.545 ;
        RECT 71.535 88.055 71.825 88.725 ;
        RECT 66.010 87.595 66.675 87.765 ;
        RECT 66.005 86.925 66.335 87.425 ;
        RECT 66.505 87.095 66.675 87.595 ;
        RECT 66.935 86.925 69.525 88.015 ;
        RECT 69.715 87.815 70.875 88.055 ;
        RECT 69.715 87.105 69.975 87.815 ;
        RECT 70.145 86.925 70.475 87.635 ;
        RECT 70.645 87.105 70.875 87.815 ;
        RECT 71.055 87.835 71.825 88.055 ;
        RECT 71.055 87.105 71.325 87.835 ;
        RECT 71.505 86.925 71.845 87.655 ;
        RECT 72.015 87.105 72.275 89.295 ;
        RECT 72.455 88.705 74.125 89.475 ;
        RECT 74.295 88.750 74.585 89.475 ;
        RECT 74.755 88.705 76.425 89.475 ;
        RECT 72.455 88.185 73.205 88.705 ;
        RECT 73.375 88.015 74.125 88.535 ;
        RECT 74.755 88.185 75.505 88.705 ;
        RECT 76.595 88.675 77.290 89.305 ;
        RECT 77.495 88.675 77.805 89.475 ;
        RECT 72.455 86.925 74.125 88.015 ;
        RECT 74.295 86.925 74.585 88.090 ;
        RECT 75.675 88.015 76.425 88.535 ;
        RECT 76.615 88.235 76.950 88.485 ;
        RECT 77.120 88.115 77.290 88.675 ;
        RECT 78.065 88.605 78.235 89.170 ;
        RECT 78.425 88.945 78.655 89.250 ;
        RECT 78.825 89.115 79.155 89.475 ;
        RECT 79.350 88.945 79.640 89.295 ;
        RECT 78.425 88.775 79.640 88.945 ;
        RECT 79.840 88.825 80.150 89.295 ;
        RECT 80.320 88.995 81.055 89.475 ;
        RECT 81.225 88.905 81.395 89.255 ;
        RECT 81.565 89.075 81.945 89.475 ;
        RECT 79.840 88.655 80.575 88.825 ;
        RECT 81.225 88.735 81.965 88.905 ;
        RECT 82.135 88.800 82.405 89.145 ;
        RECT 77.460 88.235 77.795 88.505 ;
        RECT 78.065 88.435 78.585 88.605 ;
        RECT 80.325 88.565 80.575 88.655 ;
        RECT 81.795 88.565 81.965 88.735 ;
        RECT 77.115 88.075 77.290 88.115 ;
        RECT 74.755 86.925 76.425 88.015 ;
        RECT 76.595 86.925 76.855 88.065 ;
        RECT 77.025 87.095 77.355 88.075 ;
        RECT 77.525 86.925 77.805 88.065 ;
        RECT 77.980 87.905 78.225 88.265 ;
        RECT 78.415 88.055 78.585 88.435 ;
        RECT 78.755 88.235 79.140 88.565 ;
        RECT 79.320 88.455 79.580 88.565 ;
        RECT 79.320 88.285 79.585 88.455 ;
        RECT 79.320 88.235 79.580 88.285 ;
        RECT 79.820 88.235 80.155 88.485 ;
        RECT 80.325 88.235 81.065 88.565 ;
        RECT 81.795 88.235 82.025 88.565 ;
        RECT 78.415 87.775 78.765 88.055 ;
        RECT 77.980 86.925 78.235 87.725 ;
        RECT 78.435 87.095 78.765 87.775 ;
        RECT 78.945 87.185 79.140 88.235 ;
        RECT 79.320 86.925 79.640 88.065 ;
        RECT 79.820 86.925 80.075 88.065 ;
        RECT 80.325 87.675 80.495 88.235 ;
        RECT 81.795 88.065 81.965 88.235 ;
        RECT 82.235 88.065 82.405 88.800 ;
        RECT 83.045 88.745 83.345 89.475 ;
        RECT 83.525 88.565 83.755 89.185 ;
        RECT 83.955 88.915 84.180 89.295 ;
        RECT 84.350 89.085 84.680 89.475 ;
        RECT 84.965 88.925 85.135 89.215 ;
        RECT 85.305 89.095 85.635 89.475 ;
        RECT 83.955 88.735 84.285 88.915 ;
        RECT 83.050 88.235 83.345 88.565 ;
        RECT 83.525 88.235 83.940 88.565 ;
        RECT 80.720 87.895 81.965 88.065 ;
        RECT 80.720 87.645 81.140 87.895 ;
        RECT 80.270 87.145 81.465 87.475 ;
        RECT 81.645 86.925 81.925 87.725 ;
        RECT 82.135 87.095 82.405 88.065 ;
        RECT 84.110 88.065 84.285 88.735 ;
        RECT 84.455 88.235 84.695 88.885 ;
        RECT 84.965 88.755 85.630 88.925 ;
        RECT 83.045 87.705 83.940 88.035 ;
        RECT 84.110 87.875 84.695 88.065 ;
        RECT 84.880 87.935 85.230 88.585 ;
        RECT 83.045 87.535 84.250 87.705 ;
        RECT 83.045 87.105 83.375 87.535 ;
        RECT 83.555 86.925 83.750 87.365 ;
        RECT 83.920 87.105 84.250 87.535 ;
        RECT 84.420 87.105 84.695 87.875 ;
        RECT 85.400 87.765 85.630 88.755 ;
        RECT 84.965 87.595 85.630 87.765 ;
        RECT 84.965 87.095 85.135 87.595 ;
        RECT 85.305 86.925 85.635 87.425 ;
        RECT 85.805 87.095 85.990 89.215 ;
        RECT 86.245 89.015 86.495 89.475 ;
        RECT 86.665 89.025 87.000 89.195 ;
        RECT 87.195 89.025 87.870 89.195 ;
        RECT 86.665 88.885 86.835 89.025 ;
        RECT 86.160 87.895 86.440 88.845 ;
        RECT 86.610 88.755 86.835 88.885 ;
        RECT 86.610 87.650 86.780 88.755 ;
        RECT 87.005 88.605 87.530 88.825 ;
        RECT 86.950 87.840 87.190 88.435 ;
        RECT 87.360 87.905 87.530 88.605 ;
        RECT 87.700 88.245 87.870 89.025 ;
        RECT 88.190 88.975 88.560 89.475 ;
        RECT 88.740 89.025 89.145 89.195 ;
        RECT 89.315 89.025 90.100 89.195 ;
        RECT 88.740 88.795 88.910 89.025 ;
        RECT 88.080 88.495 88.910 88.795 ;
        RECT 89.295 88.525 89.760 88.855 ;
        RECT 88.080 88.465 88.280 88.495 ;
        RECT 88.400 88.245 88.570 88.315 ;
        RECT 87.700 88.075 88.570 88.245 ;
        RECT 88.060 87.985 88.570 88.075 ;
        RECT 86.610 87.520 86.915 87.650 ;
        RECT 87.360 87.540 87.890 87.905 ;
        RECT 86.230 86.925 86.495 87.385 ;
        RECT 86.665 87.095 86.915 87.520 ;
        RECT 88.060 87.370 88.230 87.985 ;
        RECT 87.125 87.200 88.230 87.370 ;
        RECT 88.400 86.925 88.570 87.725 ;
        RECT 88.740 87.425 88.910 88.495 ;
        RECT 89.080 87.595 89.270 88.315 ;
        RECT 89.440 87.565 89.760 88.525 ;
        RECT 89.930 88.565 90.100 89.025 ;
        RECT 90.375 88.945 90.585 89.475 ;
        RECT 90.845 88.735 91.175 89.260 ;
        RECT 91.345 88.865 91.515 89.475 ;
        RECT 91.685 88.820 92.015 89.255 ;
        RECT 91.685 88.735 92.065 88.820 ;
        RECT 90.975 88.565 91.175 88.735 ;
        RECT 91.840 88.695 92.065 88.735 ;
        RECT 89.930 88.235 90.805 88.565 ;
        RECT 90.975 88.235 91.725 88.565 ;
        RECT 88.740 87.095 88.990 87.425 ;
        RECT 89.930 87.395 90.100 88.235 ;
        RECT 90.975 88.030 91.165 88.235 ;
        RECT 91.895 88.115 92.065 88.695 ;
        RECT 91.850 88.065 92.065 88.115 ;
        RECT 90.270 87.655 91.165 88.030 ;
        RECT 91.675 87.985 92.065 88.065 ;
        RECT 92.235 88.735 92.675 89.295 ;
        RECT 92.845 88.735 93.295 89.475 ;
        RECT 93.465 88.905 93.635 89.305 ;
        RECT 93.805 89.075 94.225 89.475 ;
        RECT 94.395 88.905 94.625 89.305 ;
        RECT 93.465 88.735 94.625 88.905 ;
        RECT 94.795 88.735 95.285 89.305 ;
        RECT 95.545 89.135 95.715 89.170 ;
        RECT 95.515 88.965 95.715 89.135 ;
        RECT 89.215 87.225 90.100 87.395 ;
        RECT 90.280 86.925 90.595 87.425 ;
        RECT 90.825 87.095 91.165 87.655 ;
        RECT 91.335 86.925 91.505 87.935 ;
        RECT 91.675 87.140 92.005 87.985 ;
        RECT 92.235 87.725 92.545 88.735 ;
        RECT 92.715 88.115 92.885 88.565 ;
        RECT 93.055 88.285 93.445 88.565 ;
        RECT 93.630 88.235 93.875 88.565 ;
        RECT 92.715 87.945 93.505 88.115 ;
        RECT 92.235 87.095 92.675 87.725 ;
        RECT 92.850 86.925 93.165 87.775 ;
        RECT 93.335 87.265 93.505 87.945 ;
        RECT 93.675 87.435 93.875 88.235 ;
        RECT 94.075 87.435 94.325 88.565 ;
        RECT 94.540 88.235 94.945 88.565 ;
        RECT 95.115 88.065 95.285 88.735 ;
        RECT 95.545 88.605 95.715 88.965 ;
        RECT 95.905 88.945 96.135 89.250 ;
        RECT 96.305 89.115 96.635 89.475 ;
        RECT 96.830 88.945 97.120 89.295 ;
        RECT 95.905 88.775 97.120 88.945 ;
        RECT 97.295 88.705 99.885 89.475 ;
        RECT 100.055 88.750 100.345 89.475 ;
        RECT 100.515 88.705 102.185 89.475 ;
        RECT 95.545 88.435 96.065 88.605 ;
        RECT 94.515 87.895 95.285 88.065 ;
        RECT 95.460 87.905 95.705 88.265 ;
        RECT 95.895 88.055 96.065 88.435 ;
        RECT 96.235 88.235 96.620 88.565 ;
        RECT 96.800 88.455 97.060 88.565 ;
        RECT 96.800 88.285 97.065 88.455 ;
        RECT 96.800 88.235 97.060 88.285 ;
        RECT 94.515 87.265 94.765 87.895 ;
        RECT 95.895 87.775 96.245 88.055 ;
        RECT 93.335 87.095 94.765 87.265 ;
        RECT 94.945 86.925 95.275 87.725 ;
        RECT 95.460 86.925 95.715 87.725 ;
        RECT 95.915 87.095 96.245 87.775 ;
        RECT 96.425 87.185 96.620 88.235 ;
        RECT 97.295 88.185 98.505 88.705 ;
        RECT 96.800 86.925 97.120 88.065 ;
        RECT 98.675 88.015 99.885 88.535 ;
        RECT 100.515 88.185 101.265 88.705 ;
        RECT 102.815 88.675 103.510 89.305 ;
        RECT 103.715 88.675 104.025 89.475 ;
        RECT 104.195 88.930 109.540 89.475 ;
        RECT 109.720 88.970 110.055 89.475 ;
        RECT 97.295 86.925 99.885 88.015 ;
        RECT 100.055 86.925 100.345 88.090 ;
        RECT 101.435 88.015 102.185 88.535 ;
        RECT 102.835 88.235 103.170 88.485 ;
        RECT 103.340 88.075 103.510 88.675 ;
        RECT 103.680 88.235 104.015 88.505 ;
        RECT 105.780 88.100 106.120 88.930 ;
        RECT 110.225 88.905 110.465 89.280 ;
        RECT 110.745 89.145 110.915 89.290 ;
        RECT 110.745 88.950 111.120 89.145 ;
        RECT 111.480 88.980 111.875 89.475 ;
        RECT 100.515 86.925 102.185 88.015 ;
        RECT 102.815 86.925 103.075 88.065 ;
        RECT 103.245 87.095 103.575 88.075 ;
        RECT 103.745 86.925 104.025 88.065 ;
        RECT 107.600 87.360 107.950 88.610 ;
        RECT 109.775 87.945 110.075 88.795 ;
        RECT 110.245 88.755 110.465 88.905 ;
        RECT 110.245 88.425 110.780 88.755 ;
        RECT 110.950 88.615 111.120 88.950 ;
        RECT 112.045 88.785 112.285 89.305 ;
        RECT 110.245 87.775 110.480 88.425 ;
        RECT 110.950 88.255 111.935 88.615 ;
        RECT 109.805 87.545 110.480 87.775 ;
        RECT 110.650 88.235 111.935 88.255 ;
        RECT 110.650 88.085 111.510 88.235 ;
        RECT 104.195 86.925 109.540 87.360 ;
        RECT 109.805 87.115 109.975 87.545 ;
        RECT 110.145 86.925 110.475 87.375 ;
        RECT 110.650 87.140 110.935 88.085 ;
        RECT 112.110 87.980 112.285 88.785 ;
        RECT 112.475 88.705 114.145 89.475 ;
        RECT 114.515 88.845 114.845 89.205 ;
        RECT 115.465 89.015 115.715 89.475 ;
        RECT 115.885 89.015 116.445 89.305 ;
        RECT 112.475 88.185 113.225 88.705 ;
        RECT 114.515 88.655 115.905 88.845 ;
        RECT 115.735 88.565 115.905 88.655 ;
        RECT 113.395 88.015 114.145 88.535 ;
        RECT 111.110 87.605 111.805 87.915 ;
        RECT 111.115 86.925 111.800 87.395 ;
        RECT 111.980 87.195 112.285 87.980 ;
        RECT 112.475 86.925 114.145 88.015 ;
        RECT 114.330 88.235 115.005 88.485 ;
        RECT 115.225 88.235 115.565 88.485 ;
        RECT 115.735 88.235 116.025 88.565 ;
        RECT 114.330 87.875 114.595 88.235 ;
        RECT 115.735 87.985 115.905 88.235 ;
        RECT 114.965 87.815 115.905 87.985 ;
        RECT 114.515 86.925 114.795 87.595 ;
        RECT 114.965 87.265 115.265 87.815 ;
        RECT 116.195 87.645 116.445 89.015 ;
        RECT 116.705 88.925 116.875 89.305 ;
        RECT 117.055 89.095 117.385 89.475 ;
        RECT 116.705 88.755 117.370 88.925 ;
        RECT 117.565 88.800 117.825 89.305 ;
        RECT 116.635 88.205 116.965 88.575 ;
        RECT 117.200 88.500 117.370 88.755 ;
        RECT 117.200 88.170 117.485 88.500 ;
        RECT 117.200 88.025 117.370 88.170 ;
        RECT 115.465 86.925 115.795 87.645 ;
        RECT 115.985 87.095 116.445 87.645 ;
        RECT 116.705 87.855 117.370 88.025 ;
        RECT 117.655 88.000 117.825 88.800 ;
        RECT 116.705 87.095 116.875 87.855 ;
        RECT 117.055 86.925 117.385 87.685 ;
        RECT 117.555 87.095 117.825 88.000 ;
        RECT 118.915 87.820 119.435 89.305 ;
        RECT 119.605 88.815 119.945 89.475 ;
        RECT 120.295 88.705 122.885 89.475 ;
        RECT 123.055 88.845 123.395 89.305 ;
        RECT 123.565 89.015 123.735 89.475 ;
        RECT 124.365 89.040 124.725 89.305 ;
        RECT 124.370 89.035 124.725 89.040 ;
        RECT 124.375 89.025 124.725 89.035 ;
        RECT 124.380 89.020 124.725 89.025 ;
        RECT 124.385 89.010 124.725 89.020 ;
        RECT 124.965 89.015 125.135 89.475 ;
        RECT 124.390 89.005 124.725 89.010 ;
        RECT 124.400 88.995 124.725 89.005 ;
        RECT 124.410 88.985 124.725 88.995 ;
        RECT 123.905 88.845 124.235 88.925 ;
        RECT 119.105 86.925 119.435 87.650 ;
        RECT 119.605 87.095 120.125 88.645 ;
        RECT 120.295 88.185 121.505 88.705 ;
        RECT 123.055 88.655 124.235 88.845 ;
        RECT 124.425 88.845 124.725 88.985 ;
        RECT 124.425 88.655 125.135 88.845 ;
        RECT 121.675 88.015 122.885 88.535 ;
        RECT 120.295 86.925 122.885 88.015 ;
        RECT 123.055 88.285 123.385 88.485 ;
        RECT 123.695 88.465 124.025 88.485 ;
        RECT 123.575 88.285 124.025 88.465 ;
        RECT 123.055 87.945 123.285 88.285 ;
        RECT 123.065 86.925 123.395 87.645 ;
        RECT 123.575 87.170 123.790 88.285 ;
        RECT 124.195 88.255 124.665 88.485 ;
        RECT 124.850 88.085 125.135 88.655 ;
        RECT 125.305 88.530 125.645 89.305 ;
        RECT 125.815 88.750 126.105 89.475 ;
        RECT 126.295 88.665 126.535 89.475 ;
        RECT 126.705 88.665 127.035 89.305 ;
        RECT 127.205 88.665 127.475 89.475 ;
        RECT 128.205 88.925 128.375 89.215 ;
        RECT 128.545 89.095 128.875 89.475 ;
        RECT 128.205 88.755 128.810 88.925 ;
        RECT 123.985 87.870 125.135 88.085 ;
        RECT 123.985 87.095 124.315 87.870 ;
        RECT 124.485 86.925 125.195 87.700 ;
        RECT 125.365 87.095 125.645 88.530 ;
        RECT 126.275 88.235 126.625 88.485 ;
        RECT 125.815 86.925 126.105 88.090 ;
        RECT 126.795 88.065 126.965 88.665 ;
        RECT 127.135 88.235 127.485 88.485 ;
        RECT 126.285 87.895 126.965 88.065 ;
        RECT 126.285 87.110 126.615 87.895 ;
        RECT 127.145 86.925 127.475 88.065 ;
        RECT 128.115 87.935 128.360 88.575 ;
        RECT 128.640 88.490 128.810 88.755 ;
        RECT 128.640 88.160 128.870 88.490 ;
        RECT 128.640 87.765 128.810 88.160 ;
        RECT 128.205 87.595 128.810 87.765 ;
        RECT 129.045 87.875 129.215 89.215 ;
        RECT 129.540 88.945 129.735 89.215 ;
        RECT 129.905 89.115 130.235 89.475 ;
        RECT 130.795 89.025 131.635 89.195 ;
        RECT 129.540 88.795 130.145 88.945 ;
        RECT 129.540 88.775 130.350 88.795 ;
        RECT 129.465 88.235 129.795 88.605 ;
        RECT 129.975 88.325 130.350 88.775 ;
        RECT 130.590 88.520 131.295 88.825 ;
        RECT 129.975 88.065 130.145 88.325 ;
        RECT 129.460 87.895 130.145 88.065 ;
        RECT 128.205 87.095 128.375 87.595 ;
        RECT 128.545 86.925 128.875 87.425 ;
        RECT 129.045 87.095 129.270 87.875 ;
        RECT 129.460 87.145 129.815 87.895 ;
        RECT 129.985 86.925 130.275 87.725 ;
        RECT 130.475 87.555 130.810 88.205 ;
        RECT 130.980 88.000 131.295 88.520 ;
        RECT 131.465 88.565 131.635 89.025 ;
        RECT 131.805 89.015 132.075 89.475 ;
        RECT 132.325 88.840 132.570 89.300 ;
        RECT 132.785 88.845 133.010 89.475 ;
        RECT 132.400 88.565 132.570 88.840 ;
        RECT 133.205 88.815 133.465 89.145 ;
        RECT 133.635 88.930 138.980 89.475 ;
        RECT 131.465 88.235 132.230 88.565 ;
        RECT 132.400 88.235 133.125 88.565 ;
        RECT 131.465 88.110 131.675 88.235 ;
        RECT 130.980 87.650 131.315 88.000 ;
        RECT 131.485 87.550 131.675 88.110 ;
        RECT 132.400 88.025 132.570 88.235 ;
        RECT 131.845 87.695 132.570 88.025 ;
        RECT 131.460 87.525 131.675 87.550 ;
        RECT 131.435 87.515 131.675 87.525 ;
        RECT 131.420 87.495 131.675 87.515 ;
        RECT 131.420 87.475 131.660 87.495 ;
        RECT 131.420 87.470 131.650 87.475 ;
        RECT 131.325 87.455 131.650 87.470 ;
        RECT 131.325 87.305 131.635 87.455 ;
        RECT 130.775 87.135 131.635 87.305 ;
        RECT 131.805 86.925 132.125 87.385 ;
        RECT 132.325 87.125 132.570 87.695 ;
        RECT 132.750 86.925 133.035 87.990 ;
        RECT 133.295 87.890 133.465 88.815 ;
        RECT 135.220 88.100 135.560 88.930 ;
        RECT 139.815 88.845 140.145 89.205 ;
        RECT 140.765 89.015 141.015 89.475 ;
        RECT 141.185 89.015 141.745 89.305 ;
        RECT 139.815 88.655 141.205 88.845 ;
        RECT 133.205 87.105 133.465 87.890 ;
        RECT 137.040 87.360 137.390 88.610 ;
        RECT 141.035 88.565 141.205 88.655 ;
        RECT 139.630 88.235 140.305 88.485 ;
        RECT 140.525 88.235 140.865 88.485 ;
        RECT 141.035 88.235 141.325 88.565 ;
        RECT 139.630 87.875 139.895 88.235 ;
        RECT 141.035 87.985 141.205 88.235 ;
        RECT 140.265 87.815 141.205 87.985 ;
        RECT 133.635 86.925 138.980 87.360 ;
        RECT 139.815 86.925 140.095 87.595 ;
        RECT 140.265 87.265 140.565 87.815 ;
        RECT 141.495 87.645 141.745 89.015 ;
        RECT 142.005 88.925 142.175 89.305 ;
        RECT 142.355 89.095 142.685 89.475 ;
        RECT 142.005 88.755 142.670 88.925 ;
        RECT 142.865 88.800 143.125 89.305 ;
        RECT 141.935 88.205 142.265 88.575 ;
        RECT 142.500 88.500 142.670 88.755 ;
        RECT 142.500 88.170 142.785 88.500 ;
        RECT 142.500 88.025 142.670 88.170 ;
        RECT 140.765 86.925 141.095 87.645 ;
        RECT 141.285 87.095 141.745 87.645 ;
        RECT 142.005 87.855 142.670 88.025 ;
        RECT 142.955 88.000 143.125 88.800 ;
        RECT 143.295 88.705 146.805 89.475 ;
        RECT 143.295 88.185 144.945 88.705 ;
        RECT 147.445 88.665 147.715 89.475 ;
        RECT 147.885 88.665 148.215 89.305 ;
        RECT 148.385 88.665 148.625 89.475 ;
        RECT 148.815 88.675 149.125 89.475 ;
        RECT 149.330 88.675 150.025 89.305 ;
        RECT 150.195 88.725 151.405 89.475 ;
        RECT 151.575 88.750 151.865 89.475 ;
        RECT 145.115 88.015 146.805 88.535 ;
        RECT 147.435 88.235 147.785 88.485 ;
        RECT 147.955 88.065 148.125 88.665 ;
        RECT 148.295 88.235 148.645 88.485 ;
        RECT 148.825 88.235 149.160 88.505 ;
        RECT 149.330 88.075 149.500 88.675 ;
        RECT 149.670 88.235 150.005 88.485 ;
        RECT 150.195 88.185 150.715 88.725 ;
        RECT 152.035 88.705 155.545 89.475 ;
        RECT 155.715 88.725 156.925 89.475 ;
        RECT 142.005 87.095 142.175 87.855 ;
        RECT 142.355 86.925 142.685 87.685 ;
        RECT 142.855 87.095 143.125 88.000 ;
        RECT 143.295 86.925 146.805 88.015 ;
        RECT 147.445 86.925 147.775 88.065 ;
        RECT 147.955 87.895 148.635 88.065 ;
        RECT 148.305 87.110 148.635 87.895 ;
        RECT 148.815 86.925 149.095 88.065 ;
        RECT 149.265 87.095 149.595 88.075 ;
        RECT 149.765 86.925 150.025 88.065 ;
        RECT 150.885 88.015 151.405 88.555 ;
        RECT 152.035 88.185 153.685 88.705 ;
        RECT 150.195 86.925 151.405 88.015 ;
        RECT 151.575 86.925 151.865 88.090 ;
        RECT 153.855 88.015 155.545 88.535 ;
        RECT 152.035 86.925 155.545 88.015 ;
        RECT 155.715 88.015 156.235 88.555 ;
        RECT 156.405 88.185 156.925 88.725 ;
        RECT 155.715 86.925 156.925 88.015 ;
        RECT 22.690 86.755 157.010 86.925 ;
        RECT 22.775 85.665 23.985 86.755 ;
        RECT 24.155 85.665 26.745 86.755 ;
        RECT 22.775 84.955 23.295 85.495 ;
        RECT 23.465 85.125 23.985 85.665 ;
        RECT 24.155 84.975 25.365 85.495 ;
        RECT 25.535 85.145 26.745 85.665 ;
        RECT 26.915 85.150 27.195 86.585 ;
        RECT 27.365 85.980 28.075 86.755 ;
        RECT 28.245 85.810 28.575 86.585 ;
        RECT 27.425 85.595 28.575 85.810 ;
        RECT 22.775 84.205 23.985 84.955 ;
        RECT 24.155 84.205 26.745 84.975 ;
        RECT 26.915 84.375 27.255 85.150 ;
        RECT 27.425 85.025 27.710 85.595 ;
        RECT 27.895 85.195 28.365 85.425 ;
        RECT 28.770 85.395 28.985 86.510 ;
        RECT 29.165 86.035 29.495 86.755 ;
        RECT 29.275 85.395 29.505 85.735 ;
        RECT 29.685 85.615 30.015 86.755 ;
        RECT 30.545 85.785 30.875 86.570 ;
        RECT 30.195 85.615 30.875 85.785 ;
        RECT 31.055 85.615 31.335 86.755 ;
        RECT 28.535 85.215 28.985 85.395 ;
        RECT 28.535 85.195 28.865 85.215 ;
        RECT 29.175 85.195 29.505 85.395 ;
        RECT 29.675 85.195 30.025 85.445 ;
        RECT 27.425 84.835 28.135 85.025 ;
        RECT 27.835 84.695 28.135 84.835 ;
        RECT 28.325 84.835 29.505 85.025 ;
        RECT 30.195 85.015 30.365 85.615 ;
        RECT 31.505 85.605 31.835 86.585 ;
        RECT 32.005 85.615 32.265 86.755 ;
        RECT 30.535 85.195 30.885 85.445 ;
        RECT 31.065 85.175 31.400 85.445 ;
        RECT 28.325 84.755 28.655 84.835 ;
        RECT 27.835 84.685 28.150 84.695 ;
        RECT 27.835 84.675 28.160 84.685 ;
        RECT 27.835 84.670 28.170 84.675 ;
        RECT 27.425 84.205 27.595 84.665 ;
        RECT 27.835 84.660 28.175 84.670 ;
        RECT 27.835 84.655 28.180 84.660 ;
        RECT 27.835 84.645 28.185 84.655 ;
        RECT 27.835 84.640 28.190 84.645 ;
        RECT 27.835 84.375 28.195 84.640 ;
        RECT 28.825 84.205 28.995 84.665 ;
        RECT 29.165 84.375 29.505 84.835 ;
        RECT 29.685 84.205 29.955 85.015 ;
        RECT 30.125 84.375 30.455 85.015 ;
        RECT 30.625 84.205 30.865 85.015 ;
        RECT 31.570 85.005 31.740 85.605 ;
        RECT 31.910 85.195 32.245 85.445 ;
        RECT 33.355 85.035 33.875 86.585 ;
        RECT 34.045 86.030 34.375 86.755 ;
        RECT 31.055 84.205 31.365 85.005 ;
        RECT 31.570 84.375 32.265 85.005 ;
        RECT 33.535 84.205 33.875 84.865 ;
        RECT 34.045 84.375 34.565 85.860 ;
        RECT 35.655 85.590 35.945 86.755 ;
        RECT 37.035 86.245 37.335 86.755 ;
        RECT 37.505 86.075 37.835 86.585 ;
        RECT 38.005 86.245 38.635 86.755 ;
        RECT 39.215 86.245 39.595 86.415 ;
        RECT 39.765 86.245 40.065 86.755 ;
        RECT 39.425 86.075 39.595 86.245 ;
        RECT 37.035 85.905 39.255 86.075 ;
        RECT 37.035 84.945 37.205 85.905 ;
        RECT 37.375 85.565 38.915 85.735 ;
        RECT 37.375 85.115 37.620 85.565 ;
        RECT 37.880 85.195 38.575 85.395 ;
        RECT 38.745 85.365 38.915 85.565 ;
        RECT 39.085 85.705 39.255 85.905 ;
        RECT 39.425 85.875 40.085 86.075 ;
        RECT 39.085 85.535 39.745 85.705 ;
        RECT 38.745 85.195 39.345 85.365 ;
        RECT 39.575 85.115 39.745 85.535 ;
        RECT 35.655 84.205 35.945 84.930 ;
        RECT 37.035 84.400 37.500 84.945 ;
        RECT 38.005 84.205 38.175 85.025 ;
        RECT 38.345 84.945 39.255 85.025 ;
        RECT 39.915 84.945 40.085 85.875 ;
        RECT 40.255 85.665 42.845 86.755 ;
        RECT 43.205 86.030 43.535 86.755 ;
        RECT 38.345 84.855 39.595 84.945 ;
        RECT 38.345 84.375 38.675 84.855 ;
        RECT 39.085 84.775 39.595 84.855 ;
        RECT 38.845 84.205 39.195 84.595 ;
        RECT 39.365 84.375 39.595 84.775 ;
        RECT 39.765 84.465 40.085 84.945 ;
        RECT 40.255 84.975 41.465 85.495 ;
        RECT 41.635 85.145 42.845 85.665 ;
        RECT 40.255 84.205 42.845 84.975 ;
        RECT 43.015 84.375 43.535 85.860 ;
        RECT 43.705 85.035 44.225 86.585 ;
        RECT 44.395 85.665 47.905 86.755 ;
        RECT 48.265 86.030 48.595 86.755 ;
        RECT 44.395 84.975 46.045 85.495 ;
        RECT 46.215 85.145 47.905 85.665 ;
        RECT 43.705 84.205 44.045 84.865 ;
        RECT 44.395 84.205 47.905 84.975 ;
        RECT 48.075 84.375 48.595 85.860 ;
        RECT 48.765 85.035 49.285 86.585 ;
        RECT 49.455 85.665 52.045 86.755 ;
        RECT 49.455 84.975 50.665 85.495 ;
        RECT 50.835 85.145 52.045 85.665 ;
        RECT 52.675 85.615 52.955 86.755 ;
        RECT 53.125 85.605 53.455 86.585 ;
        RECT 53.625 85.615 53.885 86.755 ;
        RECT 54.055 85.665 55.725 86.755 ;
        RECT 52.685 85.175 53.020 85.445 ;
        RECT 53.190 85.005 53.360 85.605 ;
        RECT 53.530 85.195 53.865 85.445 ;
        RECT 48.765 84.205 49.105 84.865 ;
        RECT 49.455 84.205 52.045 84.975 ;
        RECT 52.675 84.205 52.985 85.005 ;
        RECT 53.190 84.375 53.885 85.005 ;
        RECT 54.055 84.975 54.805 85.495 ;
        RECT 54.975 85.145 55.725 85.665 ;
        RECT 55.895 85.150 56.175 86.585 ;
        RECT 56.345 85.980 57.055 86.755 ;
        RECT 57.225 85.810 57.555 86.585 ;
        RECT 56.405 85.595 57.555 85.810 ;
        RECT 54.055 84.205 55.725 84.975 ;
        RECT 55.895 84.375 56.235 85.150 ;
        RECT 56.405 85.025 56.690 85.595 ;
        RECT 56.875 85.195 57.345 85.425 ;
        RECT 57.750 85.395 57.965 86.510 ;
        RECT 58.145 86.035 58.475 86.755 ;
        RECT 58.745 86.135 58.915 86.565 ;
        RECT 59.085 86.305 59.415 86.755 ;
        RECT 58.745 85.905 59.420 86.135 ;
        RECT 58.255 85.395 58.485 85.735 ;
        RECT 57.515 85.215 57.965 85.395 ;
        RECT 57.515 85.195 57.845 85.215 ;
        RECT 58.155 85.195 58.485 85.395 ;
        RECT 56.405 84.835 57.115 85.025 ;
        RECT 56.815 84.695 57.115 84.835 ;
        RECT 57.305 84.835 58.485 85.025 ;
        RECT 58.715 84.885 59.015 85.735 ;
        RECT 59.185 85.255 59.420 85.905 ;
        RECT 59.590 85.595 59.875 86.540 ;
        RECT 60.055 86.285 60.740 86.755 ;
        RECT 60.050 85.765 60.745 86.075 ;
        RECT 60.920 85.700 61.225 86.485 ;
        RECT 59.590 85.445 60.450 85.595 ;
        RECT 61.015 85.565 61.225 85.700 ;
        RECT 61.415 85.590 61.705 86.755 ;
        RECT 61.875 86.245 62.175 86.755 ;
        RECT 62.345 86.075 62.675 86.585 ;
        RECT 62.845 86.245 63.475 86.755 ;
        RECT 64.055 86.245 64.435 86.415 ;
        RECT 64.605 86.245 64.905 86.755 ;
        RECT 64.265 86.075 64.435 86.245 ;
        RECT 61.875 85.905 64.095 86.075 ;
        RECT 59.590 85.425 60.875 85.445 ;
        RECT 59.185 84.925 59.720 85.255 ;
        RECT 59.890 85.065 60.875 85.425 ;
        RECT 57.305 84.755 57.635 84.835 ;
        RECT 56.815 84.685 57.130 84.695 ;
        RECT 56.815 84.675 57.140 84.685 ;
        RECT 56.815 84.670 57.150 84.675 ;
        RECT 56.405 84.205 56.575 84.665 ;
        RECT 56.815 84.660 57.155 84.670 ;
        RECT 56.815 84.655 57.160 84.660 ;
        RECT 56.815 84.645 57.165 84.655 ;
        RECT 56.815 84.640 57.170 84.645 ;
        RECT 56.815 84.375 57.175 84.640 ;
        RECT 57.805 84.205 57.975 84.665 ;
        RECT 58.145 84.375 58.485 84.835 ;
        RECT 59.185 84.775 59.405 84.925 ;
        RECT 58.660 84.205 58.995 84.710 ;
        RECT 59.165 84.400 59.405 84.775 ;
        RECT 59.890 84.730 60.060 85.065 ;
        RECT 61.050 84.895 61.225 85.565 ;
        RECT 61.875 84.945 62.045 85.905 ;
        RECT 62.215 85.565 63.755 85.735 ;
        RECT 62.215 85.115 62.460 85.565 ;
        RECT 62.720 85.195 63.415 85.395 ;
        RECT 63.585 85.365 63.755 85.565 ;
        RECT 63.925 85.705 64.095 85.905 ;
        RECT 64.265 85.875 64.925 86.075 ;
        RECT 63.925 85.535 64.585 85.705 ;
        RECT 63.585 85.195 64.185 85.365 ;
        RECT 64.415 85.115 64.585 85.535 ;
        RECT 59.685 84.535 60.060 84.730 ;
        RECT 59.685 84.390 59.855 84.535 ;
        RECT 60.420 84.205 60.815 84.700 ;
        RECT 60.985 84.375 61.225 84.895 ;
        RECT 61.415 84.205 61.705 84.930 ;
        RECT 61.875 84.400 62.340 84.945 ;
        RECT 62.845 84.205 63.015 85.025 ;
        RECT 63.185 84.945 64.095 85.025 ;
        RECT 64.755 84.945 64.925 85.875 ;
        RECT 65.095 85.665 68.605 86.755 ;
        RECT 68.865 86.010 69.135 86.755 ;
        RECT 69.765 86.750 76.040 86.755 ;
        RECT 69.305 85.840 69.595 86.580 ;
        RECT 69.765 86.025 70.020 86.750 ;
        RECT 70.205 85.855 70.465 86.580 ;
        RECT 70.635 86.025 70.880 86.750 ;
        RECT 71.065 85.855 71.325 86.580 ;
        RECT 71.495 86.025 71.740 86.750 ;
        RECT 71.925 85.855 72.185 86.580 ;
        RECT 72.355 86.025 72.600 86.750 ;
        RECT 72.770 85.855 73.030 86.580 ;
        RECT 73.200 86.025 73.460 86.750 ;
        RECT 73.630 85.855 73.890 86.580 ;
        RECT 74.060 86.025 74.320 86.750 ;
        RECT 74.490 85.855 74.750 86.580 ;
        RECT 74.920 86.025 75.180 86.750 ;
        RECT 75.350 85.855 75.610 86.580 ;
        RECT 75.780 85.955 76.040 86.750 ;
        RECT 70.205 85.840 75.610 85.855 ;
        RECT 63.185 84.855 64.435 84.945 ;
        RECT 63.185 84.375 63.515 84.855 ;
        RECT 63.925 84.775 64.435 84.855 ;
        RECT 63.685 84.205 64.035 84.595 ;
        RECT 64.205 84.375 64.435 84.775 ;
        RECT 64.605 84.465 64.925 84.945 ;
        RECT 65.095 84.975 66.745 85.495 ;
        RECT 66.915 85.145 68.605 85.665 ;
        RECT 68.865 85.615 75.610 85.840 ;
        RECT 68.865 85.025 70.030 85.615 ;
        RECT 76.210 85.445 76.460 86.580 ;
        RECT 76.640 85.945 76.900 86.755 ;
        RECT 77.075 85.445 77.320 86.585 ;
        RECT 77.500 85.945 77.795 86.755 ;
        RECT 77.985 86.035 78.315 86.755 ;
        RECT 70.200 85.195 77.320 85.445 ;
        RECT 65.095 84.205 68.605 84.975 ;
        RECT 68.865 84.855 75.610 85.025 ;
        RECT 68.865 84.205 69.165 84.685 ;
        RECT 69.335 84.400 69.595 84.855 ;
        RECT 69.765 84.205 70.025 84.685 ;
        RECT 70.205 84.400 70.465 84.855 ;
        RECT 70.635 84.205 70.885 84.685 ;
        RECT 71.065 84.400 71.325 84.855 ;
        RECT 71.495 84.205 71.745 84.685 ;
        RECT 71.925 84.400 72.185 84.855 ;
        RECT 72.355 84.205 72.600 84.685 ;
        RECT 72.770 84.400 73.045 84.855 ;
        RECT 73.215 84.205 73.460 84.685 ;
        RECT 73.630 84.400 73.890 84.855 ;
        RECT 74.060 84.205 74.320 84.685 ;
        RECT 74.490 84.400 74.750 84.855 ;
        RECT 74.920 84.205 75.180 84.685 ;
        RECT 75.350 84.400 75.610 84.855 ;
        RECT 75.780 84.205 76.040 84.765 ;
        RECT 76.210 84.385 76.460 85.195 ;
        RECT 76.640 84.205 76.900 84.730 ;
        RECT 77.070 84.385 77.320 85.195 ;
        RECT 77.490 84.885 77.805 85.445 ;
        RECT 77.975 85.395 78.205 85.735 ;
        RECT 78.495 85.395 78.710 86.510 ;
        RECT 78.905 85.810 79.235 86.585 ;
        RECT 79.405 85.980 80.115 86.755 ;
        RECT 78.905 85.595 80.055 85.810 ;
        RECT 77.975 85.195 78.305 85.395 ;
        RECT 78.495 85.215 78.945 85.395 ;
        RECT 78.615 85.195 78.945 85.215 ;
        RECT 79.115 85.195 79.585 85.425 ;
        RECT 79.770 85.025 80.055 85.595 ;
        RECT 80.285 85.150 80.565 86.585 ;
        RECT 80.745 85.615 81.075 86.755 ;
        RECT 81.605 85.785 81.935 86.570 ;
        RECT 81.255 85.615 81.935 85.785 ;
        RECT 82.115 85.665 85.625 86.755 ;
        RECT 85.795 85.665 87.005 86.755 ;
        RECT 80.735 85.195 81.085 85.445 ;
        RECT 77.975 84.835 79.155 85.025 ;
        RECT 77.500 84.205 77.805 84.715 ;
        RECT 77.975 84.375 78.315 84.835 ;
        RECT 78.825 84.755 79.155 84.835 ;
        RECT 79.345 84.835 80.055 85.025 ;
        RECT 79.345 84.695 79.645 84.835 ;
        RECT 79.330 84.685 79.645 84.695 ;
        RECT 79.320 84.675 79.645 84.685 ;
        RECT 79.310 84.670 79.645 84.675 ;
        RECT 78.485 84.205 78.655 84.665 ;
        RECT 79.305 84.660 79.645 84.670 ;
        RECT 79.300 84.655 79.645 84.660 ;
        RECT 79.295 84.645 79.645 84.655 ;
        RECT 79.290 84.640 79.645 84.645 ;
        RECT 79.285 84.375 79.645 84.640 ;
        RECT 79.885 84.205 80.055 84.665 ;
        RECT 80.225 84.375 80.565 85.150 ;
        RECT 81.255 85.015 81.425 85.615 ;
        RECT 81.595 85.195 81.945 85.445 ;
        RECT 80.745 84.205 81.015 85.015 ;
        RECT 81.185 84.375 81.515 85.015 ;
        RECT 81.685 84.205 81.925 85.015 ;
        RECT 82.115 84.975 83.765 85.495 ;
        RECT 83.935 85.145 85.625 85.665 ;
        RECT 82.115 84.205 85.625 84.975 ;
        RECT 85.795 84.955 86.315 85.495 ;
        RECT 86.485 85.125 87.005 85.665 ;
        RECT 87.175 85.590 87.465 86.755 ;
        RECT 87.640 85.955 87.895 86.755 ;
        RECT 88.095 85.905 88.425 86.585 ;
        RECT 87.640 85.415 87.885 85.775 ;
        RECT 88.075 85.625 88.425 85.905 ;
        RECT 88.075 85.245 88.245 85.625 ;
        RECT 88.605 85.445 88.800 86.495 ;
        RECT 88.980 85.615 89.300 86.755 ;
        RECT 90.395 85.615 90.675 86.755 ;
        RECT 90.845 85.605 91.175 86.585 ;
        RECT 91.345 85.615 91.605 86.755 ;
        RECT 91.785 86.145 92.115 86.575 ;
        RECT 92.295 86.315 92.490 86.755 ;
        RECT 92.660 86.145 92.990 86.575 ;
        RECT 91.785 85.975 92.990 86.145 ;
        RECT 91.785 85.645 92.680 85.975 ;
        RECT 93.160 85.805 93.435 86.575 ;
        RECT 92.850 85.615 93.435 85.805 ;
        RECT 93.615 85.615 93.955 86.585 ;
        RECT 94.125 85.615 94.295 86.755 ;
        RECT 94.565 85.955 94.815 86.755 ;
        RECT 95.460 85.785 95.790 86.585 ;
        RECT 96.090 85.955 96.420 86.755 ;
        RECT 96.590 85.785 96.920 86.585 ;
        RECT 94.485 85.615 96.920 85.785 ;
        RECT 97.480 85.785 97.870 85.960 ;
        RECT 98.355 85.955 98.685 86.755 ;
        RECT 98.855 85.965 99.390 86.585 ;
        RECT 97.480 85.615 98.905 85.785 ;
        RECT 87.725 85.075 88.245 85.245 ;
        RECT 88.415 85.115 88.800 85.445 ;
        RECT 88.980 85.395 89.240 85.445 ;
        RECT 88.980 85.225 89.245 85.395 ;
        RECT 88.980 85.115 89.240 85.225 ;
        RECT 90.405 85.175 90.740 85.445 ;
        RECT 85.795 84.205 87.005 84.955 ;
        RECT 87.175 84.205 87.465 84.930 ;
        RECT 87.725 84.510 87.895 85.075 ;
        RECT 90.910 85.005 91.080 85.605 ;
        RECT 91.250 85.195 91.585 85.445 ;
        RECT 91.790 85.115 92.085 85.445 ;
        RECT 92.265 85.115 92.680 85.445 ;
        RECT 88.085 84.735 89.300 84.905 ;
        RECT 88.085 84.430 88.315 84.735 ;
        RECT 88.485 84.205 88.815 84.565 ;
        RECT 89.010 84.385 89.300 84.735 ;
        RECT 90.395 84.205 90.705 85.005 ;
        RECT 90.910 84.375 91.605 85.005 ;
        RECT 91.785 84.205 92.085 84.935 ;
        RECT 92.265 84.495 92.495 85.115 ;
        RECT 92.850 84.945 93.025 85.615 ;
        RECT 92.695 84.765 93.025 84.945 ;
        RECT 93.195 84.795 93.435 85.445 ;
        RECT 93.615 85.055 93.790 85.615 ;
        RECT 94.485 85.365 94.655 85.615 ;
        RECT 93.960 85.195 94.655 85.365 ;
        RECT 94.830 85.195 95.250 85.395 ;
        RECT 95.420 85.195 95.750 85.395 ;
        RECT 95.920 85.195 96.250 85.395 ;
        RECT 93.615 85.005 93.845 85.055 ;
        RECT 92.695 84.385 92.920 84.765 ;
        RECT 93.090 84.205 93.420 84.595 ;
        RECT 93.615 84.375 93.955 85.005 ;
        RECT 94.125 84.205 94.375 85.005 ;
        RECT 94.565 84.855 95.790 85.025 ;
        RECT 94.565 84.375 94.895 84.855 ;
        RECT 95.065 84.205 95.290 84.665 ;
        RECT 95.460 84.375 95.790 84.855 ;
        RECT 96.420 84.985 96.590 85.615 ;
        RECT 96.775 85.195 97.125 85.445 ;
        RECT 96.420 84.375 96.920 84.985 ;
        RECT 97.355 84.885 97.710 85.445 ;
        RECT 97.880 84.715 98.050 85.615 ;
        RECT 98.220 84.885 98.485 85.445 ;
        RECT 98.735 85.115 98.905 85.615 ;
        RECT 99.075 84.945 99.390 85.965 ;
        RECT 97.460 84.205 97.700 84.715 ;
        RECT 97.880 84.385 98.160 84.715 ;
        RECT 98.390 84.205 98.605 84.715 ;
        RECT 98.775 84.375 99.390 84.945 ;
        RECT 100.055 85.150 100.335 86.585 ;
        RECT 100.505 85.980 101.215 86.755 ;
        RECT 101.385 85.810 101.715 86.585 ;
        RECT 100.565 85.595 101.715 85.810 ;
        RECT 100.055 84.375 100.395 85.150 ;
        RECT 100.565 85.025 100.850 85.595 ;
        RECT 101.035 85.195 101.505 85.425 ;
        RECT 101.910 85.395 102.125 86.510 ;
        RECT 102.305 86.035 102.635 86.755 ;
        RECT 102.815 86.245 103.115 86.755 ;
        RECT 103.285 86.075 103.615 86.585 ;
        RECT 103.785 86.245 104.415 86.755 ;
        RECT 104.995 86.245 105.375 86.415 ;
        RECT 105.545 86.245 105.845 86.755 ;
        RECT 105.205 86.075 105.375 86.245 ;
        RECT 102.815 85.905 105.035 86.075 ;
        RECT 102.415 85.395 102.645 85.735 ;
        RECT 101.675 85.215 102.125 85.395 ;
        RECT 101.675 85.195 102.005 85.215 ;
        RECT 102.315 85.195 102.645 85.395 ;
        RECT 100.565 84.835 101.275 85.025 ;
        RECT 100.975 84.695 101.275 84.835 ;
        RECT 101.465 84.835 102.645 85.025 ;
        RECT 101.465 84.755 101.795 84.835 ;
        RECT 100.975 84.685 101.290 84.695 ;
        RECT 100.975 84.675 101.300 84.685 ;
        RECT 100.975 84.670 101.310 84.675 ;
        RECT 100.565 84.205 100.735 84.665 ;
        RECT 100.975 84.660 101.315 84.670 ;
        RECT 100.975 84.655 101.320 84.660 ;
        RECT 100.975 84.645 101.325 84.655 ;
        RECT 100.975 84.640 101.330 84.645 ;
        RECT 100.975 84.375 101.335 84.640 ;
        RECT 101.965 84.205 102.135 84.665 ;
        RECT 102.305 84.375 102.645 84.835 ;
        RECT 102.815 84.945 102.985 85.905 ;
        RECT 103.155 85.565 104.695 85.735 ;
        RECT 103.155 85.115 103.400 85.565 ;
        RECT 103.660 85.195 104.355 85.395 ;
        RECT 104.525 85.365 104.695 85.565 ;
        RECT 104.865 85.705 105.035 85.905 ;
        RECT 105.205 85.875 105.865 86.075 ;
        RECT 104.865 85.535 105.525 85.705 ;
        RECT 104.525 85.195 105.125 85.365 ;
        RECT 105.355 85.115 105.525 85.535 ;
        RECT 102.815 84.400 103.280 84.945 ;
        RECT 103.785 84.205 103.955 85.025 ;
        RECT 104.125 84.945 105.035 85.025 ;
        RECT 105.695 84.945 105.865 85.875 ;
        RECT 104.125 84.855 105.375 84.945 ;
        RECT 104.125 84.375 104.455 84.855 ;
        RECT 104.865 84.775 105.375 84.855 ;
        RECT 104.625 84.205 104.975 84.595 ;
        RECT 105.145 84.375 105.375 84.775 ;
        RECT 105.545 84.465 105.865 84.945 ;
        RECT 106.055 85.700 106.360 86.485 ;
        RECT 106.540 86.285 107.225 86.755 ;
        RECT 106.535 85.765 107.230 86.075 ;
        RECT 106.055 85.565 106.265 85.700 ;
        RECT 107.405 85.595 107.690 86.540 ;
        RECT 107.865 86.305 108.195 86.755 ;
        RECT 108.365 86.135 108.535 86.565 ;
        RECT 109.715 86.245 110.015 86.755 ;
        RECT 106.055 84.895 106.230 85.565 ;
        RECT 106.830 85.445 107.690 85.595 ;
        RECT 106.405 85.425 107.690 85.445 ;
        RECT 107.860 85.905 108.535 86.135 ;
        RECT 110.185 86.075 110.515 86.585 ;
        RECT 110.685 86.245 111.315 86.755 ;
        RECT 111.895 86.245 112.275 86.415 ;
        RECT 112.445 86.245 112.745 86.755 ;
        RECT 112.105 86.075 112.275 86.245 ;
        RECT 109.715 85.905 111.935 86.075 ;
        RECT 106.405 85.065 107.390 85.425 ;
        RECT 107.860 85.255 108.095 85.905 ;
        RECT 106.055 84.375 106.295 84.895 ;
        RECT 107.220 84.730 107.390 85.065 ;
        RECT 107.560 84.925 108.095 85.255 ;
        RECT 107.875 84.775 108.095 84.925 ;
        RECT 108.265 84.885 108.565 85.735 ;
        RECT 109.715 84.945 109.885 85.905 ;
        RECT 110.055 85.565 111.595 85.735 ;
        RECT 110.055 85.115 110.300 85.565 ;
        RECT 110.560 85.195 111.255 85.395 ;
        RECT 111.425 85.365 111.595 85.565 ;
        RECT 111.765 85.705 111.935 85.905 ;
        RECT 112.105 85.875 112.765 86.075 ;
        RECT 111.765 85.535 112.425 85.705 ;
        RECT 111.425 85.195 112.025 85.365 ;
        RECT 112.255 85.115 112.425 85.535 ;
        RECT 106.465 84.205 106.860 84.700 ;
        RECT 107.220 84.535 107.595 84.730 ;
        RECT 107.425 84.390 107.595 84.535 ;
        RECT 107.875 84.400 108.115 84.775 ;
        RECT 108.285 84.205 108.620 84.710 ;
        RECT 109.715 84.400 110.180 84.945 ;
        RECT 110.685 84.205 110.855 85.025 ;
        RECT 111.025 84.945 111.935 85.025 ;
        RECT 112.595 84.945 112.765 85.875 ;
        RECT 112.935 85.590 113.225 86.755 ;
        RECT 114.375 85.695 114.705 86.540 ;
        RECT 114.875 85.745 115.045 86.755 ;
        RECT 115.215 86.025 115.555 86.585 ;
        RECT 115.785 86.255 116.100 86.755 ;
        RECT 116.280 86.285 117.165 86.455 ;
        RECT 114.315 85.615 114.705 85.695 ;
        RECT 115.215 85.650 116.110 86.025 ;
        RECT 111.025 84.855 112.275 84.945 ;
        RECT 111.025 84.375 111.355 84.855 ;
        RECT 111.765 84.775 112.275 84.855 ;
        RECT 111.525 84.205 111.875 84.595 ;
        RECT 112.045 84.375 112.275 84.775 ;
        RECT 112.445 84.465 112.765 84.945 ;
        RECT 114.315 85.565 114.530 85.615 ;
        RECT 114.315 84.985 114.485 85.565 ;
        RECT 115.215 85.445 115.405 85.650 ;
        RECT 116.280 85.445 116.450 86.285 ;
        RECT 117.390 86.255 117.640 86.585 ;
        RECT 114.655 85.115 115.405 85.445 ;
        RECT 115.575 85.115 116.450 85.445 ;
        RECT 114.315 84.945 114.540 84.985 ;
        RECT 115.205 84.945 115.405 85.115 ;
        RECT 112.935 84.205 113.225 84.930 ;
        RECT 114.315 84.860 114.695 84.945 ;
        RECT 114.365 84.425 114.695 84.860 ;
        RECT 114.865 84.205 115.035 84.815 ;
        RECT 115.205 84.420 115.535 84.945 ;
        RECT 115.795 84.205 116.005 84.735 ;
        RECT 116.280 84.655 116.450 85.115 ;
        RECT 116.620 85.155 116.940 86.115 ;
        RECT 117.110 85.365 117.300 86.085 ;
        RECT 117.470 85.185 117.640 86.255 ;
        RECT 117.810 85.955 117.980 86.755 ;
        RECT 118.150 86.310 119.255 86.480 ;
        RECT 118.150 85.695 118.320 86.310 ;
        RECT 119.465 86.160 119.715 86.585 ;
        RECT 119.885 86.295 120.150 86.755 ;
        RECT 118.490 85.775 119.020 86.140 ;
        RECT 119.465 86.030 119.770 86.160 ;
        RECT 117.810 85.605 118.320 85.695 ;
        RECT 117.810 85.435 118.680 85.605 ;
        RECT 117.810 85.365 117.980 85.435 ;
        RECT 118.100 85.185 118.300 85.215 ;
        RECT 116.620 84.825 117.085 85.155 ;
        RECT 117.470 84.885 118.300 85.185 ;
        RECT 117.470 84.655 117.640 84.885 ;
        RECT 116.280 84.485 117.065 84.655 ;
        RECT 117.235 84.485 117.640 84.655 ;
        RECT 117.820 84.205 118.190 84.705 ;
        RECT 118.510 84.655 118.680 85.435 ;
        RECT 118.850 85.075 119.020 85.775 ;
        RECT 119.190 85.245 119.430 85.840 ;
        RECT 118.850 84.855 119.375 85.075 ;
        RECT 119.600 84.925 119.770 86.030 ;
        RECT 119.545 84.795 119.770 84.925 ;
        RECT 119.940 84.835 120.220 85.785 ;
        RECT 119.545 84.655 119.715 84.795 ;
        RECT 118.510 84.485 119.185 84.655 ;
        RECT 119.380 84.485 119.715 84.655 ;
        RECT 119.885 84.205 120.135 84.665 ;
        RECT 120.390 84.465 120.575 86.585 ;
        RECT 120.745 86.255 121.075 86.755 ;
        RECT 121.245 86.085 121.415 86.585 ;
        RECT 120.750 85.915 121.415 86.085 ;
        RECT 121.765 86.085 121.935 86.585 ;
        RECT 122.105 86.255 122.435 86.755 ;
        RECT 121.765 85.915 122.370 86.085 ;
        RECT 120.750 84.925 120.980 85.915 ;
        RECT 121.150 85.095 121.500 85.745 ;
        RECT 121.675 85.105 121.920 85.745 ;
        RECT 122.200 85.520 122.370 85.915 ;
        RECT 122.605 85.805 122.830 86.585 ;
        RECT 122.200 85.190 122.430 85.520 ;
        RECT 122.200 84.925 122.370 85.190 ;
        RECT 120.750 84.755 121.415 84.925 ;
        RECT 120.745 84.205 121.075 84.585 ;
        RECT 121.245 84.465 121.415 84.755 ;
        RECT 121.765 84.755 122.370 84.925 ;
        RECT 121.765 84.465 121.935 84.755 ;
        RECT 122.105 84.205 122.435 84.585 ;
        RECT 122.605 84.465 122.775 85.805 ;
        RECT 123.020 85.785 123.375 86.535 ;
        RECT 123.545 85.955 123.835 86.755 ;
        RECT 124.335 86.375 125.195 86.545 ;
        RECT 124.885 86.225 125.195 86.375 ;
        RECT 125.365 86.295 125.685 86.755 ;
        RECT 124.885 86.210 125.210 86.225 ;
        RECT 124.980 86.205 125.210 86.210 ;
        RECT 124.980 86.185 125.220 86.205 ;
        RECT 124.980 86.165 125.235 86.185 ;
        RECT 124.995 86.155 125.235 86.165 ;
        RECT 125.020 86.130 125.235 86.155 ;
        RECT 123.020 85.615 123.705 85.785 ;
        RECT 123.025 85.075 123.355 85.445 ;
        RECT 123.535 85.355 123.705 85.615 ;
        RECT 124.035 85.475 124.370 86.125 ;
        RECT 124.540 85.680 124.875 86.030 ;
        RECT 123.535 84.905 123.910 85.355 ;
        RECT 124.540 85.160 124.855 85.680 ;
        RECT 125.045 85.570 125.235 86.130 ;
        RECT 125.885 85.985 126.130 86.555 ;
        RECT 125.405 85.655 126.130 85.985 ;
        RECT 126.310 85.690 126.595 86.755 ;
        RECT 126.765 85.790 127.025 86.575 ;
        RECT 127.285 86.085 127.455 86.585 ;
        RECT 127.625 86.255 127.955 86.755 ;
        RECT 127.285 85.915 127.890 86.085 ;
        RECT 123.100 84.885 123.910 84.905 ;
        RECT 123.100 84.735 123.705 84.885 ;
        RECT 124.150 84.855 124.855 85.160 ;
        RECT 125.025 85.445 125.235 85.570 ;
        RECT 125.960 85.445 126.130 85.655 ;
        RECT 125.025 85.115 125.790 85.445 ;
        RECT 125.960 85.115 126.685 85.445 ;
        RECT 123.100 84.465 123.295 84.735 ;
        RECT 125.025 84.655 125.195 85.115 ;
        RECT 125.960 84.840 126.130 85.115 ;
        RECT 126.855 84.865 127.025 85.790 ;
        RECT 127.195 85.105 127.440 85.745 ;
        RECT 127.720 85.520 127.890 85.915 ;
        RECT 128.125 85.805 128.350 86.585 ;
        RECT 127.720 85.190 127.950 85.520 ;
        RECT 127.720 84.925 127.890 85.190 ;
        RECT 123.465 84.205 123.795 84.565 ;
        RECT 124.355 84.485 125.195 84.655 ;
        RECT 125.365 84.205 125.635 84.665 ;
        RECT 125.885 84.380 126.130 84.840 ;
        RECT 126.345 84.205 126.570 84.835 ;
        RECT 126.765 84.535 127.025 84.865 ;
        RECT 127.285 84.755 127.890 84.925 ;
        RECT 127.285 84.465 127.455 84.755 ;
        RECT 127.625 84.205 127.955 84.585 ;
        RECT 128.125 84.465 128.295 85.805 ;
        RECT 128.540 85.785 128.895 86.535 ;
        RECT 129.065 85.955 129.355 86.755 ;
        RECT 129.855 86.375 130.715 86.545 ;
        RECT 130.405 86.225 130.715 86.375 ;
        RECT 130.885 86.295 131.205 86.755 ;
        RECT 130.405 86.210 130.730 86.225 ;
        RECT 130.500 86.205 130.730 86.210 ;
        RECT 130.500 86.185 130.740 86.205 ;
        RECT 130.500 86.165 130.755 86.185 ;
        RECT 130.515 86.155 130.755 86.165 ;
        RECT 130.540 86.130 130.755 86.155 ;
        RECT 128.540 85.615 129.225 85.785 ;
        RECT 128.545 85.075 128.875 85.445 ;
        RECT 129.055 85.355 129.225 85.615 ;
        RECT 129.555 85.475 129.890 86.125 ;
        RECT 130.060 85.680 130.395 86.030 ;
        RECT 129.055 84.905 129.430 85.355 ;
        RECT 130.060 85.160 130.375 85.680 ;
        RECT 130.565 85.570 130.755 86.130 ;
        RECT 131.405 85.985 131.650 86.555 ;
        RECT 130.925 85.655 131.650 85.985 ;
        RECT 131.830 85.690 132.115 86.755 ;
        RECT 132.285 85.790 132.545 86.575 ;
        RECT 132.805 86.085 132.975 86.585 ;
        RECT 133.145 86.255 133.475 86.755 ;
        RECT 132.805 85.915 133.410 86.085 ;
        RECT 128.620 84.885 129.430 84.905 ;
        RECT 128.620 84.735 129.225 84.885 ;
        RECT 129.670 84.855 130.375 85.160 ;
        RECT 130.545 85.445 130.755 85.570 ;
        RECT 131.480 85.445 131.650 85.655 ;
        RECT 130.545 85.115 131.310 85.445 ;
        RECT 131.480 85.115 132.205 85.445 ;
        RECT 128.620 84.465 128.815 84.735 ;
        RECT 130.545 84.655 130.715 85.115 ;
        RECT 131.480 84.840 131.650 85.115 ;
        RECT 132.375 84.865 132.545 85.790 ;
        RECT 132.715 85.105 132.960 85.745 ;
        RECT 133.240 85.520 133.410 85.915 ;
        RECT 133.645 85.805 133.870 86.585 ;
        RECT 133.240 85.190 133.470 85.520 ;
        RECT 133.240 84.925 133.410 85.190 ;
        RECT 128.985 84.205 129.315 84.565 ;
        RECT 129.875 84.485 130.715 84.655 ;
        RECT 130.885 84.205 131.155 84.665 ;
        RECT 131.405 84.380 131.650 84.840 ;
        RECT 131.865 84.205 132.090 84.835 ;
        RECT 132.285 84.535 132.545 84.865 ;
        RECT 132.805 84.755 133.410 84.925 ;
        RECT 132.805 84.465 132.975 84.755 ;
        RECT 133.145 84.205 133.475 84.585 ;
        RECT 133.645 84.465 133.815 85.805 ;
        RECT 134.060 85.785 134.415 86.535 ;
        RECT 134.585 85.955 134.875 86.755 ;
        RECT 135.375 86.375 136.235 86.545 ;
        RECT 135.925 86.225 136.235 86.375 ;
        RECT 136.405 86.295 136.725 86.755 ;
        RECT 135.925 86.210 136.250 86.225 ;
        RECT 136.020 86.205 136.250 86.210 ;
        RECT 136.020 86.185 136.260 86.205 ;
        RECT 136.020 86.165 136.275 86.185 ;
        RECT 136.035 86.155 136.275 86.165 ;
        RECT 136.060 86.130 136.275 86.155 ;
        RECT 134.060 85.615 134.745 85.785 ;
        RECT 134.065 85.075 134.395 85.445 ;
        RECT 134.575 85.355 134.745 85.615 ;
        RECT 135.075 85.475 135.410 86.125 ;
        RECT 135.580 85.680 135.915 86.030 ;
        RECT 134.575 84.905 134.950 85.355 ;
        RECT 135.580 85.160 135.895 85.680 ;
        RECT 136.085 85.570 136.275 86.130 ;
        RECT 136.925 85.985 137.170 86.555 ;
        RECT 136.445 85.655 137.170 85.985 ;
        RECT 137.350 85.690 137.635 86.755 ;
        RECT 137.805 85.790 138.065 86.575 ;
        RECT 134.140 84.885 134.950 84.905 ;
        RECT 134.140 84.735 134.745 84.885 ;
        RECT 135.190 84.855 135.895 85.160 ;
        RECT 136.065 85.445 136.275 85.570 ;
        RECT 137.000 85.445 137.170 85.655 ;
        RECT 136.065 85.115 136.830 85.445 ;
        RECT 137.000 85.115 137.725 85.445 ;
        RECT 134.140 84.465 134.335 84.735 ;
        RECT 136.065 84.655 136.235 85.115 ;
        RECT 137.000 84.840 137.170 85.115 ;
        RECT 137.895 84.865 138.065 85.790 ;
        RECT 138.695 85.590 138.985 86.755 ;
        RECT 139.155 85.035 139.675 86.585 ;
        RECT 139.845 86.030 140.175 86.755 ;
        RECT 141.085 86.085 141.255 86.585 ;
        RECT 141.425 86.255 141.755 86.755 ;
        RECT 141.085 85.915 141.750 86.085 ;
        RECT 134.505 84.205 134.835 84.565 ;
        RECT 135.395 84.485 136.235 84.655 ;
        RECT 136.405 84.205 136.675 84.665 ;
        RECT 136.925 84.380 137.170 84.840 ;
        RECT 137.385 84.205 137.610 84.835 ;
        RECT 137.805 84.535 138.065 84.865 ;
        RECT 138.695 84.205 138.985 84.930 ;
        RECT 139.335 84.205 139.675 84.865 ;
        RECT 139.845 84.375 140.365 85.860 ;
        RECT 141.000 85.095 141.350 85.745 ;
        RECT 141.520 84.925 141.750 85.915 ;
        RECT 141.085 84.755 141.750 84.925 ;
        RECT 141.085 84.465 141.255 84.755 ;
        RECT 141.425 84.205 141.755 84.585 ;
        RECT 141.925 84.465 142.110 86.585 ;
        RECT 142.350 86.295 142.615 86.755 ;
        RECT 142.785 86.160 143.035 86.585 ;
        RECT 143.245 86.310 144.350 86.480 ;
        RECT 142.730 86.030 143.035 86.160 ;
        RECT 142.280 84.835 142.560 85.785 ;
        RECT 142.730 84.925 142.900 86.030 ;
        RECT 143.070 85.245 143.310 85.840 ;
        RECT 143.480 85.775 144.010 86.140 ;
        RECT 143.480 85.075 143.650 85.775 ;
        RECT 144.180 85.695 144.350 86.310 ;
        RECT 144.520 85.955 144.690 86.755 ;
        RECT 144.860 86.255 145.110 86.585 ;
        RECT 145.335 86.285 146.220 86.455 ;
        RECT 144.180 85.605 144.690 85.695 ;
        RECT 142.730 84.795 142.955 84.925 ;
        RECT 143.125 84.855 143.650 85.075 ;
        RECT 143.820 85.435 144.690 85.605 ;
        RECT 142.365 84.205 142.615 84.665 ;
        RECT 142.785 84.655 142.955 84.795 ;
        RECT 143.820 84.655 143.990 85.435 ;
        RECT 144.520 85.365 144.690 85.435 ;
        RECT 144.200 85.185 144.400 85.215 ;
        RECT 144.860 85.185 145.030 86.255 ;
        RECT 145.200 85.365 145.390 86.085 ;
        RECT 144.200 84.885 145.030 85.185 ;
        RECT 145.560 85.155 145.880 86.115 ;
        RECT 142.785 84.485 143.120 84.655 ;
        RECT 143.315 84.485 143.990 84.655 ;
        RECT 144.310 84.205 144.680 84.705 ;
        RECT 144.860 84.655 145.030 84.885 ;
        RECT 145.415 84.825 145.880 85.155 ;
        RECT 146.050 85.445 146.220 86.285 ;
        RECT 146.400 86.255 146.715 86.755 ;
        RECT 146.945 86.025 147.285 86.585 ;
        RECT 146.390 85.650 147.285 86.025 ;
        RECT 147.455 85.745 147.625 86.755 ;
        RECT 147.095 85.445 147.285 85.650 ;
        RECT 147.795 85.695 148.125 86.540 ;
        RECT 149.295 86.245 149.595 86.755 ;
        RECT 149.765 86.245 150.145 86.415 ;
        RECT 150.725 86.245 151.355 86.755 ;
        RECT 149.765 86.075 149.935 86.245 ;
        RECT 151.525 86.075 151.855 86.585 ;
        RECT 152.025 86.245 152.325 86.755 ;
        RECT 149.275 85.875 149.935 86.075 ;
        RECT 150.105 85.905 152.325 86.075 ;
        RECT 147.795 85.615 148.185 85.695 ;
        RECT 147.970 85.565 148.185 85.615 ;
        RECT 146.050 85.115 146.925 85.445 ;
        RECT 147.095 85.115 147.845 85.445 ;
        RECT 146.050 84.655 146.220 85.115 ;
        RECT 147.095 84.945 147.295 85.115 ;
        RECT 148.015 84.985 148.185 85.565 ;
        RECT 147.960 84.945 148.185 84.985 ;
        RECT 144.860 84.485 145.265 84.655 ;
        RECT 145.435 84.485 146.220 84.655 ;
        RECT 146.495 84.205 146.705 84.735 ;
        RECT 146.965 84.420 147.295 84.945 ;
        RECT 147.805 84.860 148.185 84.945 ;
        RECT 149.275 84.945 149.445 85.875 ;
        RECT 150.105 85.705 150.275 85.905 ;
        RECT 149.615 85.535 150.275 85.705 ;
        RECT 150.445 85.565 151.985 85.735 ;
        RECT 149.615 85.115 149.785 85.535 ;
        RECT 150.445 85.365 150.615 85.565 ;
        RECT 150.015 85.195 150.615 85.365 ;
        RECT 150.785 85.195 151.480 85.395 ;
        RECT 151.740 85.115 151.985 85.565 ;
        RECT 150.105 84.945 151.015 85.025 ;
        RECT 147.465 84.205 147.635 84.815 ;
        RECT 147.805 84.425 148.135 84.860 ;
        RECT 149.275 84.465 149.595 84.945 ;
        RECT 149.765 84.855 151.015 84.945 ;
        RECT 149.765 84.775 150.275 84.855 ;
        RECT 149.765 84.375 149.995 84.775 ;
        RECT 150.165 84.205 150.515 84.595 ;
        RECT 150.685 84.375 151.015 84.855 ;
        RECT 151.185 84.205 151.355 85.025 ;
        RECT 152.155 84.945 152.325 85.905 ;
        RECT 151.860 84.400 152.325 84.945 ;
        RECT 152.515 85.700 152.820 86.485 ;
        RECT 153.000 86.285 153.685 86.755 ;
        RECT 152.995 85.765 153.690 86.075 ;
        RECT 152.515 85.565 152.725 85.700 ;
        RECT 153.865 85.595 154.150 86.540 ;
        RECT 154.325 86.305 154.655 86.755 ;
        RECT 154.825 86.135 154.995 86.565 ;
        RECT 152.515 84.895 152.690 85.565 ;
        RECT 153.290 85.445 154.150 85.595 ;
        RECT 152.865 85.425 154.150 85.445 ;
        RECT 154.320 85.905 154.995 86.135 ;
        RECT 152.865 85.065 153.850 85.425 ;
        RECT 154.320 85.255 154.555 85.905 ;
        RECT 152.515 84.375 152.755 84.895 ;
        RECT 153.680 84.730 153.850 85.065 ;
        RECT 154.020 84.925 154.555 85.255 ;
        RECT 154.335 84.775 154.555 84.925 ;
        RECT 154.725 84.885 155.025 85.735 ;
        RECT 155.715 85.665 156.925 86.755 ;
        RECT 155.715 85.125 156.235 85.665 ;
        RECT 156.405 84.955 156.925 85.495 ;
        RECT 152.925 84.205 153.320 84.700 ;
        RECT 153.680 84.535 154.055 84.730 ;
        RECT 153.885 84.390 154.055 84.535 ;
        RECT 154.335 84.400 154.575 84.775 ;
        RECT 154.745 84.205 155.080 84.710 ;
        RECT 155.715 84.205 156.925 84.955 ;
        RECT 22.690 84.035 157.010 84.205 ;
        RECT 22.775 83.285 23.985 84.035 ;
        RECT 22.775 82.745 23.295 83.285 ;
        RECT 24.155 83.265 25.825 84.035 ;
        RECT 26.635 83.375 26.975 84.035 ;
        RECT 23.465 82.575 23.985 83.115 ;
        RECT 24.155 82.745 24.905 83.265 ;
        RECT 25.075 82.575 25.825 83.095 ;
        RECT 22.775 81.485 23.985 82.575 ;
        RECT 24.155 81.485 25.825 82.575 ;
        RECT 26.455 81.655 26.975 83.205 ;
        RECT 27.145 82.380 27.665 83.865 ;
        RECT 27.835 83.265 30.425 84.035 ;
        RECT 27.835 82.745 29.045 83.265 ;
        RECT 29.215 82.575 30.425 83.095 ;
        RECT 27.145 81.485 27.475 82.210 ;
        RECT 27.835 81.485 30.425 82.575 ;
        RECT 30.595 83.090 30.935 83.865 ;
        RECT 31.105 83.575 31.275 84.035 ;
        RECT 31.515 83.600 31.875 83.865 ;
        RECT 31.515 83.595 31.870 83.600 ;
        RECT 31.515 83.585 31.865 83.595 ;
        RECT 31.515 83.580 31.860 83.585 ;
        RECT 31.515 83.570 31.855 83.580 ;
        RECT 32.505 83.575 32.675 84.035 ;
        RECT 31.515 83.565 31.850 83.570 ;
        RECT 31.515 83.555 31.840 83.565 ;
        RECT 31.515 83.545 31.830 83.555 ;
        RECT 31.515 83.405 31.815 83.545 ;
        RECT 31.105 83.215 31.815 83.405 ;
        RECT 32.005 83.405 32.335 83.485 ;
        RECT 32.845 83.405 33.185 83.865 ;
        RECT 32.005 83.215 33.185 83.405 ;
        RECT 33.445 83.485 33.615 83.775 ;
        RECT 33.785 83.655 34.115 84.035 ;
        RECT 33.445 83.315 34.050 83.485 ;
        RECT 30.595 81.655 30.875 83.090 ;
        RECT 31.105 82.645 31.390 83.215 ;
        RECT 31.575 82.815 32.045 83.045 ;
        RECT 32.215 83.025 32.545 83.045 ;
        RECT 32.215 82.845 32.665 83.025 ;
        RECT 32.855 82.845 33.185 83.045 ;
        RECT 31.105 82.430 32.255 82.645 ;
        RECT 31.045 81.485 31.755 82.260 ;
        RECT 31.925 81.655 32.255 82.430 ;
        RECT 32.450 81.730 32.665 82.845 ;
        RECT 32.955 82.505 33.185 82.845 ;
        RECT 33.355 82.495 33.600 83.135 ;
        RECT 33.880 83.050 34.050 83.315 ;
        RECT 33.880 82.720 34.110 83.050 ;
        RECT 33.880 82.325 34.050 82.720 ;
        RECT 32.845 81.485 33.175 82.205 ;
        RECT 33.445 82.155 34.050 82.325 ;
        RECT 34.285 82.435 34.455 83.775 ;
        RECT 34.780 83.505 34.975 83.775 ;
        RECT 35.145 83.675 35.475 84.035 ;
        RECT 36.035 83.585 36.875 83.755 ;
        RECT 34.780 83.355 35.385 83.505 ;
        RECT 34.780 83.335 35.590 83.355 ;
        RECT 34.705 82.795 35.035 83.165 ;
        RECT 35.215 82.885 35.590 83.335 ;
        RECT 35.830 83.080 36.535 83.385 ;
        RECT 35.215 82.625 35.385 82.885 ;
        RECT 34.700 82.455 35.385 82.625 ;
        RECT 33.445 81.655 33.615 82.155 ;
        RECT 33.785 81.485 34.115 81.985 ;
        RECT 34.285 81.655 34.510 82.435 ;
        RECT 34.700 81.705 35.055 82.455 ;
        RECT 35.225 81.485 35.515 82.285 ;
        RECT 35.715 82.115 36.050 82.765 ;
        RECT 36.220 82.560 36.535 83.080 ;
        RECT 36.705 83.125 36.875 83.585 ;
        RECT 37.045 83.575 37.315 84.035 ;
        RECT 37.565 83.400 37.810 83.860 ;
        RECT 38.025 83.405 38.250 84.035 ;
        RECT 37.640 83.125 37.810 83.400 ;
        RECT 38.445 83.375 38.705 83.705 ;
        RECT 36.705 82.795 37.470 83.125 ;
        RECT 37.640 82.795 38.365 83.125 ;
        RECT 36.705 82.670 36.915 82.795 ;
        RECT 36.220 82.210 36.555 82.560 ;
        RECT 36.725 82.110 36.915 82.670 ;
        RECT 37.640 82.585 37.810 82.795 ;
        RECT 37.085 82.255 37.810 82.585 ;
        RECT 36.700 82.085 36.915 82.110 ;
        RECT 36.675 82.075 36.915 82.085 ;
        RECT 36.660 82.055 36.915 82.075 ;
        RECT 36.660 82.035 36.900 82.055 ;
        RECT 36.660 82.030 36.890 82.035 ;
        RECT 36.565 82.015 36.890 82.030 ;
        RECT 36.565 81.865 36.875 82.015 ;
        RECT 36.015 81.695 36.875 81.865 ;
        RECT 37.045 81.485 37.365 81.945 ;
        RECT 37.565 81.685 37.810 82.255 ;
        RECT 37.990 81.485 38.275 82.550 ;
        RECT 38.535 82.450 38.705 83.375 ;
        RECT 38.875 83.265 42.385 84.035 ;
        RECT 42.555 83.375 42.815 83.705 ;
        RECT 43.010 83.405 43.235 84.035 ;
        RECT 43.450 83.400 43.695 83.860 ;
        RECT 43.945 83.575 44.215 84.035 ;
        RECT 44.385 83.585 45.225 83.755 ;
        RECT 45.785 83.675 46.115 84.035 ;
        RECT 38.875 82.745 40.525 83.265 ;
        RECT 40.695 82.575 42.385 83.095 ;
        RECT 38.445 81.665 38.705 82.450 ;
        RECT 38.875 81.485 42.385 82.575 ;
        RECT 42.555 82.450 42.725 83.375 ;
        RECT 43.450 83.125 43.620 83.400 ;
        RECT 44.385 83.125 44.555 83.585 ;
        RECT 46.285 83.505 46.480 83.775 ;
        RECT 42.895 82.795 43.620 83.125 ;
        RECT 43.790 82.795 44.555 83.125 ;
        RECT 43.450 82.585 43.620 82.795 ;
        RECT 44.345 82.670 44.555 82.795 ;
        RECT 44.725 83.080 45.430 83.385 ;
        RECT 45.875 83.355 46.480 83.505 ;
        RECT 45.670 83.335 46.480 83.355 ;
        RECT 42.555 81.665 42.815 82.450 ;
        RECT 42.985 81.485 43.270 82.550 ;
        RECT 43.450 82.255 44.175 82.585 ;
        RECT 43.450 81.685 43.695 82.255 ;
        RECT 44.345 82.110 44.535 82.670 ;
        RECT 44.725 82.560 45.040 83.080 ;
        RECT 45.670 82.885 46.045 83.335 ;
        RECT 44.705 82.210 45.040 82.560 ;
        RECT 45.210 82.115 45.545 82.765 ;
        RECT 45.875 82.625 46.045 82.885 ;
        RECT 46.225 82.795 46.555 83.165 ;
        RECT 45.875 82.455 46.560 82.625 ;
        RECT 44.345 82.085 44.560 82.110 ;
        RECT 44.345 82.075 44.585 82.085 ;
        RECT 44.345 82.055 44.600 82.075 ;
        RECT 44.360 82.035 44.600 82.055 ;
        RECT 44.370 82.030 44.600 82.035 ;
        RECT 44.370 82.015 44.695 82.030 ;
        RECT 43.895 81.485 44.215 81.945 ;
        RECT 44.385 81.865 44.695 82.015 ;
        RECT 44.385 81.695 45.245 81.865 ;
        RECT 45.745 81.485 46.035 82.285 ;
        RECT 46.205 81.705 46.560 82.455 ;
        RECT 46.805 82.435 46.975 83.775 ;
        RECT 47.145 83.655 47.475 84.035 ;
        RECT 47.645 83.485 47.815 83.775 ;
        RECT 47.210 83.315 47.815 83.485 ;
        RECT 47.210 83.050 47.380 83.315 ;
        RECT 48.535 83.310 48.825 84.035 ;
        RECT 49.085 83.485 49.255 83.775 ;
        RECT 49.425 83.655 49.755 84.035 ;
        RECT 49.085 83.315 49.690 83.485 ;
        RECT 47.150 82.720 47.380 83.050 ;
        RECT 46.750 81.655 46.975 82.435 ;
        RECT 47.210 82.325 47.380 82.720 ;
        RECT 47.660 82.495 47.905 83.135 ;
        RECT 47.210 82.155 47.815 82.325 ;
        RECT 47.145 81.485 47.475 81.985 ;
        RECT 47.645 81.655 47.815 82.155 ;
        RECT 48.535 81.485 48.825 82.650 ;
        RECT 48.995 82.495 49.240 83.135 ;
        RECT 49.520 83.050 49.690 83.315 ;
        RECT 49.520 82.720 49.750 83.050 ;
        RECT 49.520 82.325 49.690 82.720 ;
        RECT 49.085 82.155 49.690 82.325 ;
        RECT 49.925 82.435 50.095 83.775 ;
        RECT 50.420 83.505 50.615 83.775 ;
        RECT 50.785 83.675 51.115 84.035 ;
        RECT 51.675 83.585 52.515 83.755 ;
        RECT 50.420 83.355 51.025 83.505 ;
        RECT 50.420 83.335 51.230 83.355 ;
        RECT 50.345 82.795 50.675 83.165 ;
        RECT 50.855 82.885 51.230 83.335 ;
        RECT 51.470 83.080 52.175 83.385 ;
        RECT 50.855 82.625 51.025 82.885 ;
        RECT 50.340 82.455 51.025 82.625 ;
        RECT 49.085 81.655 49.255 82.155 ;
        RECT 49.425 81.485 49.755 81.985 ;
        RECT 49.925 81.655 50.150 82.435 ;
        RECT 50.340 81.705 50.695 82.455 ;
        RECT 50.865 81.485 51.155 82.285 ;
        RECT 51.355 82.115 51.690 82.765 ;
        RECT 51.860 82.560 52.175 83.080 ;
        RECT 52.345 83.125 52.515 83.585 ;
        RECT 52.685 83.575 52.955 84.035 ;
        RECT 53.205 83.400 53.450 83.860 ;
        RECT 53.665 83.405 53.890 84.035 ;
        RECT 53.280 83.125 53.450 83.400 ;
        RECT 54.085 83.375 54.345 83.705 ;
        RECT 54.695 83.375 55.035 84.035 ;
        RECT 52.345 82.795 53.110 83.125 ;
        RECT 53.280 82.795 54.005 83.125 ;
        RECT 52.345 82.670 52.555 82.795 ;
        RECT 51.860 82.210 52.195 82.560 ;
        RECT 52.365 82.110 52.555 82.670 ;
        RECT 53.280 82.585 53.450 82.795 ;
        RECT 52.725 82.255 53.450 82.585 ;
        RECT 52.340 82.085 52.555 82.110 ;
        RECT 52.315 82.075 52.555 82.085 ;
        RECT 52.300 82.055 52.555 82.075 ;
        RECT 52.300 82.035 52.540 82.055 ;
        RECT 52.300 82.030 52.530 82.035 ;
        RECT 52.205 82.015 52.530 82.030 ;
        RECT 52.205 81.865 52.515 82.015 ;
        RECT 51.655 81.695 52.515 81.865 ;
        RECT 52.685 81.485 53.005 81.945 ;
        RECT 53.205 81.685 53.450 82.255 ;
        RECT 53.630 81.485 53.915 82.550 ;
        RECT 54.175 82.450 54.345 83.375 ;
        RECT 54.085 81.665 54.345 82.450 ;
        RECT 54.515 81.655 55.035 83.205 ;
        RECT 55.205 82.380 55.725 83.865 ;
        RECT 55.895 83.265 58.485 84.035 ;
        RECT 55.895 82.745 57.105 83.265 ;
        RECT 58.665 83.225 58.935 84.035 ;
        RECT 59.105 83.225 59.435 83.865 ;
        RECT 59.605 83.225 59.845 84.035 ;
        RECT 60.035 83.235 60.730 83.865 ;
        RECT 60.935 83.235 61.245 84.035 ;
        RECT 61.415 83.265 64.925 84.035 ;
        RECT 65.605 83.380 65.935 83.815 ;
        RECT 66.105 83.425 66.275 84.035 ;
        RECT 65.555 83.295 65.935 83.380 ;
        RECT 66.445 83.295 66.775 83.820 ;
        RECT 67.035 83.505 67.245 84.035 ;
        RECT 67.520 83.585 68.305 83.755 ;
        RECT 68.475 83.585 68.880 83.755 ;
        RECT 57.275 82.575 58.485 83.095 ;
        RECT 58.655 82.795 59.005 83.045 ;
        RECT 59.175 82.625 59.345 83.225 ;
        RECT 59.515 82.795 59.865 83.045 ;
        RECT 60.055 82.795 60.390 83.045 ;
        RECT 60.560 82.635 60.730 83.235 ;
        RECT 60.900 82.795 61.235 83.065 ;
        RECT 61.415 82.745 63.065 83.265 ;
        RECT 65.555 83.255 65.780 83.295 ;
        RECT 55.205 81.485 55.535 82.210 ;
        RECT 55.895 81.485 58.485 82.575 ;
        RECT 58.665 81.485 58.995 82.625 ;
        RECT 59.175 82.455 59.855 82.625 ;
        RECT 59.525 81.670 59.855 82.455 ;
        RECT 60.035 81.485 60.295 82.625 ;
        RECT 60.465 81.655 60.795 82.635 ;
        RECT 60.965 81.485 61.245 82.625 ;
        RECT 63.235 82.575 64.925 83.095 ;
        RECT 61.415 81.485 64.925 82.575 ;
        RECT 65.555 82.675 65.725 83.255 ;
        RECT 66.445 83.125 66.645 83.295 ;
        RECT 67.520 83.125 67.690 83.585 ;
        RECT 65.895 82.795 66.645 83.125 ;
        RECT 66.815 82.795 67.690 83.125 ;
        RECT 65.555 82.625 65.770 82.675 ;
        RECT 65.555 82.545 65.945 82.625 ;
        RECT 65.615 81.700 65.945 82.545 ;
        RECT 66.455 82.590 66.645 82.795 ;
        RECT 66.115 81.485 66.285 82.495 ;
        RECT 66.455 82.215 67.350 82.590 ;
        RECT 66.455 81.655 66.795 82.215 ;
        RECT 67.025 81.485 67.340 81.985 ;
        RECT 67.520 81.955 67.690 82.795 ;
        RECT 67.860 83.085 68.325 83.415 ;
        RECT 68.710 83.355 68.880 83.585 ;
        RECT 69.060 83.535 69.430 84.035 ;
        RECT 69.750 83.585 70.425 83.755 ;
        RECT 70.620 83.585 70.955 83.755 ;
        RECT 67.860 82.125 68.180 83.085 ;
        RECT 68.710 83.055 69.540 83.355 ;
        RECT 68.350 82.155 68.540 82.875 ;
        RECT 68.710 81.985 68.880 83.055 ;
        RECT 69.340 83.025 69.540 83.055 ;
        RECT 69.050 82.805 69.220 82.875 ;
        RECT 69.750 82.805 69.920 83.585 ;
        RECT 70.785 83.445 70.955 83.585 ;
        RECT 71.125 83.575 71.375 84.035 ;
        RECT 69.050 82.635 69.920 82.805 ;
        RECT 70.090 83.165 70.615 83.385 ;
        RECT 70.785 83.315 71.010 83.445 ;
        RECT 69.050 82.545 69.560 82.635 ;
        RECT 67.520 81.785 68.405 81.955 ;
        RECT 68.630 81.655 68.880 81.985 ;
        RECT 69.050 81.485 69.220 82.285 ;
        RECT 69.390 81.930 69.560 82.545 ;
        RECT 70.090 82.465 70.260 83.165 ;
        RECT 69.730 82.100 70.260 82.465 ;
        RECT 70.430 82.400 70.670 82.995 ;
        RECT 70.840 82.210 71.010 83.315 ;
        RECT 71.180 82.455 71.460 83.405 ;
        RECT 70.705 82.080 71.010 82.210 ;
        RECT 69.390 81.760 70.495 81.930 ;
        RECT 70.705 81.655 70.955 82.080 ;
        RECT 71.125 81.485 71.390 81.945 ;
        RECT 71.630 81.655 71.815 83.775 ;
        RECT 71.985 83.655 72.315 84.035 ;
        RECT 72.485 83.485 72.655 83.775 ;
        RECT 71.990 83.315 72.655 83.485 ;
        RECT 71.990 82.325 72.220 83.315 ;
        RECT 72.915 83.285 74.125 84.035 ;
        RECT 74.295 83.310 74.585 84.035 ;
        RECT 74.805 83.645 75.135 84.035 ;
        RECT 75.305 83.465 75.475 83.785 ;
        RECT 75.645 83.645 75.975 84.035 ;
        RECT 76.390 83.635 77.345 83.805 ;
        RECT 74.755 83.295 77.005 83.465 ;
        RECT 72.390 82.495 72.740 83.145 ;
        RECT 72.915 82.745 73.435 83.285 ;
        RECT 73.605 82.575 74.125 83.115 ;
        RECT 71.990 82.155 72.655 82.325 ;
        RECT 71.985 81.485 72.315 81.985 ;
        RECT 72.485 81.655 72.655 82.155 ;
        RECT 72.915 81.485 74.125 82.575 ;
        RECT 74.295 81.485 74.585 82.650 ;
        RECT 74.755 82.335 74.925 83.295 ;
        RECT 75.095 82.675 75.340 83.125 ;
        RECT 75.510 82.845 76.060 83.045 ;
        RECT 76.230 82.875 76.605 83.045 ;
        RECT 76.230 82.675 76.400 82.875 ;
        RECT 76.775 82.795 77.005 83.295 ;
        RECT 75.095 82.505 76.400 82.675 ;
        RECT 77.175 82.755 77.345 83.635 ;
        RECT 77.515 83.200 77.805 84.035 ;
        RECT 77.175 82.585 77.805 82.755 ;
        RECT 74.755 81.655 75.135 82.335 ;
        RECT 75.725 81.485 75.895 82.335 ;
        RECT 76.065 82.165 77.305 82.335 ;
        RECT 76.065 81.655 76.395 82.165 ;
        RECT 76.565 81.485 76.735 81.995 ;
        RECT 76.905 81.655 77.305 82.165 ;
        RECT 77.485 81.655 77.805 82.585 ;
        RECT 77.975 82.380 78.495 83.865 ;
        RECT 78.665 83.375 79.005 84.035 ;
        RECT 79.355 83.265 81.025 84.035 ;
        RECT 81.195 83.405 81.535 83.865 ;
        RECT 81.705 83.575 81.875 84.035 ;
        RECT 82.505 83.600 82.865 83.865 ;
        RECT 82.510 83.595 82.865 83.600 ;
        RECT 82.515 83.585 82.865 83.595 ;
        RECT 82.520 83.580 82.865 83.585 ;
        RECT 82.525 83.570 82.865 83.580 ;
        RECT 83.105 83.575 83.275 84.035 ;
        RECT 82.530 83.565 82.865 83.570 ;
        RECT 82.540 83.555 82.865 83.565 ;
        RECT 82.550 83.545 82.865 83.555 ;
        RECT 82.045 83.405 82.375 83.485 ;
        RECT 78.165 81.485 78.495 82.210 ;
        RECT 78.665 81.655 79.185 83.205 ;
        RECT 79.355 82.745 80.105 83.265 ;
        RECT 81.195 83.215 82.375 83.405 ;
        RECT 82.565 83.405 82.865 83.545 ;
        RECT 82.565 83.215 83.275 83.405 ;
        RECT 80.275 82.575 81.025 83.095 ;
        RECT 79.355 81.485 81.025 82.575 ;
        RECT 81.195 82.845 81.525 83.045 ;
        RECT 81.835 83.025 82.165 83.045 ;
        RECT 81.715 82.845 82.165 83.025 ;
        RECT 81.195 82.505 81.425 82.845 ;
        RECT 81.205 81.485 81.535 82.205 ;
        RECT 81.715 81.730 81.930 82.845 ;
        RECT 82.335 82.815 82.805 83.045 ;
        RECT 82.990 82.645 83.275 83.215 ;
        RECT 83.445 83.090 83.785 83.865 ;
        RECT 84.965 83.485 85.135 83.775 ;
        RECT 85.305 83.655 85.635 84.035 ;
        RECT 84.965 83.315 85.570 83.485 ;
        RECT 82.125 82.430 83.275 82.645 ;
        RECT 82.125 81.655 82.455 82.430 ;
        RECT 82.625 81.485 83.335 82.260 ;
        RECT 83.505 81.655 83.785 83.090 ;
        RECT 84.875 82.495 85.120 83.135 ;
        RECT 85.400 83.050 85.570 83.315 ;
        RECT 85.400 82.720 85.630 83.050 ;
        RECT 85.400 82.325 85.570 82.720 ;
        RECT 84.965 82.155 85.570 82.325 ;
        RECT 85.805 82.435 85.975 83.775 ;
        RECT 86.300 83.505 86.495 83.775 ;
        RECT 86.665 83.675 86.995 84.035 ;
        RECT 87.555 83.585 88.395 83.755 ;
        RECT 86.300 83.355 86.905 83.505 ;
        RECT 86.300 83.335 87.110 83.355 ;
        RECT 86.225 82.795 86.555 83.165 ;
        RECT 86.735 82.885 87.110 83.335 ;
        RECT 87.350 83.080 88.055 83.385 ;
        RECT 86.735 82.625 86.905 82.885 ;
        RECT 86.220 82.455 86.905 82.625 ;
        RECT 84.965 81.655 85.135 82.155 ;
        RECT 85.305 81.485 85.635 81.985 ;
        RECT 85.805 81.655 86.030 82.435 ;
        RECT 86.220 81.705 86.575 82.455 ;
        RECT 86.745 81.485 87.035 82.285 ;
        RECT 87.235 82.115 87.570 82.765 ;
        RECT 87.740 82.560 88.055 83.080 ;
        RECT 88.225 83.125 88.395 83.585 ;
        RECT 88.565 83.575 88.835 84.035 ;
        RECT 89.085 83.400 89.330 83.860 ;
        RECT 89.545 83.405 89.770 84.035 ;
        RECT 89.160 83.125 89.330 83.400 ;
        RECT 89.965 83.375 90.225 83.705 ;
        RECT 91.035 83.375 91.375 84.035 ;
        RECT 88.225 82.795 88.990 83.125 ;
        RECT 89.160 82.795 89.885 83.125 ;
        RECT 88.225 82.670 88.435 82.795 ;
        RECT 87.740 82.210 88.075 82.560 ;
        RECT 88.245 82.110 88.435 82.670 ;
        RECT 89.160 82.585 89.330 82.795 ;
        RECT 88.605 82.255 89.330 82.585 ;
        RECT 88.220 82.085 88.435 82.110 ;
        RECT 88.195 82.075 88.435 82.085 ;
        RECT 88.180 82.055 88.435 82.075 ;
        RECT 88.180 82.035 88.420 82.055 ;
        RECT 88.180 82.030 88.410 82.035 ;
        RECT 88.085 82.015 88.410 82.030 ;
        RECT 88.085 81.865 88.395 82.015 ;
        RECT 87.535 81.695 88.395 81.865 ;
        RECT 88.565 81.485 88.885 81.945 ;
        RECT 89.085 81.685 89.330 82.255 ;
        RECT 89.510 81.485 89.795 82.550 ;
        RECT 90.055 82.450 90.225 83.375 ;
        RECT 89.965 81.665 90.225 82.450 ;
        RECT 90.855 81.655 91.375 83.205 ;
        RECT 91.545 82.380 92.065 83.865 ;
        RECT 92.235 83.265 93.905 84.035 ;
        RECT 92.235 82.745 92.985 83.265 ;
        RECT 94.535 83.235 94.845 84.035 ;
        RECT 95.050 83.235 95.745 83.865 ;
        RECT 95.915 83.265 97.585 84.035 ;
        RECT 98.395 83.375 98.735 84.035 ;
        RECT 93.155 82.575 93.905 83.095 ;
        RECT 94.545 82.795 94.880 83.065 ;
        RECT 95.050 82.635 95.220 83.235 ;
        RECT 95.390 82.795 95.725 83.045 ;
        RECT 95.915 82.745 96.665 83.265 ;
        RECT 91.545 81.485 91.875 82.210 ;
        RECT 92.235 81.485 93.905 82.575 ;
        RECT 94.535 81.485 94.815 82.625 ;
        RECT 94.985 81.655 95.315 82.635 ;
        RECT 95.485 81.485 95.745 82.625 ;
        RECT 96.835 82.575 97.585 83.095 ;
        RECT 95.915 81.485 97.585 82.575 ;
        RECT 98.215 81.655 98.735 83.205 ;
        RECT 98.905 82.380 99.425 83.865 ;
        RECT 100.055 83.310 100.345 84.035 ;
        RECT 100.515 83.265 102.185 84.035 ;
        RECT 100.515 82.745 101.265 83.265 ;
        RECT 102.825 83.225 103.095 84.035 ;
        RECT 103.265 83.225 103.595 83.865 ;
        RECT 103.765 83.225 104.005 84.035 ;
        RECT 104.195 83.265 107.705 84.035 ;
        RECT 98.905 81.485 99.235 82.210 ;
        RECT 100.055 81.485 100.345 82.650 ;
        RECT 101.435 82.575 102.185 83.095 ;
        RECT 102.815 82.795 103.165 83.045 ;
        RECT 103.335 82.625 103.505 83.225 ;
        RECT 103.675 82.795 104.025 83.045 ;
        RECT 104.195 82.745 105.845 83.265 ;
        RECT 100.515 81.485 102.185 82.575 ;
        RECT 102.825 81.485 103.155 82.625 ;
        RECT 103.335 82.455 104.015 82.625 ;
        RECT 106.015 82.575 107.705 83.095 ;
        RECT 103.685 81.670 104.015 82.455 ;
        RECT 104.195 81.485 107.705 82.575 ;
        RECT 107.875 83.090 108.215 83.865 ;
        RECT 108.385 83.575 108.555 84.035 ;
        RECT 108.795 83.600 109.155 83.865 ;
        RECT 108.795 83.595 109.150 83.600 ;
        RECT 108.795 83.585 109.145 83.595 ;
        RECT 108.795 83.580 109.140 83.585 ;
        RECT 108.795 83.570 109.135 83.580 ;
        RECT 109.785 83.575 109.955 84.035 ;
        RECT 108.795 83.565 109.130 83.570 ;
        RECT 108.795 83.555 109.120 83.565 ;
        RECT 108.795 83.545 109.110 83.555 ;
        RECT 108.795 83.405 109.095 83.545 ;
        RECT 108.385 83.215 109.095 83.405 ;
        RECT 109.285 83.405 109.615 83.485 ;
        RECT 110.125 83.405 110.465 83.865 ;
        RECT 109.285 83.215 110.465 83.405 ;
        RECT 110.645 83.225 110.915 84.035 ;
        RECT 111.085 83.225 111.415 83.865 ;
        RECT 111.585 83.225 111.825 84.035 ;
        RECT 112.015 83.235 112.710 83.865 ;
        RECT 112.915 83.235 113.225 84.035 ;
        RECT 113.395 83.490 118.740 84.035 ;
        RECT 107.875 81.655 108.155 83.090 ;
        RECT 108.385 82.645 108.670 83.215 ;
        RECT 108.855 82.815 109.325 83.045 ;
        RECT 109.495 83.025 109.825 83.045 ;
        RECT 109.495 82.845 109.945 83.025 ;
        RECT 110.135 82.845 110.465 83.045 ;
        RECT 108.385 82.430 109.535 82.645 ;
        RECT 108.325 81.485 109.035 82.260 ;
        RECT 109.205 81.655 109.535 82.430 ;
        RECT 109.730 81.730 109.945 82.845 ;
        RECT 110.235 82.505 110.465 82.845 ;
        RECT 110.635 82.795 110.985 83.045 ;
        RECT 111.155 82.625 111.325 83.225 ;
        RECT 111.495 82.795 111.845 83.045 ;
        RECT 112.035 82.795 112.370 83.045 ;
        RECT 112.540 82.635 112.710 83.235 ;
        RECT 112.880 82.795 113.215 83.065 ;
        RECT 114.980 82.660 115.320 83.490 ;
        RECT 118.915 83.265 122.425 84.035 ;
        RECT 122.595 83.285 123.805 84.035 ;
        RECT 110.125 81.485 110.455 82.205 ;
        RECT 110.645 81.485 110.975 82.625 ;
        RECT 111.155 82.455 111.835 82.625 ;
        RECT 111.505 81.670 111.835 82.455 ;
        RECT 112.015 81.485 112.275 82.625 ;
        RECT 112.445 81.655 112.775 82.635 ;
        RECT 112.945 81.485 113.225 82.625 ;
        RECT 116.800 81.920 117.150 83.170 ;
        RECT 118.915 82.745 120.565 83.265 ;
        RECT 120.735 82.575 122.425 83.095 ;
        RECT 122.595 82.745 123.115 83.285 ;
        RECT 123.285 82.575 123.805 83.115 ;
        RECT 113.395 81.485 118.740 81.920 ;
        RECT 118.915 81.485 122.425 82.575 ;
        RECT 122.595 81.485 123.805 82.575 ;
        RECT 123.975 82.380 124.495 83.865 ;
        RECT 124.665 83.375 125.005 84.035 ;
        RECT 125.815 83.310 126.105 84.035 ;
        RECT 126.275 83.490 131.620 84.035 ;
        RECT 124.165 81.485 124.495 82.210 ;
        RECT 124.665 81.655 125.185 83.205 ;
        RECT 127.860 82.660 128.200 83.490 ;
        RECT 132.895 83.375 133.235 84.035 ;
        RECT 125.815 81.485 126.105 82.650 ;
        RECT 129.680 81.920 130.030 83.170 ;
        RECT 126.275 81.485 131.620 81.920 ;
        RECT 132.715 81.655 133.235 83.205 ;
        RECT 133.405 82.380 133.925 83.865 ;
        RECT 134.095 83.360 134.355 83.865 ;
        RECT 134.535 83.655 134.865 84.035 ;
        RECT 135.045 83.485 135.215 83.865 ;
        RECT 134.095 82.560 134.265 83.360 ;
        RECT 134.550 83.315 135.215 83.485 ;
        RECT 136.025 83.485 136.195 83.865 ;
        RECT 136.375 83.655 136.705 84.035 ;
        RECT 136.025 83.315 136.690 83.485 ;
        RECT 136.885 83.360 137.145 83.865 ;
        RECT 134.550 83.060 134.720 83.315 ;
        RECT 134.435 82.730 134.720 83.060 ;
        RECT 134.955 82.765 135.285 83.135 ;
        RECT 135.955 82.765 136.285 83.135 ;
        RECT 136.520 83.060 136.690 83.315 ;
        RECT 134.550 82.585 134.720 82.730 ;
        RECT 136.520 82.730 136.805 83.060 ;
        RECT 136.520 82.585 136.690 82.730 ;
        RECT 133.405 81.485 133.735 82.210 ;
        RECT 134.095 81.655 134.365 82.560 ;
        RECT 134.550 82.415 135.215 82.585 ;
        RECT 134.535 81.485 134.865 82.245 ;
        RECT 135.045 81.655 135.215 82.415 ;
        RECT 136.025 82.415 136.690 82.585 ;
        RECT 136.975 82.560 137.145 83.360 ;
        RECT 137.405 83.485 137.575 83.775 ;
        RECT 137.745 83.655 138.075 84.035 ;
        RECT 137.405 83.315 138.010 83.485 ;
        RECT 136.025 81.655 136.195 82.415 ;
        RECT 136.375 81.485 136.705 82.245 ;
        RECT 136.875 81.655 137.145 82.560 ;
        RECT 137.315 82.495 137.560 83.135 ;
        RECT 137.840 83.050 138.010 83.315 ;
        RECT 137.840 82.720 138.070 83.050 ;
        RECT 137.840 82.325 138.010 82.720 ;
        RECT 137.405 82.155 138.010 82.325 ;
        RECT 138.245 82.435 138.415 83.775 ;
        RECT 138.740 83.505 138.935 83.775 ;
        RECT 139.105 83.675 139.435 84.035 ;
        RECT 139.995 83.585 140.835 83.755 ;
        RECT 138.740 83.355 139.345 83.505 ;
        RECT 138.740 83.335 139.550 83.355 ;
        RECT 138.665 82.795 138.995 83.165 ;
        RECT 139.175 82.885 139.550 83.335 ;
        RECT 139.790 83.080 140.495 83.385 ;
        RECT 139.175 82.625 139.345 82.885 ;
        RECT 138.660 82.455 139.345 82.625 ;
        RECT 137.405 81.655 137.575 82.155 ;
        RECT 137.745 81.485 138.075 81.985 ;
        RECT 138.245 81.655 138.470 82.435 ;
        RECT 138.660 81.705 139.015 82.455 ;
        RECT 139.185 81.485 139.475 82.285 ;
        RECT 139.675 82.115 140.010 82.765 ;
        RECT 140.180 82.560 140.495 83.080 ;
        RECT 140.665 83.125 140.835 83.585 ;
        RECT 141.005 83.575 141.275 84.035 ;
        RECT 141.525 83.400 141.770 83.860 ;
        RECT 141.985 83.405 142.210 84.035 ;
        RECT 141.600 83.125 141.770 83.400 ;
        RECT 142.405 83.375 142.665 83.705 ;
        RECT 143.015 83.375 143.355 84.035 ;
        RECT 140.665 82.795 141.430 83.125 ;
        RECT 141.600 82.795 142.325 83.125 ;
        RECT 140.665 82.670 140.875 82.795 ;
        RECT 140.180 82.210 140.515 82.560 ;
        RECT 140.685 82.110 140.875 82.670 ;
        RECT 141.600 82.585 141.770 82.795 ;
        RECT 141.045 82.255 141.770 82.585 ;
        RECT 140.660 82.085 140.875 82.110 ;
        RECT 140.635 82.075 140.875 82.085 ;
        RECT 140.620 82.055 140.875 82.075 ;
        RECT 140.620 82.035 140.860 82.055 ;
        RECT 140.620 82.030 140.850 82.035 ;
        RECT 140.525 82.015 140.850 82.030 ;
        RECT 140.525 81.865 140.835 82.015 ;
        RECT 139.975 81.695 140.835 81.865 ;
        RECT 141.005 81.485 141.325 81.945 ;
        RECT 141.525 81.685 141.770 82.255 ;
        RECT 141.950 81.485 142.235 82.550 ;
        RECT 142.495 82.450 142.665 83.375 ;
        RECT 142.405 81.665 142.665 82.450 ;
        RECT 142.835 81.655 143.355 83.205 ;
        RECT 143.525 82.380 144.045 83.865 ;
        RECT 144.215 83.265 146.805 84.035 ;
        RECT 144.215 82.745 145.425 83.265 ;
        RECT 145.595 82.575 146.805 83.095 ;
        RECT 143.525 81.485 143.855 82.210 ;
        RECT 144.215 81.485 146.805 82.575 ;
        RECT 146.975 83.090 147.315 83.865 ;
        RECT 147.485 83.575 147.655 84.035 ;
        RECT 147.895 83.600 148.255 83.865 ;
        RECT 147.895 83.595 148.250 83.600 ;
        RECT 147.895 83.585 148.245 83.595 ;
        RECT 147.895 83.580 148.240 83.585 ;
        RECT 147.895 83.570 148.235 83.580 ;
        RECT 148.885 83.575 149.055 84.035 ;
        RECT 147.895 83.565 148.230 83.570 ;
        RECT 147.895 83.555 148.220 83.565 ;
        RECT 147.895 83.545 148.210 83.555 ;
        RECT 147.895 83.405 148.195 83.545 ;
        RECT 147.485 83.215 148.195 83.405 ;
        RECT 148.385 83.405 148.715 83.485 ;
        RECT 149.225 83.405 149.565 83.865 ;
        RECT 148.385 83.215 149.565 83.405 ;
        RECT 149.735 83.265 151.405 84.035 ;
        RECT 151.575 83.310 151.865 84.035 ;
        RECT 152.035 83.265 155.545 84.035 ;
        RECT 155.715 83.285 156.925 84.035 ;
        RECT 146.975 81.655 147.255 83.090 ;
        RECT 147.485 82.645 147.770 83.215 ;
        RECT 147.955 82.815 148.425 83.045 ;
        RECT 148.595 83.025 148.925 83.045 ;
        RECT 148.595 82.845 149.045 83.025 ;
        RECT 149.235 82.845 149.565 83.045 ;
        RECT 147.485 82.430 148.635 82.645 ;
        RECT 147.425 81.485 148.135 82.260 ;
        RECT 148.305 81.655 148.635 82.430 ;
        RECT 148.830 81.730 149.045 82.845 ;
        RECT 149.335 82.505 149.565 82.845 ;
        RECT 149.735 82.745 150.485 83.265 ;
        RECT 150.655 82.575 151.405 83.095 ;
        RECT 152.035 82.745 153.685 83.265 ;
        RECT 149.225 81.485 149.555 82.205 ;
        RECT 149.735 81.485 151.405 82.575 ;
        RECT 151.575 81.485 151.865 82.650 ;
        RECT 153.855 82.575 155.545 83.095 ;
        RECT 152.035 81.485 155.545 82.575 ;
        RECT 155.715 82.575 156.235 83.115 ;
        RECT 156.405 82.745 156.925 83.285 ;
        RECT 155.715 81.485 156.925 82.575 ;
        RECT 22.690 81.315 157.010 81.485 ;
        RECT 22.775 80.225 23.985 81.315 ;
        RECT 24.805 80.590 25.135 81.315 ;
        RECT 22.775 79.515 23.295 80.055 ;
        RECT 23.465 79.685 23.985 80.225 ;
        RECT 22.775 78.765 23.985 79.515 ;
        RECT 24.615 78.935 25.135 80.420 ;
        RECT 25.305 79.595 25.825 81.145 ;
        RECT 26.085 80.645 26.255 81.145 ;
        RECT 26.425 80.815 26.755 81.315 ;
        RECT 26.085 80.475 26.690 80.645 ;
        RECT 25.995 79.665 26.240 80.305 ;
        RECT 26.520 80.080 26.690 80.475 ;
        RECT 26.925 80.365 27.150 81.145 ;
        RECT 26.520 79.750 26.750 80.080 ;
        RECT 26.520 79.485 26.690 79.750 ;
        RECT 25.305 78.765 25.645 79.425 ;
        RECT 26.085 79.315 26.690 79.485 ;
        RECT 26.085 79.025 26.255 79.315 ;
        RECT 26.425 78.765 26.755 79.145 ;
        RECT 26.925 79.025 27.095 80.365 ;
        RECT 27.340 80.345 27.695 81.095 ;
        RECT 27.865 80.515 28.155 81.315 ;
        RECT 28.655 80.935 29.515 81.105 ;
        RECT 29.205 80.785 29.515 80.935 ;
        RECT 29.685 80.855 30.005 81.315 ;
        RECT 29.205 80.770 29.530 80.785 ;
        RECT 29.300 80.765 29.530 80.770 ;
        RECT 29.300 80.745 29.540 80.765 ;
        RECT 29.300 80.725 29.555 80.745 ;
        RECT 29.315 80.715 29.555 80.725 ;
        RECT 29.340 80.690 29.555 80.715 ;
        RECT 27.340 80.175 28.025 80.345 ;
        RECT 27.345 79.635 27.675 80.005 ;
        RECT 27.855 79.915 28.025 80.175 ;
        RECT 28.355 80.035 28.690 80.685 ;
        RECT 28.860 80.240 29.195 80.590 ;
        RECT 27.855 79.465 28.230 79.915 ;
        RECT 28.860 79.720 29.175 80.240 ;
        RECT 29.365 80.130 29.555 80.690 ;
        RECT 30.205 80.545 30.450 81.115 ;
        RECT 29.725 80.215 30.450 80.545 ;
        RECT 30.630 80.250 30.915 81.315 ;
        RECT 31.085 80.350 31.345 81.135 ;
        RECT 27.420 79.445 28.230 79.465 ;
        RECT 27.420 79.295 28.025 79.445 ;
        RECT 28.470 79.415 29.175 79.720 ;
        RECT 29.345 80.005 29.555 80.130 ;
        RECT 30.280 80.005 30.450 80.215 ;
        RECT 29.345 79.675 30.110 80.005 ;
        RECT 30.280 79.675 31.005 80.005 ;
        RECT 27.420 79.025 27.615 79.295 ;
        RECT 29.345 79.215 29.515 79.675 ;
        RECT 30.280 79.400 30.450 79.675 ;
        RECT 31.175 79.425 31.345 80.350 ;
        RECT 31.515 80.225 33.185 81.315 ;
        RECT 27.785 78.765 28.115 79.125 ;
        RECT 28.675 79.045 29.515 79.215 ;
        RECT 29.685 78.765 29.955 79.225 ;
        RECT 30.205 78.940 30.450 79.400 ;
        RECT 30.665 78.765 30.890 79.395 ;
        RECT 31.085 79.095 31.345 79.425 ;
        RECT 31.515 79.535 32.265 80.055 ;
        RECT 32.435 79.705 33.185 80.225 ;
        RECT 33.365 80.345 33.695 81.130 ;
        RECT 33.365 80.175 34.045 80.345 ;
        RECT 34.225 80.175 34.555 81.315 ;
        RECT 33.355 79.755 33.705 80.005 ;
        RECT 33.875 79.575 34.045 80.175 ;
        RECT 35.655 80.150 35.945 81.315 ;
        RECT 36.115 80.880 41.460 81.315 ;
        RECT 34.215 79.755 34.565 80.005 ;
        RECT 31.515 78.765 33.185 79.535 ;
        RECT 33.375 78.765 33.615 79.575 ;
        RECT 33.785 78.935 34.115 79.575 ;
        RECT 34.285 78.765 34.555 79.575 ;
        RECT 35.655 78.765 35.945 79.490 ;
        RECT 37.700 79.310 38.040 80.140 ;
        RECT 39.520 79.630 39.870 80.880 ;
        RECT 41.635 80.225 44.225 81.315 ;
        RECT 41.635 79.535 42.845 80.055 ;
        RECT 43.015 79.705 44.225 80.225 ;
        RECT 44.485 80.385 44.655 81.145 ;
        RECT 44.835 80.555 45.165 81.315 ;
        RECT 44.485 80.215 45.150 80.385 ;
        RECT 45.335 80.240 45.605 81.145 ;
        RECT 44.980 80.070 45.150 80.215 ;
        RECT 44.415 79.665 44.745 80.035 ;
        RECT 44.980 79.740 45.265 80.070 ;
        RECT 36.115 78.765 41.460 79.310 ;
        RECT 41.635 78.765 44.225 79.535 ;
        RECT 44.980 79.485 45.150 79.740 ;
        RECT 44.485 79.315 45.150 79.485 ;
        RECT 45.435 79.440 45.605 80.240 ;
        RECT 45.775 80.225 48.365 81.315 ;
        RECT 44.485 78.935 44.655 79.315 ;
        RECT 44.835 78.765 45.165 79.145 ;
        RECT 45.345 78.935 45.605 79.440 ;
        RECT 45.775 79.535 46.985 80.055 ;
        RECT 47.155 79.705 48.365 80.225 ;
        RECT 48.625 80.385 48.795 81.145 ;
        RECT 48.975 80.555 49.305 81.315 ;
        RECT 48.625 80.215 49.290 80.385 ;
        RECT 49.475 80.240 49.745 81.145 ;
        RECT 49.120 80.070 49.290 80.215 ;
        RECT 48.555 79.665 48.885 80.035 ;
        RECT 49.120 79.740 49.405 80.070 ;
        RECT 45.775 78.765 48.365 79.535 ;
        RECT 49.120 79.485 49.290 79.740 ;
        RECT 48.625 79.315 49.290 79.485 ;
        RECT 49.575 79.440 49.745 80.240 ;
        RECT 49.915 80.225 51.585 81.315 ;
        RECT 48.625 78.935 48.795 79.315 ;
        RECT 48.975 78.765 49.305 79.145 ;
        RECT 49.485 78.935 49.745 79.440 ;
        RECT 49.915 79.535 50.665 80.055 ;
        RECT 50.835 79.705 51.585 80.225 ;
        RECT 51.845 80.385 52.015 81.145 ;
        RECT 52.195 80.555 52.525 81.315 ;
        RECT 51.845 80.215 52.510 80.385 ;
        RECT 52.695 80.240 52.965 81.145 ;
        RECT 53.225 80.645 53.395 81.145 ;
        RECT 53.565 80.815 53.895 81.315 ;
        RECT 53.225 80.475 53.830 80.645 ;
        RECT 52.340 80.070 52.510 80.215 ;
        RECT 51.775 79.665 52.105 80.035 ;
        RECT 52.340 79.740 52.625 80.070 ;
        RECT 49.915 78.765 51.585 79.535 ;
        RECT 52.340 79.485 52.510 79.740 ;
        RECT 51.845 79.315 52.510 79.485 ;
        RECT 52.795 79.440 52.965 80.240 ;
        RECT 53.135 79.665 53.380 80.305 ;
        RECT 53.660 80.080 53.830 80.475 ;
        RECT 54.065 80.365 54.290 81.145 ;
        RECT 53.660 79.750 53.890 80.080 ;
        RECT 53.660 79.485 53.830 79.750 ;
        RECT 51.845 78.935 52.015 79.315 ;
        RECT 52.195 78.765 52.525 79.145 ;
        RECT 52.705 78.935 52.965 79.440 ;
        RECT 53.225 79.315 53.830 79.485 ;
        RECT 53.225 79.025 53.395 79.315 ;
        RECT 53.565 78.765 53.895 79.145 ;
        RECT 54.065 79.025 54.235 80.365 ;
        RECT 54.480 80.345 54.835 81.095 ;
        RECT 55.005 80.515 55.295 81.315 ;
        RECT 55.795 80.935 56.655 81.105 ;
        RECT 56.345 80.785 56.655 80.935 ;
        RECT 56.825 80.855 57.145 81.315 ;
        RECT 56.345 80.770 56.670 80.785 ;
        RECT 56.440 80.765 56.670 80.770 ;
        RECT 56.440 80.745 56.680 80.765 ;
        RECT 56.440 80.725 56.695 80.745 ;
        RECT 56.455 80.715 56.695 80.725 ;
        RECT 56.480 80.690 56.695 80.715 ;
        RECT 54.480 80.175 55.165 80.345 ;
        RECT 54.485 79.635 54.815 80.005 ;
        RECT 54.995 79.915 55.165 80.175 ;
        RECT 55.495 80.035 55.830 80.685 ;
        RECT 56.000 80.240 56.335 80.590 ;
        RECT 54.995 79.465 55.370 79.915 ;
        RECT 56.000 79.720 56.315 80.240 ;
        RECT 56.505 80.130 56.695 80.690 ;
        RECT 57.345 80.545 57.590 81.115 ;
        RECT 56.865 80.215 57.590 80.545 ;
        RECT 57.770 80.250 58.055 81.315 ;
        RECT 58.225 80.350 58.485 81.135 ;
        RECT 54.560 79.445 55.370 79.465 ;
        RECT 54.560 79.295 55.165 79.445 ;
        RECT 55.610 79.415 56.315 79.720 ;
        RECT 56.485 80.005 56.695 80.130 ;
        RECT 57.420 80.005 57.590 80.215 ;
        RECT 56.485 79.675 57.250 80.005 ;
        RECT 57.420 79.675 58.145 80.005 ;
        RECT 54.560 79.025 54.755 79.295 ;
        RECT 56.485 79.215 56.655 79.675 ;
        RECT 57.420 79.400 57.590 79.675 ;
        RECT 58.315 79.425 58.485 80.350 ;
        RECT 58.655 80.225 61.245 81.315 ;
        RECT 54.925 78.765 55.255 79.125 ;
        RECT 55.815 79.045 56.655 79.215 ;
        RECT 56.825 78.765 57.095 79.225 ;
        RECT 57.345 78.940 57.590 79.400 ;
        RECT 57.805 78.765 58.030 79.395 ;
        RECT 58.225 79.095 58.485 79.425 ;
        RECT 58.655 79.535 59.865 80.055 ;
        RECT 60.035 79.705 61.245 80.225 ;
        RECT 61.415 80.150 61.705 81.315 ;
        RECT 62.340 80.175 62.660 81.315 ;
        RECT 62.840 80.005 63.035 81.055 ;
        RECT 63.215 80.465 63.545 81.145 ;
        RECT 63.745 80.515 64.000 81.315 ;
        RECT 64.175 80.880 69.520 81.315 ;
        RECT 63.215 80.185 63.565 80.465 ;
        RECT 62.400 79.955 62.660 80.005 ;
        RECT 62.395 79.785 62.660 79.955 ;
        RECT 62.400 79.675 62.660 79.785 ;
        RECT 62.840 79.675 63.225 80.005 ;
        RECT 63.395 79.805 63.565 80.185 ;
        RECT 63.755 79.975 64.000 80.335 ;
        RECT 63.395 79.635 63.915 79.805 ;
        RECT 58.655 78.765 61.245 79.535 ;
        RECT 61.415 78.765 61.705 79.490 ;
        RECT 62.340 79.295 63.555 79.465 ;
        RECT 62.340 78.945 62.630 79.295 ;
        RECT 62.825 78.765 63.155 79.125 ;
        RECT 63.325 78.990 63.555 79.295 ;
        RECT 63.745 79.275 63.915 79.635 ;
        RECT 65.760 79.310 66.100 80.140 ;
        RECT 67.580 79.630 67.930 80.880 ;
        RECT 70.165 80.725 70.425 81.115 ;
        RECT 70.595 80.905 70.925 81.315 ;
        RECT 70.165 80.525 70.925 80.725 ;
        RECT 70.175 79.655 70.405 80.345 ;
        RECT 70.585 79.845 70.925 80.525 ;
        RECT 71.115 80.025 71.445 81.135 ;
        RECT 71.615 80.405 71.805 81.135 ;
        RECT 71.975 80.585 72.305 81.315 ;
        RECT 72.485 80.405 72.655 81.135 ;
        RECT 73.105 80.590 73.435 81.315 ;
        RECT 71.615 80.205 72.655 80.405 ;
        RECT 70.585 79.395 70.815 79.845 ;
        RECT 71.115 79.725 71.650 80.025 ;
        RECT 63.745 79.105 63.945 79.275 ;
        RECT 63.745 79.070 63.915 79.105 ;
        RECT 64.175 78.765 69.520 79.310 ;
        RECT 70.435 78.945 70.815 79.395 ;
        RECT 70.995 78.765 71.225 79.545 ;
        RECT 71.405 79.475 71.650 79.725 ;
        RECT 71.830 79.675 72.225 80.025 ;
        RECT 72.420 79.675 72.710 80.025 ;
        RECT 71.405 78.945 71.835 79.475 ;
        RECT 72.015 79.055 72.225 79.675 ;
        RECT 72.395 78.765 72.725 79.495 ;
        RECT 72.915 78.935 73.435 80.420 ;
        RECT 73.605 79.595 74.125 81.145 ;
        RECT 74.295 80.225 75.965 81.315 ;
        RECT 74.295 79.535 75.045 80.055 ;
        RECT 75.215 79.705 75.965 80.225 ;
        RECT 76.135 80.350 76.395 81.135 ;
        RECT 73.605 78.765 73.945 79.425 ;
        RECT 74.295 78.765 75.965 79.535 ;
        RECT 76.135 79.425 76.305 80.350 ;
        RECT 76.565 80.250 76.850 81.315 ;
        RECT 77.030 80.545 77.275 81.115 ;
        RECT 77.475 80.855 77.795 81.315 ;
        RECT 77.965 80.935 78.825 81.105 ;
        RECT 77.965 80.785 78.275 80.935 ;
        RECT 77.950 80.770 78.275 80.785 ;
        RECT 77.950 80.765 78.180 80.770 ;
        RECT 77.940 80.745 78.180 80.765 ;
        RECT 77.925 80.725 78.180 80.745 ;
        RECT 77.925 80.715 78.165 80.725 ;
        RECT 77.925 80.690 78.140 80.715 ;
        RECT 77.030 80.215 77.755 80.545 ;
        RECT 77.030 80.005 77.200 80.215 ;
        RECT 77.925 80.130 78.115 80.690 ;
        RECT 78.285 80.240 78.620 80.590 ;
        RECT 77.925 80.005 78.135 80.130 ;
        RECT 76.475 79.675 77.200 80.005 ;
        RECT 77.370 79.675 78.135 80.005 ;
        RECT 76.135 79.095 76.395 79.425 ;
        RECT 77.030 79.400 77.200 79.675 ;
        RECT 76.590 78.765 76.815 79.395 ;
        RECT 77.030 78.940 77.275 79.400 ;
        RECT 77.525 78.765 77.795 79.225 ;
        RECT 77.965 79.215 78.135 79.675 ;
        RECT 78.305 79.720 78.620 80.240 ;
        RECT 78.790 80.035 79.125 80.685 ;
        RECT 79.325 80.515 79.615 81.315 ;
        RECT 79.785 80.345 80.140 81.095 ;
        RECT 80.330 80.365 80.555 81.145 ;
        RECT 80.725 80.815 81.055 81.315 ;
        RECT 81.225 80.645 81.395 81.145 ;
        RECT 79.455 80.175 80.140 80.345 ;
        RECT 79.455 79.915 79.625 80.175 ;
        RECT 78.305 79.415 79.010 79.720 ;
        RECT 79.250 79.465 79.625 79.915 ;
        RECT 79.805 79.635 80.135 80.005 ;
        RECT 79.250 79.445 80.060 79.465 ;
        RECT 79.455 79.295 80.060 79.445 ;
        RECT 77.965 79.045 78.805 79.215 ;
        RECT 79.365 78.765 79.695 79.125 ;
        RECT 79.865 79.025 80.060 79.295 ;
        RECT 80.385 79.025 80.555 80.365 ;
        RECT 80.790 80.475 81.395 80.645 ;
        RECT 80.790 80.080 80.960 80.475 ;
        RECT 80.730 79.750 80.960 80.080 ;
        RECT 80.790 79.485 80.960 79.750 ;
        RECT 81.240 79.665 81.485 80.305 ;
        RECT 82.585 80.175 82.915 81.315 ;
        RECT 83.445 80.345 83.775 81.130 ;
        RECT 83.095 80.175 83.775 80.345 ;
        RECT 82.575 79.755 82.925 80.005 ;
        RECT 83.095 79.575 83.265 80.175 ;
        RECT 83.435 79.755 83.785 80.005 ;
        RECT 84.875 79.595 85.395 81.145 ;
        RECT 85.565 80.590 85.895 81.315 ;
        RECT 80.790 79.315 81.395 79.485 ;
        RECT 80.725 78.765 81.055 79.145 ;
        RECT 81.225 79.025 81.395 79.315 ;
        RECT 82.585 78.765 82.855 79.575 ;
        RECT 83.025 78.935 83.355 79.575 ;
        RECT 83.525 78.765 83.765 79.575 ;
        RECT 85.055 78.765 85.395 79.425 ;
        RECT 85.565 78.935 86.085 80.420 ;
        RECT 87.175 80.150 87.465 81.315 ;
        RECT 87.635 80.225 90.225 81.315 ;
        RECT 90.945 80.645 91.115 81.145 ;
        RECT 91.285 80.815 91.615 81.315 ;
        RECT 90.945 80.475 91.550 80.645 ;
        RECT 87.635 79.535 88.845 80.055 ;
        RECT 89.015 79.705 90.225 80.225 ;
        RECT 90.855 79.665 91.100 80.305 ;
        RECT 91.380 80.080 91.550 80.475 ;
        RECT 91.785 80.365 92.010 81.145 ;
        RECT 91.380 79.750 91.610 80.080 ;
        RECT 87.175 78.765 87.465 79.490 ;
        RECT 87.635 78.765 90.225 79.535 ;
        RECT 91.380 79.485 91.550 79.750 ;
        RECT 90.945 79.315 91.550 79.485 ;
        RECT 90.945 79.025 91.115 79.315 ;
        RECT 91.285 78.765 91.615 79.145 ;
        RECT 91.785 79.025 91.955 80.365 ;
        RECT 92.200 80.345 92.555 81.095 ;
        RECT 92.725 80.515 93.015 81.315 ;
        RECT 93.515 80.935 94.375 81.105 ;
        RECT 94.065 80.785 94.375 80.935 ;
        RECT 94.545 80.855 94.865 81.315 ;
        RECT 94.065 80.770 94.390 80.785 ;
        RECT 94.160 80.765 94.390 80.770 ;
        RECT 94.160 80.745 94.400 80.765 ;
        RECT 94.160 80.725 94.415 80.745 ;
        RECT 94.175 80.715 94.415 80.725 ;
        RECT 94.200 80.690 94.415 80.715 ;
        RECT 92.200 80.175 92.885 80.345 ;
        RECT 92.205 79.635 92.535 80.005 ;
        RECT 92.715 79.915 92.885 80.175 ;
        RECT 93.215 80.035 93.550 80.685 ;
        RECT 93.720 80.240 94.055 80.590 ;
        RECT 92.715 79.465 93.090 79.915 ;
        RECT 93.720 79.720 94.035 80.240 ;
        RECT 94.225 80.130 94.415 80.690 ;
        RECT 95.065 80.545 95.310 81.115 ;
        RECT 94.585 80.215 95.310 80.545 ;
        RECT 95.490 80.250 95.775 81.315 ;
        RECT 95.945 80.350 96.205 81.135 ;
        RECT 92.280 79.445 93.090 79.465 ;
        RECT 92.280 79.295 92.885 79.445 ;
        RECT 93.330 79.415 94.035 79.720 ;
        RECT 94.205 80.005 94.415 80.130 ;
        RECT 95.140 80.005 95.310 80.215 ;
        RECT 94.205 79.675 94.970 80.005 ;
        RECT 95.140 79.675 95.865 80.005 ;
        RECT 92.280 79.025 92.475 79.295 ;
        RECT 94.205 79.215 94.375 79.675 ;
        RECT 95.140 79.400 95.310 79.675 ;
        RECT 96.035 79.425 96.205 80.350 ;
        RECT 96.465 80.385 96.635 81.145 ;
        RECT 96.815 80.555 97.145 81.315 ;
        RECT 96.465 80.215 97.130 80.385 ;
        RECT 97.315 80.240 97.585 81.145 ;
        RECT 97.845 80.645 98.015 81.145 ;
        RECT 98.185 80.815 98.515 81.315 ;
        RECT 97.845 80.475 98.450 80.645 ;
        RECT 96.960 80.070 97.130 80.215 ;
        RECT 96.395 79.665 96.725 80.035 ;
        RECT 96.960 79.740 97.245 80.070 ;
        RECT 96.960 79.485 97.130 79.740 ;
        RECT 92.645 78.765 92.975 79.125 ;
        RECT 93.535 79.045 94.375 79.215 ;
        RECT 94.545 78.765 94.815 79.225 ;
        RECT 95.065 78.940 95.310 79.400 ;
        RECT 95.525 78.765 95.750 79.395 ;
        RECT 95.945 79.095 96.205 79.425 ;
        RECT 96.465 79.315 97.130 79.485 ;
        RECT 97.415 79.440 97.585 80.240 ;
        RECT 97.755 79.665 98.000 80.305 ;
        RECT 98.280 80.080 98.450 80.475 ;
        RECT 98.685 80.365 98.910 81.145 ;
        RECT 98.280 79.750 98.510 80.080 ;
        RECT 98.280 79.485 98.450 79.750 ;
        RECT 96.465 78.935 96.635 79.315 ;
        RECT 96.815 78.765 97.145 79.145 ;
        RECT 97.325 78.935 97.585 79.440 ;
        RECT 97.845 79.315 98.450 79.485 ;
        RECT 97.845 79.025 98.015 79.315 ;
        RECT 98.185 78.765 98.515 79.145 ;
        RECT 98.685 79.025 98.855 80.365 ;
        RECT 99.100 80.345 99.455 81.095 ;
        RECT 99.625 80.515 99.915 81.315 ;
        RECT 100.415 80.935 101.275 81.105 ;
        RECT 100.965 80.785 101.275 80.935 ;
        RECT 101.445 80.855 101.765 81.315 ;
        RECT 100.965 80.770 101.290 80.785 ;
        RECT 101.060 80.765 101.290 80.770 ;
        RECT 101.060 80.745 101.300 80.765 ;
        RECT 101.060 80.725 101.315 80.745 ;
        RECT 101.075 80.715 101.315 80.725 ;
        RECT 101.100 80.690 101.315 80.715 ;
        RECT 99.100 80.175 99.785 80.345 ;
        RECT 99.105 79.635 99.435 80.005 ;
        RECT 99.615 79.915 99.785 80.175 ;
        RECT 100.115 80.035 100.450 80.685 ;
        RECT 100.620 80.240 100.955 80.590 ;
        RECT 99.615 79.465 99.990 79.915 ;
        RECT 100.620 79.720 100.935 80.240 ;
        RECT 101.125 80.130 101.315 80.690 ;
        RECT 101.965 80.545 102.210 81.115 ;
        RECT 101.485 80.215 102.210 80.545 ;
        RECT 102.390 80.250 102.675 81.315 ;
        RECT 102.845 80.350 103.105 81.135 ;
        RECT 103.275 80.880 108.620 81.315 ;
        RECT 99.180 79.445 99.990 79.465 ;
        RECT 99.180 79.295 99.785 79.445 ;
        RECT 100.230 79.415 100.935 79.720 ;
        RECT 101.105 80.005 101.315 80.130 ;
        RECT 102.040 80.005 102.210 80.215 ;
        RECT 101.105 79.675 101.870 80.005 ;
        RECT 102.040 79.675 102.765 80.005 ;
        RECT 99.180 79.025 99.375 79.295 ;
        RECT 101.105 79.215 101.275 79.675 ;
        RECT 102.040 79.400 102.210 79.675 ;
        RECT 102.935 79.425 103.105 80.350 ;
        RECT 99.545 78.765 99.875 79.125 ;
        RECT 100.435 79.045 101.275 79.215 ;
        RECT 101.445 78.765 101.715 79.225 ;
        RECT 101.965 78.940 102.210 79.400 ;
        RECT 102.425 78.765 102.650 79.395 ;
        RECT 102.845 79.095 103.105 79.425 ;
        RECT 104.860 79.310 105.200 80.140 ;
        RECT 106.680 79.630 107.030 80.880 ;
        RECT 108.795 80.225 112.305 81.315 ;
        RECT 108.795 79.535 110.445 80.055 ;
        RECT 110.615 79.705 112.305 80.225 ;
        RECT 112.935 80.150 113.225 81.315 ;
        RECT 113.395 80.225 116.905 81.315 ;
        RECT 113.395 79.535 115.045 80.055 ;
        RECT 115.215 79.705 116.905 80.225 ;
        RECT 118.180 80.345 118.570 80.520 ;
        RECT 119.055 80.515 119.385 81.315 ;
        RECT 119.555 80.525 120.090 81.145 ;
        RECT 118.180 80.175 119.605 80.345 ;
        RECT 103.275 78.765 108.620 79.310 ;
        RECT 108.795 78.765 112.305 79.535 ;
        RECT 112.935 78.765 113.225 79.490 ;
        RECT 113.395 78.765 116.905 79.535 ;
        RECT 118.055 79.445 118.410 80.005 ;
        RECT 118.580 79.275 118.750 80.175 ;
        RECT 118.920 79.445 119.185 80.005 ;
        RECT 119.435 79.675 119.605 80.175 ;
        RECT 119.775 79.505 120.090 80.525 ;
        RECT 118.160 78.765 118.400 79.275 ;
        RECT 118.580 78.945 118.860 79.275 ;
        RECT 119.090 78.765 119.305 79.275 ;
        RECT 119.475 78.935 120.090 79.505 ;
        RECT 120.330 80.525 120.865 81.145 ;
        RECT 120.330 79.505 120.645 80.525 ;
        RECT 121.035 80.515 121.365 81.315 ;
        RECT 121.850 80.345 122.240 80.520 ;
        RECT 120.815 80.175 122.240 80.345 ;
        RECT 122.605 80.345 122.935 81.130 ;
        RECT 122.605 80.175 123.285 80.345 ;
        RECT 123.465 80.175 123.795 81.315 ;
        RECT 123.985 80.175 124.315 81.315 ;
        RECT 124.845 80.345 125.175 81.130 ;
        RECT 125.905 80.695 126.075 81.125 ;
        RECT 126.245 80.865 126.575 81.315 ;
        RECT 125.905 80.465 126.580 80.695 ;
        RECT 124.495 80.175 125.175 80.345 ;
        RECT 120.815 79.675 120.985 80.175 ;
        RECT 120.330 78.935 120.945 79.505 ;
        RECT 121.235 79.445 121.500 80.005 ;
        RECT 121.670 79.275 121.840 80.175 ;
        RECT 122.010 79.445 122.365 80.005 ;
        RECT 122.595 79.755 122.945 80.005 ;
        RECT 123.115 79.575 123.285 80.175 ;
        RECT 123.455 79.755 123.805 80.005 ;
        RECT 123.975 79.755 124.325 80.005 ;
        RECT 124.495 79.575 124.665 80.175 ;
        RECT 124.835 79.755 125.185 80.005 ;
        RECT 121.115 78.765 121.330 79.275 ;
        RECT 121.560 78.945 121.840 79.275 ;
        RECT 122.020 78.765 122.260 79.275 ;
        RECT 122.615 78.765 122.855 79.575 ;
        RECT 123.025 78.935 123.355 79.575 ;
        RECT 123.525 78.765 123.795 79.575 ;
        RECT 123.985 78.765 124.255 79.575 ;
        RECT 124.425 78.935 124.755 79.575 ;
        RECT 124.925 78.765 125.165 79.575 ;
        RECT 125.875 79.445 126.175 80.295 ;
        RECT 126.345 79.815 126.580 80.465 ;
        RECT 126.750 80.155 127.035 81.100 ;
        RECT 127.215 80.845 127.900 81.315 ;
        RECT 127.210 80.325 127.905 80.635 ;
        RECT 128.080 80.260 128.385 81.045 ;
        RECT 128.775 80.645 129.055 81.315 ;
        RECT 129.225 80.425 129.525 80.975 ;
        RECT 129.725 80.595 130.055 81.315 ;
        RECT 130.245 80.595 130.705 81.145 ;
        RECT 126.750 80.005 127.610 80.155 ;
        RECT 128.175 80.125 128.385 80.260 ;
        RECT 126.750 79.985 128.035 80.005 ;
        RECT 126.345 79.485 126.880 79.815 ;
        RECT 127.050 79.625 128.035 79.985 ;
        RECT 126.345 79.335 126.565 79.485 ;
        RECT 125.820 78.765 126.155 79.270 ;
        RECT 126.325 78.960 126.565 79.335 ;
        RECT 127.050 79.290 127.220 79.625 ;
        RECT 128.210 79.455 128.385 80.125 ;
        RECT 128.590 80.005 128.855 80.365 ;
        RECT 129.225 80.255 130.165 80.425 ;
        RECT 129.995 80.005 130.165 80.255 ;
        RECT 128.590 79.755 129.265 80.005 ;
        RECT 129.485 79.755 129.825 80.005 ;
        RECT 129.995 79.675 130.285 80.005 ;
        RECT 129.995 79.585 130.165 79.675 ;
        RECT 126.845 79.095 127.220 79.290 ;
        RECT 126.845 78.950 127.015 79.095 ;
        RECT 127.580 78.765 127.975 79.260 ;
        RECT 128.145 78.935 128.385 79.455 ;
        RECT 128.775 79.395 130.165 79.585 ;
        RECT 128.775 79.035 129.105 79.395 ;
        RECT 130.455 79.225 130.705 80.595 ;
        RECT 130.915 80.175 131.145 81.315 ;
        RECT 131.315 80.165 131.645 81.145 ;
        RECT 131.815 80.175 132.025 81.315 ;
        RECT 132.255 80.225 133.465 81.315 ;
        RECT 133.635 80.805 134.825 81.095 ;
        RECT 130.895 79.755 131.225 80.005 ;
        RECT 129.725 78.765 129.975 79.225 ;
        RECT 130.145 78.935 130.705 79.225 ;
        RECT 130.915 78.765 131.145 79.585 ;
        RECT 131.395 79.565 131.645 80.165 ;
        RECT 131.315 78.935 131.645 79.565 ;
        RECT 131.815 78.765 132.025 79.585 ;
        RECT 132.255 79.515 132.775 80.055 ;
        RECT 132.945 79.685 133.465 80.225 ;
        RECT 133.655 80.465 134.825 80.635 ;
        RECT 134.995 80.515 135.275 81.315 ;
        RECT 133.655 80.175 133.980 80.465 ;
        RECT 134.655 80.345 134.825 80.465 ;
        RECT 134.150 80.005 134.345 80.295 ;
        RECT 134.655 80.175 135.315 80.345 ;
        RECT 135.485 80.175 135.760 81.145 ;
        RECT 135.935 80.225 138.525 81.315 ;
        RECT 135.145 80.005 135.315 80.175 ;
        RECT 133.635 79.675 133.980 80.005 ;
        RECT 134.150 79.675 134.975 80.005 ;
        RECT 135.145 79.675 135.420 80.005 ;
        RECT 132.255 78.765 133.465 79.515 ;
        RECT 135.145 79.505 135.315 79.675 ;
        RECT 133.650 79.335 135.315 79.505 ;
        RECT 135.590 79.440 135.760 80.175 ;
        RECT 133.650 78.985 133.905 79.335 ;
        RECT 134.075 78.765 134.405 79.165 ;
        RECT 134.575 78.985 134.745 79.335 ;
        RECT 134.915 78.765 135.295 79.165 ;
        RECT 135.485 79.095 135.760 79.440 ;
        RECT 135.935 79.535 137.145 80.055 ;
        RECT 137.315 79.705 138.525 80.225 ;
        RECT 138.695 80.150 138.985 81.315 ;
        RECT 139.155 80.225 140.365 81.315 ;
        RECT 135.935 78.765 138.525 79.535 ;
        RECT 139.155 79.515 139.675 80.055 ;
        RECT 139.845 79.685 140.365 80.225 ;
        RECT 140.535 79.595 141.055 81.145 ;
        RECT 141.225 80.590 141.555 81.315 ;
        RECT 142.845 80.505 143.140 81.315 ;
        RECT 138.695 78.765 138.985 79.490 ;
        RECT 139.155 78.765 140.365 79.515 ;
        RECT 140.715 78.765 141.055 79.425 ;
        RECT 141.225 78.935 141.745 80.420 ;
        RECT 143.320 80.005 143.565 81.145 ;
        RECT 143.740 80.505 144.000 81.315 ;
        RECT 144.600 81.310 150.875 81.315 ;
        RECT 144.180 80.005 144.430 81.140 ;
        RECT 144.600 80.515 144.860 81.310 ;
        RECT 145.030 80.415 145.290 81.140 ;
        RECT 145.460 80.585 145.720 81.310 ;
        RECT 145.890 80.415 146.150 81.140 ;
        RECT 146.320 80.585 146.580 81.310 ;
        RECT 146.750 80.415 147.010 81.140 ;
        RECT 147.180 80.585 147.440 81.310 ;
        RECT 147.610 80.415 147.870 81.140 ;
        RECT 148.040 80.585 148.285 81.310 ;
        RECT 148.455 80.415 148.715 81.140 ;
        RECT 148.900 80.585 149.145 81.310 ;
        RECT 149.315 80.415 149.575 81.140 ;
        RECT 149.760 80.585 150.005 81.310 ;
        RECT 150.175 80.415 150.435 81.140 ;
        RECT 150.620 80.585 150.875 81.310 ;
        RECT 145.030 80.400 150.435 80.415 ;
        RECT 151.045 80.400 151.335 81.140 ;
        RECT 151.505 80.570 151.775 81.315 ;
        RECT 152.035 80.805 153.225 81.095 ;
        RECT 152.055 80.465 153.225 80.635 ;
        RECT 153.395 80.515 153.675 81.315 ;
        RECT 145.030 80.175 151.775 80.400 ;
        RECT 152.055 80.175 152.380 80.465 ;
        RECT 153.055 80.345 153.225 80.465 ;
        RECT 142.835 79.445 143.150 80.005 ;
        RECT 143.320 79.755 150.440 80.005 ;
        RECT 142.835 78.765 143.140 79.275 ;
        RECT 143.320 78.945 143.570 79.755 ;
        RECT 143.740 78.765 144.000 79.290 ;
        RECT 144.180 78.945 144.430 79.755 ;
        RECT 150.610 79.585 151.775 80.175 ;
        RECT 152.550 80.005 152.745 80.295 ;
        RECT 153.055 80.175 153.715 80.345 ;
        RECT 153.885 80.175 154.160 81.145 ;
        RECT 154.335 80.225 155.545 81.315 ;
        RECT 153.545 80.005 153.715 80.175 ;
        RECT 152.035 79.675 152.380 80.005 ;
        RECT 152.550 79.675 153.375 80.005 ;
        RECT 153.545 79.675 153.820 80.005 ;
        RECT 145.030 79.415 151.775 79.585 ;
        RECT 153.545 79.505 153.715 79.675 ;
        RECT 144.600 78.765 144.860 79.325 ;
        RECT 145.030 78.960 145.290 79.415 ;
        RECT 145.460 78.765 145.720 79.245 ;
        RECT 145.890 78.960 146.150 79.415 ;
        RECT 146.320 78.765 146.580 79.245 ;
        RECT 146.750 78.960 147.010 79.415 ;
        RECT 147.180 78.765 147.425 79.245 ;
        RECT 147.595 78.960 147.870 79.415 ;
        RECT 148.040 78.765 148.285 79.245 ;
        RECT 148.455 78.960 148.715 79.415 ;
        RECT 148.895 78.765 149.145 79.245 ;
        RECT 149.315 78.960 149.575 79.415 ;
        RECT 149.755 78.765 150.005 79.245 ;
        RECT 150.175 78.960 150.435 79.415 ;
        RECT 150.615 78.765 150.875 79.245 ;
        RECT 151.045 78.960 151.305 79.415 ;
        RECT 152.050 79.335 153.715 79.505 ;
        RECT 153.990 79.440 154.160 80.175 ;
        RECT 151.475 78.765 151.775 79.245 ;
        RECT 152.050 78.985 152.305 79.335 ;
        RECT 152.475 78.765 152.805 79.165 ;
        RECT 152.975 78.985 153.145 79.335 ;
        RECT 153.315 78.765 153.695 79.165 ;
        RECT 153.885 79.095 154.160 79.440 ;
        RECT 154.335 79.515 154.855 80.055 ;
        RECT 155.025 79.685 155.545 80.225 ;
        RECT 155.715 80.225 156.925 81.315 ;
        RECT 155.715 79.685 156.235 80.225 ;
        RECT 156.405 79.515 156.925 80.055 ;
        RECT 154.335 78.765 155.545 79.515 ;
        RECT 155.715 78.765 156.925 79.515 ;
        RECT 22.690 78.595 157.010 78.765 ;
        RECT 22.775 77.845 23.985 78.595 ;
        RECT 22.775 77.305 23.295 77.845 ;
        RECT 24.155 77.825 25.825 78.595 ;
        RECT 26.085 78.045 26.255 78.335 ;
        RECT 26.425 78.215 26.755 78.595 ;
        RECT 26.085 77.875 26.690 78.045 ;
        RECT 23.465 77.135 23.985 77.675 ;
        RECT 24.155 77.305 24.905 77.825 ;
        RECT 25.075 77.135 25.825 77.655 ;
        RECT 22.775 76.045 23.985 77.135 ;
        RECT 24.155 76.045 25.825 77.135 ;
        RECT 25.995 77.055 26.240 77.695 ;
        RECT 26.520 77.610 26.690 77.875 ;
        RECT 26.520 77.280 26.750 77.610 ;
        RECT 26.520 76.885 26.690 77.280 ;
        RECT 26.085 76.715 26.690 76.885 ;
        RECT 26.925 76.995 27.095 78.335 ;
        RECT 27.420 78.065 27.615 78.335 ;
        RECT 27.785 78.235 28.115 78.595 ;
        RECT 28.675 78.145 29.515 78.315 ;
        RECT 27.420 77.915 28.025 78.065 ;
        RECT 27.420 77.895 28.230 77.915 ;
        RECT 27.345 77.355 27.675 77.725 ;
        RECT 27.855 77.445 28.230 77.895 ;
        RECT 28.470 77.640 29.175 77.945 ;
        RECT 27.855 77.185 28.025 77.445 ;
        RECT 27.340 77.015 28.025 77.185 ;
        RECT 26.085 76.215 26.255 76.715 ;
        RECT 26.425 76.045 26.755 76.545 ;
        RECT 26.925 76.215 27.150 76.995 ;
        RECT 27.340 76.265 27.695 77.015 ;
        RECT 27.865 76.045 28.155 76.845 ;
        RECT 28.355 76.675 28.690 77.325 ;
        RECT 28.860 77.120 29.175 77.640 ;
        RECT 29.345 77.685 29.515 78.145 ;
        RECT 29.685 78.135 29.955 78.595 ;
        RECT 30.205 77.960 30.450 78.420 ;
        RECT 30.665 77.965 30.890 78.595 ;
        RECT 30.280 77.685 30.450 77.960 ;
        RECT 31.085 77.935 31.345 78.265 ;
        RECT 29.345 77.355 30.110 77.685 ;
        RECT 30.280 77.355 31.005 77.685 ;
        RECT 29.345 77.230 29.555 77.355 ;
        RECT 28.860 76.770 29.195 77.120 ;
        RECT 29.365 76.670 29.555 77.230 ;
        RECT 30.280 77.145 30.450 77.355 ;
        RECT 29.725 76.815 30.450 77.145 ;
        RECT 29.340 76.645 29.555 76.670 ;
        RECT 29.315 76.635 29.555 76.645 ;
        RECT 29.300 76.615 29.555 76.635 ;
        RECT 29.300 76.595 29.540 76.615 ;
        RECT 29.300 76.590 29.530 76.595 ;
        RECT 29.205 76.575 29.530 76.590 ;
        RECT 29.205 76.425 29.515 76.575 ;
        RECT 28.655 76.255 29.515 76.425 ;
        RECT 29.685 76.045 30.005 76.505 ;
        RECT 30.205 76.245 30.450 76.815 ;
        RECT 30.630 76.045 30.915 77.110 ;
        RECT 31.175 77.010 31.345 77.935 ;
        RECT 31.515 77.825 33.185 78.595 ;
        RECT 33.850 77.855 34.465 78.425 ;
        RECT 34.635 78.085 34.850 78.595 ;
        RECT 35.080 78.085 35.360 78.415 ;
        RECT 35.540 78.085 35.780 78.595 ;
        RECT 31.515 77.305 32.265 77.825 ;
        RECT 32.435 77.135 33.185 77.655 ;
        RECT 31.085 76.225 31.345 77.010 ;
        RECT 31.515 76.045 33.185 77.135 ;
        RECT 33.850 76.835 34.165 77.855 ;
        RECT 34.335 77.185 34.505 77.685 ;
        RECT 34.755 77.355 35.020 77.915 ;
        RECT 35.190 77.185 35.360 78.085 ;
        RECT 35.530 77.355 35.885 77.915 ;
        RECT 36.125 77.785 36.395 78.595 ;
        RECT 36.565 77.785 36.895 78.425 ;
        RECT 37.065 77.785 37.305 78.595 ;
        RECT 37.515 77.785 37.755 78.595 ;
        RECT 37.925 77.785 38.255 78.425 ;
        RECT 38.425 77.785 38.695 78.595 ;
        RECT 38.875 77.825 40.545 78.595 ;
        RECT 40.720 78.090 41.055 78.595 ;
        RECT 41.225 78.025 41.465 78.400 ;
        RECT 41.745 78.265 41.915 78.410 ;
        RECT 41.745 78.070 42.120 78.265 ;
        RECT 42.480 78.100 42.875 78.595 ;
        RECT 36.115 77.355 36.465 77.605 ;
        RECT 36.635 77.185 36.805 77.785 ;
        RECT 36.975 77.355 37.325 77.605 ;
        RECT 37.495 77.355 37.845 77.605 ;
        RECT 38.015 77.185 38.185 77.785 ;
        RECT 38.355 77.355 38.705 77.605 ;
        RECT 38.875 77.305 39.625 77.825 ;
        RECT 34.335 77.015 35.760 77.185 ;
        RECT 33.850 76.215 34.385 76.835 ;
        RECT 34.555 76.045 34.885 76.845 ;
        RECT 35.370 76.840 35.760 77.015 ;
        RECT 36.125 76.045 36.455 77.185 ;
        RECT 36.635 77.015 37.315 77.185 ;
        RECT 36.985 76.230 37.315 77.015 ;
        RECT 37.505 77.015 38.185 77.185 ;
        RECT 37.505 76.230 37.835 77.015 ;
        RECT 38.365 76.045 38.695 77.185 ;
        RECT 39.795 77.135 40.545 77.655 ;
        RECT 38.875 76.045 40.545 77.135 ;
        RECT 40.775 77.065 41.075 77.915 ;
        RECT 41.245 77.875 41.465 78.025 ;
        RECT 41.245 77.545 41.780 77.875 ;
        RECT 41.950 77.735 42.120 78.070 ;
        RECT 43.045 77.905 43.285 78.425 ;
        RECT 41.245 76.895 41.480 77.545 ;
        RECT 41.950 77.375 42.935 77.735 ;
        RECT 40.805 76.665 41.480 76.895 ;
        RECT 41.650 77.355 42.935 77.375 ;
        RECT 41.650 77.205 42.510 77.355 ;
        RECT 43.110 77.235 43.285 77.905 ;
        RECT 43.675 77.965 44.005 78.325 ;
        RECT 44.625 78.135 44.875 78.595 ;
        RECT 45.045 78.135 45.605 78.425 ;
        RECT 43.675 77.775 45.065 77.965 ;
        RECT 44.895 77.685 45.065 77.775 ;
        RECT 40.805 76.235 40.975 76.665 ;
        RECT 41.145 76.045 41.475 76.495 ;
        RECT 41.650 76.260 41.935 77.205 ;
        RECT 43.075 77.100 43.285 77.235 ;
        RECT 42.110 76.725 42.805 77.035 ;
        RECT 42.115 76.045 42.800 76.515 ;
        RECT 42.980 76.315 43.285 77.100 ;
        RECT 43.490 77.355 44.165 77.605 ;
        RECT 44.385 77.355 44.725 77.605 ;
        RECT 44.895 77.355 45.185 77.685 ;
        RECT 43.490 76.995 43.755 77.355 ;
        RECT 44.895 77.105 45.065 77.355 ;
        RECT 44.125 76.935 45.065 77.105 ;
        RECT 43.675 76.045 43.955 76.715 ;
        RECT 44.125 76.385 44.425 76.935 ;
        RECT 45.355 76.765 45.605 78.135 ;
        RECT 45.865 78.045 46.035 78.425 ;
        RECT 46.215 78.215 46.545 78.595 ;
        RECT 45.865 77.875 46.530 78.045 ;
        RECT 46.725 77.920 46.985 78.425 ;
        RECT 45.795 77.325 46.135 77.695 ;
        RECT 46.360 77.620 46.530 77.875 ;
        RECT 46.360 77.290 46.635 77.620 ;
        RECT 46.360 77.145 46.530 77.290 ;
        RECT 44.625 76.045 44.955 76.765 ;
        RECT 45.145 76.215 45.605 76.765 ;
        RECT 45.855 76.975 46.530 77.145 ;
        RECT 46.805 77.120 46.985 77.920 ;
        RECT 47.155 77.845 48.365 78.595 ;
        RECT 48.535 77.870 48.825 78.595 ;
        RECT 49.000 77.920 49.275 78.265 ;
        RECT 49.465 78.195 49.845 78.595 ;
        RECT 50.015 78.025 50.185 78.375 ;
        RECT 50.355 78.195 50.685 78.595 ;
        RECT 50.855 78.025 51.110 78.375 ;
        RECT 47.155 77.305 47.675 77.845 ;
        RECT 47.845 77.135 48.365 77.675 ;
        RECT 45.855 76.215 46.035 76.975 ;
        RECT 46.215 76.045 46.545 76.805 ;
        RECT 46.715 76.215 46.985 77.120 ;
        RECT 47.155 76.045 48.365 77.135 ;
        RECT 48.535 76.045 48.825 77.210 ;
        RECT 49.000 77.185 49.170 77.920 ;
        RECT 49.445 77.855 51.110 78.025 ;
        RECT 49.445 77.685 49.615 77.855 ;
        RECT 51.295 77.825 54.805 78.595 ;
        RECT 55.615 77.935 55.955 78.595 ;
        RECT 49.340 77.355 49.615 77.685 ;
        RECT 49.785 77.355 50.610 77.685 ;
        RECT 50.780 77.355 51.125 77.685 ;
        RECT 49.445 77.185 49.615 77.355 ;
        RECT 49.000 76.215 49.275 77.185 ;
        RECT 49.445 77.015 50.105 77.185 ;
        RECT 50.415 77.065 50.610 77.355 ;
        RECT 51.295 77.305 52.945 77.825 ;
        RECT 49.935 76.895 50.105 77.015 ;
        RECT 50.780 76.895 51.105 77.185 ;
        RECT 53.115 77.135 54.805 77.655 ;
        RECT 49.485 76.045 49.765 76.845 ;
        RECT 49.935 76.725 51.105 76.895 ;
        RECT 49.935 76.265 51.125 76.555 ;
        RECT 51.295 76.045 54.805 77.135 ;
        RECT 55.435 76.215 55.955 77.765 ;
        RECT 56.125 76.940 56.645 78.425 ;
        RECT 57.285 77.785 57.555 78.595 ;
        RECT 57.725 77.785 58.055 78.425 ;
        RECT 58.225 77.785 58.465 78.595 ;
        RECT 58.855 77.965 59.185 78.325 ;
        RECT 59.805 78.135 60.055 78.595 ;
        RECT 60.225 78.135 60.785 78.425 ;
        RECT 61.015 78.230 61.185 78.255 ;
        RECT 57.275 77.355 57.625 77.605 ;
        RECT 57.795 77.185 57.965 77.785 ;
        RECT 58.855 77.775 60.245 77.965 ;
        RECT 60.075 77.685 60.245 77.775 ;
        RECT 58.135 77.355 58.485 77.605 ;
        RECT 58.670 77.355 59.345 77.605 ;
        RECT 59.565 77.355 59.905 77.605 ;
        RECT 60.075 77.355 60.365 77.685 ;
        RECT 56.125 76.045 56.455 76.770 ;
        RECT 57.285 76.045 57.615 77.185 ;
        RECT 57.795 77.015 58.475 77.185 ;
        RECT 58.145 76.230 58.475 77.015 ;
        RECT 58.670 76.995 58.935 77.355 ;
        RECT 60.075 77.105 60.245 77.355 ;
        RECT 59.305 76.935 60.245 77.105 ;
        RECT 58.855 76.045 59.135 76.715 ;
        RECT 59.305 76.385 59.605 76.935 ;
        RECT 60.535 76.765 60.785 78.135 ;
        RECT 59.805 76.045 60.135 76.765 ;
        RECT 60.325 76.215 60.785 76.765 ;
        RECT 60.955 77.855 61.315 78.230 ;
        RECT 61.580 77.855 61.750 78.595 ;
        RECT 62.030 78.025 62.200 78.230 ;
        RECT 62.030 77.855 62.570 78.025 ;
        RECT 60.955 77.200 61.210 77.855 ;
        RECT 61.380 77.355 61.730 77.685 ;
        RECT 61.900 77.355 62.230 77.685 ;
        RECT 60.955 76.215 61.295 77.200 ;
        RECT 61.465 76.815 61.730 77.355 ;
        RECT 62.400 77.155 62.570 77.855 ;
        RECT 61.945 76.985 62.570 77.155 ;
        RECT 62.740 77.225 62.910 78.425 ;
        RECT 63.140 77.945 63.470 78.425 ;
        RECT 63.640 78.125 63.810 78.595 ;
        RECT 63.980 77.945 64.310 78.410 ;
        RECT 64.635 78.215 65.525 78.385 ;
        RECT 63.140 77.775 64.310 77.945 ;
        RECT 64.635 77.660 65.185 78.045 ;
        RECT 63.080 77.395 63.650 77.605 ;
        RECT 63.820 77.395 64.465 77.605 ;
        RECT 65.355 77.490 65.525 78.215 ;
        RECT 64.635 77.420 65.525 77.490 ;
        RECT 65.695 77.890 65.915 78.375 ;
        RECT 66.085 78.055 66.335 78.595 ;
        RECT 66.505 77.945 66.765 78.425 ;
        RECT 65.695 77.465 66.025 77.890 ;
        RECT 64.635 77.395 65.530 77.420 ;
        RECT 64.635 77.380 65.540 77.395 ;
        RECT 64.635 77.365 65.545 77.380 ;
        RECT 64.635 77.360 65.555 77.365 ;
        RECT 64.635 77.350 65.560 77.360 ;
        RECT 64.635 77.340 65.565 77.350 ;
        RECT 64.635 77.335 65.575 77.340 ;
        RECT 64.635 77.325 65.585 77.335 ;
        RECT 64.635 77.320 65.595 77.325 ;
        RECT 62.740 76.815 63.445 77.225 ;
        RECT 61.465 76.645 63.445 76.815 ;
        RECT 61.465 76.045 61.875 76.475 ;
        RECT 62.620 76.045 62.950 76.465 ;
        RECT 63.120 76.215 63.445 76.645 ;
        RECT 63.920 76.045 64.250 77.145 ;
        RECT 64.635 76.870 64.895 77.320 ;
        RECT 65.260 77.315 65.595 77.320 ;
        RECT 65.260 77.310 65.610 77.315 ;
        RECT 65.260 77.300 65.625 77.310 ;
        RECT 65.260 77.295 65.650 77.300 ;
        RECT 66.195 77.295 66.425 77.690 ;
        RECT 65.260 77.290 66.425 77.295 ;
        RECT 65.290 77.255 66.425 77.290 ;
        RECT 65.325 77.230 66.425 77.255 ;
        RECT 65.355 77.200 66.425 77.230 ;
        RECT 65.375 77.170 66.425 77.200 ;
        RECT 65.395 77.140 66.425 77.170 ;
        RECT 65.465 77.130 66.425 77.140 ;
        RECT 65.490 77.120 66.425 77.130 ;
        RECT 65.510 77.105 66.425 77.120 ;
        RECT 65.530 77.090 66.425 77.105 ;
        RECT 65.535 77.080 66.320 77.090 ;
        RECT 65.550 77.045 66.320 77.080 ;
        RECT 65.065 76.725 65.395 76.970 ;
        RECT 65.565 76.795 66.320 77.045 ;
        RECT 66.595 76.915 66.765 77.945 ;
        RECT 67.025 78.045 67.195 78.425 ;
        RECT 67.375 78.215 67.705 78.595 ;
        RECT 67.025 77.875 67.690 78.045 ;
        RECT 67.885 77.920 68.145 78.425 ;
        RECT 66.955 77.325 67.285 77.695 ;
        RECT 67.520 77.620 67.690 77.875 ;
        RECT 67.520 77.290 67.805 77.620 ;
        RECT 67.520 77.145 67.690 77.290 ;
        RECT 65.065 76.700 65.250 76.725 ;
        RECT 64.635 76.600 65.250 76.700 ;
        RECT 64.635 76.045 65.240 76.600 ;
        RECT 65.415 76.215 65.895 76.555 ;
        RECT 66.065 76.045 66.320 76.590 ;
        RECT 66.490 76.215 66.765 76.915 ;
        RECT 67.025 76.975 67.690 77.145 ;
        RECT 67.975 77.120 68.145 77.920 ;
        RECT 67.025 76.215 67.195 76.975 ;
        RECT 67.375 76.045 67.705 76.805 ;
        RECT 67.875 76.215 68.145 77.120 ;
        RECT 68.775 77.935 69.035 78.265 ;
        RECT 69.230 77.965 69.455 78.595 ;
        RECT 69.670 77.960 69.915 78.420 ;
        RECT 70.165 78.135 70.435 78.595 ;
        RECT 70.605 78.145 71.445 78.315 ;
        RECT 72.005 78.235 72.335 78.595 ;
        RECT 68.775 77.010 68.945 77.935 ;
        RECT 69.670 77.685 69.840 77.960 ;
        RECT 70.605 77.685 70.775 78.145 ;
        RECT 72.505 78.065 72.700 78.335 ;
        RECT 69.115 77.355 69.840 77.685 ;
        RECT 70.010 77.355 70.775 77.685 ;
        RECT 69.670 77.145 69.840 77.355 ;
        RECT 70.565 77.230 70.775 77.355 ;
        RECT 70.945 77.640 71.650 77.945 ;
        RECT 72.095 77.915 72.700 78.065 ;
        RECT 71.890 77.895 72.700 77.915 ;
        RECT 68.775 76.225 69.035 77.010 ;
        RECT 69.205 76.045 69.490 77.110 ;
        RECT 69.670 76.815 70.395 77.145 ;
        RECT 69.670 76.245 69.915 76.815 ;
        RECT 70.565 76.670 70.755 77.230 ;
        RECT 70.945 77.120 71.260 77.640 ;
        RECT 71.890 77.445 72.265 77.895 ;
        RECT 70.925 76.770 71.260 77.120 ;
        RECT 71.430 76.675 71.765 77.325 ;
        RECT 72.095 77.185 72.265 77.445 ;
        RECT 72.445 77.355 72.775 77.725 ;
        RECT 72.095 77.015 72.780 77.185 ;
        RECT 70.565 76.645 70.780 76.670 ;
        RECT 70.565 76.635 70.805 76.645 ;
        RECT 70.565 76.615 70.820 76.635 ;
        RECT 70.580 76.595 70.820 76.615 ;
        RECT 70.590 76.590 70.820 76.595 ;
        RECT 70.590 76.575 70.915 76.590 ;
        RECT 70.115 76.045 70.435 76.505 ;
        RECT 70.605 76.425 70.915 76.575 ;
        RECT 70.605 76.255 71.465 76.425 ;
        RECT 71.965 76.045 72.255 76.845 ;
        RECT 72.425 76.265 72.780 77.015 ;
        RECT 73.025 76.995 73.195 78.335 ;
        RECT 73.365 78.215 73.695 78.595 ;
        RECT 73.865 78.045 74.035 78.335 ;
        RECT 73.430 77.875 74.035 78.045 ;
        RECT 73.430 77.610 73.600 77.875 ;
        RECT 74.295 77.870 74.585 78.595 ;
        RECT 74.790 77.855 75.405 78.425 ;
        RECT 75.575 78.085 75.790 78.595 ;
        RECT 76.020 78.085 76.300 78.415 ;
        RECT 76.480 78.085 76.720 78.595 ;
        RECT 73.370 77.280 73.600 77.610 ;
        RECT 72.970 76.215 73.195 76.995 ;
        RECT 73.430 76.885 73.600 77.280 ;
        RECT 73.880 77.055 74.125 77.695 ;
        RECT 73.430 76.715 74.035 76.885 ;
        RECT 73.365 76.045 73.695 76.545 ;
        RECT 73.865 76.215 74.035 76.715 ;
        RECT 74.295 76.045 74.585 77.210 ;
        RECT 74.790 76.835 75.105 77.855 ;
        RECT 75.275 77.185 75.445 77.685 ;
        RECT 75.695 77.355 75.960 77.915 ;
        RECT 76.130 77.185 76.300 78.085 ;
        RECT 76.470 77.355 76.825 77.915 ;
        RECT 77.550 77.855 78.165 78.425 ;
        RECT 78.335 78.085 78.550 78.595 ;
        RECT 78.780 78.085 79.060 78.415 ;
        RECT 79.240 78.085 79.480 78.595 ;
        RECT 75.275 77.015 76.700 77.185 ;
        RECT 74.790 76.215 75.325 76.835 ;
        RECT 75.495 76.045 75.825 76.845 ;
        RECT 76.310 76.840 76.700 77.015 ;
        RECT 77.550 76.835 77.865 77.855 ;
        RECT 78.035 77.185 78.205 77.685 ;
        RECT 78.455 77.355 78.720 77.915 ;
        RECT 78.890 77.185 79.060 78.085 ;
        RECT 79.230 77.355 79.585 77.915 ;
        RECT 79.825 77.785 80.095 78.595 ;
        RECT 80.265 77.785 80.595 78.425 ;
        RECT 80.765 77.785 81.005 78.595 ;
        RECT 81.215 77.785 81.455 78.595 ;
        RECT 81.625 77.785 81.955 78.425 ;
        RECT 82.125 77.785 82.395 78.595 ;
        RECT 83.500 78.090 83.835 78.595 ;
        RECT 84.005 78.025 84.245 78.400 ;
        RECT 84.525 78.265 84.695 78.410 ;
        RECT 84.525 78.070 84.900 78.265 ;
        RECT 85.260 78.100 85.655 78.595 ;
        RECT 79.815 77.355 80.165 77.605 ;
        RECT 80.335 77.185 80.505 77.785 ;
        RECT 80.675 77.355 81.025 77.605 ;
        RECT 81.195 77.355 81.545 77.605 ;
        RECT 81.715 77.185 81.885 77.785 ;
        RECT 82.055 77.355 82.405 77.605 ;
        RECT 78.035 77.015 79.460 77.185 ;
        RECT 77.550 76.215 78.085 76.835 ;
        RECT 78.255 76.045 78.585 76.845 ;
        RECT 79.070 76.840 79.460 77.015 ;
        RECT 79.825 76.045 80.155 77.185 ;
        RECT 80.335 77.015 81.015 77.185 ;
        RECT 80.685 76.230 81.015 77.015 ;
        RECT 81.205 77.015 81.885 77.185 ;
        RECT 81.205 76.230 81.535 77.015 ;
        RECT 82.065 76.045 82.395 77.185 ;
        RECT 83.555 77.065 83.855 77.915 ;
        RECT 84.025 77.875 84.245 78.025 ;
        RECT 84.025 77.545 84.560 77.875 ;
        RECT 84.730 77.735 84.900 78.070 ;
        RECT 85.825 77.905 86.065 78.425 ;
        RECT 84.025 76.895 84.260 77.545 ;
        RECT 84.730 77.375 85.715 77.735 ;
        RECT 83.585 76.665 84.260 76.895 ;
        RECT 84.430 77.355 85.715 77.375 ;
        RECT 84.430 77.205 85.290 77.355 ;
        RECT 85.890 77.235 86.065 77.905 ;
        RECT 86.455 77.965 86.785 78.325 ;
        RECT 87.405 78.135 87.655 78.595 ;
        RECT 87.825 78.135 88.385 78.425 ;
        RECT 86.455 77.775 87.845 77.965 ;
        RECT 87.675 77.685 87.845 77.775 ;
        RECT 83.585 76.235 83.755 76.665 ;
        RECT 83.925 76.045 84.255 76.495 ;
        RECT 84.430 76.260 84.715 77.205 ;
        RECT 85.855 77.100 86.065 77.235 ;
        RECT 84.890 76.725 85.585 77.035 ;
        RECT 84.895 76.045 85.580 76.515 ;
        RECT 85.760 76.315 86.065 77.100 ;
        RECT 86.270 77.355 86.945 77.605 ;
        RECT 87.165 77.355 87.505 77.605 ;
        RECT 87.675 77.355 87.965 77.685 ;
        RECT 86.270 76.995 86.535 77.355 ;
        RECT 87.675 77.105 87.845 77.355 ;
        RECT 86.905 76.935 87.845 77.105 ;
        RECT 86.455 76.045 86.735 76.715 ;
        RECT 86.905 76.385 87.205 76.935 ;
        RECT 88.135 76.765 88.385 78.135 ;
        RECT 88.645 78.045 88.815 78.425 ;
        RECT 88.995 78.215 89.325 78.595 ;
        RECT 88.645 77.875 89.310 78.045 ;
        RECT 89.505 77.920 89.765 78.425 ;
        RECT 88.575 77.325 88.915 77.695 ;
        RECT 89.140 77.620 89.310 77.875 ;
        RECT 89.140 77.290 89.415 77.620 ;
        RECT 89.140 77.145 89.310 77.290 ;
        RECT 87.405 76.045 87.735 76.765 ;
        RECT 87.925 76.215 88.385 76.765 ;
        RECT 88.635 76.975 89.310 77.145 ;
        RECT 89.585 77.120 89.765 77.920 ;
        RECT 90.945 78.045 91.115 78.425 ;
        RECT 91.295 78.215 91.625 78.595 ;
        RECT 90.945 77.875 91.610 78.045 ;
        RECT 91.805 77.920 92.065 78.425 ;
        RECT 90.875 77.325 91.205 77.695 ;
        RECT 91.440 77.620 91.610 77.875 ;
        RECT 91.440 77.290 91.725 77.620 ;
        RECT 91.440 77.145 91.610 77.290 ;
        RECT 88.635 76.215 88.815 76.975 ;
        RECT 88.995 76.045 89.325 76.805 ;
        RECT 89.495 76.215 89.765 77.120 ;
        RECT 90.945 76.975 91.610 77.145 ;
        RECT 91.895 77.120 92.065 77.920 ;
        RECT 92.235 77.845 93.445 78.595 ;
        RECT 93.630 78.025 93.885 78.375 ;
        RECT 94.055 78.195 94.385 78.595 ;
        RECT 94.555 78.025 94.725 78.375 ;
        RECT 94.895 78.195 95.275 78.595 ;
        RECT 93.630 77.855 95.295 78.025 ;
        RECT 95.465 77.920 95.740 78.265 ;
        RECT 92.235 77.305 92.755 77.845 ;
        RECT 95.125 77.685 95.295 77.855 ;
        RECT 92.925 77.135 93.445 77.675 ;
        RECT 93.615 77.355 93.960 77.685 ;
        RECT 94.130 77.355 94.955 77.685 ;
        RECT 95.125 77.355 95.400 77.685 ;
        RECT 90.945 76.215 91.115 76.975 ;
        RECT 91.295 76.045 91.625 76.805 ;
        RECT 91.795 76.215 92.065 77.120 ;
        RECT 92.235 76.045 93.445 77.135 ;
        RECT 93.635 76.895 93.960 77.185 ;
        RECT 94.130 77.065 94.325 77.355 ;
        RECT 95.125 77.185 95.295 77.355 ;
        RECT 95.570 77.185 95.740 77.920 ;
        RECT 95.915 77.825 98.505 78.595 ;
        RECT 95.915 77.305 97.125 77.825 ;
        RECT 94.635 77.015 95.295 77.185 ;
        RECT 94.635 76.895 94.805 77.015 ;
        RECT 93.635 76.725 94.805 76.895 ;
        RECT 93.615 76.265 94.805 76.555 ;
        RECT 94.975 76.045 95.255 76.845 ;
        RECT 95.465 76.215 95.740 77.185 ;
        RECT 97.295 77.135 98.505 77.655 ;
        RECT 95.915 76.045 98.505 77.135 ;
        RECT 98.675 76.940 99.195 78.425 ;
        RECT 99.365 77.935 99.705 78.595 ;
        RECT 100.055 77.870 100.345 78.595 ;
        RECT 101.525 78.045 101.695 78.335 ;
        RECT 101.865 78.215 102.195 78.595 ;
        RECT 101.525 77.875 102.130 78.045 ;
        RECT 98.865 76.045 99.195 76.770 ;
        RECT 99.365 76.215 99.885 77.765 ;
        RECT 100.055 76.045 100.345 77.210 ;
        RECT 101.435 77.055 101.680 77.695 ;
        RECT 101.960 77.610 102.130 77.875 ;
        RECT 101.960 77.280 102.190 77.610 ;
        RECT 101.960 76.885 102.130 77.280 ;
        RECT 101.525 76.715 102.130 76.885 ;
        RECT 102.365 76.995 102.535 78.335 ;
        RECT 102.860 78.065 103.055 78.335 ;
        RECT 103.225 78.235 103.555 78.595 ;
        RECT 104.115 78.145 104.955 78.315 ;
        RECT 102.860 77.915 103.465 78.065 ;
        RECT 102.860 77.895 103.670 77.915 ;
        RECT 102.785 77.355 103.115 77.725 ;
        RECT 103.295 77.445 103.670 77.895 ;
        RECT 103.910 77.640 104.615 77.945 ;
        RECT 103.295 77.185 103.465 77.445 ;
        RECT 102.780 77.015 103.465 77.185 ;
        RECT 101.525 76.215 101.695 76.715 ;
        RECT 101.865 76.045 102.195 76.545 ;
        RECT 102.365 76.215 102.590 76.995 ;
        RECT 102.780 76.265 103.135 77.015 ;
        RECT 103.305 76.045 103.595 76.845 ;
        RECT 103.795 76.675 104.130 77.325 ;
        RECT 104.300 77.120 104.615 77.640 ;
        RECT 104.785 77.685 104.955 78.145 ;
        RECT 105.125 78.135 105.395 78.595 ;
        RECT 105.645 77.960 105.890 78.420 ;
        RECT 106.105 77.965 106.330 78.595 ;
        RECT 105.720 77.685 105.890 77.960 ;
        RECT 106.525 77.935 106.785 78.265 ;
        RECT 104.785 77.355 105.550 77.685 ;
        RECT 105.720 77.355 106.445 77.685 ;
        RECT 104.785 77.230 104.995 77.355 ;
        RECT 104.300 76.770 104.635 77.120 ;
        RECT 104.805 76.670 104.995 77.230 ;
        RECT 105.720 77.145 105.890 77.355 ;
        RECT 105.165 76.815 105.890 77.145 ;
        RECT 104.780 76.645 104.995 76.670 ;
        RECT 104.755 76.635 104.995 76.645 ;
        RECT 104.740 76.615 104.995 76.635 ;
        RECT 104.740 76.595 104.980 76.615 ;
        RECT 104.740 76.590 104.970 76.595 ;
        RECT 104.645 76.575 104.970 76.590 ;
        RECT 104.645 76.425 104.955 76.575 ;
        RECT 104.095 76.255 104.955 76.425 ;
        RECT 105.125 76.045 105.445 76.505 ;
        RECT 105.645 76.245 105.890 76.815 ;
        RECT 106.070 76.045 106.355 77.110 ;
        RECT 106.615 77.010 106.785 77.935 ;
        RECT 107.570 77.945 107.900 78.410 ;
        RECT 108.070 78.125 108.240 78.595 ;
        RECT 108.410 77.945 108.740 78.425 ;
        RECT 107.570 77.775 108.740 77.945 ;
        RECT 107.415 77.395 108.060 77.605 ;
        RECT 108.230 77.395 108.800 77.605 ;
        RECT 108.970 77.225 109.140 78.425 ;
        RECT 109.680 78.025 109.850 78.230 ;
        RECT 106.525 76.225 106.785 77.010 ;
        RECT 107.630 76.045 107.960 77.145 ;
        RECT 108.435 76.815 109.140 77.225 ;
        RECT 109.310 77.855 109.850 78.025 ;
        RECT 110.130 77.855 110.300 78.595 ;
        RECT 110.695 78.230 110.865 78.255 ;
        RECT 110.565 77.855 110.925 78.230 ;
        RECT 111.145 77.940 111.475 78.375 ;
        RECT 111.645 77.985 111.815 78.595 ;
        RECT 109.310 77.155 109.480 77.855 ;
        RECT 109.650 77.355 109.980 77.685 ;
        RECT 110.150 77.355 110.500 77.685 ;
        RECT 109.310 76.985 109.935 77.155 ;
        RECT 110.150 76.815 110.415 77.355 ;
        RECT 110.670 77.200 110.925 77.855 ;
        RECT 108.435 76.645 110.415 76.815 ;
        RECT 108.435 76.215 108.760 76.645 ;
        RECT 108.930 76.045 109.260 76.465 ;
        RECT 110.005 76.045 110.415 76.475 ;
        RECT 110.585 76.215 110.925 77.200 ;
        RECT 111.095 77.855 111.475 77.940 ;
        RECT 111.985 77.855 112.315 78.380 ;
        RECT 112.575 78.065 112.785 78.595 ;
        RECT 113.060 78.145 113.845 78.315 ;
        RECT 114.015 78.145 114.420 78.315 ;
        RECT 111.095 77.815 111.320 77.855 ;
        RECT 111.095 77.235 111.265 77.815 ;
        RECT 111.985 77.685 112.185 77.855 ;
        RECT 113.060 77.685 113.230 78.145 ;
        RECT 111.435 77.355 112.185 77.685 ;
        RECT 112.355 77.355 113.230 77.685 ;
        RECT 111.095 77.185 111.310 77.235 ;
        RECT 111.095 77.105 111.485 77.185 ;
        RECT 111.155 76.260 111.485 77.105 ;
        RECT 111.995 77.150 112.185 77.355 ;
        RECT 111.655 76.045 111.825 77.055 ;
        RECT 111.995 76.775 112.890 77.150 ;
        RECT 111.995 76.215 112.335 76.775 ;
        RECT 112.565 76.045 112.880 76.545 ;
        RECT 113.060 76.515 113.230 77.355 ;
        RECT 113.400 77.645 113.865 77.975 ;
        RECT 114.250 77.915 114.420 78.145 ;
        RECT 114.600 78.095 114.970 78.595 ;
        RECT 115.290 78.145 115.965 78.315 ;
        RECT 116.160 78.145 116.495 78.315 ;
        RECT 113.400 76.685 113.720 77.645 ;
        RECT 114.250 77.615 115.080 77.915 ;
        RECT 113.890 76.715 114.080 77.435 ;
        RECT 114.250 76.545 114.420 77.615 ;
        RECT 114.880 77.585 115.080 77.615 ;
        RECT 114.590 77.365 114.760 77.435 ;
        RECT 115.290 77.365 115.460 78.145 ;
        RECT 116.325 78.005 116.495 78.145 ;
        RECT 116.665 78.135 116.915 78.595 ;
        RECT 114.590 77.195 115.460 77.365 ;
        RECT 115.630 77.725 116.155 77.945 ;
        RECT 116.325 77.875 116.550 78.005 ;
        RECT 114.590 77.105 115.100 77.195 ;
        RECT 113.060 76.345 113.945 76.515 ;
        RECT 114.170 76.215 114.420 76.545 ;
        RECT 114.590 76.045 114.760 76.845 ;
        RECT 114.930 76.490 115.100 77.105 ;
        RECT 115.630 77.025 115.800 77.725 ;
        RECT 115.270 76.660 115.800 77.025 ;
        RECT 115.970 76.960 116.210 77.555 ;
        RECT 116.380 76.770 116.550 77.875 ;
        RECT 116.720 77.015 117.000 77.965 ;
        RECT 116.245 76.640 116.550 76.770 ;
        RECT 114.930 76.320 116.035 76.490 ;
        RECT 116.245 76.215 116.495 76.640 ;
        RECT 116.665 76.045 116.930 76.505 ;
        RECT 117.170 76.215 117.355 78.335 ;
        RECT 117.525 78.215 117.855 78.595 ;
        RECT 118.025 78.045 118.195 78.335 ;
        RECT 117.530 77.875 118.195 78.045 ;
        RECT 117.530 76.885 117.760 77.875 ;
        RECT 119.415 77.775 119.645 78.595 ;
        RECT 119.815 77.795 120.145 78.425 ;
        RECT 117.930 77.055 118.280 77.705 ;
        RECT 119.395 77.355 119.725 77.605 ;
        RECT 119.895 77.195 120.145 77.795 ;
        RECT 120.315 77.775 120.525 78.595 ;
        RECT 120.755 77.825 124.265 78.595 ;
        RECT 124.435 77.845 125.645 78.595 ;
        RECT 125.815 77.870 126.105 78.595 ;
        RECT 126.275 78.215 127.165 78.385 ;
        RECT 120.755 77.305 122.405 77.825 ;
        RECT 117.530 76.715 118.195 76.885 ;
        RECT 117.525 76.045 117.855 76.545 ;
        RECT 118.025 76.215 118.195 76.715 ;
        RECT 119.415 76.045 119.645 77.185 ;
        RECT 119.815 76.215 120.145 77.195 ;
        RECT 120.315 76.045 120.525 77.185 ;
        RECT 122.575 77.135 124.265 77.655 ;
        RECT 124.435 77.305 124.955 77.845 ;
        RECT 125.125 77.135 125.645 77.675 ;
        RECT 126.275 77.660 126.825 78.045 ;
        RECT 126.995 77.490 127.165 78.215 ;
        RECT 126.275 77.420 127.165 77.490 ;
        RECT 127.335 77.890 127.555 78.375 ;
        RECT 127.725 78.055 127.975 78.595 ;
        RECT 128.145 77.945 128.405 78.425 ;
        RECT 127.335 77.465 127.665 77.890 ;
        RECT 126.275 77.395 127.170 77.420 ;
        RECT 126.275 77.380 127.180 77.395 ;
        RECT 126.275 77.365 127.185 77.380 ;
        RECT 126.275 77.360 127.195 77.365 ;
        RECT 126.275 77.350 127.200 77.360 ;
        RECT 126.275 77.340 127.205 77.350 ;
        RECT 126.275 77.335 127.215 77.340 ;
        RECT 126.275 77.325 127.225 77.335 ;
        RECT 126.275 77.320 127.235 77.325 ;
        RECT 120.755 76.045 124.265 77.135 ;
        RECT 124.435 76.045 125.645 77.135 ;
        RECT 125.815 76.045 126.105 77.210 ;
        RECT 126.275 76.870 126.535 77.320 ;
        RECT 126.900 77.315 127.235 77.320 ;
        RECT 126.900 77.310 127.250 77.315 ;
        RECT 126.900 77.300 127.265 77.310 ;
        RECT 126.900 77.295 127.290 77.300 ;
        RECT 127.835 77.295 128.065 77.690 ;
        RECT 126.900 77.290 128.065 77.295 ;
        RECT 126.930 77.255 128.065 77.290 ;
        RECT 126.965 77.230 128.065 77.255 ;
        RECT 126.995 77.200 128.065 77.230 ;
        RECT 127.015 77.170 128.065 77.200 ;
        RECT 127.035 77.140 128.065 77.170 ;
        RECT 127.105 77.130 128.065 77.140 ;
        RECT 127.130 77.120 128.065 77.130 ;
        RECT 127.150 77.105 128.065 77.120 ;
        RECT 127.170 77.090 128.065 77.105 ;
        RECT 127.175 77.080 127.960 77.090 ;
        RECT 127.190 77.045 127.960 77.080 ;
        RECT 126.705 76.725 127.035 76.970 ;
        RECT 127.205 76.795 127.960 77.045 ;
        RECT 128.235 76.915 128.405 77.945 ;
        RECT 128.575 77.845 129.785 78.595 ;
        RECT 130.045 78.045 130.215 78.425 ;
        RECT 130.395 78.215 130.725 78.595 ;
        RECT 130.045 77.875 130.710 78.045 ;
        RECT 130.905 77.920 131.165 78.425 ;
        RECT 128.575 77.305 129.095 77.845 ;
        RECT 129.265 77.135 129.785 77.675 ;
        RECT 129.975 77.325 130.315 77.695 ;
        RECT 130.540 77.620 130.710 77.875 ;
        RECT 130.540 77.290 130.815 77.620 ;
        RECT 130.540 77.145 130.710 77.290 ;
        RECT 126.705 76.700 126.890 76.725 ;
        RECT 126.275 76.600 126.890 76.700 ;
        RECT 126.275 76.045 126.880 76.600 ;
        RECT 127.055 76.215 127.535 76.555 ;
        RECT 127.705 76.045 127.960 76.590 ;
        RECT 128.130 76.215 128.405 76.915 ;
        RECT 128.575 76.045 129.785 77.135 ;
        RECT 130.035 76.975 130.710 77.145 ;
        RECT 130.985 77.120 131.165 77.920 ;
        RECT 131.425 78.045 131.595 78.425 ;
        RECT 131.775 78.215 132.105 78.595 ;
        RECT 131.425 77.875 132.090 78.045 ;
        RECT 132.285 77.920 132.545 78.425 ;
        RECT 131.355 77.325 131.685 77.695 ;
        RECT 131.920 77.620 132.090 77.875 ;
        RECT 131.920 77.290 132.205 77.620 ;
        RECT 131.920 77.145 132.090 77.290 ;
        RECT 130.035 76.215 130.215 76.975 ;
        RECT 130.395 76.045 130.725 76.805 ;
        RECT 130.895 76.215 131.165 77.120 ;
        RECT 131.425 76.975 132.090 77.145 ;
        RECT 132.375 77.120 132.545 77.920 ;
        RECT 132.715 77.825 134.385 78.595 ;
        RECT 135.025 78.095 135.355 78.595 ;
        RECT 135.555 78.025 135.725 78.375 ;
        RECT 135.925 78.195 136.255 78.595 ;
        RECT 136.425 78.025 136.595 78.375 ;
        RECT 136.765 78.195 137.145 78.595 ;
        RECT 132.715 77.305 133.465 77.825 ;
        RECT 133.635 77.135 134.385 77.655 ;
        RECT 135.020 77.355 135.370 77.925 ;
        RECT 135.555 77.855 137.165 78.025 ;
        RECT 137.335 77.920 137.605 78.265 ;
        RECT 136.995 77.685 137.165 77.855 ;
        RECT 135.540 77.235 136.250 77.685 ;
        RECT 136.420 77.355 136.825 77.685 ;
        RECT 136.995 77.355 137.265 77.685 ;
        RECT 131.425 76.215 131.595 76.975 ;
        RECT 131.775 76.045 132.105 76.805 ;
        RECT 132.275 76.215 132.545 77.120 ;
        RECT 132.715 76.045 134.385 77.135 ;
        RECT 135.020 76.895 135.340 77.185 ;
        RECT 135.535 77.065 136.250 77.235 ;
        RECT 136.995 77.185 137.165 77.355 ;
        RECT 137.435 77.185 137.605 77.920 ;
        RECT 138.785 78.045 138.955 78.425 ;
        RECT 139.135 78.215 139.465 78.595 ;
        RECT 138.785 77.875 139.450 78.045 ;
        RECT 139.645 77.920 139.905 78.425 ;
        RECT 138.715 77.325 139.045 77.695 ;
        RECT 139.280 77.620 139.450 77.875 ;
        RECT 136.440 77.015 137.165 77.185 ;
        RECT 136.440 76.895 136.610 77.015 ;
        RECT 135.020 76.725 136.610 76.895 ;
        RECT 135.020 76.265 136.675 76.555 ;
        RECT 136.845 76.045 137.125 76.845 ;
        RECT 137.335 76.215 137.605 77.185 ;
        RECT 139.280 77.290 139.565 77.620 ;
        RECT 139.280 77.145 139.450 77.290 ;
        RECT 138.785 76.975 139.450 77.145 ;
        RECT 139.735 77.120 139.905 77.920 ;
        RECT 140.165 78.045 140.335 78.335 ;
        RECT 140.505 78.215 140.835 78.595 ;
        RECT 140.165 77.875 140.770 78.045 ;
        RECT 138.785 76.215 138.955 76.975 ;
        RECT 139.135 76.045 139.465 76.805 ;
        RECT 139.635 76.215 139.905 77.120 ;
        RECT 140.075 77.055 140.320 77.695 ;
        RECT 140.600 77.610 140.770 77.875 ;
        RECT 140.600 77.280 140.830 77.610 ;
        RECT 140.600 76.885 140.770 77.280 ;
        RECT 140.165 76.715 140.770 76.885 ;
        RECT 141.005 76.995 141.175 78.335 ;
        RECT 141.500 78.065 141.695 78.335 ;
        RECT 141.865 78.235 142.195 78.595 ;
        RECT 142.755 78.145 143.595 78.315 ;
        RECT 141.500 77.915 142.105 78.065 ;
        RECT 141.500 77.895 142.310 77.915 ;
        RECT 141.425 77.355 141.755 77.725 ;
        RECT 141.935 77.445 142.310 77.895 ;
        RECT 142.550 77.640 143.255 77.945 ;
        RECT 141.935 77.185 142.105 77.445 ;
        RECT 141.420 77.015 142.105 77.185 ;
        RECT 140.165 76.215 140.335 76.715 ;
        RECT 140.505 76.045 140.835 76.545 ;
        RECT 141.005 76.215 141.230 76.995 ;
        RECT 141.420 76.265 141.775 77.015 ;
        RECT 141.945 76.045 142.235 76.845 ;
        RECT 142.435 76.675 142.770 77.325 ;
        RECT 142.940 77.120 143.255 77.640 ;
        RECT 143.425 77.685 143.595 78.145 ;
        RECT 143.765 78.135 144.035 78.595 ;
        RECT 144.285 77.960 144.530 78.420 ;
        RECT 144.745 77.965 144.970 78.595 ;
        RECT 144.360 77.685 144.530 77.960 ;
        RECT 145.165 77.935 145.425 78.265 ;
        RECT 143.425 77.355 144.190 77.685 ;
        RECT 144.360 77.355 145.085 77.685 ;
        RECT 143.425 77.230 143.635 77.355 ;
        RECT 142.940 76.770 143.275 77.120 ;
        RECT 143.445 76.670 143.635 77.230 ;
        RECT 144.360 77.145 144.530 77.355 ;
        RECT 143.805 76.815 144.530 77.145 ;
        RECT 143.420 76.645 143.635 76.670 ;
        RECT 143.395 76.635 143.635 76.645 ;
        RECT 143.380 76.615 143.635 76.635 ;
        RECT 143.380 76.595 143.620 76.615 ;
        RECT 143.380 76.590 143.610 76.595 ;
        RECT 143.285 76.575 143.610 76.590 ;
        RECT 143.285 76.425 143.595 76.575 ;
        RECT 142.735 76.255 143.595 76.425 ;
        RECT 143.765 76.045 144.085 76.505 ;
        RECT 144.285 76.245 144.530 76.815 ;
        RECT 144.710 76.045 144.995 77.110 ;
        RECT 145.255 77.010 145.425 77.935 ;
        RECT 145.600 78.065 145.890 78.415 ;
        RECT 146.085 78.235 146.415 78.595 ;
        RECT 146.585 78.065 146.815 78.370 ;
        RECT 145.600 77.895 146.815 78.065 ;
        RECT 147.005 77.915 147.175 78.290 ;
        RECT 147.590 77.945 147.920 78.410 ;
        RECT 148.090 78.125 148.260 78.595 ;
        RECT 148.430 77.945 148.760 78.425 ;
        RECT 147.005 77.745 147.205 77.915 ;
        RECT 147.590 77.775 148.760 77.945 ;
        RECT 147.005 77.725 147.175 77.745 ;
        RECT 145.660 77.575 145.920 77.685 ;
        RECT 145.655 77.405 145.920 77.575 ;
        RECT 145.660 77.355 145.920 77.405 ;
        RECT 146.100 77.355 146.485 77.685 ;
        RECT 146.655 77.555 147.175 77.725 ;
        RECT 145.165 76.225 145.425 77.010 ;
        RECT 145.600 76.045 145.920 77.185 ;
        RECT 146.100 76.305 146.295 77.355 ;
        RECT 146.655 77.175 146.825 77.555 ;
        RECT 147.435 77.395 148.080 77.605 ;
        RECT 148.250 77.395 148.820 77.605 ;
        RECT 146.475 76.895 146.825 77.175 ;
        RECT 147.015 77.025 147.260 77.385 ;
        RECT 148.990 77.225 149.160 78.425 ;
        RECT 149.700 78.025 149.870 78.230 ;
        RECT 146.475 76.215 146.805 76.895 ;
        RECT 147.005 76.045 147.260 76.845 ;
        RECT 147.650 76.045 147.980 77.145 ;
        RECT 148.455 76.815 149.160 77.225 ;
        RECT 149.330 77.855 149.870 78.025 ;
        RECT 150.150 77.855 150.320 78.595 ;
        RECT 150.715 78.230 150.885 78.255 ;
        RECT 150.585 77.855 150.945 78.230 ;
        RECT 151.575 77.870 151.865 78.595 ;
        RECT 152.035 78.215 152.925 78.385 ;
        RECT 149.330 77.155 149.500 77.855 ;
        RECT 149.670 77.355 150.000 77.685 ;
        RECT 150.170 77.355 150.520 77.685 ;
        RECT 149.330 76.985 149.955 77.155 ;
        RECT 150.170 76.815 150.435 77.355 ;
        RECT 150.690 77.200 150.945 77.855 ;
        RECT 152.035 77.660 152.585 78.045 ;
        RECT 152.755 77.490 152.925 78.215 ;
        RECT 152.035 77.420 152.925 77.490 ;
        RECT 153.095 77.890 153.315 78.375 ;
        RECT 153.485 78.055 153.735 78.595 ;
        RECT 153.905 77.945 154.165 78.425 ;
        RECT 153.095 77.465 153.425 77.890 ;
        RECT 152.035 77.395 152.930 77.420 ;
        RECT 152.035 77.380 152.940 77.395 ;
        RECT 152.035 77.365 152.945 77.380 ;
        RECT 152.035 77.360 152.955 77.365 ;
        RECT 152.035 77.350 152.960 77.360 ;
        RECT 152.035 77.340 152.965 77.350 ;
        RECT 152.035 77.335 152.975 77.340 ;
        RECT 152.035 77.325 152.985 77.335 ;
        RECT 152.035 77.320 152.995 77.325 ;
        RECT 148.455 76.645 150.435 76.815 ;
        RECT 148.455 76.215 148.780 76.645 ;
        RECT 148.950 76.045 149.280 76.465 ;
        RECT 150.025 76.045 150.435 76.475 ;
        RECT 150.605 76.215 150.945 77.200 ;
        RECT 151.575 76.045 151.865 77.210 ;
        RECT 152.035 76.870 152.295 77.320 ;
        RECT 152.660 77.315 152.995 77.320 ;
        RECT 152.660 77.310 153.010 77.315 ;
        RECT 152.660 77.300 153.025 77.310 ;
        RECT 152.660 77.295 153.050 77.300 ;
        RECT 153.595 77.295 153.825 77.690 ;
        RECT 152.660 77.290 153.825 77.295 ;
        RECT 152.690 77.255 153.825 77.290 ;
        RECT 152.725 77.230 153.825 77.255 ;
        RECT 152.755 77.200 153.825 77.230 ;
        RECT 152.775 77.170 153.825 77.200 ;
        RECT 152.795 77.140 153.825 77.170 ;
        RECT 152.865 77.130 153.825 77.140 ;
        RECT 152.890 77.120 153.825 77.130 ;
        RECT 152.910 77.105 153.825 77.120 ;
        RECT 152.930 77.090 153.825 77.105 ;
        RECT 152.935 77.080 153.720 77.090 ;
        RECT 152.950 77.045 153.720 77.080 ;
        RECT 152.465 76.725 152.795 76.970 ;
        RECT 152.965 76.795 153.720 77.045 ;
        RECT 153.995 76.915 154.165 77.945 ;
        RECT 152.465 76.700 152.650 76.725 ;
        RECT 152.035 76.600 152.650 76.700 ;
        RECT 152.035 76.045 152.640 76.600 ;
        RECT 152.815 76.215 153.295 76.555 ;
        RECT 153.465 76.045 153.720 76.590 ;
        RECT 153.890 76.215 154.165 76.915 ;
        RECT 154.335 77.920 154.595 78.425 ;
        RECT 154.775 78.215 155.105 78.595 ;
        RECT 155.285 78.045 155.455 78.425 ;
        RECT 154.335 77.120 154.505 77.920 ;
        RECT 154.790 77.875 155.455 78.045 ;
        RECT 154.790 77.620 154.960 77.875 ;
        RECT 155.715 77.845 156.925 78.595 ;
        RECT 154.675 77.290 154.960 77.620 ;
        RECT 155.195 77.325 155.525 77.695 ;
        RECT 154.790 77.145 154.960 77.290 ;
        RECT 154.335 76.215 154.605 77.120 ;
        RECT 154.790 76.975 155.455 77.145 ;
        RECT 154.775 76.045 155.105 76.805 ;
        RECT 155.285 76.215 155.455 76.975 ;
        RECT 155.715 77.135 156.235 77.675 ;
        RECT 156.405 77.305 156.925 77.845 ;
        RECT 155.715 76.045 156.925 77.135 ;
        RECT 22.690 75.875 157.010 76.045 ;
        RECT 22.775 74.785 23.985 75.875 ;
        RECT 24.155 75.440 29.500 75.875 ;
        RECT 22.775 74.075 23.295 74.615 ;
        RECT 23.465 74.245 23.985 74.785 ;
        RECT 22.775 73.325 23.985 74.075 ;
        RECT 25.740 73.870 26.080 74.700 ;
        RECT 27.560 74.190 27.910 75.440 ;
        RECT 30.175 74.735 30.405 75.875 ;
        RECT 30.575 74.725 30.905 75.705 ;
        RECT 31.075 74.735 31.285 75.875 ;
        RECT 32.010 75.085 32.545 75.705 ;
        RECT 30.155 74.315 30.485 74.565 ;
        RECT 24.155 73.325 29.500 73.870 ;
        RECT 30.175 73.325 30.405 74.145 ;
        RECT 30.655 74.125 30.905 74.725 ;
        RECT 30.575 73.495 30.905 74.125 ;
        RECT 31.075 73.325 31.285 74.145 ;
        RECT 32.010 74.065 32.325 75.085 ;
        RECT 32.715 75.075 33.045 75.875 ;
        RECT 33.530 74.905 33.920 75.080 ;
        RECT 32.495 74.735 33.920 74.905 ;
        RECT 34.275 74.785 35.485 75.875 ;
        RECT 32.495 74.235 32.665 74.735 ;
        RECT 32.010 73.495 32.625 74.065 ;
        RECT 32.915 74.005 33.180 74.565 ;
        RECT 33.350 73.835 33.520 74.735 ;
        RECT 33.690 74.005 34.045 74.565 ;
        RECT 34.275 74.075 34.795 74.615 ;
        RECT 34.965 74.245 35.485 74.785 ;
        RECT 35.655 74.710 35.945 75.875 ;
        RECT 36.205 75.255 36.375 75.685 ;
        RECT 36.545 75.425 36.875 75.875 ;
        RECT 36.205 75.025 36.880 75.255 ;
        RECT 32.795 73.325 33.010 73.835 ;
        RECT 33.240 73.505 33.520 73.835 ;
        RECT 33.700 73.325 33.940 73.835 ;
        RECT 34.275 73.325 35.485 74.075 ;
        RECT 35.655 73.325 35.945 74.050 ;
        RECT 36.175 74.005 36.475 74.855 ;
        RECT 36.645 74.375 36.880 75.025 ;
        RECT 37.050 74.715 37.335 75.660 ;
        RECT 37.515 75.405 38.200 75.875 ;
        RECT 37.510 74.885 38.205 75.195 ;
        RECT 38.380 74.820 38.685 75.605 ;
        RECT 37.050 74.565 37.910 74.715 ;
        RECT 38.475 74.685 38.685 74.820 ;
        RECT 37.050 74.545 38.335 74.565 ;
        RECT 36.645 74.045 37.180 74.375 ;
        RECT 37.350 74.185 38.335 74.545 ;
        RECT 36.645 73.895 36.865 74.045 ;
        RECT 36.120 73.325 36.455 73.830 ;
        RECT 36.625 73.520 36.865 73.895 ;
        RECT 37.350 73.850 37.520 74.185 ;
        RECT 38.510 74.015 38.685 74.685 ;
        RECT 37.145 73.655 37.520 73.850 ;
        RECT 37.145 73.510 37.315 73.655 ;
        RECT 37.880 73.325 38.275 73.820 ;
        RECT 38.445 73.495 38.685 74.015 ;
        RECT 38.875 75.155 39.335 75.705 ;
        RECT 39.525 75.155 39.855 75.875 ;
        RECT 38.875 73.785 39.125 75.155 ;
        RECT 40.055 74.985 40.355 75.535 ;
        RECT 40.525 75.205 40.805 75.875 ;
        RECT 41.175 75.320 41.780 75.875 ;
        RECT 41.955 75.365 42.435 75.705 ;
        RECT 42.605 75.330 42.860 75.875 ;
        RECT 41.175 75.220 41.790 75.320 ;
        RECT 41.605 75.195 41.790 75.220 ;
        RECT 39.415 74.815 40.355 74.985 ;
        RECT 39.415 74.565 39.585 74.815 ;
        RECT 40.725 74.565 40.990 74.925 ;
        RECT 39.295 74.235 39.585 74.565 ;
        RECT 39.755 74.315 40.095 74.565 ;
        RECT 40.315 74.315 40.990 74.565 ;
        RECT 41.175 74.600 41.435 75.050 ;
        RECT 41.605 74.950 41.935 75.195 ;
        RECT 42.105 74.875 42.860 75.125 ;
        RECT 43.030 75.005 43.305 75.705 ;
        RECT 42.090 74.840 42.860 74.875 ;
        RECT 42.075 74.830 42.860 74.840 ;
        RECT 42.070 74.815 42.965 74.830 ;
        RECT 42.050 74.800 42.965 74.815 ;
        RECT 42.030 74.790 42.965 74.800 ;
        RECT 42.005 74.780 42.965 74.790 ;
        RECT 41.935 74.750 42.965 74.780 ;
        RECT 41.915 74.720 42.965 74.750 ;
        RECT 41.895 74.690 42.965 74.720 ;
        RECT 41.865 74.665 42.965 74.690 ;
        RECT 41.830 74.630 42.965 74.665 ;
        RECT 41.800 74.625 42.965 74.630 ;
        RECT 41.800 74.620 42.190 74.625 ;
        RECT 41.800 74.610 42.165 74.620 ;
        RECT 41.800 74.605 42.150 74.610 ;
        RECT 41.800 74.600 42.135 74.605 ;
        RECT 41.175 74.595 42.135 74.600 ;
        RECT 41.175 74.585 42.125 74.595 ;
        RECT 41.175 74.580 42.115 74.585 ;
        RECT 41.175 74.570 42.105 74.580 ;
        RECT 41.175 74.560 42.100 74.570 ;
        RECT 41.175 74.555 42.095 74.560 ;
        RECT 41.175 74.540 42.085 74.555 ;
        RECT 41.175 74.525 42.080 74.540 ;
        RECT 41.175 74.500 42.070 74.525 ;
        RECT 41.175 74.430 42.065 74.500 ;
        RECT 39.415 74.145 39.585 74.235 ;
        RECT 39.415 73.955 40.805 74.145 ;
        RECT 38.875 73.495 39.435 73.785 ;
        RECT 39.605 73.325 39.855 73.785 ;
        RECT 40.475 73.595 40.805 73.955 ;
        RECT 41.175 73.875 41.725 74.260 ;
        RECT 41.895 73.705 42.065 74.430 ;
        RECT 41.175 73.535 42.065 73.705 ;
        RECT 42.235 74.030 42.565 74.455 ;
        RECT 42.735 74.230 42.965 74.625 ;
        RECT 42.235 73.545 42.455 74.030 ;
        RECT 43.135 73.975 43.305 75.005 ;
        RECT 43.975 74.735 44.205 75.875 ;
        RECT 44.375 74.725 44.705 75.705 ;
        RECT 44.875 74.735 45.085 75.875 ;
        RECT 45.405 74.945 45.575 75.705 ;
        RECT 45.755 75.115 46.085 75.875 ;
        RECT 45.405 74.775 46.070 74.945 ;
        RECT 46.255 74.800 46.525 75.705 ;
        RECT 43.955 74.315 44.285 74.565 ;
        RECT 42.625 73.325 42.875 73.865 ;
        RECT 43.045 73.495 43.305 73.975 ;
        RECT 43.975 73.325 44.205 74.145 ;
        RECT 44.455 74.125 44.705 74.725 ;
        RECT 45.900 74.630 46.070 74.775 ;
        RECT 45.335 74.225 45.665 74.595 ;
        RECT 45.900 74.300 46.185 74.630 ;
        RECT 44.375 73.495 44.705 74.125 ;
        RECT 44.875 73.325 45.085 74.145 ;
        RECT 45.900 74.045 46.070 74.300 ;
        RECT 45.405 73.875 46.070 74.045 ;
        RECT 46.355 74.000 46.525 74.800 ;
        RECT 46.715 74.985 46.975 75.695 ;
        RECT 47.145 75.165 47.475 75.875 ;
        RECT 47.645 74.985 47.875 75.695 ;
        RECT 46.715 74.745 47.875 74.985 ;
        RECT 48.055 74.965 48.325 75.695 ;
        RECT 48.505 75.145 48.845 75.875 ;
        RECT 48.055 74.745 48.825 74.965 ;
        RECT 46.705 74.235 47.005 74.565 ;
        RECT 47.185 74.255 47.710 74.565 ;
        RECT 47.890 74.255 48.355 74.565 ;
        RECT 45.405 73.495 45.575 73.875 ;
        RECT 45.755 73.325 46.085 73.705 ;
        RECT 46.265 73.495 46.525 74.000 ;
        RECT 46.715 73.325 47.005 74.055 ;
        RECT 47.185 73.615 47.415 74.255 ;
        RECT 48.535 74.075 48.825 74.745 ;
        RECT 47.595 73.875 48.825 74.075 ;
        RECT 47.595 73.505 47.905 73.875 ;
        RECT 48.085 73.325 48.755 73.695 ;
        RECT 49.015 73.505 49.275 75.695 ;
        RECT 50.380 75.365 52.035 75.655 ;
        RECT 50.380 75.025 51.970 75.195 ;
        RECT 52.205 75.075 52.485 75.875 ;
        RECT 50.380 74.735 50.700 75.025 ;
        RECT 51.800 74.905 51.970 75.025 ;
        RECT 50.895 74.685 51.610 74.855 ;
        RECT 51.800 74.735 52.525 74.905 ;
        RECT 52.695 74.735 52.965 75.705 ;
        RECT 53.685 74.945 53.855 75.705 ;
        RECT 54.035 75.115 54.365 75.875 ;
        RECT 53.685 74.775 54.350 74.945 ;
        RECT 54.535 74.800 54.805 75.705 ;
        RECT 55.065 75.205 55.235 75.705 ;
        RECT 55.405 75.375 55.735 75.875 ;
        RECT 55.065 75.035 55.670 75.205 ;
        RECT 50.380 73.995 50.730 74.565 ;
        RECT 50.900 74.235 51.610 74.685 ;
        RECT 52.355 74.565 52.525 74.735 ;
        RECT 51.780 74.235 52.185 74.565 ;
        RECT 52.355 74.235 52.625 74.565 ;
        RECT 52.355 74.065 52.525 74.235 ;
        RECT 50.915 73.895 52.525 74.065 ;
        RECT 52.795 74.000 52.965 74.735 ;
        RECT 54.180 74.630 54.350 74.775 ;
        RECT 53.615 74.225 53.945 74.595 ;
        RECT 54.180 74.300 54.465 74.630 ;
        RECT 54.180 74.045 54.350 74.300 ;
        RECT 50.385 73.325 50.715 73.825 ;
        RECT 50.915 73.545 51.085 73.895 ;
        RECT 51.285 73.325 51.615 73.725 ;
        RECT 51.785 73.545 51.955 73.895 ;
        RECT 52.125 73.325 52.505 73.725 ;
        RECT 52.695 73.655 52.965 74.000 ;
        RECT 53.685 73.875 54.350 74.045 ;
        RECT 54.635 74.000 54.805 74.800 ;
        RECT 54.975 74.225 55.220 74.865 ;
        RECT 55.500 74.640 55.670 75.035 ;
        RECT 55.905 74.925 56.130 75.705 ;
        RECT 55.500 74.310 55.730 74.640 ;
        RECT 55.500 74.045 55.670 74.310 ;
        RECT 53.685 73.495 53.855 73.875 ;
        RECT 54.035 73.325 54.365 73.705 ;
        RECT 54.545 73.495 54.805 74.000 ;
        RECT 55.065 73.875 55.670 74.045 ;
        RECT 55.065 73.585 55.235 73.875 ;
        RECT 55.405 73.325 55.735 73.705 ;
        RECT 55.905 73.585 56.075 74.925 ;
        RECT 56.320 74.905 56.675 75.655 ;
        RECT 56.845 75.075 57.135 75.875 ;
        RECT 57.635 75.495 58.495 75.665 ;
        RECT 58.185 75.345 58.495 75.495 ;
        RECT 58.665 75.415 58.985 75.875 ;
        RECT 58.185 75.330 58.510 75.345 ;
        RECT 58.280 75.325 58.510 75.330 ;
        RECT 58.280 75.305 58.520 75.325 ;
        RECT 58.280 75.285 58.535 75.305 ;
        RECT 58.295 75.275 58.535 75.285 ;
        RECT 58.320 75.250 58.535 75.275 ;
        RECT 56.320 74.735 57.005 74.905 ;
        RECT 56.325 74.195 56.655 74.565 ;
        RECT 56.835 74.475 57.005 74.735 ;
        RECT 57.335 74.595 57.670 75.245 ;
        RECT 57.840 74.800 58.175 75.150 ;
        RECT 56.835 74.025 57.210 74.475 ;
        RECT 57.840 74.280 58.155 74.800 ;
        RECT 58.345 74.690 58.535 75.250 ;
        RECT 59.185 75.105 59.430 75.675 ;
        RECT 58.705 74.775 59.430 75.105 ;
        RECT 59.610 74.810 59.895 75.875 ;
        RECT 60.065 74.910 60.325 75.695 ;
        RECT 56.400 74.005 57.210 74.025 ;
        RECT 56.400 73.855 57.005 74.005 ;
        RECT 57.450 73.975 58.155 74.280 ;
        RECT 58.325 74.565 58.535 74.690 ;
        RECT 59.260 74.565 59.430 74.775 ;
        RECT 58.325 74.235 59.090 74.565 ;
        RECT 59.260 74.235 59.985 74.565 ;
        RECT 56.400 73.585 56.595 73.855 ;
        RECT 58.325 73.775 58.495 74.235 ;
        RECT 59.260 73.960 59.430 74.235 ;
        RECT 60.155 73.985 60.325 74.910 ;
        RECT 61.415 74.710 61.705 75.875 ;
        RECT 62.795 75.365 63.985 75.655 ;
        RECT 62.815 75.025 63.985 75.195 ;
        RECT 64.155 75.075 64.435 75.875 ;
        RECT 62.815 74.735 63.140 75.025 ;
        RECT 63.815 74.905 63.985 75.025 ;
        RECT 63.310 74.565 63.505 74.855 ;
        RECT 63.815 74.735 64.475 74.905 ;
        RECT 64.645 74.735 64.920 75.705 ;
        RECT 65.615 74.815 65.945 75.660 ;
        RECT 66.115 74.865 66.285 75.875 ;
        RECT 66.455 75.145 66.795 75.705 ;
        RECT 67.025 75.375 67.340 75.875 ;
        RECT 67.520 75.405 68.405 75.575 ;
        RECT 64.305 74.565 64.475 74.735 ;
        RECT 62.795 74.235 63.140 74.565 ;
        RECT 63.310 74.235 64.135 74.565 ;
        RECT 64.305 74.235 64.580 74.565 ;
        RECT 64.305 74.065 64.475 74.235 ;
        RECT 56.765 73.325 57.095 73.685 ;
        RECT 57.655 73.605 58.495 73.775 ;
        RECT 58.665 73.325 58.935 73.785 ;
        RECT 59.185 73.500 59.430 73.960 ;
        RECT 59.645 73.325 59.870 73.955 ;
        RECT 60.065 73.655 60.325 73.985 ;
        RECT 61.415 73.325 61.705 74.050 ;
        RECT 62.810 73.895 64.475 74.065 ;
        RECT 64.750 74.000 64.920 74.735 ;
        RECT 62.810 73.545 63.065 73.895 ;
        RECT 63.235 73.325 63.565 73.725 ;
        RECT 63.735 73.545 63.905 73.895 ;
        RECT 64.075 73.325 64.455 73.725 ;
        RECT 64.645 73.655 64.920 74.000 ;
        RECT 65.555 74.735 65.945 74.815 ;
        RECT 66.455 74.770 67.350 75.145 ;
        RECT 65.555 74.685 65.770 74.735 ;
        RECT 65.555 74.105 65.725 74.685 ;
        RECT 66.455 74.565 66.645 74.770 ;
        RECT 67.520 74.565 67.690 75.405 ;
        RECT 68.630 75.375 68.880 75.705 ;
        RECT 65.895 74.235 66.645 74.565 ;
        RECT 66.815 74.235 67.690 74.565 ;
        RECT 65.555 74.065 65.780 74.105 ;
        RECT 66.445 74.065 66.645 74.235 ;
        RECT 65.555 73.980 65.935 74.065 ;
        RECT 65.605 73.545 65.935 73.980 ;
        RECT 66.105 73.325 66.275 73.935 ;
        RECT 66.445 73.540 66.775 74.065 ;
        RECT 67.035 73.325 67.245 73.855 ;
        RECT 67.520 73.775 67.690 74.235 ;
        RECT 67.860 74.275 68.180 75.235 ;
        RECT 68.350 74.485 68.540 75.205 ;
        RECT 68.710 74.305 68.880 75.375 ;
        RECT 69.050 75.075 69.220 75.875 ;
        RECT 69.390 75.430 70.495 75.600 ;
        RECT 69.390 74.815 69.560 75.430 ;
        RECT 70.705 75.280 70.955 75.705 ;
        RECT 71.125 75.415 71.390 75.875 ;
        RECT 69.730 74.895 70.260 75.260 ;
        RECT 70.705 75.150 71.010 75.280 ;
        RECT 69.050 74.725 69.560 74.815 ;
        RECT 69.050 74.555 69.920 74.725 ;
        RECT 69.050 74.485 69.220 74.555 ;
        RECT 69.340 74.305 69.540 74.335 ;
        RECT 67.860 73.945 68.325 74.275 ;
        RECT 68.710 74.005 69.540 74.305 ;
        RECT 68.710 73.775 68.880 74.005 ;
        RECT 67.520 73.605 68.305 73.775 ;
        RECT 68.475 73.605 68.880 73.775 ;
        RECT 69.060 73.325 69.430 73.825 ;
        RECT 69.750 73.775 69.920 74.555 ;
        RECT 70.090 74.195 70.260 74.895 ;
        RECT 70.430 74.365 70.670 74.960 ;
        RECT 70.090 73.975 70.615 74.195 ;
        RECT 70.840 74.045 71.010 75.150 ;
        RECT 70.785 73.915 71.010 74.045 ;
        RECT 71.180 73.955 71.460 74.905 ;
        RECT 70.785 73.775 70.955 73.915 ;
        RECT 69.750 73.605 70.425 73.775 ;
        RECT 70.620 73.605 70.955 73.775 ;
        RECT 71.125 73.325 71.375 73.785 ;
        RECT 71.630 73.585 71.815 75.705 ;
        RECT 71.985 75.375 72.315 75.875 ;
        RECT 72.485 75.205 72.655 75.705 ;
        RECT 71.990 75.035 72.655 75.205 ;
        RECT 71.990 74.045 72.220 75.035 ;
        RECT 72.390 74.215 72.740 74.865 ;
        RECT 72.955 74.735 73.185 75.875 ;
        RECT 73.355 74.725 73.685 75.705 ;
        RECT 73.855 74.735 74.065 75.875 ;
        RECT 74.295 74.785 77.805 75.875 ;
        RECT 72.935 74.315 73.265 74.565 ;
        RECT 71.990 73.875 72.655 74.045 ;
        RECT 71.985 73.325 72.315 73.705 ;
        RECT 72.485 73.585 72.655 73.875 ;
        RECT 72.955 73.325 73.185 74.145 ;
        RECT 73.435 74.125 73.685 74.725 ;
        RECT 73.355 73.495 73.685 74.125 ;
        RECT 73.855 73.325 74.065 74.145 ;
        RECT 74.295 74.095 75.945 74.615 ;
        RECT 76.115 74.265 77.805 74.785 ;
        RECT 78.445 74.735 78.775 75.875 ;
        RECT 79.305 74.905 79.635 75.690 ;
        RECT 78.955 74.735 79.635 74.905 ;
        RECT 79.815 74.785 83.325 75.875 ;
        RECT 84.415 75.320 85.020 75.875 ;
        RECT 85.195 75.365 85.675 75.705 ;
        RECT 85.845 75.330 86.100 75.875 ;
        RECT 84.415 75.220 85.030 75.320 ;
        RECT 84.845 75.195 85.030 75.220 ;
        RECT 78.435 74.315 78.785 74.565 ;
        RECT 78.955 74.135 79.125 74.735 ;
        RECT 79.295 74.315 79.645 74.565 ;
        RECT 74.295 73.325 77.805 74.095 ;
        RECT 78.445 73.325 78.715 74.135 ;
        RECT 78.885 73.495 79.215 74.135 ;
        RECT 79.385 73.325 79.625 74.135 ;
        RECT 79.815 74.095 81.465 74.615 ;
        RECT 81.635 74.265 83.325 74.785 ;
        RECT 84.415 74.600 84.675 75.050 ;
        RECT 84.845 74.950 85.175 75.195 ;
        RECT 85.345 74.875 86.100 75.125 ;
        RECT 86.270 75.005 86.545 75.705 ;
        RECT 85.330 74.840 86.100 74.875 ;
        RECT 85.315 74.830 86.100 74.840 ;
        RECT 85.310 74.815 86.205 74.830 ;
        RECT 85.290 74.800 86.205 74.815 ;
        RECT 85.270 74.790 86.205 74.800 ;
        RECT 85.245 74.780 86.205 74.790 ;
        RECT 85.175 74.750 86.205 74.780 ;
        RECT 85.155 74.720 86.205 74.750 ;
        RECT 85.135 74.690 86.205 74.720 ;
        RECT 85.105 74.665 86.205 74.690 ;
        RECT 85.070 74.630 86.205 74.665 ;
        RECT 85.040 74.625 86.205 74.630 ;
        RECT 85.040 74.620 85.430 74.625 ;
        RECT 85.040 74.610 85.405 74.620 ;
        RECT 85.040 74.605 85.390 74.610 ;
        RECT 85.040 74.600 85.375 74.605 ;
        RECT 84.415 74.595 85.375 74.600 ;
        RECT 84.415 74.585 85.365 74.595 ;
        RECT 84.415 74.580 85.355 74.585 ;
        RECT 84.415 74.570 85.345 74.580 ;
        RECT 84.415 74.560 85.340 74.570 ;
        RECT 84.415 74.555 85.335 74.560 ;
        RECT 84.415 74.540 85.325 74.555 ;
        RECT 84.415 74.525 85.320 74.540 ;
        RECT 84.415 74.500 85.310 74.525 ;
        RECT 84.415 74.430 85.305 74.500 ;
        RECT 79.815 73.325 83.325 74.095 ;
        RECT 84.415 73.875 84.965 74.260 ;
        RECT 85.135 73.705 85.305 74.430 ;
        RECT 84.415 73.535 85.305 73.705 ;
        RECT 85.475 74.030 85.805 74.455 ;
        RECT 85.975 74.230 86.205 74.625 ;
        RECT 85.475 74.005 85.725 74.030 ;
        RECT 85.475 73.545 85.695 74.005 ;
        RECT 86.375 73.975 86.545 75.005 ;
        RECT 87.175 74.710 87.465 75.875 ;
        RECT 87.675 74.735 87.905 75.875 ;
        RECT 88.075 74.725 88.405 75.705 ;
        RECT 88.575 74.735 88.785 75.875 ;
        RECT 89.565 74.945 89.735 75.705 ;
        RECT 89.915 75.115 90.245 75.875 ;
        RECT 89.565 74.775 90.230 74.945 ;
        RECT 90.415 74.800 90.685 75.705 ;
        RECT 90.855 75.440 96.200 75.875 ;
        RECT 87.655 74.315 87.985 74.565 ;
        RECT 85.865 73.325 86.115 73.865 ;
        RECT 86.285 73.495 86.545 73.975 ;
        RECT 87.175 73.325 87.465 74.050 ;
        RECT 87.675 73.325 87.905 74.145 ;
        RECT 88.155 74.125 88.405 74.725 ;
        RECT 90.060 74.630 90.230 74.775 ;
        RECT 89.495 74.225 89.825 74.595 ;
        RECT 90.060 74.300 90.345 74.630 ;
        RECT 88.075 73.495 88.405 74.125 ;
        RECT 88.575 73.325 88.785 74.145 ;
        RECT 90.060 74.045 90.230 74.300 ;
        RECT 89.565 73.875 90.230 74.045 ;
        RECT 90.515 74.000 90.685 74.800 ;
        RECT 89.565 73.495 89.735 73.875 ;
        RECT 89.915 73.325 90.245 73.705 ;
        RECT 90.425 73.495 90.685 74.000 ;
        RECT 92.440 73.870 92.780 74.700 ;
        RECT 94.260 74.190 94.610 75.440 ;
        RECT 96.465 74.945 96.635 75.705 ;
        RECT 96.815 75.115 97.145 75.875 ;
        RECT 96.465 74.775 97.130 74.945 ;
        RECT 97.315 74.800 97.585 75.705 ;
        RECT 96.960 74.630 97.130 74.775 ;
        RECT 96.395 74.225 96.725 74.595 ;
        RECT 96.960 74.300 97.245 74.630 ;
        RECT 96.960 74.045 97.130 74.300 ;
        RECT 96.465 73.875 97.130 74.045 ;
        RECT 97.415 74.000 97.585 74.800 ;
        RECT 97.845 74.945 98.015 75.705 ;
        RECT 98.195 75.115 98.525 75.875 ;
        RECT 97.845 74.775 98.510 74.945 ;
        RECT 98.695 74.800 98.965 75.705 ;
        RECT 99.325 75.150 99.655 75.875 ;
        RECT 98.340 74.630 98.510 74.775 ;
        RECT 97.775 74.225 98.105 74.595 ;
        RECT 98.340 74.300 98.625 74.630 ;
        RECT 98.340 74.045 98.510 74.300 ;
        RECT 90.855 73.325 96.200 73.870 ;
        RECT 96.465 73.495 96.635 73.875 ;
        RECT 96.815 73.325 97.145 73.705 ;
        RECT 97.325 73.495 97.585 74.000 ;
        RECT 97.845 73.875 98.510 74.045 ;
        RECT 98.795 74.000 98.965 74.800 ;
        RECT 97.845 73.495 98.015 73.875 ;
        RECT 98.195 73.325 98.525 73.705 ;
        RECT 98.705 73.495 98.965 74.000 ;
        RECT 99.135 73.495 99.655 74.980 ;
        RECT 99.825 74.155 100.345 75.705 ;
        RECT 100.605 75.205 100.775 75.705 ;
        RECT 100.945 75.375 101.275 75.875 ;
        RECT 100.605 75.035 101.210 75.205 ;
        RECT 100.515 74.225 100.760 74.865 ;
        RECT 101.040 74.640 101.210 75.035 ;
        RECT 101.445 74.925 101.670 75.705 ;
        RECT 101.040 74.310 101.270 74.640 ;
        RECT 101.040 74.045 101.210 74.310 ;
        RECT 99.825 73.325 100.165 73.985 ;
        RECT 100.605 73.875 101.210 74.045 ;
        RECT 100.605 73.585 100.775 73.875 ;
        RECT 100.945 73.325 101.275 73.705 ;
        RECT 101.445 73.585 101.615 74.925 ;
        RECT 101.860 74.905 102.215 75.655 ;
        RECT 102.385 75.075 102.675 75.875 ;
        RECT 103.175 75.495 104.035 75.665 ;
        RECT 103.725 75.345 104.035 75.495 ;
        RECT 104.205 75.415 104.525 75.875 ;
        RECT 103.725 75.330 104.050 75.345 ;
        RECT 103.820 75.325 104.050 75.330 ;
        RECT 103.820 75.305 104.060 75.325 ;
        RECT 103.820 75.285 104.075 75.305 ;
        RECT 103.835 75.275 104.075 75.285 ;
        RECT 103.860 75.250 104.075 75.275 ;
        RECT 101.860 74.735 102.545 74.905 ;
        RECT 101.865 74.195 102.195 74.565 ;
        RECT 102.375 74.475 102.545 74.735 ;
        RECT 102.875 74.595 103.210 75.245 ;
        RECT 103.380 74.800 103.715 75.150 ;
        RECT 102.375 74.025 102.750 74.475 ;
        RECT 103.380 74.280 103.695 74.800 ;
        RECT 103.885 74.690 104.075 75.250 ;
        RECT 104.725 75.105 104.970 75.675 ;
        RECT 104.245 74.775 104.970 75.105 ;
        RECT 105.150 74.810 105.435 75.875 ;
        RECT 105.605 74.910 105.865 75.695 ;
        RECT 101.940 74.005 102.750 74.025 ;
        RECT 101.940 73.855 102.545 74.005 ;
        RECT 102.990 73.975 103.695 74.280 ;
        RECT 103.865 74.565 104.075 74.690 ;
        RECT 104.800 74.565 104.970 74.775 ;
        RECT 103.865 74.235 104.630 74.565 ;
        RECT 104.800 74.235 105.525 74.565 ;
        RECT 101.940 73.585 102.135 73.855 ;
        RECT 103.865 73.775 104.035 74.235 ;
        RECT 104.800 73.960 104.970 74.235 ;
        RECT 105.695 73.985 105.865 74.910 ;
        RECT 106.505 74.735 106.835 75.875 ;
        RECT 107.365 74.905 107.695 75.690 ;
        RECT 108.075 75.205 108.355 75.875 ;
        RECT 108.525 74.985 108.825 75.535 ;
        RECT 109.025 75.155 109.355 75.875 ;
        RECT 109.545 75.155 110.005 75.705 ;
        RECT 110.175 75.365 111.365 75.655 ;
        RECT 107.015 74.735 107.695 74.905 ;
        RECT 106.495 74.315 106.845 74.565 ;
        RECT 107.015 74.135 107.185 74.735 ;
        RECT 107.890 74.565 108.155 74.925 ;
        RECT 108.525 74.815 109.465 74.985 ;
        RECT 109.295 74.565 109.465 74.815 ;
        RECT 107.355 74.315 107.705 74.565 ;
        RECT 107.890 74.315 108.565 74.565 ;
        RECT 108.785 74.315 109.125 74.565 ;
        RECT 109.295 74.235 109.585 74.565 ;
        RECT 109.295 74.145 109.465 74.235 ;
        RECT 102.305 73.325 102.635 73.685 ;
        RECT 103.195 73.605 104.035 73.775 ;
        RECT 104.205 73.325 104.475 73.785 ;
        RECT 104.725 73.500 104.970 73.960 ;
        RECT 105.185 73.325 105.410 73.955 ;
        RECT 105.605 73.655 105.865 73.985 ;
        RECT 106.505 73.325 106.775 74.135 ;
        RECT 106.945 73.495 107.275 74.135 ;
        RECT 107.445 73.325 107.685 74.135 ;
        RECT 108.075 73.955 109.465 74.145 ;
        RECT 108.075 73.595 108.405 73.955 ;
        RECT 109.755 73.785 110.005 75.155 ;
        RECT 110.195 75.025 111.365 75.195 ;
        RECT 111.535 75.075 111.815 75.875 ;
        RECT 110.195 74.735 110.520 75.025 ;
        RECT 111.195 74.905 111.365 75.025 ;
        RECT 110.690 74.565 110.885 74.855 ;
        RECT 111.195 74.735 111.855 74.905 ;
        RECT 112.025 74.735 112.300 75.705 ;
        RECT 111.685 74.565 111.855 74.735 ;
        RECT 110.175 74.235 110.520 74.565 ;
        RECT 110.690 74.235 111.515 74.565 ;
        RECT 111.685 74.235 111.960 74.565 ;
        RECT 111.685 74.065 111.855 74.235 ;
        RECT 109.025 73.325 109.275 73.785 ;
        RECT 109.445 73.495 110.005 73.785 ;
        RECT 110.190 73.895 111.855 74.065 ;
        RECT 112.130 74.000 112.300 74.735 ;
        RECT 112.935 74.710 113.225 75.875 ;
        RECT 113.395 75.320 114.000 75.875 ;
        RECT 114.175 75.365 114.655 75.705 ;
        RECT 114.825 75.330 115.080 75.875 ;
        RECT 113.395 75.220 114.010 75.320 ;
        RECT 113.825 75.195 114.010 75.220 ;
        RECT 113.395 74.600 113.655 75.050 ;
        RECT 113.825 74.950 114.155 75.195 ;
        RECT 114.325 74.875 115.080 75.125 ;
        RECT 115.250 75.005 115.525 75.705 ;
        RECT 114.310 74.840 115.080 74.875 ;
        RECT 114.295 74.830 115.080 74.840 ;
        RECT 114.290 74.815 115.185 74.830 ;
        RECT 114.270 74.800 115.185 74.815 ;
        RECT 114.250 74.790 115.185 74.800 ;
        RECT 114.225 74.780 115.185 74.790 ;
        RECT 114.155 74.750 115.185 74.780 ;
        RECT 114.135 74.720 115.185 74.750 ;
        RECT 114.115 74.690 115.185 74.720 ;
        RECT 114.085 74.665 115.185 74.690 ;
        RECT 114.050 74.630 115.185 74.665 ;
        RECT 114.020 74.625 115.185 74.630 ;
        RECT 114.020 74.620 114.410 74.625 ;
        RECT 114.020 74.610 114.385 74.620 ;
        RECT 114.020 74.605 114.370 74.610 ;
        RECT 114.020 74.600 114.355 74.605 ;
        RECT 113.395 74.595 114.355 74.600 ;
        RECT 113.395 74.585 114.345 74.595 ;
        RECT 113.395 74.580 114.335 74.585 ;
        RECT 113.395 74.570 114.325 74.580 ;
        RECT 113.395 74.560 114.320 74.570 ;
        RECT 113.395 74.555 114.315 74.560 ;
        RECT 113.395 74.540 114.305 74.555 ;
        RECT 113.395 74.525 114.300 74.540 ;
        RECT 113.395 74.500 114.290 74.525 ;
        RECT 113.395 74.430 114.285 74.500 ;
        RECT 110.190 73.545 110.445 73.895 ;
        RECT 110.615 73.325 110.945 73.725 ;
        RECT 111.115 73.545 111.285 73.895 ;
        RECT 111.455 73.325 111.835 73.725 ;
        RECT 112.025 73.655 112.300 74.000 ;
        RECT 112.935 73.325 113.225 74.050 ;
        RECT 113.395 73.875 113.945 74.260 ;
        RECT 114.115 73.705 114.285 74.430 ;
        RECT 113.395 73.535 114.285 73.705 ;
        RECT 114.455 74.030 114.785 74.455 ;
        RECT 114.955 74.230 115.185 74.625 ;
        RECT 114.455 73.545 114.675 74.030 ;
        RECT 115.355 73.975 115.525 75.005 ;
        RECT 115.785 74.945 115.955 75.705 ;
        RECT 116.135 75.115 116.465 75.875 ;
        RECT 115.785 74.775 116.450 74.945 ;
        RECT 116.635 74.800 116.905 75.705 ;
        RECT 116.280 74.630 116.450 74.775 ;
        RECT 115.715 74.225 116.045 74.595 ;
        RECT 116.280 74.300 116.565 74.630 ;
        RECT 116.280 74.045 116.450 74.300 ;
        RECT 114.845 73.325 115.095 73.865 ;
        RECT 115.265 73.495 115.525 73.975 ;
        RECT 115.785 73.875 116.450 74.045 ;
        RECT 116.735 74.000 116.905 74.800 ;
        RECT 117.075 74.785 118.285 75.875 ;
        RECT 115.785 73.495 115.955 73.875 ;
        RECT 116.135 73.325 116.465 73.705 ;
        RECT 116.645 73.495 116.905 74.000 ;
        RECT 117.075 74.075 117.595 74.615 ;
        RECT 117.765 74.245 118.285 74.785 ;
        RECT 118.465 74.735 118.795 75.875 ;
        RECT 119.325 74.905 119.655 75.690 ;
        RECT 120.385 75.255 120.555 75.685 ;
        RECT 120.725 75.425 121.055 75.875 ;
        RECT 120.385 75.025 121.060 75.255 ;
        RECT 118.975 74.735 119.655 74.905 ;
        RECT 118.455 74.315 118.805 74.565 ;
        RECT 118.975 74.135 119.145 74.735 ;
        RECT 119.315 74.315 119.665 74.565 ;
        RECT 117.075 73.325 118.285 74.075 ;
        RECT 118.465 73.325 118.735 74.135 ;
        RECT 118.905 73.495 119.235 74.135 ;
        RECT 119.405 73.325 119.645 74.135 ;
        RECT 120.355 74.005 120.655 74.855 ;
        RECT 120.825 74.375 121.060 75.025 ;
        RECT 121.230 74.715 121.515 75.660 ;
        RECT 121.695 75.405 122.380 75.875 ;
        RECT 121.690 74.885 122.385 75.195 ;
        RECT 122.560 74.820 122.865 75.605 ;
        RECT 121.230 74.565 122.090 74.715 ;
        RECT 122.655 74.685 122.865 74.820 ;
        RECT 121.230 74.545 122.515 74.565 ;
        RECT 120.825 74.045 121.360 74.375 ;
        RECT 121.530 74.185 122.515 74.545 ;
        RECT 120.825 73.895 121.045 74.045 ;
        RECT 120.300 73.325 120.635 73.830 ;
        RECT 120.805 73.520 121.045 73.895 ;
        RECT 121.530 73.850 121.700 74.185 ;
        RECT 122.690 74.015 122.865 74.685 ;
        RECT 121.325 73.655 121.700 73.850 ;
        RECT 121.325 73.510 121.495 73.655 ;
        RECT 122.060 73.325 122.455 73.820 ;
        RECT 122.625 73.495 122.865 74.015 ;
        RECT 123.055 75.155 123.515 75.705 ;
        RECT 123.705 75.155 124.035 75.875 ;
        RECT 123.055 73.785 123.305 75.155 ;
        RECT 124.235 74.985 124.535 75.535 ;
        RECT 124.705 75.205 124.985 75.875 ;
        RECT 125.855 75.415 126.070 75.875 ;
        RECT 126.240 75.245 126.570 75.705 ;
        RECT 123.595 74.815 124.535 74.985 ;
        RECT 125.400 75.075 126.570 75.245 ;
        RECT 126.740 75.075 126.990 75.875 ;
        RECT 123.595 74.565 123.765 74.815 ;
        RECT 124.905 74.565 125.170 74.925 ;
        RECT 123.475 74.235 123.765 74.565 ;
        RECT 123.935 74.315 124.275 74.565 ;
        RECT 124.495 74.315 125.170 74.565 ;
        RECT 123.595 74.145 123.765 74.235 ;
        RECT 123.595 73.955 124.985 74.145 ;
        RECT 123.055 73.495 123.615 73.785 ;
        RECT 123.785 73.325 124.035 73.785 ;
        RECT 124.655 73.595 124.985 73.955 ;
        RECT 125.400 73.785 125.770 75.075 ;
        RECT 127.200 74.905 127.480 75.065 ;
        RECT 126.145 74.735 127.480 74.905 ;
        RECT 127.665 74.905 127.995 75.690 ;
        RECT 127.665 74.735 128.345 74.905 ;
        RECT 128.525 74.735 128.855 75.875 ;
        RECT 129.055 74.985 129.315 75.695 ;
        RECT 129.485 75.165 129.815 75.875 ;
        RECT 129.985 74.985 130.215 75.695 ;
        RECT 129.055 74.745 130.215 74.985 ;
        RECT 130.395 74.965 130.665 75.695 ;
        RECT 130.845 75.145 131.185 75.875 ;
        RECT 130.395 74.745 131.165 74.965 ;
        RECT 126.145 74.565 126.315 74.735 ;
        RECT 125.940 74.315 126.315 74.565 ;
        RECT 126.485 74.315 126.960 74.555 ;
        RECT 127.130 74.315 127.480 74.555 ;
        RECT 127.655 74.315 128.005 74.565 ;
        RECT 126.145 74.145 126.315 74.315 ;
        RECT 126.145 73.975 127.480 74.145 ;
        RECT 128.175 74.135 128.345 74.735 ;
        RECT 128.515 74.315 128.865 74.565 ;
        RECT 129.045 74.235 129.345 74.565 ;
        RECT 129.525 74.255 130.050 74.565 ;
        RECT 130.230 74.255 130.695 74.565 ;
        RECT 125.400 73.495 126.150 73.785 ;
        RECT 126.660 73.325 126.990 73.785 ;
        RECT 127.210 73.765 127.480 73.975 ;
        RECT 127.675 73.325 127.915 74.135 ;
        RECT 128.085 73.495 128.415 74.135 ;
        RECT 128.585 73.325 128.855 74.135 ;
        RECT 129.055 73.325 129.345 74.055 ;
        RECT 129.525 73.615 129.755 74.255 ;
        RECT 130.875 74.075 131.165 74.745 ;
        RECT 129.935 73.875 131.165 74.075 ;
        RECT 129.935 73.505 130.245 73.875 ;
        RECT 130.425 73.325 131.095 73.695 ;
        RECT 131.355 73.505 131.615 75.695 ;
        RECT 132.275 74.985 132.535 75.695 ;
        RECT 132.705 75.165 133.035 75.875 ;
        RECT 133.205 74.985 133.435 75.695 ;
        RECT 132.275 74.745 133.435 74.985 ;
        RECT 133.615 74.965 133.885 75.695 ;
        RECT 134.065 75.145 134.405 75.875 ;
        RECT 133.615 74.745 134.385 74.965 ;
        RECT 132.265 74.235 132.565 74.565 ;
        RECT 132.745 74.255 133.270 74.565 ;
        RECT 133.450 74.255 133.915 74.565 ;
        RECT 132.275 73.325 132.565 74.055 ;
        RECT 132.745 73.615 132.975 74.255 ;
        RECT 134.095 74.075 134.385 74.745 ;
        RECT 133.155 73.875 134.385 74.075 ;
        RECT 133.155 73.505 133.465 73.875 ;
        RECT 133.645 73.325 134.315 73.695 ;
        RECT 134.575 73.505 134.835 75.695 ;
        RECT 135.020 75.365 136.675 75.655 ;
        RECT 135.020 75.025 136.610 75.195 ;
        RECT 136.845 75.075 137.125 75.875 ;
        RECT 135.020 74.735 135.340 75.025 ;
        RECT 136.440 74.905 136.610 75.025 ;
        RECT 135.535 74.685 136.250 74.855 ;
        RECT 136.440 74.735 137.165 74.905 ;
        RECT 137.335 74.735 137.605 75.705 ;
        RECT 135.020 73.995 135.370 74.565 ;
        RECT 135.540 74.235 136.250 74.685 ;
        RECT 136.995 74.565 137.165 74.735 ;
        RECT 136.420 74.235 136.825 74.565 ;
        RECT 136.995 74.235 137.265 74.565 ;
        RECT 136.995 74.065 137.165 74.235 ;
        RECT 135.555 73.895 137.165 74.065 ;
        RECT 137.435 74.000 137.605 74.735 ;
        RECT 138.695 74.710 138.985 75.875 ;
        RECT 139.705 75.205 139.875 75.705 ;
        RECT 140.045 75.375 140.375 75.875 ;
        RECT 139.705 75.035 140.310 75.205 ;
        RECT 139.615 74.225 139.860 74.865 ;
        RECT 140.140 74.640 140.310 75.035 ;
        RECT 140.545 74.925 140.770 75.705 ;
        RECT 140.140 74.310 140.370 74.640 ;
        RECT 135.025 73.325 135.355 73.825 ;
        RECT 135.555 73.545 135.725 73.895 ;
        RECT 135.925 73.325 136.255 73.725 ;
        RECT 136.425 73.545 136.595 73.895 ;
        RECT 136.765 73.325 137.145 73.725 ;
        RECT 137.335 73.655 137.605 74.000 ;
        RECT 138.695 73.325 138.985 74.050 ;
        RECT 140.140 74.045 140.310 74.310 ;
        RECT 139.705 73.875 140.310 74.045 ;
        RECT 139.705 73.585 139.875 73.875 ;
        RECT 140.045 73.325 140.375 73.705 ;
        RECT 140.545 73.585 140.715 74.925 ;
        RECT 140.960 74.905 141.315 75.655 ;
        RECT 141.485 75.075 141.775 75.875 ;
        RECT 142.275 75.495 143.135 75.665 ;
        RECT 142.825 75.345 143.135 75.495 ;
        RECT 143.305 75.415 143.625 75.875 ;
        RECT 142.825 75.330 143.150 75.345 ;
        RECT 142.920 75.325 143.150 75.330 ;
        RECT 142.920 75.305 143.160 75.325 ;
        RECT 142.920 75.285 143.175 75.305 ;
        RECT 142.935 75.275 143.175 75.285 ;
        RECT 142.960 75.250 143.175 75.275 ;
        RECT 140.960 74.735 141.645 74.905 ;
        RECT 140.965 74.195 141.295 74.565 ;
        RECT 141.475 74.475 141.645 74.735 ;
        RECT 141.975 74.595 142.310 75.245 ;
        RECT 142.480 74.800 142.815 75.150 ;
        RECT 141.475 74.025 141.850 74.475 ;
        RECT 142.480 74.280 142.795 74.800 ;
        RECT 142.985 74.690 143.175 75.250 ;
        RECT 143.825 75.105 144.070 75.675 ;
        RECT 143.345 74.775 144.070 75.105 ;
        RECT 144.250 74.810 144.535 75.875 ;
        RECT 144.705 74.910 144.965 75.695 ;
        RECT 145.335 75.205 145.615 75.875 ;
        RECT 145.785 74.985 146.085 75.535 ;
        RECT 146.285 75.155 146.615 75.875 ;
        RECT 146.805 75.155 147.265 75.705 ;
        RECT 141.040 74.005 141.850 74.025 ;
        RECT 141.040 73.855 141.645 74.005 ;
        RECT 142.090 73.975 142.795 74.280 ;
        RECT 142.965 74.565 143.175 74.690 ;
        RECT 143.900 74.565 144.070 74.775 ;
        RECT 142.965 74.235 143.730 74.565 ;
        RECT 143.900 74.235 144.625 74.565 ;
        RECT 141.040 73.585 141.235 73.855 ;
        RECT 142.965 73.775 143.135 74.235 ;
        RECT 143.900 73.960 144.070 74.235 ;
        RECT 144.795 73.985 144.965 74.910 ;
        RECT 145.150 74.565 145.415 74.925 ;
        RECT 145.785 74.815 146.725 74.985 ;
        RECT 146.555 74.565 146.725 74.815 ;
        RECT 145.150 74.315 145.825 74.565 ;
        RECT 146.045 74.315 146.385 74.565 ;
        RECT 146.555 74.235 146.845 74.565 ;
        RECT 146.555 74.145 146.725 74.235 ;
        RECT 141.405 73.325 141.735 73.685 ;
        RECT 142.295 73.605 143.135 73.775 ;
        RECT 143.305 73.325 143.575 73.785 ;
        RECT 143.825 73.500 144.070 73.960 ;
        RECT 144.285 73.325 144.510 73.955 ;
        RECT 144.705 73.655 144.965 73.985 ;
        RECT 145.335 73.955 146.725 74.145 ;
        RECT 145.335 73.595 145.665 73.955 ;
        RECT 147.015 73.785 147.265 75.155 ;
        RECT 148.415 74.815 148.745 75.660 ;
        RECT 148.915 74.865 149.085 75.875 ;
        RECT 149.255 75.145 149.595 75.705 ;
        RECT 149.825 75.375 150.140 75.875 ;
        RECT 150.320 75.405 151.205 75.575 ;
        RECT 148.355 74.735 148.745 74.815 ;
        RECT 149.255 74.770 150.150 75.145 ;
        RECT 148.355 74.685 148.570 74.735 ;
        RECT 148.355 74.105 148.525 74.685 ;
        RECT 149.255 74.565 149.445 74.770 ;
        RECT 150.320 74.565 150.490 75.405 ;
        RECT 151.430 75.375 151.680 75.705 ;
        RECT 148.695 74.235 149.445 74.565 ;
        RECT 149.615 74.235 150.490 74.565 ;
        RECT 148.355 74.065 148.580 74.105 ;
        RECT 149.245 74.065 149.445 74.235 ;
        RECT 148.355 73.980 148.735 74.065 ;
        RECT 146.285 73.325 146.535 73.785 ;
        RECT 146.705 73.495 147.265 73.785 ;
        RECT 148.405 73.545 148.735 73.980 ;
        RECT 148.905 73.325 149.075 73.935 ;
        RECT 149.245 73.540 149.575 74.065 ;
        RECT 149.835 73.325 150.045 73.855 ;
        RECT 150.320 73.775 150.490 74.235 ;
        RECT 150.660 74.275 150.980 75.235 ;
        RECT 151.150 74.485 151.340 75.205 ;
        RECT 151.510 74.305 151.680 75.375 ;
        RECT 151.850 75.075 152.020 75.875 ;
        RECT 152.190 75.430 153.295 75.600 ;
        RECT 152.190 74.815 152.360 75.430 ;
        RECT 153.505 75.280 153.755 75.705 ;
        RECT 153.925 75.415 154.190 75.875 ;
        RECT 152.530 74.895 153.060 75.260 ;
        RECT 153.505 75.150 153.810 75.280 ;
        RECT 151.850 74.725 152.360 74.815 ;
        RECT 151.850 74.555 152.720 74.725 ;
        RECT 151.850 74.485 152.020 74.555 ;
        RECT 152.140 74.305 152.340 74.335 ;
        RECT 150.660 73.945 151.125 74.275 ;
        RECT 151.510 74.005 152.340 74.305 ;
        RECT 151.510 73.775 151.680 74.005 ;
        RECT 150.320 73.605 151.105 73.775 ;
        RECT 151.275 73.605 151.680 73.775 ;
        RECT 151.860 73.325 152.230 73.825 ;
        RECT 152.550 73.775 152.720 74.555 ;
        RECT 152.890 74.195 153.060 74.895 ;
        RECT 153.230 74.365 153.470 74.960 ;
        RECT 152.890 73.975 153.415 74.195 ;
        RECT 153.640 74.045 153.810 75.150 ;
        RECT 153.585 73.915 153.810 74.045 ;
        RECT 153.980 73.955 154.260 74.905 ;
        RECT 153.585 73.775 153.755 73.915 ;
        RECT 152.550 73.605 153.225 73.775 ;
        RECT 153.420 73.605 153.755 73.775 ;
        RECT 153.925 73.325 154.175 73.785 ;
        RECT 154.430 73.585 154.615 75.705 ;
        RECT 154.785 75.375 155.115 75.875 ;
        RECT 155.285 75.205 155.455 75.705 ;
        RECT 154.790 75.035 155.455 75.205 ;
        RECT 154.790 74.045 155.020 75.035 ;
        RECT 155.190 74.215 155.540 74.865 ;
        RECT 155.715 74.785 156.925 75.875 ;
        RECT 155.715 74.245 156.235 74.785 ;
        RECT 156.405 74.075 156.925 74.615 ;
        RECT 154.790 73.875 155.455 74.045 ;
        RECT 154.785 73.325 155.115 73.705 ;
        RECT 155.285 73.585 155.455 73.875 ;
        RECT 155.715 73.325 156.925 74.075 ;
        RECT 22.690 73.155 157.010 73.325 ;
        RECT 22.775 72.405 23.985 73.155 ;
        RECT 24.155 72.610 29.500 73.155 ;
        RECT 22.775 71.865 23.295 72.405 ;
        RECT 23.465 71.695 23.985 72.235 ;
        RECT 25.740 71.780 26.080 72.610 ;
        RECT 29.675 72.385 33.185 73.155 ;
        RECT 33.355 72.405 34.565 73.155 ;
        RECT 22.775 70.605 23.985 71.695 ;
        RECT 27.560 71.040 27.910 72.290 ;
        RECT 29.675 71.865 31.325 72.385 ;
        RECT 31.495 71.695 33.185 72.215 ;
        RECT 33.355 71.865 33.875 72.405 ;
        RECT 34.755 72.345 34.995 73.155 ;
        RECT 35.165 72.345 35.495 72.985 ;
        RECT 35.665 72.345 35.935 73.155 ;
        RECT 36.580 72.505 36.850 72.715 ;
        RECT 37.070 72.695 37.400 73.155 ;
        RECT 37.910 72.695 38.660 72.985 ;
        RECT 34.045 71.695 34.565 72.235 ;
        RECT 34.735 71.915 35.085 72.165 ;
        RECT 35.255 71.745 35.425 72.345 ;
        RECT 36.580 72.335 37.915 72.505 ;
        RECT 37.745 72.165 37.915 72.335 ;
        RECT 35.595 71.915 35.945 72.165 ;
        RECT 36.580 71.925 36.930 72.165 ;
        RECT 37.100 71.925 37.575 72.165 ;
        RECT 37.745 71.915 38.120 72.165 ;
        RECT 37.745 71.745 37.915 71.915 ;
        RECT 24.155 70.605 29.500 71.040 ;
        RECT 29.675 70.605 33.185 71.695 ;
        RECT 33.355 70.605 34.565 71.695 ;
        RECT 34.745 71.575 35.425 71.745 ;
        RECT 34.745 70.790 35.075 71.575 ;
        RECT 35.605 70.605 35.935 71.745 ;
        RECT 36.580 71.575 37.915 71.745 ;
        RECT 36.580 71.415 36.860 71.575 ;
        RECT 38.290 71.405 38.660 72.695 ;
        RECT 38.875 72.405 40.085 73.155 ;
        RECT 38.875 71.865 39.395 72.405 ;
        RECT 40.255 72.355 40.565 73.155 ;
        RECT 40.770 72.355 41.465 72.985 ;
        RECT 39.565 71.695 40.085 72.235 ;
        RECT 40.265 71.915 40.600 72.185 ;
        RECT 40.770 71.755 40.940 72.355 ;
        RECT 41.645 72.345 41.915 73.155 ;
        RECT 42.085 72.345 42.415 72.985 ;
        RECT 42.585 72.345 42.825 73.155 ;
        RECT 43.490 72.585 43.745 72.935 ;
        RECT 43.915 72.755 44.245 73.155 ;
        RECT 44.415 72.585 44.585 72.935 ;
        RECT 44.755 72.755 45.135 73.155 ;
        RECT 43.490 72.415 45.155 72.585 ;
        RECT 45.325 72.480 45.600 72.825 ;
        RECT 41.110 71.915 41.445 72.165 ;
        RECT 41.635 71.915 41.985 72.165 ;
        RECT 37.070 70.605 37.320 71.405 ;
        RECT 37.490 71.235 38.660 71.405 ;
        RECT 37.490 70.775 37.820 71.235 ;
        RECT 37.990 70.605 38.205 71.065 ;
        RECT 38.875 70.605 40.085 71.695 ;
        RECT 40.255 70.605 40.535 71.745 ;
        RECT 40.705 70.775 41.035 71.755 ;
        RECT 42.155 71.745 42.325 72.345 ;
        RECT 44.985 72.245 45.155 72.415 ;
        RECT 42.495 71.915 42.845 72.165 ;
        RECT 43.475 71.915 43.820 72.245 ;
        RECT 43.990 71.915 44.815 72.245 ;
        RECT 44.985 71.915 45.260 72.245 ;
        RECT 41.205 70.605 41.465 71.745 ;
        RECT 41.645 70.605 41.975 71.745 ;
        RECT 42.155 71.575 42.835 71.745 ;
        RECT 42.505 70.790 42.835 71.575 ;
        RECT 43.495 71.455 43.820 71.745 ;
        RECT 43.990 71.625 44.185 71.915 ;
        RECT 44.985 71.745 45.155 71.915 ;
        RECT 45.430 71.745 45.600 72.480 ;
        RECT 45.795 72.425 46.085 73.155 ;
        RECT 45.785 71.915 46.085 72.245 ;
        RECT 46.265 72.225 46.495 72.865 ;
        RECT 46.675 72.605 46.985 72.975 ;
        RECT 47.165 72.785 47.835 73.155 ;
        RECT 46.675 72.405 47.905 72.605 ;
        RECT 46.265 71.915 46.790 72.225 ;
        RECT 46.970 71.915 47.435 72.225 ;
        RECT 44.495 71.575 45.155 71.745 ;
        RECT 44.495 71.455 44.665 71.575 ;
        RECT 43.495 71.285 44.665 71.455 ;
        RECT 43.475 70.825 44.665 71.115 ;
        RECT 44.835 70.605 45.115 71.405 ;
        RECT 45.325 70.775 45.600 71.745 ;
        RECT 47.615 71.735 47.905 72.405 ;
        RECT 45.795 71.495 46.955 71.735 ;
        RECT 45.795 70.785 46.055 71.495 ;
        RECT 46.225 70.605 46.555 71.315 ;
        RECT 46.725 70.785 46.955 71.495 ;
        RECT 47.135 71.515 47.905 71.735 ;
        RECT 47.135 70.785 47.405 71.515 ;
        RECT 47.585 70.605 47.925 71.335 ;
        RECT 48.095 70.785 48.355 72.975 ;
        RECT 48.535 72.430 48.825 73.155 ;
        RECT 48.995 72.405 50.205 73.155 ;
        RECT 50.385 72.655 50.715 73.155 ;
        RECT 50.915 72.585 51.085 72.935 ;
        RECT 51.285 72.755 51.615 73.155 ;
        RECT 51.785 72.585 51.955 72.935 ;
        RECT 52.125 72.755 52.505 73.155 ;
        RECT 48.995 71.865 49.515 72.405 ;
        RECT 48.535 70.605 48.825 71.770 ;
        RECT 49.685 71.695 50.205 72.235 ;
        RECT 50.380 71.915 50.730 72.485 ;
        RECT 50.915 72.415 52.525 72.585 ;
        RECT 52.695 72.480 52.965 72.825 ;
        RECT 52.355 72.245 52.525 72.415 ;
        RECT 50.900 71.795 51.610 72.245 ;
        RECT 51.780 71.915 52.185 72.245 ;
        RECT 52.355 71.915 52.625 72.245 ;
        RECT 48.995 70.605 50.205 71.695 ;
        RECT 50.380 71.455 50.700 71.745 ;
        RECT 50.895 71.625 51.610 71.795 ;
        RECT 52.355 71.745 52.525 71.915 ;
        RECT 52.795 71.745 52.965 72.480 ;
        RECT 53.150 72.585 53.405 72.935 ;
        RECT 53.575 72.755 53.905 73.155 ;
        RECT 54.075 72.585 54.245 72.935 ;
        RECT 54.415 72.755 54.795 73.155 ;
        RECT 53.150 72.415 54.815 72.585 ;
        RECT 54.985 72.480 55.260 72.825 ;
        RECT 54.645 72.245 54.815 72.415 ;
        RECT 53.135 71.915 53.480 72.245 ;
        RECT 53.650 71.915 54.475 72.245 ;
        RECT 54.645 71.915 54.920 72.245 ;
        RECT 51.800 71.575 52.525 71.745 ;
        RECT 51.800 71.455 51.970 71.575 ;
        RECT 50.380 71.285 51.970 71.455 ;
        RECT 50.380 70.825 52.035 71.115 ;
        RECT 52.205 70.605 52.485 71.405 ;
        RECT 52.695 70.775 52.965 71.745 ;
        RECT 53.155 71.455 53.480 71.745 ;
        RECT 53.650 71.625 53.845 71.915 ;
        RECT 54.645 71.745 54.815 71.915 ;
        RECT 55.090 71.745 55.260 72.480 ;
        RECT 55.525 72.605 55.695 72.985 ;
        RECT 55.875 72.775 56.205 73.155 ;
        RECT 55.525 72.435 56.190 72.605 ;
        RECT 56.385 72.480 56.645 72.985 ;
        RECT 57.455 72.495 57.795 73.155 ;
        RECT 55.455 71.885 55.785 72.255 ;
        RECT 56.020 72.180 56.190 72.435 ;
        RECT 54.155 71.575 54.815 71.745 ;
        RECT 54.155 71.455 54.325 71.575 ;
        RECT 53.155 71.285 54.325 71.455 ;
        RECT 53.135 70.825 54.325 71.115 ;
        RECT 54.495 70.605 54.775 71.405 ;
        RECT 54.985 70.775 55.260 71.745 ;
        RECT 56.020 71.850 56.305 72.180 ;
        RECT 56.020 71.705 56.190 71.850 ;
        RECT 55.525 71.535 56.190 71.705 ;
        RECT 56.475 71.680 56.645 72.480 ;
        RECT 55.525 70.775 55.695 71.535 ;
        RECT 55.875 70.605 56.205 71.365 ;
        RECT 56.375 70.775 56.645 71.680 ;
        RECT 57.275 70.775 57.795 72.325 ;
        RECT 57.965 71.500 58.485 72.985 ;
        RECT 58.655 72.385 62.165 73.155 ;
        RECT 63.420 72.645 63.660 73.155 ;
        RECT 63.840 72.645 64.120 72.975 ;
        RECT 64.350 72.645 64.565 73.155 ;
        RECT 58.655 71.865 60.305 72.385 ;
        RECT 60.475 71.695 62.165 72.215 ;
        RECT 63.315 71.915 63.670 72.475 ;
        RECT 63.840 71.745 64.010 72.645 ;
        RECT 64.180 71.915 64.445 72.475 ;
        RECT 64.735 72.415 65.350 72.985 ;
        RECT 64.695 71.745 64.865 72.245 ;
        RECT 57.965 70.605 58.295 71.330 ;
        RECT 58.655 70.605 62.165 71.695 ;
        RECT 63.440 71.575 64.865 71.745 ;
        RECT 63.440 71.400 63.830 71.575 ;
        RECT 64.315 70.605 64.645 71.405 ;
        RECT 65.035 71.395 65.350 72.415 ;
        RECT 65.555 72.355 66.250 72.985 ;
        RECT 66.455 72.355 66.765 73.155 ;
        RECT 66.935 72.610 72.280 73.155 ;
        RECT 65.575 71.915 65.910 72.165 ;
        RECT 66.080 71.755 66.250 72.355 ;
        RECT 66.420 71.915 66.755 72.185 ;
        RECT 68.520 71.780 68.860 72.610 ;
        RECT 72.925 72.345 73.195 73.155 ;
        RECT 73.365 72.345 73.695 72.985 ;
        RECT 73.865 72.345 74.105 73.155 ;
        RECT 74.295 72.430 74.585 73.155 ;
        RECT 74.755 72.405 75.965 73.155 ;
        RECT 76.180 72.695 76.930 72.985 ;
        RECT 77.440 72.695 77.770 73.155 ;
        RECT 64.815 70.775 65.350 71.395 ;
        RECT 65.555 70.605 65.815 71.745 ;
        RECT 65.985 70.775 66.315 71.755 ;
        RECT 66.485 70.605 66.765 71.745 ;
        RECT 70.340 71.040 70.690 72.290 ;
        RECT 72.915 71.915 73.265 72.165 ;
        RECT 73.435 71.745 73.605 72.345 ;
        RECT 73.775 71.915 74.125 72.165 ;
        RECT 74.755 71.865 75.275 72.405 ;
        RECT 66.935 70.605 72.280 71.040 ;
        RECT 72.925 70.605 73.255 71.745 ;
        RECT 73.435 71.575 74.115 71.745 ;
        RECT 73.785 70.790 74.115 71.575 ;
        RECT 74.295 70.605 74.585 71.770 ;
        RECT 75.445 71.695 75.965 72.235 ;
        RECT 74.755 70.605 75.965 71.695 ;
        RECT 76.180 71.405 76.550 72.695 ;
        RECT 77.990 72.505 78.260 72.715 ;
        RECT 78.440 72.650 78.775 73.155 ;
        RECT 78.945 72.585 79.185 72.960 ;
        RECT 79.465 72.825 79.635 72.970 ;
        RECT 79.465 72.630 79.840 72.825 ;
        RECT 80.200 72.660 80.595 73.155 ;
        RECT 76.925 72.335 78.260 72.505 ;
        RECT 76.925 72.165 77.095 72.335 ;
        RECT 76.720 71.915 77.095 72.165 ;
        RECT 77.265 71.925 77.740 72.165 ;
        RECT 77.910 71.925 78.260 72.165 ;
        RECT 76.925 71.745 77.095 71.915 ;
        RECT 76.925 71.575 78.260 71.745 ;
        RECT 78.495 71.625 78.795 72.475 ;
        RECT 78.965 72.435 79.185 72.585 ;
        RECT 78.965 72.105 79.500 72.435 ;
        RECT 79.670 72.295 79.840 72.630 ;
        RECT 80.765 72.465 81.005 72.985 ;
        RECT 77.980 71.415 78.260 71.575 ;
        RECT 78.965 71.455 79.200 72.105 ;
        RECT 79.670 71.935 80.655 72.295 ;
        RECT 76.180 71.235 77.350 71.405 ;
        RECT 76.635 70.605 76.850 71.065 ;
        RECT 77.020 70.775 77.350 71.235 ;
        RECT 77.520 70.605 77.770 71.405 ;
        RECT 78.525 71.225 79.200 71.455 ;
        RECT 79.370 71.915 80.655 71.935 ;
        RECT 79.370 71.765 80.230 71.915 ;
        RECT 80.830 71.795 81.005 72.465 ;
        RECT 78.525 70.795 78.695 71.225 ;
        RECT 78.865 70.605 79.195 71.055 ;
        RECT 79.370 70.820 79.655 71.765 ;
        RECT 80.795 71.660 81.005 71.795 ;
        RECT 79.830 71.285 80.525 71.595 ;
        RECT 79.835 70.605 80.520 71.075 ;
        RECT 80.700 70.875 81.005 71.660 ;
        RECT 81.195 72.695 81.755 72.985 ;
        RECT 81.925 72.695 82.175 73.155 ;
        RECT 81.195 71.325 81.445 72.695 ;
        RECT 82.795 72.525 83.125 72.885 ;
        RECT 81.735 72.335 83.125 72.525 ;
        RECT 84.435 72.345 84.675 73.155 ;
        RECT 84.845 72.345 85.175 72.985 ;
        RECT 85.345 72.345 85.615 73.155 ;
        RECT 85.795 72.355 86.105 73.155 ;
        RECT 86.310 72.355 87.005 72.985 ;
        RECT 87.655 72.425 87.945 73.155 ;
        RECT 81.735 72.245 81.905 72.335 ;
        RECT 81.615 71.915 81.905 72.245 ;
        RECT 82.075 71.915 82.415 72.165 ;
        RECT 82.635 71.915 83.310 72.165 ;
        RECT 84.415 71.915 84.765 72.165 ;
        RECT 81.735 71.665 81.905 71.915 ;
        RECT 81.735 71.495 82.675 71.665 ;
        RECT 83.045 71.555 83.310 71.915 ;
        RECT 84.935 71.745 85.105 72.345 ;
        RECT 86.310 72.305 86.485 72.355 ;
        RECT 85.275 71.915 85.625 72.165 ;
        RECT 85.805 71.915 86.140 72.185 ;
        RECT 86.310 71.755 86.480 72.305 ;
        RECT 86.650 71.915 86.985 72.165 ;
        RECT 87.645 71.915 87.945 72.245 ;
        RECT 88.125 72.225 88.355 72.865 ;
        RECT 88.535 72.605 88.845 72.975 ;
        RECT 89.025 72.785 89.695 73.155 ;
        RECT 88.535 72.405 89.765 72.605 ;
        RECT 88.125 71.915 88.650 72.225 ;
        RECT 88.830 71.915 89.295 72.225 ;
        RECT 84.425 71.575 85.105 71.745 ;
        RECT 81.195 70.775 81.655 71.325 ;
        RECT 81.845 70.605 82.175 71.325 ;
        RECT 82.375 70.945 82.675 71.495 ;
        RECT 82.845 70.605 83.125 71.275 ;
        RECT 84.425 70.790 84.755 71.575 ;
        RECT 85.285 70.605 85.615 71.745 ;
        RECT 85.795 70.605 86.075 71.745 ;
        RECT 86.245 70.775 86.575 71.755 ;
        RECT 86.745 70.605 87.005 71.745 ;
        RECT 89.475 71.735 89.765 72.405 ;
        RECT 87.655 71.495 88.815 71.735 ;
        RECT 87.655 70.785 87.915 71.495 ;
        RECT 88.085 70.605 88.415 71.315 ;
        RECT 88.585 70.785 88.815 71.495 ;
        RECT 88.995 71.515 89.765 71.735 ;
        RECT 88.995 70.785 89.265 71.515 ;
        RECT 89.445 70.605 89.785 71.335 ;
        RECT 89.955 70.785 90.215 72.975 ;
        RECT 90.395 72.385 92.065 73.155 ;
        RECT 92.255 72.425 92.545 73.155 ;
        RECT 90.395 71.865 91.145 72.385 ;
        RECT 91.315 71.695 92.065 72.215 ;
        RECT 92.245 71.915 92.545 72.245 ;
        RECT 92.725 72.225 92.955 72.865 ;
        RECT 93.135 72.605 93.445 72.975 ;
        RECT 93.625 72.785 94.295 73.155 ;
        RECT 93.135 72.405 94.365 72.605 ;
        RECT 92.725 71.915 93.250 72.225 ;
        RECT 93.430 71.915 93.895 72.225 ;
        RECT 94.075 71.735 94.365 72.405 ;
        RECT 90.395 70.605 92.065 71.695 ;
        RECT 92.255 71.495 93.415 71.735 ;
        RECT 92.255 70.785 92.515 71.495 ;
        RECT 92.685 70.605 93.015 71.315 ;
        RECT 93.185 70.785 93.415 71.495 ;
        RECT 93.595 71.515 94.365 71.735 ;
        RECT 93.595 70.785 93.865 71.515 ;
        RECT 94.045 70.605 94.385 71.335 ;
        RECT 94.555 70.785 94.815 72.975 ;
        RECT 95.005 72.655 95.335 73.155 ;
        RECT 95.535 72.585 95.705 72.935 ;
        RECT 95.905 72.755 96.235 73.155 ;
        RECT 96.405 72.585 96.575 72.935 ;
        RECT 96.745 72.755 97.125 73.155 ;
        RECT 95.000 71.915 95.350 72.485 ;
        RECT 95.535 72.415 97.145 72.585 ;
        RECT 97.315 72.480 97.585 72.825 ;
        RECT 97.920 72.645 98.160 73.155 ;
        RECT 98.340 72.645 98.620 72.975 ;
        RECT 98.850 72.645 99.065 73.155 ;
        RECT 96.975 72.245 97.145 72.415 ;
        RECT 95.520 71.795 96.230 72.245 ;
        RECT 96.400 71.915 96.805 72.245 ;
        RECT 96.975 71.915 97.245 72.245 ;
        RECT 95.000 71.455 95.320 71.745 ;
        RECT 95.515 71.625 96.230 71.795 ;
        RECT 96.975 71.745 97.145 71.915 ;
        RECT 97.415 71.745 97.585 72.480 ;
        RECT 97.815 71.915 98.170 72.475 ;
        RECT 98.340 71.745 98.510 72.645 ;
        RECT 98.680 71.915 98.945 72.475 ;
        RECT 99.235 72.415 99.850 72.985 ;
        RECT 100.055 72.430 100.345 73.155 ;
        RECT 100.530 72.585 100.785 72.935 ;
        RECT 100.955 72.755 101.285 73.155 ;
        RECT 101.455 72.585 101.625 72.935 ;
        RECT 101.795 72.755 102.175 73.155 ;
        RECT 100.530 72.415 102.195 72.585 ;
        RECT 102.365 72.480 102.640 72.825 ;
        RECT 102.815 72.610 108.160 73.155 ;
        RECT 108.800 72.625 109.090 72.975 ;
        RECT 109.285 72.795 109.615 73.155 ;
        RECT 109.785 72.625 110.015 72.930 ;
        RECT 99.195 71.745 99.365 72.245 ;
        RECT 96.420 71.575 97.145 71.745 ;
        RECT 96.420 71.455 96.590 71.575 ;
        RECT 95.000 71.285 96.590 71.455 ;
        RECT 95.000 70.825 96.655 71.115 ;
        RECT 96.825 70.605 97.105 71.405 ;
        RECT 97.315 70.775 97.585 71.745 ;
        RECT 97.940 71.575 99.365 71.745 ;
        RECT 97.940 71.400 98.330 71.575 ;
        RECT 98.815 70.605 99.145 71.405 ;
        RECT 99.535 71.395 99.850 72.415 ;
        RECT 102.025 72.245 102.195 72.415 ;
        RECT 100.515 71.915 100.860 72.245 ;
        RECT 101.030 71.915 101.855 72.245 ;
        RECT 102.025 71.915 102.300 72.245 ;
        RECT 99.315 70.775 99.850 71.395 ;
        RECT 100.055 70.605 100.345 71.770 ;
        RECT 100.535 71.455 100.860 71.745 ;
        RECT 101.030 71.625 101.225 71.915 ;
        RECT 102.025 71.745 102.195 71.915 ;
        RECT 102.470 71.745 102.640 72.480 ;
        RECT 104.400 71.780 104.740 72.610 ;
        RECT 108.800 72.455 110.015 72.625 ;
        RECT 110.205 72.815 110.375 72.850 ;
        RECT 110.205 72.645 110.405 72.815 ;
        RECT 101.535 71.575 102.195 71.745 ;
        RECT 101.535 71.455 101.705 71.575 ;
        RECT 100.535 71.285 101.705 71.455 ;
        RECT 100.515 70.825 101.705 71.115 ;
        RECT 101.875 70.605 102.155 71.405 ;
        RECT 102.365 70.775 102.640 71.745 ;
        RECT 106.220 71.040 106.570 72.290 ;
        RECT 110.205 72.285 110.375 72.645 ;
        RECT 110.635 72.610 115.980 73.155 ;
        RECT 108.860 72.135 109.120 72.245 ;
        RECT 108.855 71.965 109.120 72.135 ;
        RECT 108.860 71.915 109.120 71.965 ;
        RECT 109.300 71.915 109.685 72.245 ;
        RECT 109.855 72.115 110.375 72.285 ;
        RECT 102.815 70.605 108.160 71.040 ;
        RECT 108.800 70.605 109.120 71.745 ;
        RECT 109.300 70.865 109.495 71.915 ;
        RECT 109.855 71.735 110.025 72.115 ;
        RECT 109.675 71.455 110.025 71.735 ;
        RECT 110.215 71.585 110.460 71.945 ;
        RECT 112.220 71.780 112.560 72.610 ;
        RECT 116.155 72.405 117.365 73.155 ;
        RECT 109.675 70.775 110.005 71.455 ;
        RECT 110.205 70.605 110.460 71.405 ;
        RECT 114.040 71.040 114.390 72.290 ;
        RECT 116.155 71.865 116.675 72.405 ;
        RECT 117.535 72.355 117.845 73.155 ;
        RECT 118.050 72.355 118.745 72.985 ;
        RECT 118.915 72.610 124.260 73.155 ;
        RECT 116.845 71.695 117.365 72.235 ;
        RECT 117.545 71.915 117.880 72.185 ;
        RECT 118.050 71.755 118.220 72.355 ;
        RECT 118.390 71.915 118.725 72.165 ;
        RECT 120.500 71.780 120.840 72.610 ;
        RECT 124.435 72.405 125.645 73.155 ;
        RECT 125.815 72.430 126.105 73.155 ;
        RECT 110.635 70.605 115.980 71.040 ;
        RECT 116.155 70.605 117.365 71.695 ;
        RECT 117.535 70.605 117.815 71.745 ;
        RECT 117.985 70.775 118.315 71.755 ;
        RECT 118.485 70.605 118.745 71.745 ;
        RECT 122.320 71.040 122.670 72.290 ;
        RECT 124.435 71.865 124.955 72.405 ;
        RECT 126.735 72.355 127.430 72.985 ;
        RECT 127.635 72.355 127.945 73.155 ;
        RECT 128.115 72.355 128.425 73.155 ;
        RECT 128.630 72.355 129.325 72.985 ;
        RECT 130.430 72.585 130.685 72.935 ;
        RECT 130.855 72.755 131.185 73.155 ;
        RECT 131.355 72.585 131.525 72.935 ;
        RECT 131.695 72.755 132.075 73.155 ;
        RECT 130.430 72.415 132.095 72.585 ;
        RECT 132.265 72.480 132.540 72.825 ;
        RECT 133.340 72.645 133.580 73.155 ;
        RECT 133.760 72.645 134.040 72.975 ;
        RECT 134.270 72.645 134.485 73.155 ;
        RECT 125.125 71.695 125.645 72.235 ;
        RECT 126.755 71.915 127.090 72.165 ;
        RECT 118.915 70.605 124.260 71.040 ;
        RECT 124.435 70.605 125.645 71.695 ;
        RECT 125.815 70.605 126.105 71.770 ;
        RECT 127.260 71.755 127.430 72.355 ;
        RECT 127.600 71.915 127.935 72.185 ;
        RECT 128.125 71.915 128.460 72.185 ;
        RECT 128.630 71.755 128.800 72.355 ;
        RECT 131.925 72.245 132.095 72.415 ;
        RECT 128.970 71.915 129.305 72.165 ;
        RECT 130.415 71.915 130.760 72.245 ;
        RECT 130.930 71.915 131.755 72.245 ;
        RECT 131.925 71.915 132.200 72.245 ;
        RECT 126.735 70.605 126.995 71.745 ;
        RECT 127.165 70.775 127.495 71.755 ;
        RECT 127.665 70.605 127.945 71.745 ;
        RECT 128.115 70.605 128.395 71.745 ;
        RECT 128.565 70.775 128.895 71.755 ;
        RECT 129.065 70.605 129.325 71.745 ;
        RECT 130.435 71.455 130.760 71.745 ;
        RECT 130.930 71.625 131.125 71.915 ;
        RECT 131.925 71.745 132.095 71.915 ;
        RECT 132.370 71.745 132.540 72.480 ;
        RECT 133.235 71.915 133.590 72.475 ;
        RECT 133.760 71.745 133.930 72.645 ;
        RECT 134.100 71.915 134.365 72.475 ;
        RECT 134.655 72.415 135.270 72.985 ;
        RECT 135.490 72.585 135.745 72.935 ;
        RECT 135.915 72.755 136.245 73.155 ;
        RECT 136.415 72.585 136.585 72.935 ;
        RECT 136.755 72.755 137.135 73.155 ;
        RECT 135.490 72.415 137.155 72.585 ;
        RECT 137.325 72.480 137.600 72.825 ;
        RECT 134.615 71.745 134.785 72.245 ;
        RECT 131.435 71.575 132.095 71.745 ;
        RECT 131.435 71.455 131.605 71.575 ;
        RECT 130.435 71.285 131.605 71.455 ;
        RECT 130.415 70.825 131.605 71.115 ;
        RECT 131.775 70.605 132.055 71.405 ;
        RECT 132.265 70.775 132.540 71.745 ;
        RECT 133.360 71.575 134.785 71.745 ;
        RECT 133.360 71.400 133.750 71.575 ;
        RECT 134.235 70.605 134.565 71.405 ;
        RECT 134.955 71.395 135.270 72.415 ;
        RECT 136.985 72.245 137.155 72.415 ;
        RECT 135.475 71.915 135.820 72.245 ;
        RECT 135.990 71.915 136.815 72.245 ;
        RECT 136.985 71.915 137.260 72.245 ;
        RECT 134.735 70.775 135.270 71.395 ;
        RECT 135.495 71.455 135.820 71.745 ;
        RECT 135.990 71.625 136.185 71.915 ;
        RECT 136.985 71.745 137.155 71.915 ;
        RECT 137.430 71.745 137.600 72.480 ;
        RECT 138.325 72.605 138.495 72.985 ;
        RECT 138.675 72.775 139.005 73.155 ;
        RECT 138.325 72.435 138.990 72.605 ;
        RECT 139.185 72.480 139.445 72.985 ;
        RECT 138.255 71.885 138.585 72.255 ;
        RECT 138.820 72.180 138.990 72.435 ;
        RECT 136.495 71.575 137.155 71.745 ;
        RECT 136.495 71.455 136.665 71.575 ;
        RECT 135.495 71.285 136.665 71.455 ;
        RECT 135.475 70.825 136.665 71.115 ;
        RECT 136.835 70.605 137.115 71.405 ;
        RECT 137.325 70.775 137.600 71.745 ;
        RECT 138.820 71.850 139.105 72.180 ;
        RECT 138.820 71.705 138.990 71.850 ;
        RECT 138.325 71.535 138.990 71.705 ;
        RECT 139.275 71.680 139.445 72.480 ;
        RECT 139.705 72.605 139.875 72.985 ;
        RECT 140.055 72.775 140.385 73.155 ;
        RECT 139.705 72.435 140.370 72.605 ;
        RECT 140.565 72.480 140.825 72.985 ;
        RECT 141.175 72.495 141.515 73.155 ;
        RECT 139.635 71.885 139.965 72.255 ;
        RECT 140.200 72.180 140.370 72.435 ;
        RECT 140.200 71.850 140.485 72.180 ;
        RECT 140.200 71.705 140.370 71.850 ;
        RECT 138.325 70.775 138.495 71.535 ;
        RECT 138.675 70.605 139.005 71.365 ;
        RECT 139.175 70.775 139.445 71.680 ;
        RECT 139.705 71.535 140.370 71.705 ;
        RECT 140.655 71.680 140.825 72.480 ;
        RECT 139.705 70.775 139.875 71.535 ;
        RECT 140.055 70.605 140.385 71.365 ;
        RECT 140.555 70.775 140.825 71.680 ;
        RECT 140.995 70.775 141.515 72.325 ;
        RECT 141.685 71.500 142.205 72.985 ;
        RECT 142.375 72.385 145.885 73.155 ;
        RECT 142.375 71.865 144.025 72.385 ;
        RECT 146.985 72.345 147.255 73.155 ;
        RECT 147.425 72.345 147.755 72.985 ;
        RECT 147.925 72.345 148.165 73.155 ;
        RECT 148.355 72.385 150.945 73.155 ;
        RECT 151.575 72.430 151.865 73.155 ;
        RECT 152.035 72.385 155.545 73.155 ;
        RECT 155.715 72.405 156.925 73.155 ;
        RECT 144.195 71.695 145.885 72.215 ;
        RECT 146.975 71.915 147.325 72.165 ;
        RECT 147.495 71.745 147.665 72.345 ;
        RECT 147.835 71.915 148.185 72.165 ;
        RECT 148.355 71.865 149.565 72.385 ;
        RECT 141.685 70.605 142.015 71.330 ;
        RECT 142.375 70.605 145.885 71.695 ;
        RECT 146.985 70.605 147.315 71.745 ;
        RECT 147.495 71.575 148.175 71.745 ;
        RECT 149.735 71.695 150.945 72.215 ;
        RECT 152.035 71.865 153.685 72.385 ;
        RECT 147.845 70.790 148.175 71.575 ;
        RECT 148.355 70.605 150.945 71.695 ;
        RECT 151.575 70.605 151.865 71.770 ;
        RECT 153.855 71.695 155.545 72.215 ;
        RECT 152.035 70.605 155.545 71.695 ;
        RECT 155.715 71.695 156.235 72.235 ;
        RECT 156.405 71.865 156.925 72.405 ;
        RECT 155.715 70.605 156.925 71.695 ;
        RECT 22.690 70.435 157.010 70.605 ;
        RECT 22.775 69.345 23.985 70.435 ;
        RECT 24.155 69.345 27.665 70.435 ;
        RECT 22.775 68.635 23.295 69.175 ;
        RECT 23.465 68.805 23.985 69.345 ;
        RECT 24.155 68.655 25.805 69.175 ;
        RECT 25.975 68.825 27.665 69.345 ;
        RECT 28.305 69.465 28.635 70.250 ;
        RECT 28.305 69.295 28.985 69.465 ;
        RECT 29.165 69.295 29.495 70.435 ;
        RECT 29.685 69.295 30.015 70.435 ;
        RECT 30.545 69.465 30.875 70.250 ;
        RECT 30.195 69.295 30.875 69.465 ;
        RECT 31.065 69.295 31.395 70.435 ;
        RECT 31.925 69.465 32.255 70.250 ;
        RECT 31.575 69.295 32.255 69.465 ;
        RECT 33.355 69.295 33.635 70.435 ;
        RECT 28.295 68.875 28.645 69.125 ;
        RECT 28.815 68.695 28.985 69.295 ;
        RECT 29.155 68.875 29.505 69.125 ;
        RECT 29.675 68.875 30.025 69.125 ;
        RECT 30.195 68.695 30.365 69.295 ;
        RECT 30.535 68.875 30.885 69.125 ;
        RECT 31.055 68.875 31.405 69.125 ;
        RECT 31.575 68.695 31.745 69.295 ;
        RECT 33.805 69.285 34.135 70.265 ;
        RECT 34.305 69.295 34.565 70.435 ;
        RECT 31.915 68.875 32.265 69.125 ;
        RECT 33.365 68.855 33.700 69.125 ;
        RECT 22.775 67.885 23.985 68.635 ;
        RECT 24.155 67.885 27.665 68.655 ;
        RECT 28.315 67.885 28.555 68.695 ;
        RECT 28.725 68.055 29.055 68.695 ;
        RECT 29.225 67.885 29.495 68.695 ;
        RECT 29.685 67.885 29.955 68.695 ;
        RECT 30.125 68.055 30.455 68.695 ;
        RECT 30.625 67.885 30.865 68.695 ;
        RECT 31.065 67.885 31.335 68.695 ;
        RECT 31.505 68.055 31.835 68.695 ;
        RECT 32.005 67.885 32.245 68.695 ;
        RECT 33.870 68.685 34.040 69.285 ;
        RECT 35.655 69.270 35.945 70.435 ;
        RECT 37.220 69.465 37.610 69.640 ;
        RECT 38.095 69.635 38.425 70.435 ;
        RECT 38.595 69.645 39.130 70.265 ;
        RECT 39.335 70.000 44.680 70.435 ;
        RECT 37.220 69.295 38.645 69.465 ;
        RECT 34.210 68.875 34.545 69.125 ;
        RECT 33.355 67.885 33.665 68.685 ;
        RECT 33.870 68.055 34.565 68.685 ;
        RECT 35.655 67.885 35.945 68.610 ;
        RECT 37.095 68.565 37.450 69.125 ;
        RECT 37.620 68.395 37.790 69.295 ;
        RECT 37.960 68.565 38.225 69.125 ;
        RECT 38.475 68.795 38.645 69.295 ;
        RECT 38.815 68.625 39.130 69.645 ;
        RECT 37.200 67.885 37.440 68.395 ;
        RECT 37.620 68.065 37.900 68.395 ;
        RECT 38.130 67.885 38.345 68.395 ;
        RECT 38.515 68.055 39.130 68.625 ;
        RECT 40.920 68.430 41.260 69.260 ;
        RECT 42.740 68.750 43.090 70.000 ;
        RECT 44.855 69.345 47.445 70.435 ;
        RECT 44.855 68.655 46.065 69.175 ;
        RECT 46.235 68.825 47.445 69.345 ;
        RECT 48.260 69.465 48.650 69.640 ;
        RECT 49.135 69.635 49.465 70.435 ;
        RECT 49.635 69.645 50.170 70.265 ;
        RECT 48.260 69.295 49.685 69.465 ;
        RECT 39.335 67.885 44.680 68.430 ;
        RECT 44.855 67.885 47.445 68.655 ;
        RECT 48.135 68.565 48.490 69.125 ;
        RECT 48.660 68.395 48.830 69.295 ;
        RECT 49.000 68.565 49.265 69.125 ;
        RECT 49.515 68.795 49.685 69.295 ;
        RECT 49.855 68.625 50.170 69.645 ;
        RECT 50.845 69.465 51.175 70.250 ;
        RECT 50.845 69.295 51.525 69.465 ;
        RECT 51.705 69.295 52.035 70.435 ;
        RECT 52.225 69.295 52.555 70.435 ;
        RECT 53.085 69.465 53.415 70.250 ;
        RECT 52.735 69.295 53.415 69.465 ;
        RECT 53.595 69.295 53.855 70.435 ;
        RECT 50.835 68.875 51.185 69.125 ;
        RECT 51.355 68.695 51.525 69.295 ;
        RECT 51.695 68.875 52.045 69.125 ;
        RECT 52.215 68.875 52.565 69.125 ;
        RECT 52.735 68.695 52.905 69.295 ;
        RECT 54.025 69.285 54.355 70.265 ;
        RECT 54.525 69.295 54.805 70.435 ;
        RECT 55.985 69.765 56.155 70.265 ;
        RECT 56.325 69.935 56.655 70.435 ;
        RECT 55.985 69.595 56.590 69.765 ;
        RECT 53.075 68.875 53.425 69.125 ;
        RECT 53.615 68.875 53.950 69.125 ;
        RECT 54.120 68.735 54.290 69.285 ;
        RECT 54.460 68.855 54.795 69.125 ;
        RECT 55.895 68.785 56.140 69.425 ;
        RECT 56.420 69.200 56.590 69.595 ;
        RECT 56.825 69.485 57.050 70.265 ;
        RECT 56.420 68.870 56.650 69.200 ;
        RECT 48.240 67.885 48.480 68.395 ;
        RECT 48.660 68.065 48.940 68.395 ;
        RECT 49.170 67.885 49.385 68.395 ;
        RECT 49.555 68.055 50.170 68.625 ;
        RECT 50.855 67.885 51.095 68.695 ;
        RECT 51.265 68.055 51.595 68.695 ;
        RECT 51.765 67.885 52.035 68.695 ;
        RECT 52.225 67.885 52.495 68.695 ;
        RECT 52.665 68.055 52.995 68.695 ;
        RECT 53.165 67.885 53.405 68.695 ;
        RECT 54.115 68.685 54.290 68.735 ;
        RECT 53.595 68.055 54.290 68.685 ;
        RECT 54.495 67.885 54.805 68.685 ;
        RECT 56.420 68.605 56.590 68.870 ;
        RECT 55.985 68.435 56.590 68.605 ;
        RECT 55.985 68.145 56.155 68.435 ;
        RECT 56.325 67.885 56.655 68.265 ;
        RECT 56.825 68.145 56.995 69.485 ;
        RECT 57.240 69.465 57.595 70.215 ;
        RECT 57.765 69.635 58.055 70.435 ;
        RECT 58.555 70.055 59.415 70.225 ;
        RECT 59.105 69.905 59.415 70.055 ;
        RECT 59.585 69.975 59.905 70.435 ;
        RECT 59.105 69.890 59.430 69.905 ;
        RECT 59.200 69.885 59.430 69.890 ;
        RECT 59.200 69.865 59.440 69.885 ;
        RECT 59.200 69.845 59.455 69.865 ;
        RECT 59.215 69.835 59.455 69.845 ;
        RECT 59.240 69.810 59.455 69.835 ;
        RECT 57.240 69.295 57.925 69.465 ;
        RECT 57.245 68.755 57.575 69.125 ;
        RECT 57.755 69.035 57.925 69.295 ;
        RECT 58.255 69.155 58.590 69.805 ;
        RECT 58.760 69.360 59.095 69.710 ;
        RECT 57.755 68.585 58.130 69.035 ;
        RECT 58.760 68.840 59.075 69.360 ;
        RECT 59.265 69.250 59.455 69.810 ;
        RECT 60.105 69.665 60.350 70.235 ;
        RECT 59.625 69.335 60.350 69.665 ;
        RECT 60.530 69.370 60.815 70.435 ;
        RECT 60.985 69.470 61.245 70.255 ;
        RECT 57.320 68.565 58.130 68.585 ;
        RECT 57.320 68.415 57.925 68.565 ;
        RECT 58.370 68.535 59.075 68.840 ;
        RECT 59.245 69.125 59.455 69.250 ;
        RECT 60.180 69.125 60.350 69.335 ;
        RECT 59.245 68.795 60.010 69.125 ;
        RECT 60.180 68.795 60.905 69.125 ;
        RECT 57.320 68.145 57.515 68.415 ;
        RECT 59.245 68.335 59.415 68.795 ;
        RECT 60.180 68.520 60.350 68.795 ;
        RECT 61.075 68.545 61.245 69.470 ;
        RECT 61.415 69.270 61.705 70.435 ;
        RECT 62.855 69.375 63.185 70.220 ;
        RECT 63.355 69.425 63.525 70.435 ;
        RECT 63.695 69.705 64.035 70.265 ;
        RECT 64.265 69.935 64.580 70.435 ;
        RECT 64.760 69.965 65.645 70.135 ;
        RECT 62.795 69.295 63.185 69.375 ;
        RECT 63.695 69.330 64.590 69.705 ;
        RECT 62.795 69.245 63.010 69.295 ;
        RECT 62.795 68.665 62.965 69.245 ;
        RECT 63.695 69.125 63.885 69.330 ;
        RECT 64.760 69.125 64.930 69.965 ;
        RECT 65.870 69.935 66.120 70.265 ;
        RECT 63.135 68.795 63.885 69.125 ;
        RECT 64.055 68.795 64.930 69.125 ;
        RECT 62.795 68.625 63.020 68.665 ;
        RECT 63.685 68.625 63.885 68.795 ;
        RECT 57.685 67.885 58.015 68.245 ;
        RECT 58.575 68.165 59.415 68.335 ;
        RECT 59.585 67.885 59.855 68.345 ;
        RECT 60.105 68.060 60.350 68.520 ;
        RECT 60.565 67.885 60.790 68.515 ;
        RECT 60.985 68.215 61.245 68.545 ;
        RECT 61.415 67.885 61.705 68.610 ;
        RECT 62.795 68.540 63.175 68.625 ;
        RECT 62.845 68.105 63.175 68.540 ;
        RECT 63.345 67.885 63.515 68.495 ;
        RECT 63.685 68.100 64.015 68.625 ;
        RECT 64.275 67.885 64.485 68.415 ;
        RECT 64.760 68.335 64.930 68.795 ;
        RECT 65.100 68.835 65.420 69.795 ;
        RECT 65.590 69.045 65.780 69.765 ;
        RECT 65.950 68.865 66.120 69.935 ;
        RECT 66.290 69.635 66.460 70.435 ;
        RECT 66.630 69.990 67.735 70.160 ;
        RECT 66.630 69.375 66.800 69.990 ;
        RECT 67.945 69.840 68.195 70.265 ;
        RECT 68.365 69.975 68.630 70.435 ;
        RECT 66.970 69.455 67.500 69.820 ;
        RECT 67.945 69.710 68.250 69.840 ;
        RECT 66.290 69.285 66.800 69.375 ;
        RECT 66.290 69.115 67.160 69.285 ;
        RECT 66.290 69.045 66.460 69.115 ;
        RECT 66.580 68.865 66.780 68.895 ;
        RECT 65.100 68.505 65.565 68.835 ;
        RECT 65.950 68.565 66.780 68.865 ;
        RECT 65.950 68.335 66.120 68.565 ;
        RECT 64.760 68.165 65.545 68.335 ;
        RECT 65.715 68.165 66.120 68.335 ;
        RECT 66.300 67.885 66.670 68.385 ;
        RECT 66.990 68.335 67.160 69.115 ;
        RECT 67.330 68.755 67.500 69.455 ;
        RECT 67.670 68.925 67.910 69.520 ;
        RECT 67.330 68.535 67.855 68.755 ;
        RECT 68.080 68.605 68.250 69.710 ;
        RECT 68.025 68.475 68.250 68.605 ;
        RECT 68.420 68.515 68.700 69.465 ;
        RECT 68.025 68.335 68.195 68.475 ;
        RECT 66.990 68.165 67.665 68.335 ;
        RECT 67.860 68.165 68.195 68.335 ;
        RECT 68.365 67.885 68.615 68.345 ;
        RECT 68.870 68.145 69.055 70.265 ;
        RECT 69.225 69.935 69.555 70.435 ;
        RECT 69.725 69.765 69.895 70.265 ;
        RECT 69.230 69.595 69.895 69.765 ;
        RECT 69.230 68.605 69.460 69.595 ;
        RECT 71.085 69.465 71.415 70.250 ;
        RECT 69.630 68.775 69.980 69.425 ;
        RECT 71.085 69.295 71.765 69.465 ;
        RECT 71.945 69.295 72.275 70.435 ;
        RECT 72.465 69.295 72.795 70.435 ;
        RECT 73.325 69.465 73.655 70.250 ;
        RECT 72.975 69.295 73.655 69.465 ;
        RECT 73.845 69.295 74.175 70.435 ;
        RECT 74.705 69.465 75.035 70.250 ;
        RECT 74.355 69.295 75.035 69.465 ;
        RECT 75.215 69.295 75.475 70.435 ;
        RECT 71.075 68.875 71.425 69.125 ;
        RECT 71.595 68.695 71.765 69.295 ;
        RECT 71.935 68.875 72.285 69.125 ;
        RECT 72.455 68.875 72.805 69.125 ;
        RECT 72.975 68.695 73.145 69.295 ;
        RECT 73.315 68.875 73.665 69.125 ;
        RECT 73.835 68.875 74.185 69.125 ;
        RECT 74.355 68.695 74.525 69.295 ;
        RECT 75.645 69.285 75.975 70.265 ;
        RECT 76.145 69.295 76.425 70.435 ;
        RECT 77.700 69.465 78.090 69.640 ;
        RECT 78.575 69.635 78.905 70.435 ;
        RECT 79.075 69.645 79.610 70.265 ;
        RECT 77.700 69.295 79.125 69.465 ;
        RECT 75.735 69.245 75.910 69.285 ;
        RECT 74.695 68.875 75.045 69.125 ;
        RECT 75.235 68.875 75.570 69.125 ;
        RECT 69.230 68.435 69.895 68.605 ;
        RECT 69.225 67.885 69.555 68.265 ;
        RECT 69.725 68.145 69.895 68.435 ;
        RECT 71.095 67.885 71.335 68.695 ;
        RECT 71.505 68.055 71.835 68.695 ;
        RECT 72.005 67.885 72.275 68.695 ;
        RECT 72.465 67.885 72.735 68.695 ;
        RECT 72.905 68.055 73.235 68.695 ;
        RECT 73.405 67.885 73.645 68.695 ;
        RECT 73.845 67.885 74.115 68.695 ;
        RECT 74.285 68.055 74.615 68.695 ;
        RECT 74.785 67.885 75.025 68.695 ;
        RECT 75.740 68.685 75.910 69.245 ;
        RECT 76.080 68.855 76.415 69.125 ;
        RECT 75.215 68.055 75.910 68.685 ;
        RECT 76.115 67.885 76.425 68.685 ;
        RECT 77.575 68.565 77.930 69.125 ;
        RECT 78.100 68.395 78.270 69.295 ;
        RECT 78.440 68.565 78.705 69.125 ;
        RECT 78.955 68.795 79.125 69.295 ;
        RECT 79.295 68.625 79.610 69.645 ;
        RECT 79.815 69.345 82.405 70.435 ;
        RECT 77.680 67.885 77.920 68.395 ;
        RECT 78.100 68.065 78.380 68.395 ;
        RECT 78.610 67.885 78.825 68.395 ;
        RECT 78.995 68.055 79.610 68.625 ;
        RECT 79.815 68.655 81.025 69.175 ;
        RECT 81.195 68.825 82.405 69.345 ;
        RECT 82.575 69.295 82.855 70.435 ;
        RECT 83.025 69.285 83.355 70.265 ;
        RECT 83.525 69.295 83.785 70.435 ;
        RECT 83.955 69.295 84.235 70.435 ;
        RECT 84.405 69.285 84.735 70.265 ;
        RECT 84.905 69.295 85.165 70.435 ;
        RECT 85.335 69.345 87.005 70.435 ;
        RECT 82.585 68.855 82.920 69.125 ;
        RECT 83.090 68.685 83.260 69.285 ;
        RECT 83.430 68.875 83.765 69.125 ;
        RECT 83.965 68.855 84.300 69.125 ;
        RECT 84.470 68.685 84.640 69.285 ;
        RECT 84.810 68.875 85.145 69.125 ;
        RECT 79.815 67.885 82.405 68.655 ;
        RECT 82.575 67.885 82.885 68.685 ;
        RECT 83.090 68.055 83.785 68.685 ;
        RECT 83.955 67.885 84.265 68.685 ;
        RECT 84.470 68.055 85.165 68.685 ;
        RECT 85.335 68.655 86.085 69.175 ;
        RECT 86.255 68.825 87.005 69.345 ;
        RECT 87.175 69.270 87.465 70.435 ;
        RECT 87.635 69.345 88.845 70.435 ;
        RECT 89.015 69.925 90.205 70.215 ;
        RECT 85.335 67.885 87.005 68.655 ;
        RECT 87.635 68.635 88.155 69.175 ;
        RECT 88.325 68.805 88.845 69.345 ;
        RECT 89.035 69.585 90.205 69.755 ;
        RECT 90.375 69.635 90.655 70.435 ;
        RECT 89.035 69.295 89.360 69.585 ;
        RECT 90.035 69.465 90.205 69.585 ;
        RECT 89.530 69.125 89.725 69.415 ;
        RECT 90.035 69.295 90.695 69.465 ;
        RECT 90.865 69.295 91.140 70.265 ;
        RECT 91.325 69.465 91.655 70.250 ;
        RECT 91.325 69.295 92.005 69.465 ;
        RECT 92.185 69.295 92.515 70.435 ;
        RECT 92.705 69.295 93.035 70.435 ;
        RECT 93.565 69.465 93.895 70.250 ;
        RECT 93.215 69.295 93.895 69.465 ;
        RECT 94.075 69.345 95.745 70.435 ;
        RECT 95.920 69.925 97.575 70.215 ;
        RECT 90.525 69.125 90.695 69.295 ;
        RECT 89.015 68.795 89.360 69.125 ;
        RECT 89.530 68.795 90.355 69.125 ;
        RECT 90.525 68.795 90.800 69.125 ;
        RECT 87.175 67.885 87.465 68.610 ;
        RECT 87.635 67.885 88.845 68.635 ;
        RECT 90.525 68.625 90.695 68.795 ;
        RECT 89.030 68.455 90.695 68.625 ;
        RECT 90.970 68.560 91.140 69.295 ;
        RECT 91.315 68.875 91.665 69.125 ;
        RECT 91.835 68.695 92.005 69.295 ;
        RECT 92.175 68.875 92.525 69.125 ;
        RECT 92.695 68.875 93.045 69.125 ;
        RECT 93.215 68.695 93.385 69.295 ;
        RECT 93.555 68.875 93.905 69.125 ;
        RECT 89.030 68.105 89.285 68.455 ;
        RECT 89.455 67.885 89.785 68.285 ;
        RECT 89.955 68.105 90.125 68.455 ;
        RECT 90.295 67.885 90.675 68.285 ;
        RECT 90.865 68.215 91.140 68.560 ;
        RECT 91.335 67.885 91.575 68.695 ;
        RECT 91.745 68.055 92.075 68.695 ;
        RECT 92.245 67.885 92.515 68.695 ;
        RECT 92.705 67.885 92.975 68.695 ;
        RECT 93.145 68.055 93.475 68.695 ;
        RECT 93.645 67.885 93.885 68.695 ;
        RECT 94.075 68.655 94.825 69.175 ;
        RECT 94.995 68.825 95.745 69.345 ;
        RECT 95.920 69.585 97.510 69.755 ;
        RECT 97.745 69.635 98.025 70.435 ;
        RECT 95.920 69.295 96.240 69.585 ;
        RECT 97.340 69.465 97.510 69.585 ;
        RECT 96.435 69.245 97.150 69.415 ;
        RECT 97.340 69.295 98.065 69.465 ;
        RECT 98.235 69.295 98.505 70.265 ;
        RECT 99.685 69.505 99.855 70.265 ;
        RECT 100.035 69.675 100.365 70.435 ;
        RECT 99.685 69.335 100.350 69.505 ;
        RECT 100.535 69.360 100.805 70.265 ;
        RECT 101.065 69.765 101.235 70.265 ;
        RECT 101.405 69.935 101.735 70.435 ;
        RECT 101.065 69.595 101.670 69.765 ;
        RECT 94.075 67.885 95.745 68.655 ;
        RECT 95.920 68.555 96.270 69.125 ;
        RECT 96.440 68.795 97.150 69.245 ;
        RECT 97.895 69.125 98.065 69.295 ;
        RECT 97.320 68.795 97.725 69.125 ;
        RECT 97.895 68.795 98.165 69.125 ;
        RECT 97.895 68.625 98.065 68.795 ;
        RECT 96.455 68.455 98.065 68.625 ;
        RECT 98.335 68.560 98.505 69.295 ;
        RECT 100.180 69.190 100.350 69.335 ;
        RECT 99.615 68.785 99.945 69.155 ;
        RECT 100.180 68.860 100.465 69.190 ;
        RECT 100.180 68.605 100.350 68.860 ;
        RECT 95.925 67.885 96.255 68.385 ;
        RECT 96.455 68.105 96.625 68.455 ;
        RECT 96.825 67.885 97.155 68.285 ;
        RECT 97.325 68.105 97.495 68.455 ;
        RECT 97.665 67.885 98.045 68.285 ;
        RECT 98.235 68.215 98.505 68.560 ;
        RECT 99.685 68.435 100.350 68.605 ;
        RECT 100.635 68.560 100.805 69.360 ;
        RECT 100.975 68.785 101.220 69.425 ;
        RECT 101.500 69.200 101.670 69.595 ;
        RECT 101.905 69.485 102.130 70.265 ;
        RECT 101.500 68.870 101.730 69.200 ;
        RECT 101.500 68.605 101.670 68.870 ;
        RECT 99.685 68.055 99.855 68.435 ;
        RECT 100.035 67.885 100.365 68.265 ;
        RECT 100.545 68.055 100.805 68.560 ;
        RECT 101.065 68.435 101.670 68.605 ;
        RECT 101.065 68.145 101.235 68.435 ;
        RECT 101.405 67.885 101.735 68.265 ;
        RECT 101.905 68.145 102.075 69.485 ;
        RECT 102.320 69.465 102.675 70.215 ;
        RECT 102.845 69.635 103.135 70.435 ;
        RECT 103.635 70.055 104.495 70.225 ;
        RECT 104.185 69.905 104.495 70.055 ;
        RECT 104.665 69.975 104.985 70.435 ;
        RECT 104.185 69.890 104.510 69.905 ;
        RECT 104.280 69.885 104.510 69.890 ;
        RECT 104.280 69.865 104.520 69.885 ;
        RECT 104.280 69.845 104.535 69.865 ;
        RECT 104.295 69.835 104.535 69.845 ;
        RECT 104.320 69.810 104.535 69.835 ;
        RECT 102.320 69.295 103.005 69.465 ;
        RECT 102.325 68.755 102.655 69.125 ;
        RECT 102.835 69.035 103.005 69.295 ;
        RECT 103.335 69.155 103.670 69.805 ;
        RECT 103.840 69.360 104.175 69.710 ;
        RECT 102.835 68.585 103.210 69.035 ;
        RECT 103.840 68.840 104.155 69.360 ;
        RECT 104.345 69.250 104.535 69.810 ;
        RECT 105.185 69.665 105.430 70.235 ;
        RECT 104.705 69.335 105.430 69.665 ;
        RECT 105.610 69.370 105.895 70.435 ;
        RECT 106.065 69.470 106.325 70.255 ;
        RECT 102.400 68.565 103.210 68.585 ;
        RECT 102.400 68.415 103.005 68.565 ;
        RECT 103.450 68.535 104.155 68.840 ;
        RECT 104.325 69.125 104.535 69.250 ;
        RECT 105.260 69.125 105.430 69.335 ;
        RECT 104.325 68.795 105.090 69.125 ;
        RECT 105.260 68.795 105.985 69.125 ;
        RECT 102.400 68.145 102.595 68.415 ;
        RECT 104.325 68.335 104.495 68.795 ;
        RECT 105.260 68.520 105.430 68.795 ;
        RECT 106.155 68.545 106.325 69.470 ;
        RECT 106.495 69.345 108.165 70.435 ;
        RECT 102.765 67.885 103.095 68.245 ;
        RECT 103.655 68.165 104.495 68.335 ;
        RECT 104.665 67.885 104.935 68.345 ;
        RECT 105.185 68.060 105.430 68.520 ;
        RECT 105.645 67.885 105.870 68.515 ;
        RECT 106.065 68.215 106.325 68.545 ;
        RECT 106.495 68.655 107.245 69.175 ;
        RECT 107.415 68.825 108.165 69.345 ;
        RECT 108.335 69.565 108.610 70.265 ;
        RECT 108.780 69.890 109.035 70.435 ;
        RECT 109.205 69.925 109.685 70.265 ;
        RECT 109.860 69.880 110.465 70.435 ;
        RECT 109.850 69.780 110.465 69.880 ;
        RECT 109.850 69.755 110.035 69.780 ;
        RECT 106.495 67.885 108.165 68.655 ;
        RECT 108.335 68.535 108.505 69.565 ;
        RECT 108.780 69.435 109.535 69.685 ;
        RECT 109.705 69.510 110.035 69.755 ;
        RECT 108.780 69.400 109.550 69.435 ;
        RECT 108.780 69.390 109.565 69.400 ;
        RECT 108.675 69.375 109.570 69.390 ;
        RECT 108.675 69.360 109.590 69.375 ;
        RECT 108.675 69.350 109.610 69.360 ;
        RECT 108.675 69.340 109.635 69.350 ;
        RECT 108.675 69.310 109.705 69.340 ;
        RECT 108.675 69.280 109.725 69.310 ;
        RECT 108.675 69.250 109.745 69.280 ;
        RECT 108.675 69.225 109.775 69.250 ;
        RECT 108.675 69.190 109.810 69.225 ;
        RECT 108.675 69.185 109.840 69.190 ;
        RECT 108.675 68.790 108.905 69.185 ;
        RECT 109.450 69.180 109.840 69.185 ;
        RECT 109.475 69.170 109.840 69.180 ;
        RECT 109.490 69.165 109.840 69.170 ;
        RECT 109.505 69.160 109.840 69.165 ;
        RECT 110.205 69.160 110.465 69.610 ;
        RECT 110.635 69.295 110.895 70.435 ;
        RECT 111.065 69.285 111.395 70.265 ;
        RECT 111.565 69.295 111.845 70.435 ;
        RECT 109.505 69.155 110.465 69.160 ;
        RECT 109.515 69.145 110.465 69.155 ;
        RECT 109.525 69.140 110.465 69.145 ;
        RECT 109.535 69.130 110.465 69.140 ;
        RECT 109.540 69.120 110.465 69.130 ;
        RECT 109.545 69.115 110.465 69.120 ;
        RECT 109.555 69.100 110.465 69.115 ;
        RECT 109.560 69.085 110.465 69.100 ;
        RECT 109.570 69.060 110.465 69.085 ;
        RECT 109.075 68.590 109.405 69.015 ;
        RECT 108.335 68.055 108.595 68.535 ;
        RECT 108.765 67.885 109.015 68.425 ;
        RECT 109.185 68.105 109.405 68.590 ;
        RECT 109.575 68.990 110.465 69.060 ;
        RECT 109.575 68.265 109.745 68.990 ;
        RECT 110.655 68.875 110.990 69.125 ;
        RECT 109.915 68.435 110.465 68.820 ;
        RECT 111.160 68.685 111.330 69.285 ;
        RECT 112.935 69.270 113.225 70.435 ;
        RECT 113.395 69.345 115.065 70.435 ;
        RECT 111.500 68.855 111.835 69.125 ;
        RECT 109.575 68.095 110.465 68.265 ;
        RECT 110.635 68.055 111.330 68.685 ;
        RECT 111.535 67.885 111.845 68.685 ;
        RECT 113.395 68.655 114.145 69.175 ;
        RECT 114.315 68.825 115.065 69.345 ;
        RECT 115.245 69.465 115.575 70.250 ;
        RECT 115.245 69.295 115.925 69.465 ;
        RECT 116.105 69.295 116.435 70.435 ;
        RECT 116.625 69.295 116.955 70.435 ;
        RECT 117.485 69.465 117.815 70.250 ;
        RECT 117.135 69.295 117.815 69.465 ;
        RECT 118.005 69.295 118.335 70.435 ;
        RECT 118.865 69.465 119.195 70.250 ;
        RECT 118.515 69.295 119.195 69.465 ;
        RECT 119.385 69.465 119.715 70.250 ;
        RECT 119.385 69.295 120.065 69.465 ;
        RECT 120.245 69.295 120.575 70.435 ;
        RECT 121.675 69.295 121.955 70.435 ;
        RECT 115.235 68.875 115.585 69.125 ;
        RECT 115.755 68.695 115.925 69.295 ;
        RECT 116.095 68.875 116.445 69.125 ;
        RECT 116.615 68.875 116.965 69.125 ;
        RECT 117.135 68.695 117.305 69.295 ;
        RECT 117.475 68.875 117.825 69.125 ;
        RECT 117.995 68.875 118.345 69.125 ;
        RECT 118.515 68.695 118.685 69.295 ;
        RECT 118.855 68.875 119.205 69.125 ;
        RECT 119.375 68.875 119.725 69.125 ;
        RECT 119.895 68.695 120.065 69.295 ;
        RECT 122.125 69.285 122.455 70.265 ;
        RECT 122.625 69.295 122.885 70.435 ;
        RECT 123.550 69.645 124.085 70.265 ;
        RECT 122.190 69.245 122.365 69.285 ;
        RECT 120.235 68.875 120.585 69.125 ;
        RECT 121.685 68.855 122.020 69.125 ;
        RECT 112.935 67.885 113.225 68.610 ;
        RECT 113.395 67.885 115.065 68.655 ;
        RECT 115.255 67.885 115.495 68.695 ;
        RECT 115.665 68.055 115.995 68.695 ;
        RECT 116.165 67.885 116.435 68.695 ;
        RECT 116.625 67.885 116.895 68.695 ;
        RECT 117.065 68.055 117.395 68.695 ;
        RECT 117.565 67.885 117.805 68.695 ;
        RECT 118.005 67.885 118.275 68.695 ;
        RECT 118.445 68.055 118.775 68.695 ;
        RECT 118.945 67.885 119.185 68.695 ;
        RECT 119.395 67.885 119.635 68.695 ;
        RECT 119.805 68.055 120.135 68.695 ;
        RECT 120.305 67.885 120.575 68.695 ;
        RECT 122.190 68.685 122.360 69.245 ;
        RECT 122.530 68.875 122.865 69.125 ;
        RECT 121.675 67.885 121.985 68.685 ;
        RECT 122.190 68.055 122.885 68.685 ;
        RECT 123.550 68.625 123.865 69.645 ;
        RECT 124.255 69.635 124.585 70.435 ;
        RECT 125.070 69.465 125.460 69.640 ;
        RECT 124.035 69.295 125.460 69.465 ;
        RECT 125.815 69.345 129.325 70.435 ;
        RECT 124.035 68.795 124.205 69.295 ;
        RECT 123.550 68.055 124.165 68.625 ;
        RECT 124.455 68.565 124.720 69.125 ;
        RECT 124.890 68.395 125.060 69.295 ;
        RECT 125.230 68.565 125.585 69.125 ;
        RECT 125.815 68.655 127.465 69.175 ;
        RECT 127.635 68.825 129.325 69.345 ;
        RECT 129.965 69.465 130.295 70.250 ;
        RECT 129.965 69.295 130.645 69.465 ;
        RECT 130.825 69.295 131.155 70.435 ;
        RECT 131.345 69.465 131.675 70.250 ;
        RECT 131.345 69.295 132.025 69.465 ;
        RECT 132.205 69.295 132.535 70.435 ;
        RECT 132.725 69.295 133.055 70.435 ;
        RECT 133.585 69.465 133.915 70.250 ;
        RECT 133.235 69.295 133.915 69.465 ;
        RECT 134.095 69.345 136.685 70.435 ;
        RECT 129.955 68.875 130.305 69.125 ;
        RECT 130.475 68.695 130.645 69.295 ;
        RECT 130.815 68.875 131.165 69.125 ;
        RECT 131.335 68.875 131.685 69.125 ;
        RECT 131.855 68.695 132.025 69.295 ;
        RECT 132.195 68.875 132.545 69.125 ;
        RECT 132.715 68.875 133.065 69.125 ;
        RECT 133.235 68.695 133.405 69.295 ;
        RECT 133.575 68.875 133.925 69.125 ;
        RECT 124.335 67.885 124.550 68.395 ;
        RECT 124.780 68.065 125.060 68.395 ;
        RECT 125.240 67.885 125.480 68.395 ;
        RECT 125.815 67.885 129.325 68.655 ;
        RECT 129.975 67.885 130.215 68.695 ;
        RECT 130.385 68.055 130.715 68.695 ;
        RECT 130.885 67.885 131.155 68.695 ;
        RECT 131.355 67.885 131.595 68.695 ;
        RECT 131.765 68.055 132.095 68.695 ;
        RECT 132.265 67.885 132.535 68.695 ;
        RECT 132.725 67.885 132.995 68.695 ;
        RECT 133.165 68.055 133.495 68.695 ;
        RECT 133.665 67.885 133.905 68.695 ;
        RECT 134.095 68.655 135.305 69.175 ;
        RECT 135.475 68.825 136.685 69.345 ;
        RECT 136.855 68.715 137.375 70.265 ;
        RECT 137.545 69.710 137.875 70.435 ;
        RECT 134.095 67.885 136.685 68.655 ;
        RECT 137.035 67.885 137.375 68.545 ;
        RECT 137.545 68.055 138.065 69.540 ;
        RECT 138.695 69.270 138.985 70.435 ;
        RECT 139.705 69.765 139.875 70.265 ;
        RECT 140.045 69.935 140.375 70.435 ;
        RECT 139.705 69.595 140.310 69.765 ;
        RECT 139.615 68.785 139.860 69.425 ;
        RECT 140.140 69.200 140.310 69.595 ;
        RECT 140.545 69.485 140.770 70.265 ;
        RECT 140.140 68.870 140.370 69.200 ;
        RECT 138.695 67.885 138.985 68.610 ;
        RECT 140.140 68.605 140.310 68.870 ;
        RECT 139.705 68.435 140.310 68.605 ;
        RECT 139.705 68.145 139.875 68.435 ;
        RECT 140.045 67.885 140.375 68.265 ;
        RECT 140.545 68.145 140.715 69.485 ;
        RECT 140.960 69.465 141.315 70.215 ;
        RECT 141.485 69.635 141.775 70.435 ;
        RECT 142.275 70.055 143.135 70.225 ;
        RECT 142.825 69.905 143.135 70.055 ;
        RECT 143.305 69.975 143.625 70.435 ;
        RECT 142.825 69.890 143.150 69.905 ;
        RECT 142.920 69.885 143.150 69.890 ;
        RECT 142.920 69.865 143.160 69.885 ;
        RECT 142.920 69.845 143.175 69.865 ;
        RECT 142.935 69.835 143.175 69.845 ;
        RECT 142.960 69.810 143.175 69.835 ;
        RECT 140.960 69.295 141.645 69.465 ;
        RECT 140.965 68.755 141.295 69.125 ;
        RECT 141.475 69.035 141.645 69.295 ;
        RECT 141.975 69.155 142.310 69.805 ;
        RECT 142.480 69.360 142.815 69.710 ;
        RECT 141.475 68.585 141.850 69.035 ;
        RECT 142.480 68.840 142.795 69.360 ;
        RECT 142.985 69.250 143.175 69.810 ;
        RECT 143.825 69.665 144.070 70.235 ;
        RECT 143.345 69.335 144.070 69.665 ;
        RECT 144.250 69.370 144.535 70.435 ;
        RECT 144.705 69.470 144.965 70.255 ;
        RECT 141.040 68.565 141.850 68.585 ;
        RECT 141.040 68.415 141.645 68.565 ;
        RECT 142.090 68.535 142.795 68.840 ;
        RECT 142.965 69.125 143.175 69.250 ;
        RECT 143.900 69.125 144.070 69.335 ;
        RECT 142.965 68.795 143.730 69.125 ;
        RECT 143.900 68.795 144.625 69.125 ;
        RECT 141.040 68.145 141.235 68.415 ;
        RECT 142.965 68.335 143.135 68.795 ;
        RECT 143.900 68.520 144.070 68.795 ;
        RECT 144.795 68.545 144.965 69.470 ;
        RECT 141.405 67.885 141.735 68.245 ;
        RECT 142.295 68.165 143.135 68.335 ;
        RECT 143.305 67.885 143.575 68.345 ;
        RECT 143.825 68.060 144.070 68.520 ;
        RECT 144.285 67.885 144.510 68.515 ;
        RECT 144.705 68.215 144.965 68.545 ;
        RECT 145.135 69.360 145.405 70.265 ;
        RECT 145.575 69.675 145.905 70.435 ;
        RECT 146.085 69.505 146.255 70.265 ;
        RECT 145.135 68.560 145.305 69.360 ;
        RECT 145.590 69.335 146.255 69.505 ;
        RECT 146.515 69.565 146.790 70.265 ;
        RECT 146.960 69.890 147.215 70.435 ;
        RECT 147.385 69.925 147.865 70.265 ;
        RECT 148.040 69.880 148.645 70.435 ;
        RECT 148.030 69.780 148.645 69.880 ;
        RECT 148.030 69.755 148.215 69.780 ;
        RECT 145.590 69.190 145.760 69.335 ;
        RECT 145.475 68.860 145.760 69.190 ;
        RECT 145.590 68.605 145.760 68.860 ;
        RECT 145.995 68.785 146.325 69.155 ;
        RECT 145.135 68.055 145.395 68.560 ;
        RECT 145.590 68.435 146.255 68.605 ;
        RECT 145.575 67.885 145.905 68.265 ;
        RECT 146.085 68.055 146.255 68.435 ;
        RECT 146.515 68.535 146.685 69.565 ;
        RECT 146.960 69.435 147.715 69.685 ;
        RECT 147.885 69.510 148.215 69.755 ;
        RECT 148.850 69.645 149.385 70.265 ;
        RECT 146.960 69.400 147.730 69.435 ;
        RECT 146.960 69.390 147.745 69.400 ;
        RECT 146.855 69.375 147.750 69.390 ;
        RECT 146.855 69.360 147.770 69.375 ;
        RECT 146.855 69.350 147.790 69.360 ;
        RECT 146.855 69.340 147.815 69.350 ;
        RECT 146.855 69.310 147.885 69.340 ;
        RECT 146.855 69.280 147.905 69.310 ;
        RECT 146.855 69.250 147.925 69.280 ;
        RECT 146.855 69.225 147.955 69.250 ;
        RECT 146.855 69.190 147.990 69.225 ;
        RECT 146.855 69.185 148.020 69.190 ;
        RECT 146.855 68.790 147.085 69.185 ;
        RECT 147.630 69.180 148.020 69.185 ;
        RECT 147.655 69.170 148.020 69.180 ;
        RECT 147.670 69.165 148.020 69.170 ;
        RECT 147.685 69.160 148.020 69.165 ;
        RECT 148.385 69.160 148.645 69.610 ;
        RECT 147.685 69.155 148.645 69.160 ;
        RECT 147.695 69.145 148.645 69.155 ;
        RECT 147.705 69.140 148.645 69.145 ;
        RECT 147.715 69.130 148.645 69.140 ;
        RECT 147.720 69.120 148.645 69.130 ;
        RECT 147.725 69.115 148.645 69.120 ;
        RECT 147.735 69.100 148.645 69.115 ;
        RECT 147.740 69.085 148.645 69.100 ;
        RECT 147.750 69.060 148.645 69.085 ;
        RECT 147.255 68.590 147.585 69.015 ;
        RECT 146.515 68.055 146.775 68.535 ;
        RECT 146.945 67.885 147.195 68.425 ;
        RECT 147.365 68.105 147.585 68.590 ;
        RECT 147.755 68.990 148.645 69.060 ;
        RECT 147.755 68.265 147.925 68.990 ;
        RECT 148.095 68.435 148.645 68.820 ;
        RECT 148.850 68.625 149.165 69.645 ;
        RECT 149.555 69.635 149.885 70.435 ;
        RECT 150.370 69.465 150.760 69.640 ;
        RECT 149.335 69.295 150.760 69.465 ;
        RECT 151.115 69.295 151.395 70.435 ;
        RECT 149.335 68.795 149.505 69.295 ;
        RECT 147.755 68.095 148.645 68.265 ;
        RECT 148.850 68.055 149.465 68.625 ;
        RECT 149.755 68.565 150.020 69.125 ;
        RECT 150.190 68.395 150.360 69.295 ;
        RECT 151.565 69.285 151.895 70.265 ;
        RECT 152.065 69.295 152.325 70.435 ;
        RECT 152.495 69.345 155.085 70.435 ;
        RECT 150.530 68.565 150.885 69.125 ;
        RECT 151.125 68.855 151.460 69.125 ;
        RECT 151.630 68.685 151.800 69.285 ;
        RECT 151.970 68.875 152.305 69.125 ;
        RECT 149.635 67.885 149.850 68.395 ;
        RECT 150.080 68.065 150.360 68.395 ;
        RECT 150.540 67.885 150.780 68.395 ;
        RECT 151.115 67.885 151.425 68.685 ;
        RECT 151.630 68.055 152.325 68.685 ;
        RECT 152.495 68.655 153.705 69.175 ;
        RECT 153.875 68.825 155.085 69.345 ;
        RECT 155.715 69.345 156.925 70.435 ;
        RECT 155.715 68.805 156.235 69.345 ;
        RECT 152.495 67.885 155.085 68.655 ;
        RECT 156.405 68.635 156.925 69.175 ;
        RECT 155.715 67.885 156.925 68.635 ;
        RECT 22.690 67.715 157.010 67.885 ;
        RECT 22.775 66.965 23.985 67.715 ;
        RECT 24.155 67.170 29.500 67.715 ;
        RECT 22.775 66.425 23.295 66.965 ;
        RECT 23.465 66.255 23.985 66.795 ;
        RECT 25.740 66.340 26.080 67.170 ;
        RECT 29.675 66.945 32.265 67.715 ;
        RECT 22.775 65.165 23.985 66.255 ;
        RECT 27.560 65.600 27.910 66.850 ;
        RECT 29.675 66.425 30.885 66.945 ;
        RECT 32.445 66.905 32.715 67.715 ;
        RECT 32.885 66.905 33.215 67.545 ;
        RECT 33.385 66.905 33.625 67.715 ;
        RECT 33.815 66.945 36.405 67.715 ;
        RECT 31.055 66.255 32.265 66.775 ;
        RECT 32.435 66.475 32.785 66.725 ;
        RECT 32.955 66.305 33.125 66.905 ;
        RECT 33.295 66.475 33.645 66.725 ;
        RECT 33.815 66.425 35.025 66.945 ;
        RECT 37.045 66.905 37.315 67.715 ;
        RECT 37.485 66.905 37.815 67.545 ;
        RECT 37.985 66.905 38.225 67.715 ;
        RECT 38.415 66.945 40.085 67.715 ;
        RECT 40.435 67.055 40.775 67.715 ;
        RECT 24.155 65.165 29.500 65.600 ;
        RECT 29.675 65.165 32.265 66.255 ;
        RECT 32.445 65.165 32.775 66.305 ;
        RECT 32.955 66.135 33.635 66.305 ;
        RECT 35.195 66.255 36.405 66.775 ;
        RECT 37.035 66.475 37.385 66.725 ;
        RECT 37.555 66.305 37.725 66.905 ;
        RECT 37.895 66.475 38.245 66.725 ;
        RECT 38.415 66.425 39.165 66.945 ;
        RECT 33.305 65.350 33.635 66.135 ;
        RECT 33.815 65.165 36.405 66.255 ;
        RECT 37.045 65.165 37.375 66.305 ;
        RECT 37.555 66.135 38.235 66.305 ;
        RECT 39.335 66.255 40.085 66.775 ;
        RECT 37.905 65.350 38.235 66.135 ;
        RECT 38.415 65.165 40.085 66.255 ;
        RECT 40.255 65.335 40.775 66.885 ;
        RECT 40.945 66.060 41.465 67.545 ;
        RECT 41.645 66.905 41.915 67.715 ;
        RECT 42.085 66.905 42.415 67.545 ;
        RECT 42.585 66.905 42.825 67.715 ;
        RECT 43.025 66.905 43.295 67.715 ;
        RECT 43.465 66.905 43.795 67.545 ;
        RECT 43.965 66.905 44.205 67.715 ;
        RECT 44.875 66.905 45.115 67.715 ;
        RECT 45.285 66.905 45.615 67.545 ;
        RECT 45.785 66.905 46.055 67.715 ;
        RECT 46.705 66.905 46.975 67.715 ;
        RECT 47.145 66.905 47.475 67.545 ;
        RECT 47.645 66.905 47.885 67.715 ;
        RECT 48.535 66.990 48.825 67.715 ;
        RECT 49.160 67.205 49.400 67.715 ;
        RECT 49.580 67.205 49.860 67.535 ;
        RECT 50.090 67.205 50.305 67.715 ;
        RECT 41.635 66.475 41.985 66.725 ;
        RECT 42.155 66.305 42.325 66.905 ;
        RECT 42.495 66.475 42.845 66.725 ;
        RECT 43.015 66.475 43.365 66.725 ;
        RECT 43.535 66.305 43.705 66.905 ;
        RECT 43.875 66.475 44.225 66.725 ;
        RECT 44.855 66.475 45.205 66.725 ;
        RECT 45.375 66.305 45.545 66.905 ;
        RECT 45.715 66.475 46.065 66.725 ;
        RECT 46.695 66.475 47.045 66.725 ;
        RECT 47.215 66.305 47.385 66.905 ;
        RECT 47.555 66.475 47.905 66.725 ;
        RECT 49.055 66.475 49.410 67.035 ;
        RECT 40.945 65.165 41.275 65.890 ;
        RECT 41.645 65.165 41.975 66.305 ;
        RECT 42.155 66.135 42.835 66.305 ;
        RECT 42.505 65.350 42.835 66.135 ;
        RECT 43.025 65.165 43.355 66.305 ;
        RECT 43.535 66.135 44.215 66.305 ;
        RECT 43.885 65.350 44.215 66.135 ;
        RECT 44.865 66.135 45.545 66.305 ;
        RECT 44.865 65.350 45.195 66.135 ;
        RECT 45.725 65.165 46.055 66.305 ;
        RECT 46.705 65.165 47.035 66.305 ;
        RECT 47.215 66.135 47.895 66.305 ;
        RECT 47.565 65.350 47.895 66.135 ;
        RECT 48.535 65.165 48.825 66.330 ;
        RECT 49.580 66.305 49.750 67.205 ;
        RECT 49.920 66.475 50.185 67.035 ;
        RECT 50.475 66.975 51.090 67.545 ;
        RECT 50.435 66.305 50.605 66.805 ;
        RECT 49.180 66.135 50.605 66.305 ;
        RECT 49.180 65.960 49.570 66.135 ;
        RECT 50.055 65.165 50.385 65.965 ;
        RECT 50.775 65.955 51.090 66.975 ;
        RECT 51.305 66.905 51.575 67.715 ;
        RECT 51.745 66.905 52.075 67.545 ;
        RECT 52.245 66.905 52.485 67.715 ;
        RECT 53.595 66.915 54.290 67.545 ;
        RECT 54.495 66.915 54.805 67.715 ;
        RECT 55.155 67.055 55.495 67.715 ;
        RECT 51.295 66.475 51.645 66.725 ;
        RECT 51.815 66.305 51.985 66.905 ;
        RECT 52.155 66.475 52.505 66.725 ;
        RECT 53.615 66.475 53.950 66.725 ;
        RECT 54.120 66.315 54.290 66.915 ;
        RECT 54.460 66.475 54.795 66.745 ;
        RECT 50.555 65.335 51.090 65.955 ;
        RECT 51.305 65.165 51.635 66.305 ;
        RECT 51.815 66.135 52.495 66.305 ;
        RECT 52.165 65.350 52.495 66.135 ;
        RECT 53.595 65.165 53.855 66.305 ;
        RECT 54.025 65.335 54.355 66.315 ;
        RECT 54.525 65.165 54.805 66.305 ;
        RECT 54.975 65.335 55.495 66.885 ;
        RECT 55.665 66.060 56.185 67.545 ;
        RECT 56.355 67.170 61.700 67.715 ;
        RECT 57.940 66.340 58.280 67.170 ;
        RECT 61.875 66.965 63.085 67.715 ;
        RECT 63.255 67.335 64.145 67.505 ;
        RECT 55.665 65.165 55.995 65.890 ;
        RECT 59.760 65.600 60.110 66.850 ;
        RECT 61.875 66.425 62.395 66.965 ;
        RECT 62.565 66.255 63.085 66.795 ;
        RECT 63.255 66.780 63.805 67.165 ;
        RECT 63.975 66.610 64.145 67.335 ;
        RECT 56.355 65.165 61.700 65.600 ;
        RECT 61.875 65.165 63.085 66.255 ;
        RECT 63.255 66.540 64.145 66.610 ;
        RECT 64.315 67.010 64.535 67.495 ;
        RECT 64.705 67.175 64.955 67.715 ;
        RECT 65.125 67.065 65.385 67.545 ;
        RECT 64.315 66.585 64.645 67.010 ;
        RECT 63.255 66.515 64.150 66.540 ;
        RECT 63.255 66.500 64.160 66.515 ;
        RECT 63.255 66.485 64.165 66.500 ;
        RECT 63.255 66.480 64.175 66.485 ;
        RECT 63.255 66.470 64.180 66.480 ;
        RECT 63.255 66.460 64.185 66.470 ;
        RECT 63.255 66.455 64.195 66.460 ;
        RECT 63.255 66.445 64.205 66.455 ;
        RECT 63.255 66.440 64.215 66.445 ;
        RECT 63.255 65.990 63.515 66.440 ;
        RECT 63.880 66.435 64.215 66.440 ;
        RECT 63.880 66.430 64.230 66.435 ;
        RECT 63.880 66.420 64.245 66.430 ;
        RECT 63.880 66.415 64.270 66.420 ;
        RECT 64.815 66.415 65.045 66.810 ;
        RECT 63.880 66.410 65.045 66.415 ;
        RECT 63.910 66.375 65.045 66.410 ;
        RECT 63.945 66.350 65.045 66.375 ;
        RECT 63.975 66.320 65.045 66.350 ;
        RECT 63.995 66.290 65.045 66.320 ;
        RECT 64.015 66.260 65.045 66.290 ;
        RECT 64.085 66.250 65.045 66.260 ;
        RECT 64.110 66.240 65.045 66.250 ;
        RECT 64.130 66.225 65.045 66.240 ;
        RECT 64.150 66.210 65.045 66.225 ;
        RECT 64.155 66.200 64.940 66.210 ;
        RECT 64.170 66.165 64.940 66.200 ;
        RECT 63.685 65.845 64.015 66.090 ;
        RECT 64.185 65.915 64.940 66.165 ;
        RECT 65.215 66.035 65.385 67.065 ;
        RECT 65.645 67.165 65.815 67.545 ;
        RECT 65.995 67.335 66.325 67.715 ;
        RECT 65.645 66.995 66.310 67.165 ;
        RECT 66.505 67.040 66.765 67.545 ;
        RECT 65.575 66.445 65.905 66.815 ;
        RECT 66.140 66.740 66.310 66.995 ;
        RECT 66.140 66.410 66.425 66.740 ;
        RECT 66.140 66.265 66.310 66.410 ;
        RECT 63.685 65.820 63.870 65.845 ;
        RECT 63.255 65.720 63.870 65.820 ;
        RECT 63.255 65.165 63.860 65.720 ;
        RECT 64.035 65.335 64.515 65.675 ;
        RECT 64.685 65.165 64.940 65.710 ;
        RECT 65.110 65.335 65.385 66.035 ;
        RECT 65.645 66.095 66.310 66.265 ;
        RECT 66.595 66.240 66.765 67.040 ;
        RECT 66.935 66.945 70.445 67.715 ;
        RECT 66.935 66.425 68.585 66.945 ;
        RECT 68.755 66.255 70.445 66.775 ;
        RECT 65.645 65.335 65.815 66.095 ;
        RECT 65.995 65.165 66.325 65.925 ;
        RECT 66.495 65.335 66.765 66.240 ;
        RECT 66.935 65.165 70.445 66.255 ;
        RECT 70.615 66.060 71.135 67.545 ;
        RECT 71.305 67.055 71.645 67.715 ;
        RECT 71.995 66.945 73.665 67.715 ;
        RECT 74.295 66.990 74.585 67.715 ;
        RECT 74.755 66.945 78.265 67.715 ;
        RECT 70.805 65.165 71.135 65.890 ;
        RECT 71.305 65.335 71.825 66.885 ;
        RECT 71.995 66.425 72.745 66.945 ;
        RECT 72.915 66.255 73.665 66.775 ;
        RECT 74.755 66.425 76.405 66.945 ;
        RECT 78.445 66.905 78.715 67.715 ;
        RECT 78.885 66.905 79.215 67.545 ;
        RECT 79.385 66.905 79.625 67.715 ;
        RECT 79.815 67.040 80.075 67.545 ;
        RECT 80.255 67.335 80.585 67.715 ;
        RECT 80.765 67.165 80.935 67.545 ;
        RECT 71.995 65.165 73.665 66.255 ;
        RECT 74.295 65.165 74.585 66.330 ;
        RECT 76.575 66.255 78.265 66.775 ;
        RECT 78.435 66.475 78.785 66.725 ;
        RECT 78.955 66.305 79.125 66.905 ;
        RECT 79.295 66.475 79.645 66.725 ;
        RECT 74.755 65.165 78.265 66.255 ;
        RECT 78.445 65.165 78.775 66.305 ;
        RECT 78.955 66.135 79.635 66.305 ;
        RECT 79.305 65.350 79.635 66.135 ;
        RECT 79.815 66.240 79.985 67.040 ;
        RECT 80.270 66.995 80.935 67.165 ;
        RECT 80.270 66.740 80.440 66.995 ;
        RECT 81.195 66.965 82.405 67.715 ;
        RECT 80.155 66.410 80.440 66.740 ;
        RECT 80.675 66.445 81.005 66.815 ;
        RECT 81.195 66.425 81.715 66.965 ;
        RECT 82.585 66.905 82.855 67.715 ;
        RECT 83.025 66.905 83.355 67.545 ;
        RECT 83.525 66.905 83.765 67.715 ;
        RECT 83.975 66.905 84.215 67.715 ;
        RECT 84.385 66.905 84.715 67.545 ;
        RECT 84.885 66.905 85.155 67.715 ;
        RECT 85.335 66.945 87.925 67.715 ;
        RECT 80.270 66.265 80.440 66.410 ;
        RECT 79.815 65.335 80.085 66.240 ;
        RECT 80.270 66.095 80.935 66.265 ;
        RECT 81.885 66.255 82.405 66.795 ;
        RECT 82.575 66.475 82.925 66.725 ;
        RECT 83.095 66.305 83.265 66.905 ;
        RECT 83.435 66.475 83.785 66.725 ;
        RECT 83.955 66.475 84.305 66.725 ;
        RECT 84.475 66.305 84.645 66.905 ;
        RECT 84.815 66.475 85.165 66.725 ;
        RECT 85.335 66.425 86.545 66.945 ;
        RECT 88.105 66.905 88.375 67.715 ;
        RECT 88.545 66.905 88.875 67.545 ;
        RECT 89.045 66.905 89.285 67.715 ;
        RECT 89.475 66.945 91.145 67.715 ;
        RECT 80.255 65.165 80.585 65.925 ;
        RECT 80.765 65.335 80.935 66.095 ;
        RECT 81.195 65.165 82.405 66.255 ;
        RECT 82.585 65.165 82.915 66.305 ;
        RECT 83.095 66.135 83.775 66.305 ;
        RECT 83.445 65.350 83.775 66.135 ;
        RECT 83.965 66.135 84.645 66.305 ;
        RECT 83.965 65.350 84.295 66.135 ;
        RECT 84.825 65.165 85.155 66.305 ;
        RECT 86.715 66.255 87.925 66.775 ;
        RECT 88.095 66.475 88.445 66.725 ;
        RECT 88.615 66.305 88.785 66.905 ;
        RECT 88.955 66.475 89.305 66.725 ;
        RECT 89.475 66.425 90.225 66.945 ;
        RECT 91.335 66.905 91.575 67.715 ;
        RECT 91.745 66.905 92.075 67.545 ;
        RECT 92.245 66.905 92.515 67.715 ;
        RECT 92.705 66.905 92.975 67.715 ;
        RECT 93.145 66.905 93.475 67.545 ;
        RECT 93.645 66.905 93.885 67.715 ;
        RECT 94.700 67.205 94.940 67.715 ;
        RECT 95.120 67.205 95.400 67.535 ;
        RECT 95.630 67.205 95.845 67.715 ;
        RECT 85.335 65.165 87.925 66.255 ;
        RECT 88.105 65.165 88.435 66.305 ;
        RECT 88.615 66.135 89.295 66.305 ;
        RECT 90.395 66.255 91.145 66.775 ;
        RECT 91.315 66.475 91.665 66.725 ;
        RECT 91.835 66.305 92.005 66.905 ;
        RECT 92.175 66.475 92.525 66.725 ;
        RECT 92.695 66.475 93.045 66.725 ;
        RECT 93.215 66.305 93.385 66.905 ;
        RECT 93.555 66.475 93.905 66.725 ;
        RECT 94.595 66.475 94.950 67.035 ;
        RECT 95.120 66.305 95.290 67.205 ;
        RECT 95.460 66.475 95.725 67.035 ;
        RECT 96.015 66.975 96.630 67.545 ;
        RECT 95.975 66.305 96.145 66.805 ;
        RECT 88.965 65.350 89.295 66.135 ;
        RECT 89.475 65.165 91.145 66.255 ;
        RECT 91.325 66.135 92.005 66.305 ;
        RECT 91.325 65.350 91.655 66.135 ;
        RECT 92.185 65.165 92.515 66.305 ;
        RECT 92.705 65.165 93.035 66.305 ;
        RECT 93.215 66.135 93.895 66.305 ;
        RECT 93.565 65.350 93.895 66.135 ;
        RECT 94.720 66.135 96.145 66.305 ;
        RECT 94.720 65.960 95.110 66.135 ;
        RECT 95.595 65.165 95.925 65.965 ;
        RECT 96.315 65.955 96.630 66.975 ;
        RECT 96.835 66.945 99.425 67.715 ;
        RECT 100.055 66.990 100.345 67.715 ;
        RECT 101.155 67.055 101.495 67.715 ;
        RECT 96.835 66.425 98.045 66.945 ;
        RECT 98.215 66.255 99.425 66.775 ;
        RECT 96.095 65.335 96.630 65.955 ;
        RECT 96.835 65.165 99.425 66.255 ;
        RECT 100.055 65.165 100.345 66.330 ;
        RECT 100.975 65.335 101.495 66.885 ;
        RECT 101.665 66.060 102.185 67.545 ;
        RECT 102.355 66.945 104.025 67.715 ;
        RECT 104.285 67.165 104.455 67.455 ;
        RECT 104.625 67.335 104.955 67.715 ;
        RECT 104.285 66.995 104.950 67.165 ;
        RECT 102.355 66.425 103.105 66.945 ;
        RECT 103.275 66.255 104.025 66.775 ;
        RECT 101.665 65.165 101.995 65.890 ;
        RECT 102.355 65.165 104.025 66.255 ;
        RECT 104.200 66.175 104.550 66.825 ;
        RECT 104.720 66.005 104.950 66.995 ;
        RECT 104.285 65.835 104.950 66.005 ;
        RECT 104.285 65.335 104.455 65.835 ;
        RECT 104.625 65.165 104.955 65.665 ;
        RECT 105.125 65.335 105.310 67.455 ;
        RECT 105.565 67.255 105.815 67.715 ;
        RECT 105.985 67.265 106.320 67.435 ;
        RECT 106.515 67.265 107.190 67.435 ;
        RECT 105.985 67.125 106.155 67.265 ;
        RECT 105.480 66.135 105.760 67.085 ;
        RECT 105.930 66.995 106.155 67.125 ;
        RECT 105.930 65.890 106.100 66.995 ;
        RECT 106.325 66.845 106.850 67.065 ;
        RECT 106.270 66.080 106.510 66.675 ;
        RECT 106.680 66.145 106.850 66.845 ;
        RECT 107.020 66.485 107.190 67.265 ;
        RECT 107.510 67.215 107.880 67.715 ;
        RECT 108.060 67.265 108.465 67.435 ;
        RECT 108.635 67.265 109.420 67.435 ;
        RECT 108.060 67.035 108.230 67.265 ;
        RECT 107.400 66.735 108.230 67.035 ;
        RECT 108.615 66.765 109.080 67.095 ;
        RECT 107.400 66.705 107.600 66.735 ;
        RECT 107.720 66.485 107.890 66.555 ;
        RECT 107.020 66.315 107.890 66.485 ;
        RECT 107.380 66.225 107.890 66.315 ;
        RECT 105.930 65.760 106.235 65.890 ;
        RECT 106.680 65.780 107.210 66.145 ;
        RECT 105.550 65.165 105.815 65.625 ;
        RECT 105.985 65.335 106.235 65.760 ;
        RECT 107.380 65.610 107.550 66.225 ;
        RECT 106.445 65.440 107.550 65.610 ;
        RECT 107.720 65.165 107.890 65.965 ;
        RECT 108.060 65.665 108.230 66.735 ;
        RECT 108.400 65.835 108.590 66.555 ;
        RECT 108.760 65.805 109.080 66.765 ;
        RECT 109.250 66.805 109.420 67.265 ;
        RECT 109.695 67.185 109.905 67.715 ;
        RECT 110.165 66.975 110.495 67.500 ;
        RECT 110.665 67.105 110.835 67.715 ;
        RECT 111.005 67.060 111.335 67.495 ;
        RECT 111.720 67.205 111.960 67.715 ;
        RECT 112.140 67.205 112.420 67.535 ;
        RECT 112.650 67.205 112.865 67.715 ;
        RECT 111.005 66.975 111.385 67.060 ;
        RECT 110.295 66.805 110.495 66.975 ;
        RECT 111.160 66.935 111.385 66.975 ;
        RECT 109.250 66.475 110.125 66.805 ;
        RECT 110.295 66.475 111.045 66.805 ;
        RECT 108.060 65.335 108.310 65.665 ;
        RECT 109.250 65.635 109.420 66.475 ;
        RECT 110.295 66.270 110.485 66.475 ;
        RECT 111.215 66.355 111.385 66.935 ;
        RECT 111.615 66.475 111.970 67.035 ;
        RECT 111.170 66.305 111.385 66.355 ;
        RECT 112.140 66.305 112.310 67.205 ;
        RECT 112.480 66.475 112.745 67.035 ;
        RECT 113.035 66.975 113.650 67.545 ;
        RECT 113.855 67.170 119.200 67.715 ;
        RECT 112.995 66.305 113.165 66.805 ;
        RECT 109.590 65.895 110.485 66.270 ;
        RECT 110.995 66.225 111.385 66.305 ;
        RECT 108.535 65.465 109.420 65.635 ;
        RECT 109.600 65.165 109.915 65.665 ;
        RECT 110.145 65.335 110.485 65.895 ;
        RECT 110.655 65.165 110.825 66.175 ;
        RECT 110.995 65.380 111.325 66.225 ;
        RECT 111.740 66.135 113.165 66.305 ;
        RECT 111.740 65.960 112.130 66.135 ;
        RECT 112.615 65.165 112.945 65.965 ;
        RECT 113.335 65.955 113.650 66.975 ;
        RECT 115.440 66.340 115.780 67.170 ;
        RECT 119.375 66.945 121.045 67.715 ;
        RECT 121.305 67.165 121.475 67.545 ;
        RECT 121.655 67.335 121.985 67.715 ;
        RECT 121.305 66.995 121.970 67.165 ;
        RECT 122.165 67.040 122.425 67.545 ;
        RECT 113.115 65.335 113.650 65.955 ;
        RECT 117.260 65.600 117.610 66.850 ;
        RECT 119.375 66.425 120.125 66.945 ;
        RECT 120.295 66.255 121.045 66.775 ;
        RECT 121.235 66.445 121.565 66.815 ;
        RECT 121.800 66.740 121.970 66.995 ;
        RECT 121.800 66.410 122.085 66.740 ;
        RECT 121.800 66.265 121.970 66.410 ;
        RECT 113.855 65.165 119.200 65.600 ;
        RECT 119.375 65.165 121.045 66.255 ;
        RECT 121.305 66.095 121.970 66.265 ;
        RECT 122.255 66.240 122.425 67.040 ;
        RECT 122.615 66.905 122.855 67.715 ;
        RECT 123.025 66.905 123.355 67.545 ;
        RECT 123.525 66.905 123.795 67.715 ;
        RECT 123.985 66.905 124.255 67.715 ;
        RECT 124.425 66.905 124.755 67.545 ;
        RECT 124.925 66.905 125.165 67.715 ;
        RECT 125.815 66.990 126.105 67.715 ;
        RECT 126.295 66.905 126.535 67.715 ;
        RECT 126.705 66.905 127.035 67.545 ;
        RECT 127.205 66.905 127.475 67.715 ;
        RECT 127.655 66.945 130.245 67.715 ;
        RECT 122.595 66.475 122.945 66.725 ;
        RECT 123.115 66.305 123.285 66.905 ;
        RECT 123.455 66.475 123.805 66.725 ;
        RECT 123.975 66.475 124.325 66.725 ;
        RECT 124.495 66.305 124.665 66.905 ;
        RECT 124.835 66.475 125.185 66.725 ;
        RECT 126.275 66.475 126.625 66.725 ;
        RECT 121.305 65.335 121.475 66.095 ;
        RECT 121.655 65.165 121.985 65.925 ;
        RECT 122.155 65.335 122.425 66.240 ;
        RECT 122.605 66.135 123.285 66.305 ;
        RECT 122.605 65.350 122.935 66.135 ;
        RECT 123.465 65.165 123.795 66.305 ;
        RECT 123.985 65.165 124.315 66.305 ;
        RECT 124.495 66.135 125.175 66.305 ;
        RECT 124.845 65.350 125.175 66.135 ;
        RECT 125.815 65.165 126.105 66.330 ;
        RECT 126.795 66.305 126.965 66.905 ;
        RECT 127.135 66.475 127.485 66.725 ;
        RECT 127.655 66.425 128.865 66.945 ;
        RECT 130.435 66.905 130.675 67.715 ;
        RECT 130.845 66.905 131.175 67.545 ;
        RECT 131.345 66.905 131.615 67.715 ;
        RECT 131.805 66.905 132.075 67.715 ;
        RECT 132.245 66.905 132.575 67.545 ;
        RECT 132.745 66.905 132.985 67.715 ;
        RECT 134.260 67.205 134.500 67.715 ;
        RECT 134.680 67.205 134.960 67.535 ;
        RECT 135.190 67.205 135.405 67.715 ;
        RECT 126.285 66.135 126.965 66.305 ;
        RECT 126.285 65.350 126.615 66.135 ;
        RECT 127.145 65.165 127.475 66.305 ;
        RECT 129.035 66.255 130.245 66.775 ;
        RECT 130.415 66.475 130.765 66.725 ;
        RECT 130.935 66.305 131.105 66.905 ;
        RECT 131.275 66.475 131.625 66.725 ;
        RECT 131.795 66.475 132.145 66.725 ;
        RECT 132.315 66.305 132.485 66.905 ;
        RECT 132.655 66.475 133.005 66.725 ;
        RECT 134.155 66.475 134.510 67.035 ;
        RECT 134.680 66.305 134.850 67.205 ;
        RECT 135.020 66.475 135.285 67.035 ;
        RECT 135.575 66.975 136.190 67.545 ;
        RECT 136.485 67.165 136.655 67.455 ;
        RECT 136.825 67.335 137.155 67.715 ;
        RECT 136.485 66.995 137.090 67.165 ;
        RECT 135.535 66.305 135.705 66.805 ;
        RECT 127.655 65.165 130.245 66.255 ;
        RECT 130.425 66.135 131.105 66.305 ;
        RECT 130.425 65.350 130.755 66.135 ;
        RECT 131.285 65.165 131.615 66.305 ;
        RECT 131.805 65.165 132.135 66.305 ;
        RECT 132.315 66.135 132.995 66.305 ;
        RECT 132.665 65.350 132.995 66.135 ;
        RECT 134.280 66.135 135.705 66.305 ;
        RECT 134.280 65.960 134.670 66.135 ;
        RECT 135.155 65.165 135.485 65.965 ;
        RECT 135.875 65.955 136.190 66.975 ;
        RECT 136.395 66.175 136.640 66.815 ;
        RECT 136.920 66.730 137.090 66.995 ;
        RECT 136.920 66.400 137.150 66.730 ;
        RECT 136.920 66.005 137.090 66.400 ;
        RECT 135.655 65.335 136.190 65.955 ;
        RECT 136.485 65.835 137.090 66.005 ;
        RECT 137.325 66.115 137.495 67.455 ;
        RECT 137.865 67.185 138.035 67.455 ;
        RECT 138.205 67.355 138.535 67.715 ;
        RECT 139.170 67.265 139.830 67.435 ;
        RECT 137.865 67.035 138.470 67.185 ;
        RECT 137.865 67.015 138.670 67.035 ;
        RECT 137.790 66.475 138.120 66.845 ;
        RECT 138.300 66.705 138.670 67.015 ;
        RECT 139.045 66.765 139.425 67.095 ;
        RECT 138.300 66.305 138.470 66.705 ;
        RECT 137.785 66.135 138.470 66.305 ;
        RECT 136.485 65.335 136.655 65.835 ;
        RECT 136.825 65.165 137.155 65.665 ;
        RECT 137.325 65.335 137.550 66.115 ;
        RECT 137.785 65.385 138.115 66.135 ;
        RECT 138.285 65.165 138.600 65.965 ;
        RECT 138.800 65.795 139.085 66.445 ;
        RECT 139.255 66.385 139.425 66.765 ;
        RECT 139.660 66.805 139.830 67.265 ;
        RECT 140.070 66.975 140.400 67.715 ;
        RECT 140.670 66.975 140.890 67.385 ;
        RECT 141.070 66.975 141.355 67.715 ;
        RECT 141.525 67.115 141.775 67.385 ;
        RECT 141.945 67.250 142.205 67.715 ;
        RECT 142.465 67.165 142.635 67.455 ;
        RECT 142.805 67.335 143.135 67.715 ;
        RECT 141.525 66.975 141.810 67.115 ;
        RECT 142.465 66.995 143.130 67.165 ;
        RECT 140.720 66.805 140.890 66.975 ;
        RECT 141.640 66.805 141.810 66.975 ;
        RECT 139.660 66.635 140.530 66.805 ;
        RECT 139.810 66.475 140.530 66.635 ;
        RECT 140.720 66.475 141.470 66.805 ;
        RECT 141.640 66.475 142.205 66.805 ;
        RECT 139.255 65.805 139.595 66.385 ;
        RECT 139.810 65.545 139.980 66.475 ;
        RECT 140.720 66.265 140.890 66.475 ;
        RECT 141.640 66.305 141.810 66.475 ;
        RECT 140.170 65.935 140.890 66.265 ;
        RECT 139.230 65.375 139.980 65.545 ;
        RECT 140.150 65.165 140.450 65.665 ;
        RECT 140.670 65.365 140.890 65.935 ;
        RECT 141.070 65.165 141.355 66.305 ;
        RECT 141.525 66.160 141.810 66.305 ;
        RECT 142.380 66.175 142.730 66.825 ;
        RECT 141.525 65.345 141.775 66.160 ;
        RECT 141.945 65.165 142.205 66.045 ;
        RECT 142.900 66.005 143.130 66.995 ;
        RECT 142.465 65.835 143.130 66.005 ;
        RECT 142.465 65.335 142.635 65.835 ;
        RECT 142.805 65.165 143.135 65.665 ;
        RECT 143.305 65.335 143.490 67.455 ;
        RECT 143.745 67.255 143.995 67.715 ;
        RECT 144.165 67.265 144.500 67.435 ;
        RECT 144.695 67.265 145.370 67.435 ;
        RECT 144.165 67.125 144.335 67.265 ;
        RECT 143.660 66.135 143.940 67.085 ;
        RECT 144.110 66.995 144.335 67.125 ;
        RECT 144.110 65.890 144.280 66.995 ;
        RECT 144.505 66.845 145.030 67.065 ;
        RECT 144.450 66.080 144.690 66.675 ;
        RECT 144.860 66.145 145.030 66.845 ;
        RECT 145.200 66.485 145.370 67.265 ;
        RECT 145.690 67.215 146.060 67.715 ;
        RECT 146.240 67.265 146.645 67.435 ;
        RECT 146.815 67.265 147.600 67.435 ;
        RECT 146.240 67.035 146.410 67.265 ;
        RECT 145.580 66.735 146.410 67.035 ;
        RECT 146.795 66.765 147.260 67.095 ;
        RECT 145.580 66.705 145.780 66.735 ;
        RECT 145.900 66.485 146.070 66.555 ;
        RECT 145.200 66.315 146.070 66.485 ;
        RECT 145.560 66.225 146.070 66.315 ;
        RECT 144.110 65.760 144.415 65.890 ;
        RECT 144.860 65.780 145.390 66.145 ;
        RECT 143.730 65.165 143.995 65.625 ;
        RECT 144.165 65.335 144.415 65.760 ;
        RECT 145.560 65.610 145.730 66.225 ;
        RECT 144.625 65.440 145.730 65.610 ;
        RECT 145.900 65.165 146.070 65.965 ;
        RECT 146.240 65.665 146.410 66.735 ;
        RECT 146.580 65.835 146.770 66.555 ;
        RECT 146.940 65.805 147.260 66.765 ;
        RECT 147.430 66.805 147.600 67.265 ;
        RECT 147.875 67.185 148.085 67.715 ;
        RECT 148.345 66.975 148.675 67.500 ;
        RECT 148.845 67.105 149.015 67.715 ;
        RECT 149.185 67.060 149.515 67.495 ;
        RECT 149.185 66.975 149.565 67.060 ;
        RECT 148.475 66.805 148.675 66.975 ;
        RECT 149.340 66.935 149.565 66.975 ;
        RECT 147.430 66.475 148.305 66.805 ;
        RECT 148.475 66.475 149.225 66.805 ;
        RECT 146.240 65.335 146.490 65.665 ;
        RECT 147.430 65.635 147.600 66.475 ;
        RECT 148.475 66.270 148.665 66.475 ;
        RECT 149.395 66.355 149.565 66.935 ;
        RECT 149.735 66.945 151.405 67.715 ;
        RECT 151.575 66.990 151.865 67.715 ;
        RECT 152.035 66.945 155.545 67.715 ;
        RECT 155.715 66.965 156.925 67.715 ;
        RECT 149.735 66.425 150.485 66.945 ;
        RECT 149.350 66.305 149.565 66.355 ;
        RECT 147.770 65.895 148.665 66.270 ;
        RECT 149.175 66.225 149.565 66.305 ;
        RECT 150.655 66.255 151.405 66.775 ;
        RECT 152.035 66.425 153.685 66.945 ;
        RECT 146.715 65.465 147.600 65.635 ;
        RECT 147.780 65.165 148.095 65.665 ;
        RECT 148.325 65.335 148.665 65.895 ;
        RECT 148.835 65.165 149.005 66.175 ;
        RECT 149.175 65.380 149.505 66.225 ;
        RECT 149.735 65.165 151.405 66.255 ;
        RECT 151.575 65.165 151.865 66.330 ;
        RECT 153.855 66.255 155.545 66.775 ;
        RECT 152.035 65.165 155.545 66.255 ;
        RECT 155.715 66.255 156.235 66.795 ;
        RECT 156.405 66.425 156.925 66.965 ;
        RECT 155.715 65.165 156.925 66.255 ;
        RECT 22.690 64.995 157.010 65.165 ;
        RECT 22.775 63.905 23.985 64.995 ;
        RECT 22.775 63.195 23.295 63.735 ;
        RECT 23.465 63.365 23.985 63.905 ;
        RECT 24.615 63.275 25.135 64.825 ;
        RECT 25.305 64.270 25.635 64.995 ;
        RECT 22.775 62.445 23.985 63.195 ;
        RECT 24.795 62.445 25.135 63.105 ;
        RECT 25.305 62.615 25.825 64.100 ;
        RECT 26.455 63.275 26.975 64.825 ;
        RECT 27.145 64.270 27.475 64.995 ;
        RECT 28.025 64.270 28.355 64.995 ;
        RECT 26.635 62.445 26.975 63.105 ;
        RECT 27.145 62.615 27.665 64.100 ;
        RECT 27.835 62.615 28.355 64.100 ;
        RECT 28.525 63.275 29.045 64.825 ;
        RECT 29.305 64.325 29.475 64.825 ;
        RECT 29.645 64.495 29.975 64.995 ;
        RECT 29.305 64.155 29.910 64.325 ;
        RECT 29.215 63.345 29.460 63.985 ;
        RECT 29.740 63.760 29.910 64.155 ;
        RECT 30.145 64.045 30.370 64.825 ;
        RECT 29.740 63.430 29.970 63.760 ;
        RECT 29.740 63.165 29.910 63.430 ;
        RECT 28.525 62.445 28.865 63.105 ;
        RECT 29.305 62.995 29.910 63.165 ;
        RECT 29.305 62.705 29.475 62.995 ;
        RECT 29.645 62.445 29.975 62.825 ;
        RECT 30.145 62.705 30.315 64.045 ;
        RECT 30.605 64.025 30.935 64.775 ;
        RECT 31.105 64.195 31.420 64.995 ;
        RECT 32.050 64.615 32.800 64.785 ;
        RECT 30.605 63.855 31.290 64.025 ;
        RECT 30.610 63.315 30.940 63.685 ;
        RECT 31.120 63.455 31.290 63.855 ;
        RECT 31.620 63.715 31.905 64.365 ;
        RECT 32.075 63.775 32.415 64.355 ;
        RECT 31.120 63.145 31.490 63.455 ;
        RECT 32.075 63.395 32.245 63.775 ;
        RECT 32.630 63.685 32.800 64.615 ;
        RECT 32.970 64.495 33.270 64.995 ;
        RECT 33.490 64.225 33.710 64.795 ;
        RECT 32.990 63.895 33.710 64.225 ;
        RECT 33.540 63.685 33.710 63.895 ;
        RECT 33.890 63.855 34.175 64.995 ;
        RECT 34.345 64.000 34.595 64.815 ;
        RECT 34.765 64.115 35.025 64.995 ;
        RECT 34.345 63.855 34.630 64.000 ;
        RECT 34.460 63.685 34.630 63.855 ;
        RECT 35.655 63.830 35.945 64.995 ;
        RECT 32.630 63.525 33.350 63.685 ;
        RECT 30.685 63.125 31.490 63.145 ;
        RECT 30.685 62.975 31.290 63.125 ;
        RECT 31.865 63.065 32.245 63.395 ;
        RECT 32.480 63.355 33.350 63.525 ;
        RECT 33.540 63.355 34.290 63.685 ;
        RECT 34.460 63.355 35.025 63.685 ;
        RECT 30.685 62.705 30.855 62.975 ;
        RECT 32.480 62.895 32.650 63.355 ;
        RECT 33.540 63.185 33.710 63.355 ;
        RECT 34.460 63.185 34.630 63.355 ;
        RECT 36.115 63.275 36.635 64.825 ;
        RECT 36.805 64.270 37.135 64.995 ;
        RECT 31.025 62.445 31.355 62.805 ;
        RECT 31.990 62.725 32.650 62.895 ;
        RECT 32.890 62.445 33.220 63.185 ;
        RECT 33.490 62.775 33.710 63.185 ;
        RECT 33.890 62.445 34.175 63.185 ;
        RECT 34.345 63.045 34.630 63.185 ;
        RECT 34.345 62.775 34.595 63.045 ;
        RECT 34.765 62.445 35.025 62.910 ;
        RECT 35.655 62.445 35.945 63.170 ;
        RECT 36.295 62.445 36.635 63.105 ;
        RECT 36.805 62.615 37.325 64.100 ;
        RECT 37.495 63.920 37.765 64.825 ;
        RECT 37.935 64.235 38.265 64.995 ;
        RECT 38.445 64.065 38.615 64.825 ;
        RECT 39.065 64.270 39.395 64.995 ;
        RECT 37.495 63.120 37.665 63.920 ;
        RECT 37.950 63.895 38.615 64.065 ;
        RECT 37.950 63.750 38.120 63.895 ;
        RECT 37.835 63.420 38.120 63.750 ;
        RECT 37.950 63.165 38.120 63.420 ;
        RECT 38.355 63.345 38.685 63.715 ;
        RECT 37.495 62.615 37.755 63.120 ;
        RECT 37.950 62.995 38.615 63.165 ;
        RECT 37.935 62.445 38.265 62.825 ;
        RECT 38.445 62.615 38.615 62.995 ;
        RECT 38.875 62.615 39.395 64.100 ;
        RECT 39.565 63.275 40.085 64.825 ;
        RECT 40.345 64.325 40.515 64.825 ;
        RECT 40.685 64.495 41.015 64.995 ;
        RECT 40.345 64.155 40.950 64.325 ;
        RECT 40.255 63.345 40.500 63.985 ;
        RECT 40.780 63.760 40.950 64.155 ;
        RECT 41.185 64.045 41.410 64.825 ;
        RECT 40.780 63.430 41.010 63.760 ;
        RECT 40.780 63.165 40.950 63.430 ;
        RECT 39.565 62.445 39.905 63.105 ;
        RECT 40.345 62.995 40.950 63.165 ;
        RECT 40.345 62.705 40.515 62.995 ;
        RECT 40.685 62.445 41.015 62.825 ;
        RECT 41.185 62.705 41.355 64.045 ;
        RECT 41.645 64.025 41.975 64.775 ;
        RECT 42.145 64.195 42.460 64.995 ;
        RECT 43.090 64.615 43.840 64.785 ;
        RECT 41.645 63.855 42.330 64.025 ;
        RECT 41.650 63.315 41.980 63.685 ;
        RECT 42.160 63.455 42.330 63.855 ;
        RECT 42.660 63.715 42.945 64.365 ;
        RECT 43.115 63.775 43.455 64.355 ;
        RECT 42.160 63.145 42.530 63.455 ;
        RECT 43.115 63.395 43.285 63.775 ;
        RECT 43.670 63.685 43.840 64.615 ;
        RECT 44.010 64.495 44.310 64.995 ;
        RECT 44.530 64.225 44.750 64.795 ;
        RECT 44.030 63.895 44.750 64.225 ;
        RECT 44.580 63.685 44.750 63.895 ;
        RECT 44.930 63.855 45.215 64.995 ;
        RECT 45.385 64.000 45.635 64.815 ;
        RECT 45.805 64.115 46.065 64.995 ;
        RECT 45.385 63.855 45.670 64.000 ;
        RECT 45.500 63.685 45.670 63.855 ;
        RECT 43.670 63.525 44.390 63.685 ;
        RECT 41.725 63.125 42.530 63.145 ;
        RECT 41.725 62.975 42.330 63.125 ;
        RECT 42.905 63.065 43.285 63.395 ;
        RECT 43.520 63.355 44.390 63.525 ;
        RECT 44.580 63.355 45.330 63.685 ;
        RECT 45.500 63.355 46.065 63.685 ;
        RECT 41.725 62.705 41.895 62.975 ;
        RECT 43.520 62.895 43.690 63.355 ;
        RECT 44.580 63.185 44.750 63.355 ;
        RECT 45.500 63.185 45.670 63.355 ;
        RECT 46.235 63.275 46.755 64.825 ;
        RECT 46.925 64.270 47.255 64.995 ;
        RECT 47.705 64.325 47.875 64.825 ;
        RECT 48.045 64.495 48.375 64.995 ;
        RECT 47.705 64.155 48.310 64.325 ;
        RECT 42.065 62.445 42.395 62.805 ;
        RECT 43.030 62.725 43.690 62.895 ;
        RECT 43.930 62.445 44.260 63.185 ;
        RECT 44.530 62.775 44.750 63.185 ;
        RECT 44.930 62.445 45.215 63.185 ;
        RECT 45.385 63.045 45.670 63.185 ;
        RECT 45.385 62.775 45.635 63.045 ;
        RECT 45.805 62.445 46.065 62.910 ;
        RECT 46.415 62.445 46.755 63.105 ;
        RECT 46.925 62.615 47.445 64.100 ;
        RECT 47.615 63.345 47.860 63.985 ;
        RECT 48.140 63.760 48.310 64.155 ;
        RECT 48.545 64.045 48.770 64.825 ;
        RECT 48.140 63.430 48.370 63.760 ;
        RECT 48.140 63.165 48.310 63.430 ;
        RECT 47.705 62.995 48.310 63.165 ;
        RECT 47.705 62.705 47.875 62.995 ;
        RECT 48.045 62.445 48.375 62.825 ;
        RECT 48.545 62.705 48.715 64.045 ;
        RECT 49.005 64.025 49.335 64.775 ;
        RECT 49.505 64.195 49.820 64.995 ;
        RECT 50.450 64.615 51.200 64.785 ;
        RECT 49.005 63.855 49.690 64.025 ;
        RECT 49.010 63.315 49.340 63.685 ;
        RECT 49.520 63.455 49.690 63.855 ;
        RECT 50.020 63.715 50.305 64.365 ;
        RECT 50.475 63.775 50.815 64.355 ;
        RECT 49.520 63.145 49.890 63.455 ;
        RECT 50.475 63.395 50.645 63.775 ;
        RECT 51.030 63.685 51.200 64.615 ;
        RECT 51.370 64.495 51.670 64.995 ;
        RECT 51.890 64.225 52.110 64.795 ;
        RECT 51.390 63.895 52.110 64.225 ;
        RECT 51.940 63.685 52.110 63.895 ;
        RECT 52.290 63.855 52.575 64.995 ;
        RECT 52.745 64.000 52.995 64.815 ;
        RECT 53.165 64.115 53.425 64.995 ;
        RECT 53.685 64.325 53.855 64.825 ;
        RECT 54.025 64.495 54.355 64.995 ;
        RECT 53.685 64.155 54.290 64.325 ;
        RECT 52.745 63.855 53.030 64.000 ;
        RECT 52.860 63.685 53.030 63.855 ;
        RECT 51.030 63.525 51.750 63.685 ;
        RECT 49.085 63.125 49.890 63.145 ;
        RECT 49.085 62.975 49.690 63.125 ;
        RECT 50.265 63.065 50.645 63.395 ;
        RECT 50.880 63.355 51.750 63.525 ;
        RECT 51.940 63.355 52.690 63.685 ;
        RECT 52.860 63.355 53.425 63.685 ;
        RECT 49.085 62.705 49.255 62.975 ;
        RECT 50.880 62.895 51.050 63.355 ;
        RECT 51.940 63.185 52.110 63.355 ;
        RECT 52.860 63.185 53.030 63.355 ;
        RECT 53.595 63.345 53.840 63.985 ;
        RECT 54.120 63.760 54.290 64.155 ;
        RECT 54.525 64.045 54.750 64.825 ;
        RECT 54.120 63.430 54.350 63.760 ;
        RECT 49.425 62.445 49.755 62.805 ;
        RECT 50.390 62.725 51.050 62.895 ;
        RECT 51.290 62.445 51.620 63.185 ;
        RECT 51.890 62.775 52.110 63.185 ;
        RECT 52.290 62.445 52.575 63.185 ;
        RECT 52.745 63.045 53.030 63.185 ;
        RECT 54.120 63.165 54.290 63.430 ;
        RECT 52.745 62.775 52.995 63.045 ;
        RECT 53.685 62.995 54.290 63.165 ;
        RECT 53.165 62.445 53.425 62.910 ;
        RECT 53.685 62.705 53.855 62.995 ;
        RECT 54.025 62.445 54.355 62.825 ;
        RECT 54.525 62.705 54.695 64.045 ;
        RECT 54.985 64.025 55.315 64.775 ;
        RECT 55.485 64.195 55.800 64.995 ;
        RECT 56.430 64.615 57.180 64.785 ;
        RECT 54.985 63.855 55.670 64.025 ;
        RECT 54.990 63.315 55.320 63.685 ;
        RECT 55.500 63.455 55.670 63.855 ;
        RECT 56.000 63.715 56.285 64.365 ;
        RECT 56.455 63.775 56.795 64.355 ;
        RECT 55.500 63.145 55.870 63.455 ;
        RECT 56.455 63.395 56.625 63.775 ;
        RECT 57.010 63.685 57.180 64.615 ;
        RECT 57.350 64.495 57.650 64.995 ;
        RECT 57.870 64.225 58.090 64.795 ;
        RECT 57.370 63.895 58.090 64.225 ;
        RECT 57.920 63.685 58.090 63.895 ;
        RECT 58.270 63.855 58.555 64.995 ;
        RECT 58.725 64.000 58.975 64.815 ;
        RECT 59.145 64.115 59.405 64.995 ;
        RECT 58.725 63.855 59.010 64.000 ;
        RECT 58.840 63.685 59.010 63.855 ;
        RECT 57.010 63.525 57.730 63.685 ;
        RECT 55.065 63.125 55.870 63.145 ;
        RECT 55.065 62.975 55.670 63.125 ;
        RECT 56.245 63.065 56.625 63.395 ;
        RECT 56.860 63.355 57.730 63.525 ;
        RECT 57.920 63.355 58.670 63.685 ;
        RECT 58.840 63.355 59.405 63.685 ;
        RECT 55.065 62.705 55.235 62.975 ;
        RECT 56.860 62.895 57.030 63.355 ;
        RECT 57.920 63.185 58.090 63.355 ;
        RECT 58.840 63.185 59.010 63.355 ;
        RECT 59.575 63.275 60.095 64.825 ;
        RECT 60.265 64.270 60.595 64.995 ;
        RECT 55.405 62.445 55.735 62.805 ;
        RECT 56.370 62.725 57.030 62.895 ;
        RECT 57.270 62.445 57.600 63.185 ;
        RECT 57.870 62.775 58.090 63.185 ;
        RECT 58.270 62.445 58.555 63.185 ;
        RECT 58.725 63.045 59.010 63.185 ;
        RECT 58.725 62.775 58.975 63.045 ;
        RECT 59.145 62.445 59.405 62.910 ;
        RECT 59.755 62.445 60.095 63.105 ;
        RECT 60.265 62.615 60.785 64.100 ;
        RECT 61.415 63.830 61.705 64.995 ;
        RECT 61.875 63.905 64.465 64.995 ;
        RECT 65.285 64.270 65.615 64.995 ;
        RECT 61.875 63.215 63.085 63.735 ;
        RECT 63.255 63.385 64.465 63.905 ;
        RECT 61.415 62.445 61.705 63.170 ;
        RECT 61.875 62.445 64.465 63.215 ;
        RECT 65.095 62.615 65.615 64.100 ;
        RECT 65.785 63.275 66.305 64.825 ;
        RECT 66.475 64.115 66.735 64.995 ;
        RECT 66.905 64.000 67.155 64.815 ;
        RECT 66.870 63.855 67.155 64.000 ;
        RECT 67.325 63.855 67.610 64.995 ;
        RECT 67.790 64.225 68.010 64.795 ;
        RECT 68.230 64.495 68.530 64.995 ;
        RECT 68.700 64.615 69.450 64.785 ;
        RECT 67.790 63.895 68.510 64.225 ;
        RECT 66.870 63.685 67.040 63.855 ;
        RECT 67.790 63.685 67.960 63.895 ;
        RECT 68.700 63.685 68.870 64.615 ;
        RECT 69.085 63.775 69.425 64.355 ;
        RECT 66.475 63.355 67.040 63.685 ;
        RECT 67.210 63.355 67.960 63.685 ;
        RECT 68.150 63.525 68.870 63.685 ;
        RECT 68.150 63.355 69.020 63.525 ;
        RECT 66.870 63.185 67.040 63.355 ;
        RECT 67.790 63.185 67.960 63.355 ;
        RECT 65.785 62.445 66.125 63.105 ;
        RECT 66.870 63.045 67.155 63.185 ;
        RECT 66.475 62.445 66.735 62.910 ;
        RECT 66.905 62.775 67.155 63.045 ;
        RECT 67.325 62.445 67.610 63.185 ;
        RECT 67.790 62.775 68.010 63.185 ;
        RECT 68.280 62.445 68.610 63.185 ;
        RECT 68.850 62.895 69.020 63.355 ;
        RECT 69.255 63.395 69.425 63.775 ;
        RECT 69.595 63.715 69.880 64.365 ;
        RECT 70.080 64.195 70.395 64.995 ;
        RECT 70.565 64.025 70.895 64.775 ;
        RECT 71.130 64.045 71.355 64.825 ;
        RECT 71.525 64.495 71.855 64.995 ;
        RECT 72.025 64.325 72.195 64.825 ;
        RECT 70.210 63.855 70.895 64.025 ;
        RECT 70.210 63.455 70.380 63.855 ;
        RECT 69.255 63.065 69.635 63.395 ;
        RECT 70.010 63.145 70.380 63.455 ;
        RECT 70.560 63.315 70.890 63.685 ;
        RECT 70.010 63.125 70.815 63.145 ;
        RECT 70.210 62.975 70.815 63.125 ;
        RECT 68.850 62.725 69.510 62.895 ;
        RECT 70.145 62.445 70.475 62.805 ;
        RECT 70.645 62.705 70.815 62.975 ;
        RECT 71.185 62.705 71.355 64.045 ;
        RECT 71.590 64.155 72.195 64.325 ;
        RECT 72.545 64.325 72.715 64.825 ;
        RECT 72.885 64.495 73.215 64.995 ;
        RECT 72.545 64.155 73.150 64.325 ;
        RECT 71.590 63.760 71.760 64.155 ;
        RECT 71.530 63.430 71.760 63.760 ;
        RECT 71.590 63.165 71.760 63.430 ;
        RECT 72.040 63.345 72.285 63.985 ;
        RECT 72.455 63.345 72.700 63.985 ;
        RECT 72.980 63.760 73.150 64.155 ;
        RECT 73.385 64.045 73.610 64.825 ;
        RECT 72.980 63.430 73.210 63.760 ;
        RECT 72.980 63.165 73.150 63.430 ;
        RECT 71.590 62.995 72.195 63.165 ;
        RECT 71.525 62.445 71.855 62.825 ;
        RECT 72.025 62.705 72.195 62.995 ;
        RECT 72.545 62.995 73.150 63.165 ;
        RECT 72.545 62.705 72.715 62.995 ;
        RECT 72.885 62.445 73.215 62.825 ;
        RECT 73.385 62.705 73.555 64.045 ;
        RECT 73.845 64.025 74.175 64.775 ;
        RECT 74.345 64.195 74.660 64.995 ;
        RECT 75.290 64.615 76.040 64.785 ;
        RECT 73.845 63.855 74.530 64.025 ;
        RECT 73.850 63.315 74.180 63.685 ;
        RECT 74.360 63.455 74.530 63.855 ;
        RECT 74.860 63.715 75.145 64.365 ;
        RECT 75.315 63.775 75.655 64.355 ;
        RECT 74.360 63.145 74.730 63.455 ;
        RECT 75.315 63.395 75.485 63.775 ;
        RECT 75.870 63.685 76.040 64.615 ;
        RECT 76.210 64.495 76.510 64.995 ;
        RECT 76.730 64.225 76.950 64.795 ;
        RECT 76.230 63.895 76.950 64.225 ;
        RECT 76.780 63.685 76.950 63.895 ;
        RECT 77.130 63.855 77.415 64.995 ;
        RECT 77.585 64.000 77.835 64.815 ;
        RECT 78.005 64.115 78.265 64.995 ;
        RECT 78.525 64.325 78.695 64.825 ;
        RECT 78.865 64.495 79.195 64.995 ;
        RECT 78.525 64.155 79.130 64.325 ;
        RECT 77.585 63.855 77.870 64.000 ;
        RECT 77.700 63.685 77.870 63.855 ;
        RECT 75.870 63.525 76.590 63.685 ;
        RECT 73.925 63.125 74.730 63.145 ;
        RECT 73.925 62.975 74.530 63.125 ;
        RECT 75.105 63.065 75.485 63.395 ;
        RECT 75.720 63.355 76.590 63.525 ;
        RECT 76.780 63.355 77.530 63.685 ;
        RECT 77.700 63.355 78.265 63.685 ;
        RECT 73.925 62.705 74.095 62.975 ;
        RECT 75.720 62.895 75.890 63.355 ;
        RECT 76.780 63.185 76.950 63.355 ;
        RECT 77.700 63.185 77.870 63.355 ;
        RECT 78.435 63.345 78.680 63.985 ;
        RECT 78.960 63.760 79.130 64.155 ;
        RECT 79.365 64.045 79.590 64.825 ;
        RECT 78.960 63.430 79.190 63.760 ;
        RECT 74.265 62.445 74.595 62.805 ;
        RECT 75.230 62.725 75.890 62.895 ;
        RECT 76.130 62.445 76.460 63.185 ;
        RECT 76.730 62.775 76.950 63.185 ;
        RECT 77.130 62.445 77.415 63.185 ;
        RECT 77.585 63.045 77.870 63.185 ;
        RECT 78.960 63.165 79.130 63.430 ;
        RECT 77.585 62.775 77.835 63.045 ;
        RECT 78.525 62.995 79.130 63.165 ;
        RECT 78.005 62.445 78.265 62.910 ;
        RECT 78.525 62.705 78.695 62.995 ;
        RECT 78.865 62.445 79.195 62.825 ;
        RECT 79.365 62.705 79.535 64.045 ;
        RECT 79.825 64.025 80.155 64.775 ;
        RECT 80.325 64.195 80.640 64.995 ;
        RECT 81.270 64.615 82.020 64.785 ;
        RECT 79.825 63.855 80.510 64.025 ;
        RECT 79.830 63.315 80.160 63.685 ;
        RECT 80.340 63.455 80.510 63.855 ;
        RECT 80.840 63.715 81.125 64.365 ;
        RECT 81.295 63.775 81.635 64.355 ;
        RECT 80.340 63.145 80.710 63.455 ;
        RECT 81.295 63.395 81.465 63.775 ;
        RECT 81.850 63.685 82.020 64.615 ;
        RECT 82.190 64.495 82.490 64.995 ;
        RECT 82.710 64.225 82.930 64.795 ;
        RECT 82.210 63.895 82.930 64.225 ;
        RECT 82.760 63.685 82.930 63.895 ;
        RECT 83.110 63.855 83.395 64.995 ;
        RECT 83.565 64.000 83.815 64.815 ;
        RECT 83.985 64.115 84.245 64.995 ;
        RECT 83.565 63.855 83.850 64.000 ;
        RECT 83.680 63.685 83.850 63.855 ;
        RECT 81.850 63.525 82.570 63.685 ;
        RECT 79.905 63.125 80.710 63.145 ;
        RECT 79.905 62.975 80.510 63.125 ;
        RECT 81.085 63.065 81.465 63.395 ;
        RECT 81.700 63.355 82.570 63.525 ;
        RECT 82.760 63.355 83.510 63.685 ;
        RECT 83.680 63.355 84.245 63.685 ;
        RECT 79.905 62.705 80.075 62.975 ;
        RECT 81.700 62.895 81.870 63.355 ;
        RECT 82.760 63.185 82.930 63.355 ;
        RECT 83.680 63.185 83.850 63.355 ;
        RECT 84.415 63.275 84.935 64.825 ;
        RECT 85.105 64.270 85.435 64.995 ;
        RECT 80.245 62.445 80.575 62.805 ;
        RECT 81.210 62.725 81.870 62.895 ;
        RECT 82.110 62.445 82.440 63.185 ;
        RECT 82.710 62.775 82.930 63.185 ;
        RECT 83.110 62.445 83.395 63.185 ;
        RECT 83.565 63.045 83.850 63.185 ;
        RECT 83.565 62.775 83.815 63.045 ;
        RECT 83.985 62.445 84.245 62.910 ;
        RECT 84.595 62.445 84.935 63.105 ;
        RECT 85.105 62.615 85.625 64.100 ;
        RECT 85.795 63.275 86.315 64.825 ;
        RECT 86.485 64.270 86.815 64.995 ;
        RECT 85.975 62.445 86.315 63.105 ;
        RECT 86.485 62.615 87.005 64.100 ;
        RECT 87.175 63.830 87.465 64.995 ;
        RECT 87.635 63.905 90.225 64.995 ;
        RECT 87.635 63.215 88.845 63.735 ;
        RECT 89.015 63.385 90.225 63.905 ;
        RECT 90.855 63.275 91.375 64.825 ;
        RECT 91.545 64.270 91.875 64.995 ;
        RECT 87.175 62.445 87.465 63.170 ;
        RECT 87.635 62.445 90.225 63.215 ;
        RECT 91.035 62.445 91.375 63.105 ;
        RECT 91.545 62.615 92.065 64.100 ;
        RECT 93.155 63.275 93.675 64.825 ;
        RECT 93.845 64.270 94.175 64.995 ;
        RECT 94.725 64.270 95.055 64.995 ;
        RECT 93.335 62.445 93.675 63.105 ;
        RECT 93.845 62.615 94.365 64.100 ;
        RECT 94.535 62.615 95.055 64.100 ;
        RECT 95.225 63.275 95.745 64.825 ;
        RECT 96.005 64.325 96.175 64.825 ;
        RECT 96.345 64.495 96.675 64.995 ;
        RECT 96.005 64.155 96.610 64.325 ;
        RECT 95.915 63.345 96.160 63.985 ;
        RECT 96.440 63.760 96.610 64.155 ;
        RECT 96.845 64.045 97.070 64.825 ;
        RECT 96.440 63.430 96.670 63.760 ;
        RECT 96.440 63.165 96.610 63.430 ;
        RECT 95.225 62.445 95.565 63.105 ;
        RECT 96.005 62.995 96.610 63.165 ;
        RECT 96.005 62.705 96.175 62.995 ;
        RECT 96.345 62.445 96.675 62.825 ;
        RECT 96.845 62.705 97.015 64.045 ;
        RECT 97.305 64.025 97.635 64.775 ;
        RECT 97.805 64.195 98.120 64.995 ;
        RECT 98.750 64.615 99.500 64.785 ;
        RECT 97.305 63.855 97.990 64.025 ;
        RECT 97.310 63.315 97.640 63.685 ;
        RECT 97.820 63.455 97.990 63.855 ;
        RECT 98.320 63.715 98.605 64.365 ;
        RECT 98.775 63.775 99.115 64.355 ;
        RECT 97.820 63.145 98.190 63.455 ;
        RECT 98.775 63.395 98.945 63.775 ;
        RECT 99.330 63.685 99.500 64.615 ;
        RECT 99.670 64.495 99.970 64.995 ;
        RECT 100.190 64.225 100.410 64.795 ;
        RECT 99.690 63.895 100.410 64.225 ;
        RECT 100.240 63.685 100.410 63.895 ;
        RECT 100.590 63.855 100.875 64.995 ;
        RECT 101.045 64.000 101.295 64.815 ;
        RECT 101.465 64.115 101.725 64.995 ;
        RECT 101.045 63.855 101.330 64.000 ;
        RECT 101.160 63.685 101.330 63.855 ;
        RECT 99.330 63.525 100.050 63.685 ;
        RECT 97.385 63.125 98.190 63.145 ;
        RECT 97.385 62.975 97.990 63.125 ;
        RECT 98.565 63.065 98.945 63.395 ;
        RECT 99.180 63.355 100.050 63.525 ;
        RECT 100.240 63.355 100.990 63.685 ;
        RECT 101.160 63.355 101.725 63.685 ;
        RECT 97.385 62.705 97.555 62.975 ;
        RECT 99.180 62.895 99.350 63.355 ;
        RECT 100.240 63.185 100.410 63.355 ;
        RECT 101.160 63.185 101.330 63.355 ;
        RECT 101.895 63.275 102.415 64.825 ;
        RECT 102.585 64.270 102.915 64.995 ;
        RECT 103.465 64.270 103.795 64.995 ;
        RECT 97.725 62.445 98.055 62.805 ;
        RECT 98.690 62.725 99.350 62.895 ;
        RECT 99.590 62.445 99.920 63.185 ;
        RECT 100.190 62.775 100.410 63.185 ;
        RECT 100.590 62.445 100.875 63.185 ;
        RECT 101.045 63.045 101.330 63.185 ;
        RECT 101.045 62.775 101.295 63.045 ;
        RECT 101.465 62.445 101.725 62.910 ;
        RECT 102.075 62.445 102.415 63.105 ;
        RECT 102.585 62.615 103.105 64.100 ;
        RECT 103.275 62.615 103.795 64.100 ;
        RECT 103.965 63.275 104.485 64.825 ;
        RECT 104.655 63.905 107.245 64.995 ;
        RECT 104.655 63.215 105.865 63.735 ;
        RECT 106.035 63.385 107.245 63.905 ;
        RECT 107.415 63.920 107.685 64.825 ;
        RECT 107.855 64.235 108.185 64.995 ;
        RECT 108.365 64.065 108.535 64.825 ;
        RECT 103.965 62.445 104.305 63.105 ;
        RECT 104.655 62.445 107.245 63.215 ;
        RECT 107.415 63.120 107.585 63.920 ;
        RECT 107.870 63.895 108.535 64.065 ;
        RECT 108.795 63.905 112.305 64.995 ;
        RECT 107.870 63.750 108.040 63.895 ;
        RECT 107.755 63.420 108.040 63.750 ;
        RECT 107.870 63.165 108.040 63.420 ;
        RECT 108.275 63.345 108.605 63.715 ;
        RECT 108.795 63.215 110.445 63.735 ;
        RECT 110.615 63.385 112.305 63.905 ;
        RECT 112.935 63.830 113.225 64.995 ;
        RECT 113.585 64.270 113.915 64.995 ;
        RECT 107.415 62.615 107.675 63.120 ;
        RECT 107.870 62.995 108.535 63.165 ;
        RECT 107.855 62.445 108.185 62.825 ;
        RECT 108.365 62.615 108.535 62.995 ;
        RECT 108.795 62.445 112.305 63.215 ;
        RECT 112.935 62.445 113.225 63.170 ;
        RECT 113.395 62.615 113.915 64.100 ;
        RECT 114.085 63.275 114.605 64.825 ;
        RECT 114.865 64.325 115.035 64.825 ;
        RECT 115.205 64.495 115.535 64.995 ;
        RECT 114.865 64.155 115.470 64.325 ;
        RECT 114.775 63.345 115.020 63.985 ;
        RECT 115.300 63.760 115.470 64.155 ;
        RECT 115.705 64.045 115.930 64.825 ;
        RECT 115.300 63.430 115.530 63.760 ;
        RECT 115.300 63.165 115.470 63.430 ;
        RECT 114.085 62.445 114.425 63.105 ;
        RECT 114.865 62.995 115.470 63.165 ;
        RECT 114.865 62.705 115.035 62.995 ;
        RECT 115.205 62.445 115.535 62.825 ;
        RECT 115.705 62.705 115.875 64.045 ;
        RECT 116.165 64.025 116.495 64.775 ;
        RECT 116.665 64.195 116.980 64.995 ;
        RECT 117.610 64.615 118.360 64.785 ;
        RECT 116.165 63.855 116.850 64.025 ;
        RECT 116.170 63.315 116.500 63.685 ;
        RECT 116.680 63.455 116.850 63.855 ;
        RECT 117.180 63.715 117.465 64.365 ;
        RECT 117.635 63.775 117.975 64.355 ;
        RECT 116.680 63.145 117.050 63.455 ;
        RECT 117.635 63.395 117.805 63.775 ;
        RECT 118.190 63.685 118.360 64.615 ;
        RECT 118.530 64.495 118.830 64.995 ;
        RECT 119.050 64.225 119.270 64.795 ;
        RECT 118.550 63.895 119.270 64.225 ;
        RECT 119.100 63.685 119.270 63.895 ;
        RECT 119.450 63.855 119.735 64.995 ;
        RECT 119.905 64.000 120.155 64.815 ;
        RECT 120.325 64.115 120.585 64.995 ;
        RECT 120.845 64.325 121.015 64.825 ;
        RECT 121.185 64.495 121.515 64.995 ;
        RECT 120.845 64.155 121.450 64.325 ;
        RECT 119.905 63.855 120.190 64.000 ;
        RECT 120.020 63.685 120.190 63.855 ;
        RECT 118.190 63.525 118.910 63.685 ;
        RECT 116.245 63.125 117.050 63.145 ;
        RECT 116.245 62.975 116.850 63.125 ;
        RECT 117.425 63.065 117.805 63.395 ;
        RECT 118.040 63.355 118.910 63.525 ;
        RECT 119.100 63.355 119.850 63.685 ;
        RECT 120.020 63.355 120.585 63.685 ;
        RECT 116.245 62.705 116.415 62.975 ;
        RECT 118.040 62.895 118.210 63.355 ;
        RECT 119.100 63.185 119.270 63.355 ;
        RECT 120.020 63.185 120.190 63.355 ;
        RECT 120.755 63.345 121.000 63.985 ;
        RECT 121.280 63.760 121.450 64.155 ;
        RECT 121.685 64.045 121.910 64.825 ;
        RECT 121.280 63.430 121.510 63.760 ;
        RECT 116.585 62.445 116.915 62.805 ;
        RECT 117.550 62.725 118.210 62.895 ;
        RECT 118.450 62.445 118.780 63.185 ;
        RECT 119.050 62.775 119.270 63.185 ;
        RECT 119.450 62.445 119.735 63.185 ;
        RECT 119.905 63.045 120.190 63.185 ;
        RECT 121.280 63.165 121.450 63.430 ;
        RECT 119.905 62.775 120.155 63.045 ;
        RECT 120.845 62.995 121.450 63.165 ;
        RECT 120.325 62.445 120.585 62.910 ;
        RECT 120.845 62.705 121.015 62.995 ;
        RECT 121.185 62.445 121.515 62.825 ;
        RECT 121.685 62.705 121.855 64.045 ;
        RECT 122.145 64.025 122.475 64.775 ;
        RECT 122.645 64.195 122.960 64.995 ;
        RECT 123.590 64.615 124.340 64.785 ;
        RECT 122.145 63.855 122.830 64.025 ;
        RECT 122.150 63.315 122.480 63.685 ;
        RECT 122.660 63.455 122.830 63.855 ;
        RECT 123.160 63.715 123.445 64.365 ;
        RECT 123.615 63.775 123.955 64.355 ;
        RECT 122.660 63.145 123.030 63.455 ;
        RECT 123.615 63.395 123.785 63.775 ;
        RECT 124.170 63.685 124.340 64.615 ;
        RECT 124.510 64.495 124.810 64.995 ;
        RECT 125.030 64.225 125.250 64.795 ;
        RECT 124.530 63.895 125.250 64.225 ;
        RECT 125.080 63.685 125.250 63.895 ;
        RECT 125.430 63.855 125.715 64.995 ;
        RECT 125.885 64.000 126.135 64.815 ;
        RECT 126.305 64.115 126.565 64.995 ;
        RECT 125.885 63.855 126.170 64.000 ;
        RECT 126.000 63.685 126.170 63.855 ;
        RECT 124.170 63.525 124.890 63.685 ;
        RECT 122.225 63.125 123.030 63.145 ;
        RECT 122.225 62.975 122.830 63.125 ;
        RECT 123.405 63.065 123.785 63.395 ;
        RECT 124.020 63.355 124.890 63.525 ;
        RECT 125.080 63.355 125.830 63.685 ;
        RECT 126.000 63.355 126.565 63.685 ;
        RECT 122.225 62.705 122.395 62.975 ;
        RECT 124.020 62.895 124.190 63.355 ;
        RECT 125.080 63.185 125.250 63.355 ;
        RECT 126.000 63.185 126.170 63.355 ;
        RECT 126.735 63.275 127.255 64.825 ;
        RECT 127.425 64.270 127.755 64.995 ;
        RECT 122.565 62.445 122.895 62.805 ;
        RECT 123.530 62.725 124.190 62.895 ;
        RECT 124.430 62.445 124.760 63.185 ;
        RECT 125.030 62.775 125.250 63.185 ;
        RECT 125.430 62.445 125.715 63.185 ;
        RECT 125.885 63.045 126.170 63.185 ;
        RECT 125.885 62.775 126.135 63.045 ;
        RECT 126.305 62.445 126.565 62.910 ;
        RECT 126.915 62.445 127.255 63.105 ;
        RECT 127.425 62.615 127.945 64.100 ;
        RECT 128.115 63.275 128.635 64.825 ;
        RECT 128.805 64.270 129.135 64.995 ;
        RECT 128.295 62.445 128.635 63.105 ;
        RECT 128.805 62.615 129.325 64.100 ;
        RECT 129.495 63.275 130.015 64.825 ;
        RECT 130.185 64.270 130.515 64.995 ;
        RECT 131.885 64.325 132.055 64.825 ;
        RECT 132.225 64.495 132.555 64.995 ;
        RECT 131.885 64.155 132.490 64.325 ;
        RECT 129.675 62.445 130.015 63.105 ;
        RECT 130.185 62.615 130.705 64.100 ;
        RECT 131.795 63.345 132.040 63.985 ;
        RECT 132.320 63.760 132.490 64.155 ;
        RECT 132.725 64.045 132.950 64.825 ;
        RECT 132.320 63.430 132.550 63.760 ;
        RECT 132.320 63.165 132.490 63.430 ;
        RECT 131.885 62.995 132.490 63.165 ;
        RECT 131.885 62.705 132.055 62.995 ;
        RECT 132.225 62.445 132.555 62.825 ;
        RECT 132.725 62.705 132.895 64.045 ;
        RECT 133.185 64.025 133.515 64.775 ;
        RECT 133.685 64.195 134.000 64.995 ;
        RECT 134.630 64.615 135.380 64.785 ;
        RECT 133.185 63.855 133.870 64.025 ;
        RECT 133.190 63.315 133.520 63.685 ;
        RECT 133.700 63.455 133.870 63.855 ;
        RECT 134.200 63.715 134.485 64.365 ;
        RECT 134.655 63.775 134.995 64.355 ;
        RECT 133.700 63.145 134.070 63.455 ;
        RECT 134.655 63.395 134.825 63.775 ;
        RECT 135.210 63.685 135.380 64.615 ;
        RECT 135.550 64.495 135.850 64.995 ;
        RECT 136.070 64.225 136.290 64.795 ;
        RECT 135.570 63.895 136.290 64.225 ;
        RECT 136.120 63.685 136.290 63.895 ;
        RECT 136.470 63.855 136.755 64.995 ;
        RECT 136.925 64.000 137.175 64.815 ;
        RECT 137.345 64.115 137.605 64.995 ;
        RECT 136.925 63.855 137.210 64.000 ;
        RECT 137.040 63.685 137.210 63.855 ;
        RECT 138.695 63.830 138.985 64.995 ;
        RECT 135.210 63.525 135.930 63.685 ;
        RECT 133.265 63.125 134.070 63.145 ;
        RECT 133.265 62.975 133.870 63.125 ;
        RECT 134.445 63.065 134.825 63.395 ;
        RECT 135.060 63.355 135.930 63.525 ;
        RECT 136.120 63.355 136.870 63.685 ;
        RECT 137.040 63.355 137.605 63.685 ;
        RECT 133.265 62.705 133.435 62.975 ;
        RECT 135.060 62.895 135.230 63.355 ;
        RECT 136.120 63.185 136.290 63.355 ;
        RECT 137.040 63.185 137.210 63.355 ;
        RECT 139.155 63.275 139.675 64.825 ;
        RECT 139.845 64.270 140.175 64.995 ;
        RECT 133.605 62.445 133.935 62.805 ;
        RECT 134.570 62.725 135.230 62.895 ;
        RECT 135.470 62.445 135.800 63.185 ;
        RECT 136.070 62.775 136.290 63.185 ;
        RECT 136.470 62.445 136.755 63.185 ;
        RECT 136.925 63.045 137.210 63.185 ;
        RECT 136.925 62.775 137.175 63.045 ;
        RECT 137.345 62.445 137.605 62.910 ;
        RECT 138.695 62.445 138.985 63.170 ;
        RECT 139.335 62.445 139.675 63.105 ;
        RECT 139.845 62.615 140.365 64.100 ;
        RECT 140.535 63.905 142.205 64.995 ;
        RECT 142.925 64.325 143.095 64.825 ;
        RECT 143.265 64.495 143.595 64.995 ;
        RECT 142.925 64.155 143.530 64.325 ;
        RECT 140.535 63.215 141.285 63.735 ;
        RECT 141.455 63.385 142.205 63.905 ;
        RECT 142.835 63.345 143.080 63.985 ;
        RECT 143.360 63.760 143.530 64.155 ;
        RECT 143.765 64.045 143.990 64.825 ;
        RECT 143.360 63.430 143.590 63.760 ;
        RECT 140.535 62.445 142.205 63.215 ;
        RECT 143.360 63.165 143.530 63.430 ;
        RECT 142.925 62.995 143.530 63.165 ;
        RECT 142.925 62.705 143.095 62.995 ;
        RECT 143.265 62.445 143.595 62.825 ;
        RECT 143.765 62.705 143.935 64.045 ;
        RECT 144.225 64.025 144.555 64.775 ;
        RECT 144.725 64.195 145.040 64.995 ;
        RECT 145.670 64.615 146.420 64.785 ;
        RECT 144.225 63.855 144.910 64.025 ;
        RECT 144.230 63.315 144.560 63.685 ;
        RECT 144.740 63.455 144.910 63.855 ;
        RECT 145.240 63.715 145.525 64.365 ;
        RECT 145.695 63.775 146.035 64.355 ;
        RECT 144.740 63.145 145.110 63.455 ;
        RECT 145.695 63.395 145.865 63.775 ;
        RECT 146.250 63.685 146.420 64.615 ;
        RECT 146.590 64.495 146.890 64.995 ;
        RECT 147.110 64.225 147.330 64.795 ;
        RECT 146.610 63.895 147.330 64.225 ;
        RECT 147.160 63.685 147.330 63.895 ;
        RECT 147.510 63.855 147.795 64.995 ;
        RECT 147.965 64.000 148.215 64.815 ;
        RECT 148.385 64.115 148.645 64.995 ;
        RECT 148.815 64.560 154.160 64.995 ;
        RECT 147.965 63.855 148.250 64.000 ;
        RECT 148.080 63.685 148.250 63.855 ;
        RECT 146.250 63.525 146.970 63.685 ;
        RECT 144.305 63.125 145.110 63.145 ;
        RECT 144.305 62.975 144.910 63.125 ;
        RECT 145.485 63.065 145.865 63.395 ;
        RECT 146.100 63.355 146.970 63.525 ;
        RECT 147.160 63.355 147.910 63.685 ;
        RECT 148.080 63.355 148.645 63.685 ;
        RECT 144.305 62.705 144.475 62.975 ;
        RECT 146.100 62.895 146.270 63.355 ;
        RECT 147.160 63.185 147.330 63.355 ;
        RECT 148.080 63.185 148.250 63.355 ;
        RECT 144.645 62.445 144.975 62.805 ;
        RECT 145.610 62.725 146.270 62.895 ;
        RECT 146.510 62.445 146.840 63.185 ;
        RECT 147.110 62.775 147.330 63.185 ;
        RECT 147.510 62.445 147.795 63.185 ;
        RECT 147.965 63.045 148.250 63.185 ;
        RECT 147.965 62.775 148.215 63.045 ;
        RECT 150.400 62.990 150.740 63.820 ;
        RECT 152.220 63.310 152.570 64.560 ;
        RECT 154.335 63.905 155.545 64.995 ;
        RECT 154.335 63.195 154.855 63.735 ;
        RECT 155.025 63.365 155.545 63.905 ;
        RECT 155.715 63.905 156.925 64.995 ;
        RECT 155.715 63.365 156.235 63.905 ;
        RECT 156.405 63.195 156.925 63.735 ;
        RECT 148.385 62.445 148.645 62.910 ;
        RECT 148.815 62.445 154.160 62.990 ;
        RECT 154.335 62.445 155.545 63.195 ;
        RECT 155.715 62.445 156.925 63.195 ;
        RECT 22.690 62.275 157.010 62.445 ;
        RECT 22.775 61.525 23.985 62.275 ;
        RECT 24.705 61.725 24.875 62.015 ;
        RECT 25.045 61.895 25.375 62.275 ;
        RECT 24.705 61.555 25.310 61.725 ;
        RECT 22.775 60.985 23.295 61.525 ;
        RECT 23.465 60.815 23.985 61.355 ;
        RECT 22.775 59.725 23.985 60.815 ;
        RECT 24.615 60.735 24.860 61.375 ;
        RECT 25.140 61.290 25.310 61.555 ;
        RECT 25.140 60.960 25.370 61.290 ;
        RECT 25.140 60.565 25.310 60.960 ;
        RECT 24.705 60.395 25.310 60.565 ;
        RECT 25.545 60.675 25.715 62.015 ;
        RECT 26.085 61.745 26.255 62.015 ;
        RECT 26.425 61.915 26.755 62.275 ;
        RECT 27.390 61.825 28.050 61.995 ;
        RECT 26.085 61.595 26.690 61.745 ;
        RECT 26.085 61.575 26.890 61.595 ;
        RECT 26.010 61.035 26.340 61.405 ;
        RECT 26.520 61.265 26.890 61.575 ;
        RECT 27.265 61.325 27.645 61.655 ;
        RECT 26.520 60.865 26.690 61.265 ;
        RECT 26.005 60.695 26.690 60.865 ;
        RECT 24.705 59.895 24.875 60.395 ;
        RECT 25.045 59.725 25.375 60.225 ;
        RECT 25.545 59.895 25.770 60.675 ;
        RECT 26.005 59.945 26.335 60.695 ;
        RECT 26.505 59.725 26.820 60.525 ;
        RECT 27.020 60.355 27.305 61.005 ;
        RECT 27.475 60.945 27.645 61.325 ;
        RECT 27.880 61.365 28.050 61.825 ;
        RECT 28.290 61.535 28.620 62.275 ;
        RECT 28.890 61.535 29.110 61.945 ;
        RECT 29.290 61.535 29.575 62.275 ;
        RECT 29.745 61.675 29.995 61.945 ;
        RECT 30.165 61.810 30.425 62.275 ;
        RECT 30.685 61.725 30.855 62.015 ;
        RECT 31.025 61.895 31.355 62.275 ;
        RECT 29.745 61.535 30.030 61.675 ;
        RECT 30.685 61.555 31.290 61.725 ;
        RECT 28.940 61.365 29.110 61.535 ;
        RECT 29.860 61.365 30.030 61.535 ;
        RECT 27.880 61.195 28.750 61.365 ;
        RECT 28.030 61.035 28.750 61.195 ;
        RECT 28.940 61.035 29.690 61.365 ;
        RECT 29.860 61.035 30.425 61.365 ;
        RECT 27.475 60.365 27.815 60.945 ;
        RECT 28.030 60.105 28.200 61.035 ;
        RECT 28.940 60.825 29.110 61.035 ;
        RECT 29.860 60.865 30.030 61.035 ;
        RECT 28.390 60.495 29.110 60.825 ;
        RECT 27.450 59.935 28.200 60.105 ;
        RECT 28.370 59.725 28.670 60.225 ;
        RECT 28.890 59.925 29.110 60.495 ;
        RECT 29.290 59.725 29.575 60.865 ;
        RECT 29.745 60.720 30.030 60.865 ;
        RECT 30.595 60.735 30.840 61.375 ;
        RECT 31.120 61.290 31.290 61.555 ;
        RECT 31.120 60.960 31.350 61.290 ;
        RECT 29.745 59.905 29.995 60.720 ;
        RECT 30.165 59.725 30.425 60.605 ;
        RECT 31.120 60.565 31.290 60.960 ;
        RECT 30.685 60.395 31.290 60.565 ;
        RECT 31.525 60.675 31.695 62.015 ;
        RECT 32.065 61.745 32.235 62.015 ;
        RECT 32.405 61.915 32.735 62.275 ;
        RECT 33.370 61.825 34.030 61.995 ;
        RECT 32.065 61.595 32.670 61.745 ;
        RECT 32.065 61.575 32.870 61.595 ;
        RECT 31.990 61.035 32.320 61.405 ;
        RECT 32.500 61.265 32.870 61.575 ;
        RECT 33.245 61.325 33.625 61.655 ;
        RECT 32.500 60.865 32.670 61.265 ;
        RECT 31.985 60.695 32.670 60.865 ;
        RECT 30.685 59.895 30.855 60.395 ;
        RECT 31.025 59.725 31.355 60.225 ;
        RECT 31.525 59.895 31.750 60.675 ;
        RECT 31.985 59.945 32.315 60.695 ;
        RECT 32.485 59.725 32.800 60.525 ;
        RECT 33.000 60.355 33.285 61.005 ;
        RECT 33.455 60.945 33.625 61.325 ;
        RECT 33.860 61.365 34.030 61.825 ;
        RECT 34.270 61.535 34.600 62.275 ;
        RECT 34.870 61.535 35.090 61.945 ;
        RECT 35.270 61.535 35.555 62.275 ;
        RECT 35.725 61.675 35.975 61.945 ;
        RECT 36.145 61.810 36.405 62.275 ;
        RECT 36.665 61.725 36.835 62.015 ;
        RECT 37.005 61.895 37.335 62.275 ;
        RECT 35.725 61.535 36.010 61.675 ;
        RECT 36.665 61.555 37.270 61.725 ;
        RECT 34.920 61.365 35.090 61.535 ;
        RECT 35.840 61.365 36.010 61.535 ;
        RECT 33.860 61.195 34.730 61.365 ;
        RECT 34.010 61.035 34.730 61.195 ;
        RECT 34.920 61.035 35.670 61.365 ;
        RECT 35.840 61.035 36.405 61.365 ;
        RECT 33.455 60.365 33.795 60.945 ;
        RECT 34.010 60.105 34.180 61.035 ;
        RECT 34.920 60.825 35.090 61.035 ;
        RECT 35.840 60.865 36.010 61.035 ;
        RECT 34.370 60.495 35.090 60.825 ;
        RECT 33.430 59.935 34.180 60.105 ;
        RECT 34.350 59.725 34.650 60.225 ;
        RECT 34.870 59.925 35.090 60.495 ;
        RECT 35.270 59.725 35.555 60.865 ;
        RECT 35.725 60.720 36.010 60.865 ;
        RECT 36.575 60.735 36.820 61.375 ;
        RECT 37.100 61.290 37.270 61.555 ;
        RECT 37.100 60.960 37.330 61.290 ;
        RECT 35.725 59.905 35.975 60.720 ;
        RECT 36.145 59.725 36.405 60.605 ;
        RECT 37.100 60.565 37.270 60.960 ;
        RECT 36.665 60.395 37.270 60.565 ;
        RECT 37.505 60.675 37.675 62.015 ;
        RECT 38.045 61.745 38.215 62.015 ;
        RECT 38.385 61.915 38.715 62.275 ;
        RECT 39.350 61.825 40.010 61.995 ;
        RECT 38.045 61.595 38.650 61.745 ;
        RECT 38.045 61.575 38.850 61.595 ;
        RECT 37.970 61.035 38.300 61.405 ;
        RECT 38.480 61.265 38.850 61.575 ;
        RECT 39.225 61.325 39.605 61.655 ;
        RECT 38.480 60.865 38.650 61.265 ;
        RECT 37.965 60.695 38.650 60.865 ;
        RECT 36.665 59.895 36.835 60.395 ;
        RECT 37.005 59.725 37.335 60.225 ;
        RECT 37.505 59.895 37.730 60.675 ;
        RECT 37.965 59.945 38.295 60.695 ;
        RECT 38.465 59.725 38.780 60.525 ;
        RECT 38.980 60.355 39.265 61.005 ;
        RECT 39.435 60.945 39.605 61.325 ;
        RECT 39.840 61.365 40.010 61.825 ;
        RECT 40.250 61.535 40.580 62.275 ;
        RECT 40.850 61.535 41.070 61.945 ;
        RECT 41.250 61.535 41.535 62.275 ;
        RECT 41.705 61.675 41.955 61.945 ;
        RECT 42.125 61.810 42.385 62.275 ;
        RECT 42.645 61.725 42.815 62.015 ;
        RECT 42.985 61.895 43.315 62.275 ;
        RECT 41.705 61.535 41.990 61.675 ;
        RECT 42.645 61.555 43.250 61.725 ;
        RECT 40.900 61.365 41.070 61.535 ;
        RECT 41.820 61.365 41.990 61.535 ;
        RECT 39.840 61.195 40.710 61.365 ;
        RECT 39.990 61.035 40.710 61.195 ;
        RECT 40.900 61.035 41.650 61.365 ;
        RECT 41.820 61.035 42.385 61.365 ;
        RECT 39.435 60.365 39.775 60.945 ;
        RECT 39.990 60.105 40.160 61.035 ;
        RECT 40.900 60.825 41.070 61.035 ;
        RECT 41.820 60.865 41.990 61.035 ;
        RECT 40.350 60.495 41.070 60.825 ;
        RECT 39.410 59.935 40.160 60.105 ;
        RECT 40.330 59.725 40.630 60.225 ;
        RECT 40.850 59.925 41.070 60.495 ;
        RECT 41.250 59.725 41.535 60.865 ;
        RECT 41.705 60.720 41.990 60.865 ;
        RECT 42.555 60.735 42.800 61.375 ;
        RECT 43.080 61.290 43.250 61.555 ;
        RECT 43.080 60.960 43.310 61.290 ;
        RECT 41.705 59.905 41.955 60.720 ;
        RECT 42.125 59.725 42.385 60.605 ;
        RECT 43.080 60.565 43.250 60.960 ;
        RECT 42.645 60.395 43.250 60.565 ;
        RECT 43.485 60.675 43.655 62.015 ;
        RECT 44.025 61.745 44.195 62.015 ;
        RECT 44.365 61.915 44.695 62.275 ;
        RECT 45.330 61.825 45.990 61.995 ;
        RECT 44.025 61.595 44.630 61.745 ;
        RECT 44.025 61.575 44.830 61.595 ;
        RECT 43.950 61.035 44.280 61.405 ;
        RECT 44.460 61.265 44.830 61.575 ;
        RECT 45.205 61.325 45.585 61.655 ;
        RECT 44.460 60.865 44.630 61.265 ;
        RECT 43.945 60.695 44.630 60.865 ;
        RECT 42.645 59.895 42.815 60.395 ;
        RECT 42.985 59.725 43.315 60.225 ;
        RECT 43.485 59.895 43.710 60.675 ;
        RECT 43.945 59.945 44.275 60.695 ;
        RECT 44.445 59.725 44.760 60.525 ;
        RECT 44.960 60.355 45.245 61.005 ;
        RECT 45.415 60.945 45.585 61.325 ;
        RECT 45.820 61.365 45.990 61.825 ;
        RECT 46.230 61.535 46.560 62.275 ;
        RECT 46.830 61.535 47.050 61.945 ;
        RECT 47.230 61.535 47.515 62.275 ;
        RECT 47.685 61.675 47.935 61.945 ;
        RECT 48.105 61.810 48.365 62.275 ;
        RECT 47.685 61.535 47.970 61.675 ;
        RECT 48.535 61.550 48.825 62.275 ;
        RECT 49.175 61.615 49.515 62.275 ;
        RECT 46.880 61.365 47.050 61.535 ;
        RECT 47.800 61.365 47.970 61.535 ;
        RECT 45.820 61.195 46.690 61.365 ;
        RECT 45.970 61.035 46.690 61.195 ;
        RECT 46.880 61.035 47.630 61.365 ;
        RECT 47.800 61.035 48.365 61.365 ;
        RECT 45.415 60.365 45.755 60.945 ;
        RECT 45.970 60.105 46.140 61.035 ;
        RECT 46.880 60.825 47.050 61.035 ;
        RECT 47.800 60.865 47.970 61.035 ;
        RECT 46.330 60.495 47.050 60.825 ;
        RECT 45.390 59.935 46.140 60.105 ;
        RECT 46.310 59.725 46.610 60.225 ;
        RECT 46.830 59.925 47.050 60.495 ;
        RECT 47.230 59.725 47.515 60.865 ;
        RECT 47.685 60.720 47.970 60.865 ;
        RECT 47.685 59.905 47.935 60.720 ;
        RECT 48.105 59.725 48.365 60.605 ;
        RECT 48.535 59.725 48.825 60.890 ;
        RECT 48.995 59.895 49.515 61.445 ;
        RECT 49.685 60.620 50.205 62.105 ;
        RECT 51.475 61.615 51.815 62.275 ;
        RECT 49.685 59.725 50.015 60.450 ;
        RECT 51.295 59.895 51.815 61.445 ;
        RECT 51.985 60.620 52.505 62.105 ;
        RECT 52.675 60.620 53.195 62.105 ;
        RECT 53.365 61.615 53.705 62.275 ;
        RECT 54.145 61.725 54.315 62.015 ;
        RECT 54.485 61.895 54.815 62.275 ;
        RECT 54.145 61.555 54.750 61.725 ;
        RECT 51.985 59.725 52.315 60.450 ;
        RECT 52.865 59.725 53.195 60.450 ;
        RECT 53.365 59.895 53.885 61.445 ;
        RECT 54.055 60.735 54.300 61.375 ;
        RECT 54.580 61.290 54.750 61.555 ;
        RECT 54.580 60.960 54.810 61.290 ;
        RECT 54.580 60.565 54.750 60.960 ;
        RECT 54.145 60.395 54.750 60.565 ;
        RECT 54.985 60.675 55.155 62.015 ;
        RECT 55.525 61.745 55.695 62.015 ;
        RECT 55.865 61.915 56.195 62.275 ;
        RECT 56.830 61.825 57.490 61.995 ;
        RECT 55.525 61.595 56.130 61.745 ;
        RECT 55.525 61.575 56.330 61.595 ;
        RECT 55.450 61.035 55.780 61.405 ;
        RECT 55.960 61.265 56.330 61.575 ;
        RECT 56.705 61.325 57.085 61.655 ;
        RECT 55.960 60.865 56.130 61.265 ;
        RECT 55.445 60.695 56.130 60.865 ;
        RECT 54.145 59.895 54.315 60.395 ;
        RECT 54.485 59.725 54.815 60.225 ;
        RECT 54.985 59.895 55.210 60.675 ;
        RECT 55.445 59.945 55.775 60.695 ;
        RECT 55.945 59.725 56.260 60.525 ;
        RECT 56.460 60.355 56.745 61.005 ;
        RECT 56.915 60.945 57.085 61.325 ;
        RECT 57.320 61.365 57.490 61.825 ;
        RECT 57.730 61.535 58.060 62.275 ;
        RECT 58.330 61.535 58.550 61.945 ;
        RECT 58.730 61.535 59.015 62.275 ;
        RECT 59.185 61.675 59.435 61.945 ;
        RECT 59.605 61.810 59.865 62.275 ;
        RECT 60.125 61.725 60.295 62.015 ;
        RECT 60.465 61.895 60.795 62.275 ;
        RECT 59.185 61.535 59.470 61.675 ;
        RECT 60.125 61.555 60.730 61.725 ;
        RECT 58.380 61.365 58.550 61.535 ;
        RECT 59.300 61.365 59.470 61.535 ;
        RECT 57.320 61.195 58.190 61.365 ;
        RECT 57.470 61.035 58.190 61.195 ;
        RECT 58.380 61.035 59.130 61.365 ;
        RECT 59.300 61.035 59.865 61.365 ;
        RECT 56.915 60.365 57.255 60.945 ;
        RECT 57.470 60.105 57.640 61.035 ;
        RECT 58.380 60.825 58.550 61.035 ;
        RECT 59.300 60.865 59.470 61.035 ;
        RECT 57.830 60.495 58.550 60.825 ;
        RECT 56.890 59.935 57.640 60.105 ;
        RECT 57.810 59.725 58.110 60.225 ;
        RECT 58.330 59.925 58.550 60.495 ;
        RECT 58.730 59.725 59.015 60.865 ;
        RECT 59.185 60.720 59.470 60.865 ;
        RECT 60.035 60.735 60.280 61.375 ;
        RECT 60.560 61.290 60.730 61.555 ;
        RECT 60.560 60.960 60.790 61.290 ;
        RECT 59.185 59.905 59.435 60.720 ;
        RECT 59.605 59.725 59.865 60.605 ;
        RECT 60.560 60.565 60.730 60.960 ;
        RECT 60.125 60.395 60.730 60.565 ;
        RECT 60.965 60.675 61.135 62.015 ;
        RECT 61.505 61.745 61.675 62.015 ;
        RECT 61.845 61.915 62.175 62.275 ;
        RECT 62.810 61.825 63.470 61.995 ;
        RECT 61.505 61.595 62.110 61.745 ;
        RECT 61.505 61.575 62.310 61.595 ;
        RECT 61.430 61.035 61.760 61.405 ;
        RECT 61.940 61.265 62.310 61.575 ;
        RECT 62.685 61.325 63.065 61.655 ;
        RECT 61.940 60.865 62.110 61.265 ;
        RECT 61.425 60.695 62.110 60.865 ;
        RECT 60.125 59.895 60.295 60.395 ;
        RECT 60.465 59.725 60.795 60.225 ;
        RECT 60.965 59.895 61.190 60.675 ;
        RECT 61.425 59.945 61.755 60.695 ;
        RECT 61.925 59.725 62.240 60.525 ;
        RECT 62.440 60.355 62.725 61.005 ;
        RECT 62.895 60.945 63.065 61.325 ;
        RECT 63.300 61.365 63.470 61.825 ;
        RECT 63.710 61.535 64.040 62.275 ;
        RECT 64.310 61.535 64.530 61.945 ;
        RECT 64.710 61.535 64.995 62.275 ;
        RECT 65.165 61.675 65.415 61.945 ;
        RECT 65.585 61.810 65.845 62.275 ;
        RECT 65.165 61.535 65.450 61.675 ;
        RECT 64.360 61.365 64.530 61.535 ;
        RECT 65.280 61.365 65.450 61.535 ;
        RECT 63.300 61.195 64.170 61.365 ;
        RECT 63.450 61.035 64.170 61.195 ;
        RECT 64.360 61.035 65.110 61.365 ;
        RECT 65.280 61.035 65.845 61.365 ;
        RECT 62.895 60.365 63.235 60.945 ;
        RECT 63.450 60.105 63.620 61.035 ;
        RECT 64.360 60.825 64.530 61.035 ;
        RECT 65.280 60.865 65.450 61.035 ;
        RECT 63.810 60.495 64.530 60.825 ;
        RECT 62.870 59.935 63.620 60.105 ;
        RECT 63.790 59.725 64.090 60.225 ;
        RECT 64.310 59.925 64.530 60.495 ;
        RECT 64.710 59.725 64.995 60.865 ;
        RECT 65.165 60.720 65.450 60.865 ;
        RECT 65.165 59.905 65.415 60.720 ;
        RECT 66.475 60.620 66.995 62.105 ;
        RECT 67.165 61.615 67.505 62.275 ;
        RECT 67.945 61.725 68.115 62.015 ;
        RECT 68.285 61.895 68.615 62.275 ;
        RECT 67.945 61.555 68.550 61.725 ;
        RECT 65.585 59.725 65.845 60.605 ;
        RECT 66.665 59.725 66.995 60.450 ;
        RECT 67.165 59.895 67.685 61.445 ;
        RECT 67.855 60.735 68.100 61.375 ;
        RECT 68.380 61.290 68.550 61.555 ;
        RECT 68.380 60.960 68.610 61.290 ;
        RECT 68.380 60.565 68.550 60.960 ;
        RECT 67.945 60.395 68.550 60.565 ;
        RECT 68.785 60.675 68.955 62.015 ;
        RECT 69.325 61.745 69.495 62.015 ;
        RECT 69.665 61.915 69.995 62.275 ;
        RECT 70.630 61.825 71.290 61.995 ;
        RECT 69.325 61.595 69.930 61.745 ;
        RECT 69.325 61.575 70.130 61.595 ;
        RECT 69.250 61.035 69.580 61.405 ;
        RECT 69.760 61.265 70.130 61.575 ;
        RECT 70.505 61.325 70.885 61.655 ;
        RECT 69.760 60.865 69.930 61.265 ;
        RECT 69.245 60.695 69.930 60.865 ;
        RECT 67.945 59.895 68.115 60.395 ;
        RECT 68.285 59.725 68.615 60.225 ;
        RECT 68.785 59.895 69.010 60.675 ;
        RECT 69.245 59.945 69.575 60.695 ;
        RECT 69.745 59.725 70.060 60.525 ;
        RECT 70.260 60.355 70.545 61.005 ;
        RECT 70.715 60.945 70.885 61.325 ;
        RECT 71.120 61.365 71.290 61.825 ;
        RECT 71.530 61.535 71.860 62.275 ;
        RECT 72.130 61.535 72.350 61.945 ;
        RECT 72.530 61.535 72.815 62.275 ;
        RECT 72.985 61.675 73.235 61.945 ;
        RECT 73.405 61.810 73.665 62.275 ;
        RECT 72.985 61.535 73.270 61.675 ;
        RECT 74.295 61.550 74.585 62.275 ;
        RECT 75.305 61.725 75.475 62.015 ;
        RECT 75.645 61.895 75.975 62.275 ;
        RECT 75.305 61.555 75.910 61.725 ;
        RECT 72.180 61.365 72.350 61.535 ;
        RECT 73.100 61.365 73.270 61.535 ;
        RECT 71.120 61.195 71.990 61.365 ;
        RECT 71.270 61.035 71.990 61.195 ;
        RECT 72.180 61.035 72.930 61.365 ;
        RECT 73.100 61.035 73.665 61.365 ;
        RECT 70.715 60.365 71.055 60.945 ;
        RECT 71.270 60.105 71.440 61.035 ;
        RECT 72.180 60.825 72.350 61.035 ;
        RECT 73.100 60.865 73.270 61.035 ;
        RECT 71.630 60.495 72.350 60.825 ;
        RECT 70.690 59.935 71.440 60.105 ;
        RECT 71.610 59.725 71.910 60.225 ;
        RECT 72.130 59.925 72.350 60.495 ;
        RECT 72.530 59.725 72.815 60.865 ;
        RECT 72.985 60.720 73.270 60.865 ;
        RECT 72.985 59.905 73.235 60.720 ;
        RECT 73.405 59.725 73.665 60.605 ;
        RECT 74.295 59.725 74.585 60.890 ;
        RECT 75.215 60.735 75.460 61.375 ;
        RECT 75.740 61.290 75.910 61.555 ;
        RECT 75.740 60.960 75.970 61.290 ;
        RECT 75.740 60.565 75.910 60.960 ;
        RECT 75.305 60.395 75.910 60.565 ;
        RECT 76.145 60.675 76.315 62.015 ;
        RECT 76.685 61.745 76.855 62.015 ;
        RECT 77.025 61.915 77.355 62.275 ;
        RECT 77.990 61.825 78.650 61.995 ;
        RECT 76.685 61.595 77.290 61.745 ;
        RECT 76.685 61.575 77.490 61.595 ;
        RECT 76.610 61.035 76.940 61.405 ;
        RECT 77.120 61.265 77.490 61.575 ;
        RECT 77.865 61.325 78.245 61.655 ;
        RECT 77.120 60.865 77.290 61.265 ;
        RECT 76.605 60.695 77.290 60.865 ;
        RECT 75.305 59.895 75.475 60.395 ;
        RECT 75.645 59.725 75.975 60.225 ;
        RECT 76.145 59.895 76.370 60.675 ;
        RECT 76.605 59.945 76.935 60.695 ;
        RECT 77.105 59.725 77.420 60.525 ;
        RECT 77.620 60.355 77.905 61.005 ;
        RECT 78.075 60.945 78.245 61.325 ;
        RECT 78.480 61.365 78.650 61.825 ;
        RECT 78.890 61.535 79.220 62.275 ;
        RECT 79.490 61.535 79.710 61.945 ;
        RECT 79.890 61.535 80.175 62.275 ;
        RECT 80.345 61.675 80.595 61.945 ;
        RECT 80.765 61.810 81.025 62.275 ;
        RECT 81.285 61.725 81.455 62.015 ;
        RECT 81.625 61.895 81.955 62.275 ;
        RECT 80.345 61.535 80.630 61.675 ;
        RECT 81.285 61.555 81.890 61.725 ;
        RECT 79.540 61.365 79.710 61.535 ;
        RECT 80.460 61.365 80.630 61.535 ;
        RECT 78.480 61.195 79.350 61.365 ;
        RECT 78.630 61.035 79.350 61.195 ;
        RECT 79.540 61.035 80.290 61.365 ;
        RECT 80.460 61.035 81.025 61.365 ;
        RECT 78.075 60.365 78.415 60.945 ;
        RECT 78.630 60.105 78.800 61.035 ;
        RECT 79.540 60.825 79.710 61.035 ;
        RECT 80.460 60.865 80.630 61.035 ;
        RECT 78.990 60.495 79.710 60.825 ;
        RECT 78.050 59.935 78.800 60.105 ;
        RECT 78.970 59.725 79.270 60.225 ;
        RECT 79.490 59.925 79.710 60.495 ;
        RECT 79.890 59.725 80.175 60.865 ;
        RECT 80.345 60.720 80.630 60.865 ;
        RECT 81.195 60.735 81.440 61.375 ;
        RECT 81.720 61.290 81.890 61.555 ;
        RECT 81.720 60.960 81.950 61.290 ;
        RECT 80.345 59.905 80.595 60.720 ;
        RECT 80.765 59.725 81.025 60.605 ;
        RECT 81.720 60.565 81.890 60.960 ;
        RECT 81.285 60.395 81.890 60.565 ;
        RECT 82.125 60.675 82.295 62.015 ;
        RECT 82.665 61.745 82.835 62.015 ;
        RECT 83.005 61.915 83.335 62.275 ;
        RECT 83.970 61.825 84.630 61.995 ;
        RECT 82.665 61.595 83.270 61.745 ;
        RECT 82.665 61.575 83.470 61.595 ;
        RECT 82.590 61.035 82.920 61.405 ;
        RECT 83.100 61.265 83.470 61.575 ;
        RECT 83.845 61.325 84.225 61.655 ;
        RECT 83.100 60.865 83.270 61.265 ;
        RECT 82.585 60.695 83.270 60.865 ;
        RECT 81.285 59.895 81.455 60.395 ;
        RECT 81.625 59.725 81.955 60.225 ;
        RECT 82.125 59.895 82.350 60.675 ;
        RECT 82.585 59.945 82.915 60.695 ;
        RECT 83.085 59.725 83.400 60.525 ;
        RECT 83.600 60.355 83.885 61.005 ;
        RECT 84.055 60.945 84.225 61.325 ;
        RECT 84.460 61.365 84.630 61.825 ;
        RECT 84.870 61.535 85.200 62.275 ;
        RECT 85.470 61.535 85.690 61.945 ;
        RECT 85.870 61.535 86.155 62.275 ;
        RECT 86.325 61.675 86.575 61.945 ;
        RECT 86.745 61.810 87.005 62.275 ;
        RECT 87.265 61.725 87.435 62.015 ;
        RECT 87.605 61.895 87.935 62.275 ;
        RECT 86.325 61.535 86.610 61.675 ;
        RECT 87.265 61.555 87.870 61.725 ;
        RECT 85.520 61.365 85.690 61.535 ;
        RECT 86.440 61.365 86.610 61.535 ;
        RECT 84.460 61.195 85.330 61.365 ;
        RECT 84.610 61.035 85.330 61.195 ;
        RECT 85.520 61.035 86.270 61.365 ;
        RECT 86.440 61.035 87.005 61.365 ;
        RECT 84.055 60.365 84.395 60.945 ;
        RECT 84.610 60.105 84.780 61.035 ;
        RECT 85.520 60.825 85.690 61.035 ;
        RECT 86.440 60.865 86.610 61.035 ;
        RECT 84.970 60.495 85.690 60.825 ;
        RECT 84.030 59.935 84.780 60.105 ;
        RECT 84.950 59.725 85.250 60.225 ;
        RECT 85.470 59.925 85.690 60.495 ;
        RECT 85.870 59.725 86.155 60.865 ;
        RECT 86.325 60.720 86.610 60.865 ;
        RECT 87.175 60.735 87.420 61.375 ;
        RECT 87.700 61.290 87.870 61.555 ;
        RECT 87.700 60.960 87.930 61.290 ;
        RECT 86.325 59.905 86.575 60.720 ;
        RECT 86.745 59.725 87.005 60.605 ;
        RECT 87.700 60.565 87.870 60.960 ;
        RECT 87.265 60.395 87.870 60.565 ;
        RECT 88.105 60.675 88.275 62.015 ;
        RECT 88.645 61.745 88.815 62.015 ;
        RECT 88.985 61.915 89.315 62.275 ;
        RECT 89.950 61.825 90.610 61.995 ;
        RECT 88.645 61.595 89.250 61.745 ;
        RECT 88.645 61.575 89.450 61.595 ;
        RECT 88.570 61.035 88.900 61.405 ;
        RECT 89.080 61.265 89.450 61.575 ;
        RECT 89.825 61.325 90.205 61.655 ;
        RECT 89.080 60.865 89.250 61.265 ;
        RECT 88.565 60.695 89.250 60.865 ;
        RECT 87.265 59.895 87.435 60.395 ;
        RECT 87.605 59.725 87.935 60.225 ;
        RECT 88.105 59.895 88.330 60.675 ;
        RECT 88.565 59.945 88.895 60.695 ;
        RECT 89.065 59.725 89.380 60.525 ;
        RECT 89.580 60.355 89.865 61.005 ;
        RECT 90.035 60.945 90.205 61.325 ;
        RECT 90.440 61.365 90.610 61.825 ;
        RECT 90.850 61.535 91.180 62.275 ;
        RECT 91.450 61.535 91.670 61.945 ;
        RECT 91.850 61.535 92.135 62.275 ;
        RECT 92.305 61.675 92.555 61.945 ;
        RECT 92.725 61.810 92.985 62.275 ;
        RECT 93.245 61.725 93.415 62.015 ;
        RECT 93.585 61.895 93.915 62.275 ;
        RECT 92.305 61.535 92.590 61.675 ;
        RECT 93.245 61.555 93.850 61.725 ;
        RECT 91.500 61.365 91.670 61.535 ;
        RECT 92.420 61.365 92.590 61.535 ;
        RECT 90.440 61.195 91.310 61.365 ;
        RECT 90.590 61.035 91.310 61.195 ;
        RECT 91.500 61.035 92.250 61.365 ;
        RECT 92.420 61.035 92.985 61.365 ;
        RECT 90.035 60.365 90.375 60.945 ;
        RECT 90.590 60.105 90.760 61.035 ;
        RECT 91.500 60.825 91.670 61.035 ;
        RECT 92.420 60.865 92.590 61.035 ;
        RECT 90.950 60.495 91.670 60.825 ;
        RECT 90.010 59.935 90.760 60.105 ;
        RECT 90.930 59.725 91.230 60.225 ;
        RECT 91.450 59.925 91.670 60.495 ;
        RECT 91.850 59.725 92.135 60.865 ;
        RECT 92.305 60.720 92.590 60.865 ;
        RECT 93.155 60.735 93.400 61.375 ;
        RECT 93.680 61.290 93.850 61.555 ;
        RECT 93.680 60.960 93.910 61.290 ;
        RECT 92.305 59.905 92.555 60.720 ;
        RECT 92.725 59.725 92.985 60.605 ;
        RECT 93.680 60.565 93.850 60.960 ;
        RECT 93.245 60.395 93.850 60.565 ;
        RECT 94.085 60.675 94.255 62.015 ;
        RECT 94.625 61.745 94.795 62.015 ;
        RECT 94.965 61.915 95.295 62.275 ;
        RECT 95.930 61.825 96.590 61.995 ;
        RECT 94.625 61.595 95.230 61.745 ;
        RECT 94.625 61.575 95.430 61.595 ;
        RECT 94.550 61.035 94.880 61.405 ;
        RECT 95.060 61.265 95.430 61.575 ;
        RECT 95.805 61.325 96.185 61.655 ;
        RECT 95.060 60.865 95.230 61.265 ;
        RECT 94.545 60.695 95.230 60.865 ;
        RECT 93.245 59.895 93.415 60.395 ;
        RECT 93.585 59.725 93.915 60.225 ;
        RECT 94.085 59.895 94.310 60.675 ;
        RECT 94.545 59.945 94.875 60.695 ;
        RECT 95.045 59.725 95.360 60.525 ;
        RECT 95.560 60.355 95.845 61.005 ;
        RECT 96.015 60.945 96.185 61.325 ;
        RECT 96.420 61.365 96.590 61.825 ;
        RECT 96.830 61.535 97.160 62.275 ;
        RECT 97.430 61.535 97.650 61.945 ;
        RECT 97.830 61.535 98.115 62.275 ;
        RECT 98.285 61.675 98.535 61.945 ;
        RECT 98.705 61.810 98.965 62.275 ;
        RECT 98.285 61.535 98.570 61.675 ;
        RECT 100.055 61.550 100.345 62.275 ;
        RECT 100.605 61.725 100.775 62.015 ;
        RECT 100.945 61.895 101.275 62.275 ;
        RECT 100.605 61.555 101.210 61.725 ;
        RECT 97.480 61.365 97.650 61.535 ;
        RECT 98.400 61.365 98.570 61.535 ;
        RECT 96.420 61.195 97.290 61.365 ;
        RECT 96.570 61.035 97.290 61.195 ;
        RECT 97.480 61.035 98.230 61.365 ;
        RECT 98.400 61.035 98.965 61.365 ;
        RECT 96.015 60.365 96.355 60.945 ;
        RECT 96.570 60.105 96.740 61.035 ;
        RECT 97.480 60.825 97.650 61.035 ;
        RECT 98.400 60.865 98.570 61.035 ;
        RECT 96.930 60.495 97.650 60.825 ;
        RECT 95.990 59.935 96.740 60.105 ;
        RECT 96.910 59.725 97.210 60.225 ;
        RECT 97.430 59.925 97.650 60.495 ;
        RECT 97.830 59.725 98.115 60.865 ;
        RECT 98.285 60.720 98.570 60.865 ;
        RECT 98.285 59.905 98.535 60.720 ;
        RECT 98.705 59.725 98.965 60.605 ;
        RECT 100.055 59.725 100.345 60.890 ;
        RECT 100.515 60.735 100.760 61.375 ;
        RECT 101.040 61.290 101.210 61.555 ;
        RECT 101.040 60.960 101.270 61.290 ;
        RECT 101.040 60.565 101.210 60.960 ;
        RECT 100.605 60.395 101.210 60.565 ;
        RECT 101.445 60.675 101.615 62.015 ;
        RECT 101.985 61.745 102.155 62.015 ;
        RECT 102.325 61.915 102.655 62.275 ;
        RECT 103.290 61.825 103.950 61.995 ;
        RECT 101.985 61.595 102.590 61.745 ;
        RECT 101.985 61.575 102.790 61.595 ;
        RECT 101.910 61.035 102.240 61.405 ;
        RECT 102.420 61.265 102.790 61.575 ;
        RECT 103.165 61.325 103.545 61.655 ;
        RECT 102.420 60.865 102.590 61.265 ;
        RECT 101.905 60.695 102.590 60.865 ;
        RECT 100.605 59.895 100.775 60.395 ;
        RECT 100.945 59.725 101.275 60.225 ;
        RECT 101.445 59.895 101.670 60.675 ;
        RECT 101.905 59.945 102.235 60.695 ;
        RECT 102.405 59.725 102.720 60.525 ;
        RECT 102.920 60.355 103.205 61.005 ;
        RECT 103.375 60.945 103.545 61.325 ;
        RECT 103.780 61.365 103.950 61.825 ;
        RECT 104.190 61.535 104.520 62.275 ;
        RECT 104.790 61.535 105.010 61.945 ;
        RECT 105.190 61.535 105.475 62.275 ;
        RECT 105.645 61.675 105.895 61.945 ;
        RECT 106.065 61.810 106.325 62.275 ;
        RECT 106.585 61.725 106.755 62.015 ;
        RECT 106.925 61.895 107.255 62.275 ;
        RECT 105.645 61.535 105.930 61.675 ;
        RECT 106.585 61.555 107.190 61.725 ;
        RECT 104.840 61.365 105.010 61.535 ;
        RECT 105.760 61.365 105.930 61.535 ;
        RECT 103.780 61.195 104.650 61.365 ;
        RECT 103.930 61.035 104.650 61.195 ;
        RECT 104.840 61.035 105.590 61.365 ;
        RECT 105.760 61.035 106.325 61.365 ;
        RECT 103.375 60.365 103.715 60.945 ;
        RECT 103.930 60.105 104.100 61.035 ;
        RECT 104.840 60.825 105.010 61.035 ;
        RECT 105.760 60.865 105.930 61.035 ;
        RECT 104.290 60.495 105.010 60.825 ;
        RECT 103.350 59.935 104.100 60.105 ;
        RECT 104.270 59.725 104.570 60.225 ;
        RECT 104.790 59.925 105.010 60.495 ;
        RECT 105.190 59.725 105.475 60.865 ;
        RECT 105.645 60.720 105.930 60.865 ;
        RECT 106.495 60.735 106.740 61.375 ;
        RECT 107.020 61.290 107.190 61.555 ;
        RECT 107.020 60.960 107.250 61.290 ;
        RECT 105.645 59.905 105.895 60.720 ;
        RECT 106.065 59.725 106.325 60.605 ;
        RECT 107.020 60.565 107.190 60.960 ;
        RECT 106.585 60.395 107.190 60.565 ;
        RECT 107.425 60.675 107.595 62.015 ;
        RECT 107.965 61.745 108.135 62.015 ;
        RECT 108.305 61.915 108.635 62.275 ;
        RECT 109.270 61.825 109.930 61.995 ;
        RECT 107.965 61.595 108.570 61.745 ;
        RECT 107.965 61.575 108.770 61.595 ;
        RECT 107.890 61.035 108.220 61.405 ;
        RECT 108.400 61.265 108.770 61.575 ;
        RECT 109.145 61.325 109.525 61.655 ;
        RECT 108.400 60.865 108.570 61.265 ;
        RECT 107.885 60.695 108.570 60.865 ;
        RECT 106.585 59.895 106.755 60.395 ;
        RECT 106.925 59.725 107.255 60.225 ;
        RECT 107.425 59.895 107.650 60.675 ;
        RECT 107.885 59.945 108.215 60.695 ;
        RECT 108.385 59.725 108.700 60.525 ;
        RECT 108.900 60.355 109.185 61.005 ;
        RECT 109.355 60.945 109.525 61.325 ;
        RECT 109.760 61.365 109.930 61.825 ;
        RECT 110.170 61.535 110.500 62.275 ;
        RECT 110.770 61.535 110.990 61.945 ;
        RECT 111.170 61.535 111.455 62.275 ;
        RECT 111.625 61.675 111.875 61.945 ;
        RECT 112.045 61.810 112.305 62.275 ;
        RECT 112.475 61.810 112.735 62.275 ;
        RECT 112.905 61.675 113.155 61.945 ;
        RECT 111.625 61.535 111.910 61.675 ;
        RECT 110.820 61.365 110.990 61.535 ;
        RECT 111.740 61.365 111.910 61.535 ;
        RECT 112.870 61.535 113.155 61.675 ;
        RECT 113.325 61.535 113.610 62.275 ;
        RECT 113.790 61.535 114.010 61.945 ;
        RECT 114.280 61.535 114.610 62.275 ;
        RECT 114.850 61.825 115.510 61.995 ;
        RECT 116.145 61.915 116.475 62.275 ;
        RECT 112.870 61.365 113.040 61.535 ;
        RECT 113.790 61.365 113.960 61.535 ;
        RECT 114.850 61.365 115.020 61.825 ;
        RECT 116.645 61.745 116.815 62.015 ;
        RECT 109.760 61.195 110.630 61.365 ;
        RECT 109.910 61.035 110.630 61.195 ;
        RECT 110.820 61.035 111.570 61.365 ;
        RECT 111.740 61.035 112.305 61.365 ;
        RECT 112.475 61.035 113.040 61.365 ;
        RECT 113.210 61.035 113.960 61.365 ;
        RECT 114.150 61.195 115.020 61.365 ;
        RECT 115.255 61.325 115.635 61.655 ;
        RECT 116.210 61.595 116.815 61.745 ;
        RECT 116.010 61.575 116.815 61.595 ;
        RECT 114.150 61.035 114.870 61.195 ;
        RECT 109.355 60.365 109.695 60.945 ;
        RECT 109.910 60.105 110.080 61.035 ;
        RECT 110.820 60.825 110.990 61.035 ;
        RECT 111.740 60.865 111.910 61.035 ;
        RECT 110.270 60.495 110.990 60.825 ;
        RECT 109.330 59.935 110.080 60.105 ;
        RECT 110.250 59.725 110.550 60.225 ;
        RECT 110.770 59.925 110.990 60.495 ;
        RECT 111.170 59.725 111.455 60.865 ;
        RECT 111.625 60.720 111.910 60.865 ;
        RECT 112.870 60.865 113.040 61.035 ;
        RECT 112.870 60.720 113.155 60.865 ;
        RECT 111.625 59.905 111.875 60.720 ;
        RECT 112.045 59.725 112.305 60.605 ;
        RECT 112.475 59.725 112.735 60.605 ;
        RECT 112.905 59.905 113.155 60.720 ;
        RECT 113.325 59.725 113.610 60.865 ;
        RECT 113.790 60.825 113.960 61.035 ;
        RECT 113.790 60.495 114.510 60.825 ;
        RECT 113.790 59.925 114.010 60.495 ;
        RECT 114.230 59.725 114.530 60.225 ;
        RECT 114.700 60.105 114.870 61.035 ;
        RECT 115.255 60.945 115.425 61.325 ;
        RECT 116.010 61.265 116.380 61.575 ;
        RECT 115.085 60.365 115.425 60.945 ;
        RECT 115.595 60.355 115.880 61.005 ;
        RECT 116.210 60.865 116.380 61.265 ;
        RECT 116.560 61.035 116.890 61.405 ;
        RECT 116.210 60.695 116.895 60.865 ;
        RECT 114.700 59.935 115.450 60.105 ;
        RECT 116.080 59.725 116.395 60.525 ;
        RECT 116.565 59.945 116.895 60.695 ;
        RECT 117.185 60.675 117.355 62.015 ;
        RECT 117.525 61.895 117.855 62.275 ;
        RECT 118.025 61.725 118.195 62.015 ;
        RECT 117.590 61.555 118.195 61.725 ;
        RECT 118.545 61.725 118.715 62.015 ;
        RECT 118.885 61.895 119.215 62.275 ;
        RECT 118.545 61.555 119.150 61.725 ;
        RECT 117.590 61.290 117.760 61.555 ;
        RECT 117.530 60.960 117.760 61.290 ;
        RECT 117.130 59.895 117.355 60.675 ;
        RECT 117.590 60.565 117.760 60.960 ;
        RECT 118.040 60.735 118.285 61.375 ;
        RECT 118.455 60.735 118.700 61.375 ;
        RECT 118.980 61.290 119.150 61.555 ;
        RECT 118.980 60.960 119.210 61.290 ;
        RECT 118.980 60.565 119.150 60.960 ;
        RECT 117.590 60.395 118.195 60.565 ;
        RECT 117.525 59.725 117.855 60.225 ;
        RECT 118.025 59.895 118.195 60.395 ;
        RECT 118.545 60.395 119.150 60.565 ;
        RECT 119.385 60.675 119.555 62.015 ;
        RECT 119.925 61.745 120.095 62.015 ;
        RECT 120.265 61.915 120.595 62.275 ;
        RECT 121.230 61.825 121.890 61.995 ;
        RECT 119.925 61.595 120.530 61.745 ;
        RECT 119.925 61.575 120.730 61.595 ;
        RECT 119.850 61.035 120.180 61.405 ;
        RECT 120.360 61.265 120.730 61.575 ;
        RECT 121.105 61.325 121.485 61.655 ;
        RECT 120.360 60.865 120.530 61.265 ;
        RECT 119.845 60.695 120.530 60.865 ;
        RECT 118.545 59.895 118.715 60.395 ;
        RECT 118.885 59.725 119.215 60.225 ;
        RECT 119.385 59.895 119.610 60.675 ;
        RECT 119.845 59.945 120.175 60.695 ;
        RECT 120.345 59.725 120.660 60.525 ;
        RECT 120.860 60.355 121.145 61.005 ;
        RECT 121.315 60.945 121.485 61.325 ;
        RECT 121.720 61.365 121.890 61.825 ;
        RECT 122.130 61.535 122.460 62.275 ;
        RECT 122.730 61.535 122.950 61.945 ;
        RECT 123.130 61.535 123.415 62.275 ;
        RECT 123.585 61.675 123.835 61.945 ;
        RECT 124.005 61.810 124.265 62.275 ;
        RECT 123.585 61.535 123.870 61.675 ;
        RECT 122.780 61.365 122.950 61.535 ;
        RECT 123.700 61.365 123.870 61.535 ;
        RECT 121.720 61.195 122.590 61.365 ;
        RECT 121.870 61.035 122.590 61.195 ;
        RECT 122.780 61.035 123.530 61.365 ;
        RECT 123.700 61.035 124.265 61.365 ;
        RECT 121.315 60.365 121.655 60.945 ;
        RECT 121.870 60.105 122.040 61.035 ;
        RECT 122.780 60.825 122.950 61.035 ;
        RECT 123.700 60.865 123.870 61.035 ;
        RECT 122.230 60.495 122.950 60.825 ;
        RECT 121.290 59.935 122.040 60.105 ;
        RECT 122.210 59.725 122.510 60.225 ;
        RECT 122.730 59.925 122.950 60.495 ;
        RECT 123.130 59.725 123.415 60.865 ;
        RECT 123.585 60.720 123.870 60.865 ;
        RECT 123.585 59.905 123.835 60.720 ;
        RECT 124.435 60.620 124.955 62.105 ;
        RECT 125.125 61.615 125.465 62.275 ;
        RECT 125.815 61.550 126.105 62.275 ;
        RECT 126.365 61.725 126.535 62.015 ;
        RECT 126.705 61.895 127.035 62.275 ;
        RECT 126.365 61.555 126.970 61.725 ;
        RECT 124.005 59.725 124.265 60.605 ;
        RECT 124.625 59.725 124.955 60.450 ;
        RECT 125.125 59.895 125.645 61.445 ;
        RECT 125.815 59.725 126.105 60.890 ;
        RECT 126.275 60.735 126.520 61.375 ;
        RECT 126.800 61.290 126.970 61.555 ;
        RECT 126.800 60.960 127.030 61.290 ;
        RECT 126.800 60.565 126.970 60.960 ;
        RECT 126.365 60.395 126.970 60.565 ;
        RECT 127.205 60.675 127.375 62.015 ;
        RECT 127.745 61.745 127.915 62.015 ;
        RECT 128.085 61.915 128.415 62.275 ;
        RECT 129.050 61.825 129.710 61.995 ;
        RECT 127.745 61.595 128.350 61.745 ;
        RECT 127.745 61.575 128.550 61.595 ;
        RECT 127.670 61.035 128.000 61.405 ;
        RECT 128.180 61.265 128.550 61.575 ;
        RECT 128.925 61.325 129.305 61.655 ;
        RECT 128.180 60.865 128.350 61.265 ;
        RECT 127.665 60.695 128.350 60.865 ;
        RECT 126.365 59.895 126.535 60.395 ;
        RECT 126.705 59.725 127.035 60.225 ;
        RECT 127.205 59.895 127.430 60.675 ;
        RECT 127.665 59.945 127.995 60.695 ;
        RECT 128.165 59.725 128.480 60.525 ;
        RECT 128.680 60.355 128.965 61.005 ;
        RECT 129.135 60.945 129.305 61.325 ;
        RECT 129.540 61.365 129.710 61.825 ;
        RECT 129.950 61.535 130.280 62.275 ;
        RECT 130.550 61.535 130.770 61.945 ;
        RECT 130.950 61.535 131.235 62.275 ;
        RECT 131.405 61.675 131.655 61.945 ;
        RECT 131.825 61.810 132.085 62.275 ;
        RECT 132.345 61.725 132.515 62.015 ;
        RECT 132.685 61.895 133.015 62.275 ;
        RECT 131.405 61.535 131.690 61.675 ;
        RECT 132.345 61.555 132.950 61.725 ;
        RECT 130.600 61.365 130.770 61.535 ;
        RECT 131.520 61.365 131.690 61.535 ;
        RECT 129.540 61.195 130.410 61.365 ;
        RECT 129.690 61.035 130.410 61.195 ;
        RECT 130.600 61.035 131.350 61.365 ;
        RECT 131.520 61.035 132.085 61.365 ;
        RECT 129.135 60.365 129.475 60.945 ;
        RECT 129.690 60.105 129.860 61.035 ;
        RECT 130.600 60.825 130.770 61.035 ;
        RECT 131.520 60.865 131.690 61.035 ;
        RECT 130.050 60.495 130.770 60.825 ;
        RECT 129.110 59.935 129.860 60.105 ;
        RECT 130.030 59.725 130.330 60.225 ;
        RECT 130.550 59.925 130.770 60.495 ;
        RECT 130.950 59.725 131.235 60.865 ;
        RECT 131.405 60.720 131.690 60.865 ;
        RECT 132.255 60.735 132.500 61.375 ;
        RECT 132.780 61.290 132.950 61.555 ;
        RECT 132.780 60.960 133.010 61.290 ;
        RECT 131.405 59.905 131.655 60.720 ;
        RECT 131.825 59.725 132.085 60.605 ;
        RECT 132.780 60.565 132.950 60.960 ;
        RECT 132.345 60.395 132.950 60.565 ;
        RECT 133.185 60.675 133.355 62.015 ;
        RECT 133.725 61.745 133.895 62.015 ;
        RECT 134.065 61.915 134.395 62.275 ;
        RECT 135.030 61.825 135.690 61.995 ;
        RECT 133.725 61.595 134.330 61.745 ;
        RECT 133.725 61.575 134.530 61.595 ;
        RECT 133.650 61.035 133.980 61.405 ;
        RECT 134.160 61.265 134.530 61.575 ;
        RECT 134.905 61.325 135.285 61.655 ;
        RECT 134.160 60.865 134.330 61.265 ;
        RECT 133.645 60.695 134.330 60.865 ;
        RECT 132.345 59.895 132.515 60.395 ;
        RECT 132.685 59.725 133.015 60.225 ;
        RECT 133.185 59.895 133.410 60.675 ;
        RECT 133.645 59.945 133.975 60.695 ;
        RECT 134.145 59.725 134.460 60.525 ;
        RECT 134.660 60.355 134.945 61.005 ;
        RECT 135.115 60.945 135.285 61.325 ;
        RECT 135.520 61.365 135.690 61.825 ;
        RECT 135.930 61.535 136.260 62.275 ;
        RECT 136.530 61.535 136.750 61.945 ;
        RECT 136.930 61.535 137.215 62.275 ;
        RECT 137.385 61.675 137.635 61.945 ;
        RECT 137.805 61.810 138.065 62.275 ;
        RECT 138.325 61.725 138.495 62.015 ;
        RECT 138.665 61.895 138.995 62.275 ;
        RECT 137.385 61.535 137.670 61.675 ;
        RECT 138.325 61.555 138.930 61.725 ;
        RECT 136.580 61.365 136.750 61.535 ;
        RECT 137.500 61.365 137.670 61.535 ;
        RECT 135.520 61.195 136.390 61.365 ;
        RECT 135.670 61.035 136.390 61.195 ;
        RECT 136.580 61.035 137.330 61.365 ;
        RECT 137.500 61.035 138.065 61.365 ;
        RECT 135.115 60.365 135.455 60.945 ;
        RECT 135.670 60.105 135.840 61.035 ;
        RECT 136.580 60.825 136.750 61.035 ;
        RECT 137.500 60.865 137.670 61.035 ;
        RECT 136.030 60.495 136.750 60.825 ;
        RECT 135.090 59.935 135.840 60.105 ;
        RECT 136.010 59.725 136.310 60.225 ;
        RECT 136.530 59.925 136.750 60.495 ;
        RECT 136.930 59.725 137.215 60.865 ;
        RECT 137.385 60.720 137.670 60.865 ;
        RECT 138.235 60.735 138.480 61.375 ;
        RECT 138.760 61.290 138.930 61.555 ;
        RECT 138.760 60.960 138.990 61.290 ;
        RECT 137.385 59.905 137.635 60.720 ;
        RECT 137.805 59.725 138.065 60.605 ;
        RECT 138.760 60.565 138.930 60.960 ;
        RECT 138.325 60.395 138.930 60.565 ;
        RECT 139.165 60.675 139.335 62.015 ;
        RECT 139.705 61.745 139.875 62.015 ;
        RECT 140.045 61.915 140.375 62.275 ;
        RECT 141.010 61.825 141.670 61.995 ;
        RECT 139.705 61.595 140.310 61.745 ;
        RECT 139.705 61.575 140.510 61.595 ;
        RECT 139.630 61.035 139.960 61.405 ;
        RECT 140.140 61.265 140.510 61.575 ;
        RECT 140.885 61.325 141.265 61.655 ;
        RECT 140.140 60.865 140.310 61.265 ;
        RECT 139.625 60.695 140.310 60.865 ;
        RECT 138.325 59.895 138.495 60.395 ;
        RECT 138.665 59.725 138.995 60.225 ;
        RECT 139.165 59.895 139.390 60.675 ;
        RECT 139.625 59.945 139.955 60.695 ;
        RECT 140.125 59.725 140.440 60.525 ;
        RECT 140.640 60.355 140.925 61.005 ;
        RECT 141.095 60.945 141.265 61.325 ;
        RECT 141.500 61.365 141.670 61.825 ;
        RECT 141.910 61.535 142.240 62.275 ;
        RECT 142.510 61.535 142.730 61.945 ;
        RECT 142.910 61.535 143.195 62.275 ;
        RECT 143.365 61.675 143.615 61.945 ;
        RECT 143.785 61.810 144.045 62.275 ;
        RECT 144.305 61.725 144.475 62.015 ;
        RECT 144.645 61.895 144.975 62.275 ;
        RECT 143.365 61.535 143.650 61.675 ;
        RECT 144.305 61.555 144.910 61.725 ;
        RECT 142.560 61.365 142.730 61.535 ;
        RECT 143.480 61.365 143.650 61.535 ;
        RECT 141.500 61.195 142.370 61.365 ;
        RECT 141.650 61.035 142.370 61.195 ;
        RECT 142.560 61.035 143.310 61.365 ;
        RECT 143.480 61.035 144.045 61.365 ;
        RECT 141.095 60.365 141.435 60.945 ;
        RECT 141.650 60.105 141.820 61.035 ;
        RECT 142.560 60.825 142.730 61.035 ;
        RECT 143.480 60.865 143.650 61.035 ;
        RECT 142.010 60.495 142.730 60.825 ;
        RECT 141.070 59.935 141.820 60.105 ;
        RECT 141.990 59.725 142.290 60.225 ;
        RECT 142.510 59.925 142.730 60.495 ;
        RECT 142.910 59.725 143.195 60.865 ;
        RECT 143.365 60.720 143.650 60.865 ;
        RECT 144.215 60.735 144.460 61.375 ;
        RECT 144.740 61.290 144.910 61.555 ;
        RECT 144.740 60.960 144.970 61.290 ;
        RECT 143.365 59.905 143.615 60.720 ;
        RECT 143.785 59.725 144.045 60.605 ;
        RECT 144.740 60.565 144.910 60.960 ;
        RECT 144.305 60.395 144.910 60.565 ;
        RECT 145.145 60.675 145.315 62.015 ;
        RECT 145.685 61.745 145.855 62.015 ;
        RECT 146.025 61.915 146.355 62.275 ;
        RECT 146.990 61.825 147.650 61.995 ;
        RECT 145.685 61.595 146.290 61.745 ;
        RECT 145.685 61.575 146.490 61.595 ;
        RECT 145.610 61.035 145.940 61.405 ;
        RECT 146.120 61.265 146.490 61.575 ;
        RECT 146.865 61.325 147.245 61.655 ;
        RECT 146.120 60.865 146.290 61.265 ;
        RECT 145.605 60.695 146.290 60.865 ;
        RECT 144.305 59.895 144.475 60.395 ;
        RECT 144.645 59.725 144.975 60.225 ;
        RECT 145.145 59.895 145.370 60.675 ;
        RECT 145.605 59.945 145.935 60.695 ;
        RECT 146.105 59.725 146.420 60.525 ;
        RECT 146.620 60.355 146.905 61.005 ;
        RECT 147.075 60.945 147.245 61.325 ;
        RECT 147.480 61.365 147.650 61.825 ;
        RECT 147.890 61.535 148.220 62.275 ;
        RECT 148.490 61.535 148.710 61.945 ;
        RECT 148.890 61.535 149.175 62.275 ;
        RECT 149.345 61.675 149.595 61.945 ;
        RECT 149.765 61.810 150.025 62.275 ;
        RECT 149.345 61.535 149.630 61.675 ;
        RECT 148.540 61.365 148.710 61.535 ;
        RECT 149.460 61.365 149.630 61.535 ;
        RECT 150.195 61.525 151.405 62.275 ;
        RECT 151.575 61.550 151.865 62.275 ;
        RECT 147.480 61.195 148.350 61.365 ;
        RECT 147.630 61.035 148.350 61.195 ;
        RECT 148.540 61.035 149.290 61.365 ;
        RECT 149.460 61.035 150.025 61.365 ;
        RECT 147.075 60.365 147.415 60.945 ;
        RECT 147.630 60.105 147.800 61.035 ;
        RECT 148.540 60.825 148.710 61.035 ;
        RECT 149.460 60.865 149.630 61.035 ;
        RECT 150.195 60.985 150.715 61.525 ;
        RECT 152.035 61.505 155.545 62.275 ;
        RECT 155.715 61.525 156.925 62.275 ;
        RECT 147.990 60.495 148.710 60.825 ;
        RECT 147.050 59.935 147.800 60.105 ;
        RECT 147.970 59.725 148.270 60.225 ;
        RECT 148.490 59.925 148.710 60.495 ;
        RECT 148.890 59.725 149.175 60.865 ;
        RECT 149.345 60.720 149.630 60.865 ;
        RECT 150.885 60.815 151.405 61.355 ;
        RECT 152.035 60.985 153.685 61.505 ;
        RECT 149.345 59.905 149.595 60.720 ;
        RECT 149.765 59.725 150.025 60.605 ;
        RECT 150.195 59.725 151.405 60.815 ;
        RECT 151.575 59.725 151.865 60.890 ;
        RECT 153.855 60.815 155.545 61.335 ;
        RECT 152.035 59.725 155.545 60.815 ;
        RECT 155.715 60.815 156.235 61.355 ;
        RECT 156.405 60.985 156.925 61.525 ;
        RECT 155.715 59.725 156.925 60.815 ;
        RECT 22.690 59.555 157.010 59.725 ;
        RECT 22.775 58.465 23.985 59.555 ;
        RECT 24.705 58.885 24.875 59.385 ;
        RECT 25.045 59.055 25.375 59.555 ;
        RECT 24.705 58.715 25.310 58.885 ;
        RECT 22.775 57.755 23.295 58.295 ;
        RECT 23.465 57.925 23.985 58.465 ;
        RECT 24.615 57.905 24.860 58.545 ;
        RECT 25.140 58.320 25.310 58.715 ;
        RECT 25.545 58.605 25.770 59.385 ;
        RECT 25.140 57.990 25.370 58.320 ;
        RECT 22.775 57.005 23.985 57.755 ;
        RECT 25.140 57.725 25.310 57.990 ;
        RECT 24.705 57.555 25.310 57.725 ;
        RECT 24.705 57.265 24.875 57.555 ;
        RECT 25.045 57.005 25.375 57.385 ;
        RECT 25.545 57.265 25.715 58.605 ;
        RECT 26.005 58.585 26.335 59.335 ;
        RECT 26.505 58.755 26.820 59.555 ;
        RECT 27.450 59.175 28.200 59.345 ;
        RECT 26.005 58.415 26.690 58.585 ;
        RECT 26.010 57.875 26.340 58.245 ;
        RECT 26.520 58.015 26.690 58.415 ;
        RECT 27.020 58.275 27.305 58.925 ;
        RECT 27.475 58.335 27.815 58.915 ;
        RECT 26.520 57.705 26.890 58.015 ;
        RECT 27.475 57.955 27.645 58.335 ;
        RECT 28.030 58.245 28.200 59.175 ;
        RECT 28.370 59.055 28.670 59.555 ;
        RECT 28.890 58.785 29.110 59.355 ;
        RECT 28.390 58.455 29.110 58.785 ;
        RECT 28.940 58.245 29.110 58.455 ;
        RECT 29.290 58.415 29.575 59.555 ;
        RECT 29.745 58.560 29.995 59.375 ;
        RECT 30.165 58.675 30.425 59.555 ;
        RECT 29.745 58.415 30.030 58.560 ;
        RECT 29.860 58.245 30.030 58.415 ;
        RECT 28.030 58.085 28.750 58.245 ;
        RECT 26.085 57.685 26.890 57.705 ;
        RECT 26.085 57.535 26.690 57.685 ;
        RECT 27.265 57.625 27.645 57.955 ;
        RECT 27.880 57.915 28.750 58.085 ;
        RECT 28.940 57.915 29.690 58.245 ;
        RECT 29.860 57.915 30.425 58.245 ;
        RECT 26.085 57.265 26.255 57.535 ;
        RECT 27.880 57.455 28.050 57.915 ;
        RECT 28.940 57.745 29.110 57.915 ;
        RECT 29.860 57.745 30.030 57.915 ;
        RECT 31.055 57.835 31.575 59.385 ;
        RECT 31.745 58.830 32.075 59.555 ;
        RECT 26.425 57.005 26.755 57.365 ;
        RECT 27.390 57.285 28.050 57.455 ;
        RECT 28.290 57.005 28.620 57.745 ;
        RECT 28.890 57.335 29.110 57.745 ;
        RECT 29.290 57.005 29.575 57.745 ;
        RECT 29.745 57.605 30.030 57.745 ;
        RECT 29.745 57.335 29.995 57.605 ;
        RECT 30.165 57.005 30.425 57.470 ;
        RECT 31.235 57.005 31.575 57.665 ;
        RECT 31.745 57.175 32.265 58.660 ;
        RECT 32.435 58.465 34.105 59.555 ;
        RECT 34.465 58.830 34.795 59.555 ;
        RECT 32.435 57.775 33.185 58.295 ;
        RECT 33.355 57.945 34.105 58.465 ;
        RECT 32.435 57.005 34.105 57.775 ;
        RECT 34.275 57.175 34.795 58.660 ;
        RECT 34.965 57.835 35.485 59.385 ;
        RECT 35.655 58.390 35.945 59.555 ;
        RECT 36.205 58.885 36.375 59.385 ;
        RECT 36.545 59.055 36.875 59.555 ;
        RECT 36.205 58.715 36.810 58.885 ;
        RECT 36.115 57.905 36.360 58.545 ;
        RECT 36.640 58.320 36.810 58.715 ;
        RECT 37.045 58.605 37.270 59.385 ;
        RECT 36.640 57.990 36.870 58.320 ;
        RECT 34.965 57.005 35.305 57.665 ;
        RECT 35.655 57.005 35.945 57.730 ;
        RECT 36.640 57.725 36.810 57.990 ;
        RECT 36.205 57.555 36.810 57.725 ;
        RECT 36.205 57.265 36.375 57.555 ;
        RECT 36.545 57.005 36.875 57.385 ;
        RECT 37.045 57.265 37.215 58.605 ;
        RECT 37.505 58.585 37.835 59.335 ;
        RECT 38.005 58.755 38.320 59.555 ;
        RECT 38.950 59.175 39.700 59.345 ;
        RECT 37.505 58.415 38.190 58.585 ;
        RECT 37.510 57.875 37.840 58.245 ;
        RECT 38.020 58.015 38.190 58.415 ;
        RECT 38.520 58.275 38.805 58.925 ;
        RECT 38.975 58.335 39.315 58.915 ;
        RECT 38.020 57.705 38.390 58.015 ;
        RECT 38.975 57.955 39.145 58.335 ;
        RECT 39.530 58.245 39.700 59.175 ;
        RECT 39.870 59.055 40.170 59.555 ;
        RECT 40.390 58.785 40.610 59.355 ;
        RECT 39.890 58.455 40.610 58.785 ;
        RECT 40.440 58.245 40.610 58.455 ;
        RECT 40.790 58.415 41.075 59.555 ;
        RECT 41.245 58.560 41.495 59.375 ;
        RECT 41.665 58.675 41.925 59.555 ;
        RECT 42.185 58.885 42.355 59.385 ;
        RECT 42.525 59.055 42.855 59.555 ;
        RECT 42.185 58.715 42.790 58.885 ;
        RECT 41.245 58.415 41.530 58.560 ;
        RECT 41.360 58.245 41.530 58.415 ;
        RECT 39.530 58.085 40.250 58.245 ;
        RECT 37.585 57.685 38.390 57.705 ;
        RECT 37.585 57.535 38.190 57.685 ;
        RECT 38.765 57.625 39.145 57.955 ;
        RECT 39.380 57.915 40.250 58.085 ;
        RECT 40.440 57.915 41.190 58.245 ;
        RECT 41.360 57.915 41.925 58.245 ;
        RECT 37.585 57.265 37.755 57.535 ;
        RECT 39.380 57.455 39.550 57.915 ;
        RECT 40.440 57.745 40.610 57.915 ;
        RECT 41.360 57.745 41.530 57.915 ;
        RECT 42.095 57.905 42.340 58.545 ;
        RECT 42.620 58.320 42.790 58.715 ;
        RECT 43.025 58.605 43.250 59.385 ;
        RECT 42.620 57.990 42.850 58.320 ;
        RECT 37.925 57.005 38.255 57.365 ;
        RECT 38.890 57.285 39.550 57.455 ;
        RECT 39.790 57.005 40.120 57.745 ;
        RECT 40.390 57.335 40.610 57.745 ;
        RECT 40.790 57.005 41.075 57.745 ;
        RECT 41.245 57.605 41.530 57.745 ;
        RECT 42.620 57.725 42.790 57.990 ;
        RECT 41.245 57.335 41.495 57.605 ;
        RECT 42.185 57.555 42.790 57.725 ;
        RECT 41.665 57.005 41.925 57.470 ;
        RECT 42.185 57.265 42.355 57.555 ;
        RECT 42.525 57.005 42.855 57.385 ;
        RECT 43.025 57.265 43.195 58.605 ;
        RECT 43.485 58.585 43.815 59.335 ;
        RECT 43.985 58.755 44.300 59.555 ;
        RECT 44.930 59.175 45.680 59.345 ;
        RECT 43.485 58.415 44.170 58.585 ;
        RECT 43.490 57.875 43.820 58.245 ;
        RECT 44.000 58.015 44.170 58.415 ;
        RECT 44.500 58.275 44.785 58.925 ;
        RECT 44.955 58.335 45.295 58.915 ;
        RECT 44.000 57.705 44.370 58.015 ;
        RECT 44.955 57.955 45.125 58.335 ;
        RECT 45.510 58.245 45.680 59.175 ;
        RECT 45.850 59.055 46.150 59.555 ;
        RECT 46.370 58.785 46.590 59.355 ;
        RECT 45.870 58.455 46.590 58.785 ;
        RECT 46.420 58.245 46.590 58.455 ;
        RECT 46.770 58.415 47.055 59.555 ;
        RECT 47.225 58.560 47.475 59.375 ;
        RECT 47.645 58.675 47.905 59.555 ;
        RECT 47.225 58.415 47.510 58.560 ;
        RECT 47.340 58.245 47.510 58.415 ;
        RECT 48.535 58.390 48.825 59.555 ;
        RECT 49.545 58.885 49.715 59.385 ;
        RECT 49.885 59.055 50.215 59.555 ;
        RECT 49.545 58.715 50.150 58.885 ;
        RECT 45.510 58.085 46.230 58.245 ;
        RECT 43.565 57.685 44.370 57.705 ;
        RECT 43.565 57.535 44.170 57.685 ;
        RECT 44.745 57.625 45.125 57.955 ;
        RECT 45.360 57.915 46.230 58.085 ;
        RECT 46.420 57.915 47.170 58.245 ;
        RECT 47.340 57.915 47.905 58.245 ;
        RECT 43.565 57.265 43.735 57.535 ;
        RECT 45.360 57.455 45.530 57.915 ;
        RECT 46.420 57.745 46.590 57.915 ;
        RECT 47.340 57.745 47.510 57.915 ;
        RECT 49.455 57.905 49.700 58.545 ;
        RECT 49.980 58.320 50.150 58.715 ;
        RECT 50.385 58.605 50.610 59.385 ;
        RECT 49.980 57.990 50.210 58.320 ;
        RECT 43.905 57.005 44.235 57.365 ;
        RECT 44.870 57.285 45.530 57.455 ;
        RECT 45.770 57.005 46.100 57.745 ;
        RECT 46.370 57.335 46.590 57.745 ;
        RECT 46.770 57.005 47.055 57.745 ;
        RECT 47.225 57.605 47.510 57.745 ;
        RECT 47.225 57.335 47.475 57.605 ;
        RECT 47.645 57.005 47.905 57.470 ;
        RECT 48.535 57.005 48.825 57.730 ;
        RECT 49.980 57.725 50.150 57.990 ;
        RECT 49.545 57.555 50.150 57.725 ;
        RECT 49.545 57.265 49.715 57.555 ;
        RECT 49.885 57.005 50.215 57.385 ;
        RECT 50.385 57.265 50.555 58.605 ;
        RECT 50.845 58.585 51.175 59.335 ;
        RECT 51.345 58.755 51.660 59.555 ;
        RECT 52.290 59.175 53.040 59.345 ;
        RECT 50.845 58.415 51.530 58.585 ;
        RECT 50.850 57.875 51.180 58.245 ;
        RECT 51.360 58.015 51.530 58.415 ;
        RECT 51.860 58.275 52.145 58.925 ;
        RECT 52.315 58.335 52.655 58.915 ;
        RECT 51.360 57.705 51.730 58.015 ;
        RECT 52.315 57.955 52.485 58.335 ;
        RECT 52.870 58.245 53.040 59.175 ;
        RECT 53.210 59.055 53.510 59.555 ;
        RECT 53.730 58.785 53.950 59.355 ;
        RECT 53.230 58.455 53.950 58.785 ;
        RECT 53.780 58.245 53.950 58.455 ;
        RECT 54.130 58.415 54.415 59.555 ;
        RECT 54.585 58.560 54.835 59.375 ;
        RECT 55.005 58.675 55.265 59.555 ;
        RECT 55.525 58.885 55.695 59.385 ;
        RECT 55.865 59.055 56.195 59.555 ;
        RECT 55.525 58.715 56.130 58.885 ;
        RECT 54.585 58.415 54.870 58.560 ;
        RECT 54.700 58.245 54.870 58.415 ;
        RECT 52.870 58.085 53.590 58.245 ;
        RECT 50.925 57.685 51.730 57.705 ;
        RECT 50.925 57.535 51.530 57.685 ;
        RECT 52.105 57.625 52.485 57.955 ;
        RECT 52.720 57.915 53.590 58.085 ;
        RECT 53.780 57.915 54.530 58.245 ;
        RECT 54.700 57.915 55.265 58.245 ;
        RECT 50.925 57.265 51.095 57.535 ;
        RECT 52.720 57.455 52.890 57.915 ;
        RECT 53.780 57.745 53.950 57.915 ;
        RECT 54.700 57.745 54.870 57.915 ;
        RECT 55.435 57.905 55.680 58.545 ;
        RECT 55.960 58.320 56.130 58.715 ;
        RECT 56.365 58.605 56.590 59.385 ;
        RECT 55.960 57.990 56.190 58.320 ;
        RECT 51.265 57.005 51.595 57.365 ;
        RECT 52.230 57.285 52.890 57.455 ;
        RECT 53.130 57.005 53.460 57.745 ;
        RECT 53.730 57.335 53.950 57.745 ;
        RECT 54.130 57.005 54.415 57.745 ;
        RECT 54.585 57.605 54.870 57.745 ;
        RECT 55.960 57.725 56.130 57.990 ;
        RECT 54.585 57.335 54.835 57.605 ;
        RECT 55.525 57.555 56.130 57.725 ;
        RECT 55.005 57.005 55.265 57.470 ;
        RECT 55.525 57.265 55.695 57.555 ;
        RECT 55.865 57.005 56.195 57.385 ;
        RECT 56.365 57.265 56.535 58.605 ;
        RECT 56.825 58.585 57.155 59.335 ;
        RECT 57.325 58.755 57.640 59.555 ;
        RECT 58.270 59.175 59.020 59.345 ;
        RECT 56.825 58.415 57.510 58.585 ;
        RECT 56.830 57.875 57.160 58.245 ;
        RECT 57.340 58.015 57.510 58.415 ;
        RECT 57.840 58.275 58.125 58.925 ;
        RECT 58.295 58.335 58.635 58.915 ;
        RECT 57.340 57.705 57.710 58.015 ;
        RECT 58.295 57.955 58.465 58.335 ;
        RECT 58.850 58.245 59.020 59.175 ;
        RECT 59.190 59.055 59.490 59.555 ;
        RECT 59.710 58.785 59.930 59.355 ;
        RECT 59.210 58.455 59.930 58.785 ;
        RECT 59.760 58.245 59.930 58.455 ;
        RECT 60.110 58.415 60.395 59.555 ;
        RECT 60.565 58.560 60.815 59.375 ;
        RECT 60.985 58.675 61.245 59.555 ;
        RECT 60.565 58.415 60.850 58.560 ;
        RECT 60.680 58.245 60.850 58.415 ;
        RECT 61.415 58.390 61.705 59.555 ;
        RECT 58.850 58.085 59.570 58.245 ;
        RECT 56.905 57.685 57.710 57.705 ;
        RECT 56.905 57.535 57.510 57.685 ;
        RECT 58.085 57.625 58.465 57.955 ;
        RECT 58.700 57.915 59.570 58.085 ;
        RECT 59.760 57.915 60.510 58.245 ;
        RECT 60.680 57.915 61.245 58.245 ;
        RECT 56.905 57.265 57.075 57.535 ;
        RECT 58.700 57.455 58.870 57.915 ;
        RECT 59.760 57.745 59.930 57.915 ;
        RECT 60.680 57.745 60.850 57.915 ;
        RECT 61.875 57.835 62.395 59.385 ;
        RECT 62.565 58.830 62.895 59.555 ;
        RECT 57.245 57.005 57.575 57.365 ;
        RECT 58.210 57.285 58.870 57.455 ;
        RECT 59.110 57.005 59.440 57.745 ;
        RECT 59.710 57.335 59.930 57.745 ;
        RECT 60.110 57.005 60.395 57.745 ;
        RECT 60.565 57.605 60.850 57.745 ;
        RECT 60.565 57.335 60.815 57.605 ;
        RECT 60.985 57.005 61.245 57.470 ;
        RECT 61.415 57.005 61.705 57.730 ;
        RECT 62.055 57.005 62.395 57.665 ;
        RECT 62.565 57.175 63.085 58.660 ;
        RECT 63.255 58.465 65.845 59.555 ;
        RECT 66.105 58.885 66.275 59.385 ;
        RECT 66.445 59.055 66.775 59.555 ;
        RECT 66.105 58.715 66.710 58.885 ;
        RECT 63.255 57.775 64.465 58.295 ;
        RECT 64.635 57.945 65.845 58.465 ;
        RECT 66.015 57.905 66.260 58.545 ;
        RECT 66.540 58.320 66.710 58.715 ;
        RECT 66.945 58.605 67.170 59.385 ;
        RECT 66.540 57.990 66.770 58.320 ;
        RECT 63.255 57.005 65.845 57.775 ;
        RECT 66.540 57.725 66.710 57.990 ;
        RECT 66.105 57.555 66.710 57.725 ;
        RECT 66.105 57.265 66.275 57.555 ;
        RECT 66.445 57.005 66.775 57.385 ;
        RECT 66.945 57.265 67.115 58.605 ;
        RECT 67.405 58.585 67.735 59.335 ;
        RECT 67.905 58.755 68.220 59.555 ;
        RECT 68.850 59.175 69.600 59.345 ;
        RECT 67.405 58.415 68.090 58.585 ;
        RECT 67.410 57.875 67.740 58.245 ;
        RECT 67.920 58.015 68.090 58.415 ;
        RECT 68.420 58.275 68.705 58.925 ;
        RECT 68.875 58.335 69.215 58.915 ;
        RECT 67.920 57.705 68.290 58.015 ;
        RECT 68.875 57.955 69.045 58.335 ;
        RECT 69.430 58.245 69.600 59.175 ;
        RECT 69.770 59.055 70.070 59.555 ;
        RECT 70.290 58.785 70.510 59.355 ;
        RECT 69.790 58.455 70.510 58.785 ;
        RECT 70.340 58.245 70.510 58.455 ;
        RECT 70.690 58.415 70.975 59.555 ;
        RECT 71.145 58.560 71.395 59.375 ;
        RECT 71.565 58.675 71.825 59.555 ;
        RECT 71.145 58.415 71.430 58.560 ;
        RECT 71.260 58.245 71.430 58.415 ;
        RECT 69.430 58.085 70.150 58.245 ;
        RECT 67.485 57.685 68.290 57.705 ;
        RECT 67.485 57.535 68.090 57.685 ;
        RECT 68.665 57.625 69.045 57.955 ;
        RECT 69.280 57.915 70.150 58.085 ;
        RECT 70.340 57.915 71.090 58.245 ;
        RECT 71.260 57.915 71.825 58.245 ;
        RECT 67.485 57.265 67.655 57.535 ;
        RECT 69.280 57.455 69.450 57.915 ;
        RECT 70.340 57.745 70.510 57.915 ;
        RECT 71.260 57.745 71.430 57.915 ;
        RECT 72.915 57.835 73.435 59.385 ;
        RECT 73.605 58.830 73.935 59.555 ;
        RECT 67.825 57.005 68.155 57.365 ;
        RECT 68.790 57.285 69.450 57.455 ;
        RECT 69.690 57.005 70.020 57.745 ;
        RECT 70.290 57.335 70.510 57.745 ;
        RECT 70.690 57.005 70.975 57.745 ;
        RECT 71.145 57.605 71.430 57.745 ;
        RECT 71.145 57.335 71.395 57.605 ;
        RECT 71.565 57.005 71.825 57.470 ;
        RECT 73.095 57.005 73.435 57.665 ;
        RECT 73.605 57.175 74.125 58.660 ;
        RECT 74.295 58.390 74.585 59.555 ;
        RECT 74.755 58.465 75.965 59.555 ;
        RECT 74.755 57.755 75.275 58.295 ;
        RECT 75.445 57.925 75.965 58.465 ;
        RECT 76.135 57.835 76.655 59.385 ;
        RECT 76.825 58.830 77.155 59.555 ;
        RECT 74.295 57.005 74.585 57.730 ;
        RECT 74.755 57.005 75.965 57.755 ;
        RECT 76.315 57.005 76.655 57.665 ;
        RECT 76.825 57.175 77.345 58.660 ;
        RECT 78.435 57.835 78.955 59.385 ;
        RECT 79.125 58.830 79.455 59.555 ;
        RECT 78.615 57.005 78.955 57.665 ;
        RECT 79.125 57.175 79.645 58.660 ;
        RECT 79.815 58.465 81.025 59.555 ;
        RECT 81.285 58.885 81.455 59.385 ;
        RECT 81.625 59.055 81.955 59.555 ;
        RECT 81.285 58.715 81.890 58.885 ;
        RECT 79.815 57.755 80.335 58.295 ;
        RECT 80.505 57.925 81.025 58.465 ;
        RECT 81.195 57.905 81.440 58.545 ;
        RECT 81.720 58.320 81.890 58.715 ;
        RECT 82.125 58.605 82.350 59.385 ;
        RECT 81.720 57.990 81.950 58.320 ;
        RECT 79.815 57.005 81.025 57.755 ;
        RECT 81.720 57.725 81.890 57.990 ;
        RECT 81.285 57.555 81.890 57.725 ;
        RECT 81.285 57.265 81.455 57.555 ;
        RECT 81.625 57.005 81.955 57.385 ;
        RECT 82.125 57.265 82.295 58.605 ;
        RECT 82.585 58.585 82.915 59.335 ;
        RECT 83.085 58.755 83.400 59.555 ;
        RECT 84.030 59.175 84.780 59.345 ;
        RECT 82.585 58.415 83.270 58.585 ;
        RECT 82.590 57.875 82.920 58.245 ;
        RECT 83.100 58.015 83.270 58.415 ;
        RECT 83.600 58.275 83.885 58.925 ;
        RECT 84.055 58.335 84.395 58.915 ;
        RECT 83.100 57.705 83.470 58.015 ;
        RECT 84.055 57.955 84.225 58.335 ;
        RECT 84.610 58.245 84.780 59.175 ;
        RECT 84.950 59.055 85.250 59.555 ;
        RECT 85.470 58.785 85.690 59.355 ;
        RECT 84.970 58.455 85.690 58.785 ;
        RECT 85.520 58.245 85.690 58.455 ;
        RECT 85.870 58.415 86.155 59.555 ;
        RECT 86.325 58.560 86.575 59.375 ;
        RECT 86.745 58.675 87.005 59.555 ;
        RECT 86.325 58.415 86.610 58.560 ;
        RECT 86.440 58.245 86.610 58.415 ;
        RECT 87.175 58.390 87.465 59.555 ;
        RECT 84.610 58.085 85.330 58.245 ;
        RECT 82.665 57.685 83.470 57.705 ;
        RECT 82.665 57.535 83.270 57.685 ;
        RECT 83.845 57.625 84.225 57.955 ;
        RECT 84.460 57.915 85.330 58.085 ;
        RECT 85.520 57.915 86.270 58.245 ;
        RECT 86.440 57.915 87.005 58.245 ;
        RECT 82.665 57.265 82.835 57.535 ;
        RECT 84.460 57.455 84.630 57.915 ;
        RECT 85.520 57.745 85.690 57.915 ;
        RECT 86.440 57.745 86.610 57.915 ;
        RECT 87.635 57.835 88.155 59.385 ;
        RECT 88.325 58.830 88.655 59.555 ;
        RECT 83.005 57.005 83.335 57.365 ;
        RECT 83.970 57.285 84.630 57.455 ;
        RECT 84.870 57.005 85.200 57.745 ;
        RECT 85.470 57.335 85.690 57.745 ;
        RECT 85.870 57.005 86.155 57.745 ;
        RECT 86.325 57.605 86.610 57.745 ;
        RECT 86.325 57.335 86.575 57.605 ;
        RECT 86.745 57.005 87.005 57.470 ;
        RECT 87.175 57.005 87.465 57.730 ;
        RECT 87.815 57.005 88.155 57.665 ;
        RECT 88.325 57.175 88.845 58.660 ;
        RECT 89.015 58.465 90.225 59.555 ;
        RECT 90.485 58.885 90.655 59.385 ;
        RECT 90.825 59.055 91.155 59.555 ;
        RECT 90.485 58.715 91.090 58.885 ;
        RECT 89.015 57.755 89.535 58.295 ;
        RECT 89.705 57.925 90.225 58.465 ;
        RECT 90.395 57.905 90.640 58.545 ;
        RECT 90.920 58.320 91.090 58.715 ;
        RECT 91.325 58.605 91.550 59.385 ;
        RECT 90.920 57.990 91.150 58.320 ;
        RECT 89.015 57.005 90.225 57.755 ;
        RECT 90.920 57.725 91.090 57.990 ;
        RECT 90.485 57.555 91.090 57.725 ;
        RECT 90.485 57.265 90.655 57.555 ;
        RECT 90.825 57.005 91.155 57.385 ;
        RECT 91.325 57.265 91.495 58.605 ;
        RECT 91.785 58.585 92.115 59.335 ;
        RECT 92.285 58.755 92.600 59.555 ;
        RECT 93.230 59.175 93.980 59.345 ;
        RECT 91.785 58.415 92.470 58.585 ;
        RECT 91.790 57.875 92.120 58.245 ;
        RECT 92.300 58.015 92.470 58.415 ;
        RECT 92.800 58.275 93.085 58.925 ;
        RECT 93.255 58.335 93.595 58.915 ;
        RECT 92.300 57.705 92.670 58.015 ;
        RECT 93.255 57.955 93.425 58.335 ;
        RECT 93.810 58.245 93.980 59.175 ;
        RECT 94.150 59.055 94.450 59.555 ;
        RECT 94.670 58.785 94.890 59.355 ;
        RECT 94.170 58.455 94.890 58.785 ;
        RECT 94.720 58.245 94.890 58.455 ;
        RECT 95.070 58.415 95.355 59.555 ;
        RECT 95.525 58.560 95.775 59.375 ;
        RECT 95.945 58.675 96.205 59.555 ;
        RECT 95.525 58.415 95.810 58.560 ;
        RECT 96.375 58.465 97.585 59.555 ;
        RECT 97.945 58.830 98.275 59.555 ;
        RECT 95.640 58.245 95.810 58.415 ;
        RECT 93.810 58.085 94.530 58.245 ;
        RECT 91.865 57.685 92.670 57.705 ;
        RECT 91.865 57.535 92.470 57.685 ;
        RECT 93.045 57.625 93.425 57.955 ;
        RECT 93.660 57.915 94.530 58.085 ;
        RECT 94.720 57.915 95.470 58.245 ;
        RECT 95.640 57.915 96.205 58.245 ;
        RECT 91.865 57.265 92.035 57.535 ;
        RECT 93.660 57.455 93.830 57.915 ;
        RECT 94.720 57.745 94.890 57.915 ;
        RECT 95.640 57.745 95.810 57.915 ;
        RECT 92.205 57.005 92.535 57.365 ;
        RECT 93.170 57.285 93.830 57.455 ;
        RECT 94.070 57.005 94.400 57.745 ;
        RECT 94.670 57.335 94.890 57.745 ;
        RECT 95.070 57.005 95.355 57.745 ;
        RECT 95.525 57.605 95.810 57.745 ;
        RECT 96.375 57.755 96.895 58.295 ;
        RECT 97.065 57.925 97.585 58.465 ;
        RECT 95.525 57.335 95.775 57.605 ;
        RECT 95.945 57.005 96.205 57.470 ;
        RECT 96.375 57.005 97.585 57.755 ;
        RECT 97.755 57.175 98.275 58.660 ;
        RECT 98.445 57.835 98.965 59.385 ;
        RECT 100.055 58.390 100.345 59.555 ;
        RECT 101.065 58.885 101.235 59.385 ;
        RECT 101.405 59.055 101.735 59.555 ;
        RECT 101.065 58.715 101.670 58.885 ;
        RECT 100.975 57.905 101.220 58.545 ;
        RECT 101.500 58.320 101.670 58.715 ;
        RECT 101.905 58.605 102.130 59.385 ;
        RECT 101.500 57.990 101.730 58.320 ;
        RECT 98.445 57.005 98.785 57.665 ;
        RECT 100.055 57.005 100.345 57.730 ;
        RECT 101.500 57.725 101.670 57.990 ;
        RECT 101.065 57.555 101.670 57.725 ;
        RECT 101.065 57.265 101.235 57.555 ;
        RECT 101.405 57.005 101.735 57.385 ;
        RECT 101.905 57.265 102.075 58.605 ;
        RECT 102.365 58.585 102.695 59.335 ;
        RECT 102.865 58.755 103.180 59.555 ;
        RECT 103.810 59.175 104.560 59.345 ;
        RECT 102.365 58.415 103.050 58.585 ;
        RECT 102.370 57.875 102.700 58.245 ;
        RECT 102.880 58.015 103.050 58.415 ;
        RECT 103.380 58.275 103.665 58.925 ;
        RECT 103.835 58.335 104.175 58.915 ;
        RECT 102.880 57.705 103.250 58.015 ;
        RECT 103.835 57.955 104.005 58.335 ;
        RECT 104.390 58.245 104.560 59.175 ;
        RECT 104.730 59.055 105.030 59.555 ;
        RECT 105.250 58.785 105.470 59.355 ;
        RECT 104.750 58.455 105.470 58.785 ;
        RECT 105.300 58.245 105.470 58.455 ;
        RECT 105.650 58.415 105.935 59.555 ;
        RECT 106.105 58.560 106.355 59.375 ;
        RECT 106.525 58.675 106.785 59.555 ;
        RECT 106.105 58.415 106.390 58.560 ;
        RECT 106.955 58.465 108.165 59.555 ;
        RECT 108.525 58.830 108.855 59.555 ;
        RECT 106.220 58.245 106.390 58.415 ;
        RECT 104.390 58.085 105.110 58.245 ;
        RECT 102.445 57.685 103.250 57.705 ;
        RECT 102.445 57.535 103.050 57.685 ;
        RECT 103.625 57.625 104.005 57.955 ;
        RECT 104.240 57.915 105.110 58.085 ;
        RECT 105.300 57.915 106.050 58.245 ;
        RECT 106.220 57.915 106.785 58.245 ;
        RECT 102.445 57.265 102.615 57.535 ;
        RECT 104.240 57.455 104.410 57.915 ;
        RECT 105.300 57.745 105.470 57.915 ;
        RECT 106.220 57.745 106.390 57.915 ;
        RECT 102.785 57.005 103.115 57.365 ;
        RECT 103.750 57.285 104.410 57.455 ;
        RECT 104.650 57.005 104.980 57.745 ;
        RECT 105.250 57.335 105.470 57.745 ;
        RECT 105.650 57.005 105.935 57.745 ;
        RECT 106.105 57.605 106.390 57.745 ;
        RECT 106.955 57.755 107.475 58.295 ;
        RECT 107.645 57.925 108.165 58.465 ;
        RECT 106.105 57.335 106.355 57.605 ;
        RECT 106.525 57.005 106.785 57.470 ;
        RECT 106.955 57.005 108.165 57.755 ;
        RECT 108.335 57.175 108.855 58.660 ;
        RECT 109.025 57.835 109.545 59.385 ;
        RECT 110.365 58.830 110.695 59.555 ;
        RECT 109.025 57.005 109.365 57.665 ;
        RECT 110.175 57.175 110.695 58.660 ;
        RECT 110.865 57.835 111.385 59.385 ;
        RECT 111.745 58.830 112.075 59.555 ;
        RECT 110.865 57.005 111.205 57.665 ;
        RECT 111.555 57.175 112.075 58.660 ;
        RECT 112.245 57.835 112.765 59.385 ;
        RECT 112.935 58.390 113.225 59.555 ;
        RECT 113.485 58.885 113.655 59.385 ;
        RECT 113.825 59.055 114.155 59.555 ;
        RECT 113.485 58.715 114.090 58.885 ;
        RECT 113.395 57.905 113.640 58.545 ;
        RECT 113.920 58.320 114.090 58.715 ;
        RECT 114.325 58.605 114.550 59.385 ;
        RECT 113.920 57.990 114.150 58.320 ;
        RECT 112.245 57.005 112.585 57.665 ;
        RECT 112.935 57.005 113.225 57.730 ;
        RECT 113.920 57.725 114.090 57.990 ;
        RECT 113.485 57.555 114.090 57.725 ;
        RECT 113.485 57.265 113.655 57.555 ;
        RECT 113.825 57.005 114.155 57.385 ;
        RECT 114.325 57.265 114.495 58.605 ;
        RECT 114.785 58.585 115.115 59.335 ;
        RECT 115.285 58.755 115.600 59.555 ;
        RECT 116.230 59.175 116.980 59.345 ;
        RECT 114.785 58.415 115.470 58.585 ;
        RECT 114.790 57.875 115.120 58.245 ;
        RECT 115.300 58.015 115.470 58.415 ;
        RECT 115.800 58.275 116.085 58.925 ;
        RECT 116.255 58.335 116.595 58.915 ;
        RECT 115.300 57.705 115.670 58.015 ;
        RECT 116.255 57.955 116.425 58.335 ;
        RECT 116.810 58.245 116.980 59.175 ;
        RECT 117.150 59.055 117.450 59.555 ;
        RECT 117.670 58.785 117.890 59.355 ;
        RECT 117.170 58.455 117.890 58.785 ;
        RECT 117.720 58.245 117.890 58.455 ;
        RECT 118.070 58.415 118.355 59.555 ;
        RECT 118.525 58.560 118.775 59.375 ;
        RECT 118.945 58.675 119.205 59.555 ;
        RECT 119.375 58.675 119.635 59.555 ;
        RECT 119.805 58.560 120.055 59.375 ;
        RECT 118.525 58.415 118.810 58.560 ;
        RECT 118.640 58.245 118.810 58.415 ;
        RECT 119.770 58.415 120.055 58.560 ;
        RECT 120.225 58.415 120.510 59.555 ;
        RECT 120.690 58.785 120.910 59.355 ;
        RECT 121.130 59.055 121.430 59.555 ;
        RECT 121.600 59.175 122.350 59.345 ;
        RECT 120.690 58.455 121.410 58.785 ;
        RECT 119.770 58.245 119.940 58.415 ;
        RECT 120.690 58.245 120.860 58.455 ;
        RECT 121.600 58.245 121.770 59.175 ;
        RECT 121.985 58.335 122.325 58.915 ;
        RECT 116.810 58.085 117.530 58.245 ;
        RECT 114.865 57.685 115.670 57.705 ;
        RECT 114.865 57.535 115.470 57.685 ;
        RECT 116.045 57.625 116.425 57.955 ;
        RECT 116.660 57.915 117.530 58.085 ;
        RECT 117.720 57.915 118.470 58.245 ;
        RECT 118.640 57.915 119.205 58.245 ;
        RECT 119.375 57.915 119.940 58.245 ;
        RECT 120.110 57.915 120.860 58.245 ;
        RECT 121.050 58.085 121.770 58.245 ;
        RECT 121.050 57.915 121.920 58.085 ;
        RECT 114.865 57.265 115.035 57.535 ;
        RECT 116.660 57.455 116.830 57.915 ;
        RECT 117.720 57.745 117.890 57.915 ;
        RECT 118.640 57.745 118.810 57.915 ;
        RECT 115.205 57.005 115.535 57.365 ;
        RECT 116.170 57.285 116.830 57.455 ;
        RECT 117.070 57.005 117.400 57.745 ;
        RECT 117.670 57.335 117.890 57.745 ;
        RECT 118.070 57.005 118.355 57.745 ;
        RECT 118.525 57.605 118.810 57.745 ;
        RECT 119.770 57.745 119.940 57.915 ;
        RECT 120.690 57.745 120.860 57.915 ;
        RECT 119.770 57.605 120.055 57.745 ;
        RECT 118.525 57.335 118.775 57.605 ;
        RECT 118.945 57.005 119.205 57.470 ;
        RECT 119.375 57.005 119.635 57.470 ;
        RECT 119.805 57.335 120.055 57.605 ;
        RECT 120.225 57.005 120.510 57.745 ;
        RECT 120.690 57.335 120.910 57.745 ;
        RECT 121.180 57.005 121.510 57.745 ;
        RECT 121.750 57.455 121.920 57.915 ;
        RECT 122.155 57.955 122.325 58.335 ;
        RECT 122.495 58.275 122.780 58.925 ;
        RECT 122.980 58.755 123.295 59.555 ;
        RECT 123.465 58.585 123.795 59.335 ;
        RECT 124.030 58.605 124.255 59.385 ;
        RECT 124.425 59.055 124.755 59.555 ;
        RECT 124.925 58.885 125.095 59.385 ;
        RECT 123.110 58.415 123.795 58.585 ;
        RECT 123.110 58.015 123.280 58.415 ;
        RECT 122.155 57.625 122.535 57.955 ;
        RECT 122.910 57.705 123.280 58.015 ;
        RECT 123.460 57.875 123.790 58.245 ;
        RECT 122.910 57.685 123.715 57.705 ;
        RECT 123.110 57.535 123.715 57.685 ;
        RECT 121.750 57.285 122.410 57.455 ;
        RECT 123.045 57.005 123.375 57.365 ;
        RECT 123.545 57.265 123.715 57.535 ;
        RECT 124.085 57.265 124.255 58.605 ;
        RECT 124.490 58.715 125.095 58.885 ;
        RECT 124.490 58.320 124.660 58.715 ;
        RECT 124.430 57.990 124.660 58.320 ;
        RECT 124.490 57.725 124.660 57.990 ;
        RECT 124.940 57.905 125.185 58.545 ;
        RECT 125.815 58.390 126.105 59.555 ;
        RECT 126.365 58.885 126.535 59.385 ;
        RECT 126.705 59.055 127.035 59.555 ;
        RECT 126.365 58.715 126.970 58.885 ;
        RECT 126.275 57.905 126.520 58.545 ;
        RECT 126.800 58.320 126.970 58.715 ;
        RECT 127.205 58.605 127.430 59.385 ;
        RECT 126.800 57.990 127.030 58.320 ;
        RECT 124.490 57.555 125.095 57.725 ;
        RECT 124.425 57.005 124.755 57.385 ;
        RECT 124.925 57.265 125.095 57.555 ;
        RECT 125.815 57.005 126.105 57.730 ;
        RECT 126.800 57.725 126.970 57.990 ;
        RECT 126.365 57.555 126.970 57.725 ;
        RECT 126.365 57.265 126.535 57.555 ;
        RECT 126.705 57.005 127.035 57.385 ;
        RECT 127.205 57.265 127.375 58.605 ;
        RECT 127.665 58.585 127.995 59.335 ;
        RECT 128.165 58.755 128.480 59.555 ;
        RECT 129.110 59.175 129.860 59.345 ;
        RECT 127.665 58.415 128.350 58.585 ;
        RECT 127.670 57.875 128.000 58.245 ;
        RECT 128.180 58.015 128.350 58.415 ;
        RECT 128.680 58.275 128.965 58.925 ;
        RECT 129.135 58.335 129.475 58.915 ;
        RECT 128.180 57.705 128.550 58.015 ;
        RECT 129.135 57.955 129.305 58.335 ;
        RECT 129.690 58.245 129.860 59.175 ;
        RECT 130.030 59.055 130.330 59.555 ;
        RECT 130.550 58.785 130.770 59.355 ;
        RECT 130.050 58.455 130.770 58.785 ;
        RECT 130.600 58.245 130.770 58.455 ;
        RECT 130.950 58.415 131.235 59.555 ;
        RECT 131.405 58.560 131.655 59.375 ;
        RECT 131.825 58.675 132.085 59.555 ;
        RECT 131.405 58.415 131.690 58.560 ;
        RECT 131.520 58.245 131.690 58.415 ;
        RECT 129.690 58.085 130.410 58.245 ;
        RECT 127.745 57.685 128.550 57.705 ;
        RECT 127.745 57.535 128.350 57.685 ;
        RECT 128.925 57.625 129.305 57.955 ;
        RECT 129.540 57.915 130.410 58.085 ;
        RECT 130.600 57.915 131.350 58.245 ;
        RECT 131.520 57.915 132.085 58.245 ;
        RECT 127.745 57.265 127.915 57.535 ;
        RECT 129.540 57.455 129.710 57.915 ;
        RECT 130.600 57.745 130.770 57.915 ;
        RECT 131.520 57.745 131.690 57.915 ;
        RECT 132.255 57.835 132.775 59.385 ;
        RECT 132.945 58.830 133.275 59.555 ;
        RECT 128.085 57.005 128.415 57.365 ;
        RECT 129.050 57.285 129.710 57.455 ;
        RECT 129.950 57.005 130.280 57.745 ;
        RECT 130.550 57.335 130.770 57.745 ;
        RECT 130.950 57.005 131.235 57.745 ;
        RECT 131.405 57.605 131.690 57.745 ;
        RECT 131.405 57.335 131.655 57.605 ;
        RECT 131.825 57.005 132.085 57.470 ;
        RECT 132.435 57.005 132.775 57.665 ;
        RECT 132.945 57.175 133.465 58.660 ;
        RECT 133.635 57.835 134.155 59.385 ;
        RECT 134.325 58.830 134.655 59.555 ;
        RECT 135.205 58.830 135.535 59.555 ;
        RECT 133.815 57.005 134.155 57.665 ;
        RECT 134.325 57.175 134.845 58.660 ;
        RECT 135.015 57.175 135.535 58.660 ;
        RECT 135.705 57.835 136.225 59.385 ;
        RECT 136.395 58.465 138.065 59.555 ;
        RECT 136.395 57.775 137.145 58.295 ;
        RECT 137.315 57.945 138.065 58.465 ;
        RECT 138.695 58.390 138.985 59.555 ;
        RECT 139.245 58.885 139.415 59.385 ;
        RECT 139.585 59.055 139.915 59.555 ;
        RECT 139.245 58.715 139.850 58.885 ;
        RECT 139.155 57.905 139.400 58.545 ;
        RECT 139.680 58.320 139.850 58.715 ;
        RECT 140.085 58.605 140.310 59.385 ;
        RECT 139.680 57.990 139.910 58.320 ;
        RECT 135.705 57.005 136.045 57.665 ;
        RECT 136.395 57.005 138.065 57.775 ;
        RECT 138.695 57.005 138.985 57.730 ;
        RECT 139.680 57.725 139.850 57.990 ;
        RECT 139.245 57.555 139.850 57.725 ;
        RECT 139.245 57.265 139.415 57.555 ;
        RECT 139.585 57.005 139.915 57.385 ;
        RECT 140.085 57.265 140.255 58.605 ;
        RECT 140.545 58.585 140.875 59.335 ;
        RECT 141.045 58.755 141.360 59.555 ;
        RECT 141.990 59.175 142.740 59.345 ;
        RECT 140.545 58.415 141.230 58.585 ;
        RECT 140.550 57.875 140.880 58.245 ;
        RECT 141.060 58.015 141.230 58.415 ;
        RECT 141.560 58.275 141.845 58.925 ;
        RECT 142.015 58.335 142.355 58.915 ;
        RECT 141.060 57.705 141.430 58.015 ;
        RECT 142.015 57.955 142.185 58.335 ;
        RECT 142.570 58.245 142.740 59.175 ;
        RECT 142.910 59.055 143.210 59.555 ;
        RECT 143.430 58.785 143.650 59.355 ;
        RECT 142.930 58.455 143.650 58.785 ;
        RECT 143.480 58.245 143.650 58.455 ;
        RECT 143.830 58.415 144.115 59.555 ;
        RECT 144.285 58.560 144.535 59.375 ;
        RECT 144.705 58.675 144.965 59.555 ;
        RECT 144.285 58.415 144.570 58.560 ;
        RECT 144.400 58.245 144.570 58.415 ;
        RECT 142.570 58.085 143.290 58.245 ;
        RECT 140.625 57.685 141.430 57.705 ;
        RECT 140.625 57.535 141.230 57.685 ;
        RECT 141.805 57.625 142.185 57.955 ;
        RECT 142.420 57.915 143.290 58.085 ;
        RECT 143.480 57.915 144.230 58.245 ;
        RECT 144.400 57.915 144.965 58.245 ;
        RECT 140.625 57.265 140.795 57.535 ;
        RECT 142.420 57.455 142.590 57.915 ;
        RECT 143.480 57.745 143.650 57.915 ;
        RECT 144.400 57.745 144.570 57.915 ;
        RECT 145.135 57.835 145.655 59.385 ;
        RECT 145.825 58.830 146.155 59.555 ;
        RECT 140.965 57.005 141.295 57.365 ;
        RECT 141.930 57.285 142.590 57.455 ;
        RECT 142.830 57.005 143.160 57.745 ;
        RECT 143.430 57.335 143.650 57.745 ;
        RECT 143.830 57.005 144.115 57.745 ;
        RECT 144.285 57.605 144.570 57.745 ;
        RECT 144.285 57.335 144.535 57.605 ;
        RECT 144.705 57.005 144.965 57.470 ;
        RECT 145.315 57.005 145.655 57.665 ;
        RECT 145.825 57.175 146.345 58.660 ;
        RECT 146.515 57.835 147.035 59.385 ;
        RECT 147.205 58.830 147.535 59.555 ;
        RECT 146.695 57.005 147.035 57.665 ;
        RECT 147.205 57.175 147.725 58.660 ;
        RECT 147.895 58.465 151.405 59.555 ;
        RECT 147.895 57.775 149.545 58.295 ;
        RECT 149.715 57.945 151.405 58.465 ;
        RECT 151.575 58.390 151.865 59.555 ;
        RECT 152.035 58.465 155.545 59.555 ;
        RECT 152.035 57.775 153.685 58.295 ;
        RECT 153.855 57.945 155.545 58.465 ;
        RECT 155.715 58.465 156.925 59.555 ;
        RECT 155.715 57.925 156.235 58.465 ;
        RECT 147.895 57.005 151.405 57.775 ;
        RECT 151.575 57.005 151.865 57.730 ;
        RECT 152.035 57.005 155.545 57.775 ;
        RECT 156.405 57.755 156.925 58.295 ;
        RECT 155.715 57.005 156.925 57.755 ;
        RECT 22.690 56.835 157.010 57.005 ;
        RECT 114.100 49.650 116.700 49.820 ;
        RECT 114.100 48.800 114.270 49.650 ;
        RECT 114.900 49.140 115.900 49.310 ;
        RECT 74.220 48.250 76.820 48.420 ;
        RECT 33.000 47.410 35.600 47.580 ;
        RECT 33.000 46.560 33.170 47.410 ;
        RECT 33.800 46.900 34.800 47.070 ;
        RECT 32.980 44.760 33.180 46.560 ;
        RECT 33.000 34.010 33.170 44.760 ;
        RECT 33.570 34.690 33.740 46.730 ;
        RECT 34.860 34.690 35.030 46.730 ;
        RECT 33.800 34.350 34.800 34.520 ;
        RECT 35.430 34.010 35.600 47.410 ;
        RECT 74.220 47.400 74.390 48.250 ;
        RECT 75.020 47.740 76.020 47.910 ;
        RECT 74.200 45.600 74.400 47.400 ;
        RECT 33.000 33.840 35.600 34.010 ;
        RECT 40.000 38.410 42.600 38.580 ;
        RECT 40.000 34.010 40.170 38.410 ;
        RECT 40.800 37.900 41.800 38.070 ;
        RECT 42.430 38.060 42.600 38.410 ;
        RECT 40.570 34.690 40.740 37.730 ;
        RECT 41.860 34.690 42.030 37.730 ;
        RECT 42.430 36.510 42.630 38.060 ;
        RECT 43.700 37.960 46.300 38.130 ;
        RECT 43.700 37.660 43.870 37.960 ;
        RECT 43.680 36.510 43.880 37.660 ;
        RECT 44.500 37.450 45.500 37.620 ;
        RECT 40.800 34.350 41.800 34.520 ;
        RECT 42.430 34.010 42.600 36.510 ;
        RECT 43.700 34.440 43.870 36.510 ;
        RECT 44.270 35.120 44.440 37.280 ;
        RECT 45.560 35.120 45.730 37.280 ;
        RECT 44.500 34.780 45.500 34.950 ;
        RECT 46.130 34.440 46.300 37.960 ;
        RECT 43.700 34.270 46.300 34.440 ;
        RECT 46.710 34.760 49.950 34.930 ;
        RECT 40.000 33.840 42.600 34.010 ;
        RECT 46.710 33.910 46.880 34.760 ;
        RECT 49.780 34.410 49.950 34.760 ;
        RECT 50.410 34.760 53.150 34.930 ;
        RECT 50.410 34.410 50.580 34.760 ;
        RECT 47.560 34.190 49.100 34.360 ;
        RECT 35.000 32.910 37.600 33.080 ;
        RECT 35.000 31.960 35.170 32.910 ;
        RECT 35.800 32.400 36.800 32.570 ;
        RECT 34.980 30.160 35.180 31.960 ;
        RECT 35.000 23.030 35.170 30.160 ;
        RECT 35.570 23.710 35.740 32.230 ;
        RECT 36.860 23.710 37.030 32.230 ;
        RECT 35.800 23.370 36.800 23.540 ;
        RECT 37.430 23.030 37.600 32.910 ;
        RECT 46.680 32.860 46.880 33.910 ;
        RECT 47.220 33.130 47.390 34.130 ;
        RECT 49.270 33.130 49.440 34.130 ;
        RECT 47.560 32.900 49.100 33.070 ;
        RECT 46.710 32.500 46.880 32.860 ;
        RECT 49.780 32.860 49.980 34.410 ;
        RECT 50.380 32.860 50.580 34.410 ;
        RECT 51.260 34.190 52.300 34.360 ;
        RECT 50.920 33.130 51.090 34.130 ;
        RECT 52.470 33.130 52.640 34.130 ;
        RECT 51.260 32.900 52.300 33.070 ;
        RECT 49.780 32.500 49.950 32.860 ;
        RECT 46.710 32.330 49.950 32.500 ;
        RECT 50.410 32.500 50.580 32.860 ;
        RECT 52.980 32.500 53.150 34.760 ;
        RECT 74.220 34.850 74.390 45.600 ;
        RECT 74.790 35.530 74.960 47.570 ;
        RECT 76.080 35.530 76.250 47.570 ;
        RECT 75.020 35.190 76.020 35.360 ;
        RECT 76.650 34.850 76.820 48.250 ;
        RECT 114.080 47.000 114.280 48.800 ;
        RECT 74.220 34.680 76.820 34.850 ;
        RECT 81.220 39.250 83.820 39.420 ;
        RECT 81.220 34.850 81.390 39.250 ;
        RECT 82.020 38.740 83.020 38.910 ;
        RECT 83.650 38.900 83.820 39.250 ;
        RECT 81.790 35.530 81.960 38.570 ;
        RECT 83.080 35.530 83.250 38.570 ;
        RECT 83.650 37.350 83.850 38.900 ;
        RECT 84.920 38.800 87.520 38.970 ;
        RECT 84.920 38.500 85.090 38.800 ;
        RECT 84.900 37.350 85.100 38.500 ;
        RECT 85.720 38.290 86.720 38.460 ;
        RECT 82.020 35.190 83.020 35.360 ;
        RECT 83.650 34.850 83.820 37.350 ;
        RECT 84.920 35.280 85.090 37.350 ;
        RECT 85.490 35.960 85.660 38.120 ;
        RECT 86.780 35.960 86.950 38.120 ;
        RECT 85.720 35.620 86.720 35.790 ;
        RECT 87.350 35.280 87.520 38.800 ;
        RECT 114.100 36.250 114.270 47.000 ;
        RECT 114.670 36.930 114.840 48.970 ;
        RECT 115.960 36.930 116.130 48.970 ;
        RECT 114.900 36.590 115.900 36.760 ;
        RECT 116.530 36.250 116.700 49.650 ;
        RECT 114.100 36.080 116.700 36.250 ;
        RECT 121.100 40.650 123.700 40.820 ;
        RECT 121.100 36.250 121.270 40.650 ;
        RECT 121.900 40.140 122.900 40.310 ;
        RECT 123.530 40.300 123.700 40.650 ;
        RECT 121.670 36.930 121.840 39.970 ;
        RECT 122.960 36.930 123.130 39.970 ;
        RECT 123.530 38.750 123.730 40.300 ;
        RECT 124.800 40.200 127.400 40.370 ;
        RECT 124.800 39.900 124.970 40.200 ;
        RECT 124.780 38.750 124.980 39.900 ;
        RECT 125.600 39.690 126.600 39.860 ;
        RECT 121.900 36.590 122.900 36.760 ;
        RECT 123.530 36.250 123.700 38.750 ;
        RECT 124.800 36.680 124.970 38.750 ;
        RECT 125.370 37.360 125.540 39.520 ;
        RECT 126.660 37.360 126.830 39.520 ;
        RECT 125.600 37.020 126.600 37.190 ;
        RECT 127.230 36.680 127.400 40.200 ;
        RECT 124.800 36.510 127.400 36.680 ;
        RECT 127.810 37.000 131.050 37.170 ;
        RECT 121.100 36.080 123.700 36.250 ;
        RECT 127.810 36.150 127.980 37.000 ;
        RECT 130.880 36.650 131.050 37.000 ;
        RECT 131.510 37.000 134.250 37.170 ;
        RECT 131.510 36.650 131.680 37.000 ;
        RECT 128.660 36.430 130.200 36.600 ;
        RECT 84.920 35.110 87.520 35.280 ;
        RECT 87.930 35.600 91.170 35.770 ;
        RECT 81.220 34.680 83.820 34.850 ;
        RECT 87.930 34.750 88.100 35.600 ;
        RECT 91.000 35.250 91.170 35.600 ;
        RECT 91.630 35.600 94.370 35.770 ;
        RECT 91.630 35.250 91.800 35.600 ;
        RECT 88.780 35.030 90.320 35.200 ;
        RECT 76.220 33.750 78.820 33.920 ;
        RECT 76.220 32.800 76.390 33.750 ;
        RECT 77.020 33.240 78.020 33.410 ;
        RECT 50.410 32.330 53.150 32.500 ;
        RECT 50.410 31.810 53.150 31.980 ;
        RECT 50.410 30.460 50.580 31.810 ;
        RECT 51.260 31.240 52.300 31.410 ;
        RECT 50.330 29.360 50.580 30.460 ;
        RECT 50.920 29.680 51.090 31.180 ;
        RECT 52.470 29.680 52.640 31.180 ;
        RECT 51.260 29.450 52.300 29.620 ;
        RECT 50.410 29.050 50.580 29.360 ;
        RECT 52.980 29.050 53.150 31.810 ;
        RECT 76.200 31.000 76.400 32.800 ;
        RECT 50.410 28.880 53.150 29.050 ;
        RECT 50.430 28.230 50.830 28.310 ;
        RECT 49.980 28.060 53.700 28.230 ;
        RECT 49.980 27.860 50.150 28.060 ;
        RECT 49.980 27.410 50.230 27.860 ;
        RECT 50.780 27.550 52.900 27.720 ;
        RECT 49.980 25.660 50.150 27.410 ;
        RECT 50.550 26.340 50.720 27.380 ;
        RECT 52.960 26.340 53.130 27.380 ;
        RECT 50.780 26.000 52.900 26.170 ;
        RECT 53.530 25.660 53.700 28.060 ;
        RECT 49.980 25.490 53.700 25.660 ;
        RECT 35.000 22.860 37.600 23.030 ;
        RECT 50.150 24.510 54.750 24.680 ;
        RECT 50.150 22.110 50.320 24.510 ;
        RECT 50.950 24.000 53.950 24.170 ;
        RECT 50.720 22.790 50.890 23.830 ;
        RECT 54.010 22.790 54.180 23.830 ;
        RECT 50.950 22.450 53.950 22.620 ;
        RECT 54.580 22.110 54.750 24.510 ;
        RECT 76.220 23.870 76.390 31.000 ;
        RECT 76.790 24.550 76.960 33.070 ;
        RECT 78.080 24.550 78.250 33.070 ;
        RECT 77.020 24.210 78.020 24.380 ;
        RECT 78.650 23.870 78.820 33.750 ;
        RECT 87.900 33.700 88.100 34.750 ;
        RECT 88.440 33.970 88.610 34.970 ;
        RECT 90.490 33.970 90.660 34.970 ;
        RECT 88.780 33.740 90.320 33.910 ;
        RECT 87.930 33.340 88.100 33.700 ;
        RECT 91.000 33.700 91.200 35.250 ;
        RECT 91.600 33.700 91.800 35.250 ;
        RECT 92.480 35.030 93.520 35.200 ;
        RECT 92.140 33.970 92.310 34.970 ;
        RECT 93.690 33.970 93.860 34.970 ;
        RECT 92.480 33.740 93.520 33.910 ;
        RECT 91.000 33.340 91.170 33.700 ;
        RECT 87.930 33.170 91.170 33.340 ;
        RECT 91.630 33.340 91.800 33.700 ;
        RECT 94.200 33.340 94.370 35.600 ;
        RECT 116.100 35.150 118.700 35.320 ;
        RECT 116.100 34.200 116.270 35.150 ;
        RECT 116.900 34.640 117.900 34.810 ;
        RECT 91.630 33.170 94.370 33.340 ;
        RECT 91.630 32.650 94.370 32.820 ;
        RECT 91.630 31.300 91.800 32.650 ;
        RECT 92.480 32.080 93.520 32.250 ;
        RECT 91.550 30.200 91.800 31.300 ;
        RECT 92.140 30.520 92.310 32.020 ;
        RECT 93.690 30.520 93.860 32.020 ;
        RECT 92.480 30.290 93.520 30.460 ;
        RECT 91.630 29.890 91.800 30.200 ;
        RECT 94.200 29.890 94.370 32.650 ;
        RECT 116.080 32.400 116.280 34.200 ;
        RECT 91.630 29.720 94.370 29.890 ;
        RECT 91.650 29.070 92.050 29.150 ;
        RECT 91.200 28.900 94.920 29.070 ;
        RECT 91.200 28.700 91.370 28.900 ;
        RECT 91.200 28.250 91.450 28.700 ;
        RECT 92.000 28.390 94.120 28.560 ;
        RECT 91.200 26.500 91.370 28.250 ;
        RECT 91.770 27.180 91.940 28.220 ;
        RECT 94.180 27.180 94.350 28.220 ;
        RECT 92.000 26.840 94.120 27.010 ;
        RECT 94.750 26.500 94.920 28.900 ;
        RECT 91.200 26.330 94.920 26.500 ;
        RECT 76.220 23.700 78.820 23.870 ;
        RECT 91.370 25.350 95.970 25.520 ;
        RECT 91.370 22.950 91.540 25.350 ;
        RECT 92.170 24.840 95.170 25.010 ;
        RECT 91.940 23.630 92.110 24.670 ;
        RECT 95.230 23.630 95.400 24.670 ;
        RECT 92.170 23.290 95.170 23.460 ;
        RECT 95.800 22.950 95.970 25.350 ;
        RECT 116.100 25.270 116.270 32.400 ;
        RECT 116.670 25.950 116.840 34.470 ;
        RECT 117.960 25.950 118.130 34.470 ;
        RECT 116.900 25.610 117.900 25.780 ;
        RECT 118.530 25.270 118.700 35.150 ;
        RECT 127.780 35.100 127.980 36.150 ;
        RECT 128.320 35.370 128.490 36.370 ;
        RECT 130.370 35.370 130.540 36.370 ;
        RECT 128.660 35.140 130.200 35.310 ;
        RECT 127.810 34.740 127.980 35.100 ;
        RECT 130.880 35.100 131.080 36.650 ;
        RECT 131.480 35.100 131.680 36.650 ;
        RECT 132.360 36.430 133.400 36.600 ;
        RECT 132.020 35.370 132.190 36.370 ;
        RECT 133.570 35.370 133.740 36.370 ;
        RECT 132.360 35.140 133.400 35.310 ;
        RECT 130.880 34.740 131.050 35.100 ;
        RECT 127.810 34.570 131.050 34.740 ;
        RECT 131.510 34.740 131.680 35.100 ;
        RECT 134.080 34.740 134.250 37.000 ;
        RECT 131.510 34.570 134.250 34.740 ;
        RECT 131.510 34.050 134.250 34.220 ;
        RECT 131.510 32.700 131.680 34.050 ;
        RECT 132.360 33.480 133.400 33.650 ;
        RECT 131.430 31.600 131.680 32.700 ;
        RECT 132.020 31.920 132.190 33.420 ;
        RECT 133.570 31.920 133.740 33.420 ;
        RECT 132.360 31.690 133.400 31.860 ;
        RECT 131.510 31.290 131.680 31.600 ;
        RECT 134.080 31.290 134.250 34.050 ;
        RECT 131.510 31.120 134.250 31.290 ;
        RECT 131.530 30.470 131.930 30.550 ;
        RECT 131.080 30.300 134.800 30.470 ;
        RECT 131.080 30.100 131.250 30.300 ;
        RECT 131.080 29.650 131.330 30.100 ;
        RECT 131.880 29.790 134.000 29.960 ;
        RECT 131.080 27.900 131.250 29.650 ;
        RECT 131.650 28.580 131.820 29.620 ;
        RECT 134.060 28.580 134.230 29.620 ;
        RECT 131.880 28.240 134.000 28.410 ;
        RECT 134.630 27.900 134.800 30.300 ;
        RECT 131.080 27.730 134.800 27.900 ;
        RECT 116.100 25.100 118.700 25.270 ;
        RECT 131.250 26.750 135.850 26.920 ;
        RECT 131.250 24.350 131.420 26.750 ;
        RECT 132.050 26.240 135.050 26.410 ;
        RECT 131.820 25.030 131.990 26.070 ;
        RECT 135.110 25.030 135.280 26.070 ;
        RECT 132.050 24.690 135.050 24.860 ;
        RECT 135.680 24.350 135.850 26.750 ;
        RECT 117.600 24.150 120.200 24.320 ;
        RECT 131.250 24.180 135.850 24.350 ;
        RECT 131.560 24.150 134.320 24.180 ;
        RECT 117.600 23.200 117.770 24.150 ;
        RECT 118.400 23.640 119.400 23.810 ;
        RECT 36.500 21.910 39.100 22.080 ;
        RECT 50.150 21.940 54.750 22.110 ;
        RECT 77.720 22.750 80.320 22.920 ;
        RECT 91.370 22.780 95.970 22.950 ;
        RECT 91.680 22.750 94.440 22.780 ;
        RECT 50.460 21.910 53.220 21.940 ;
        RECT 36.500 20.960 36.670 21.910 ;
        RECT 37.300 21.400 38.300 21.570 ;
        RECT 36.480 19.060 36.680 20.960 ;
        RECT 36.500 14.510 36.670 19.060 ;
        RECT 37.070 15.190 37.240 21.230 ;
        RECT 38.360 15.190 38.530 21.230 ;
        RECT 37.300 14.850 38.300 15.020 ;
        RECT 38.930 14.510 39.100 21.910 ;
        RECT 77.720 21.800 77.890 22.750 ;
        RECT 78.520 22.240 79.520 22.410 ;
        RECT 50.120 20.930 55.960 21.100 ;
        RECT 50.120 18.530 50.290 20.930 ;
        RECT 50.920 20.420 55.160 20.590 ;
        RECT 50.690 19.210 50.860 20.250 ;
        RECT 55.220 19.210 55.390 20.250 ;
        RECT 50.920 18.870 55.160 19.040 ;
        RECT 55.790 18.530 55.960 20.930 ;
        RECT 77.700 19.900 77.900 21.800 ;
        RECT 50.120 18.360 55.960 18.530 ;
        RECT 50.460 18.330 53.220 18.360 ;
        RECT 49.990 17.350 57.590 17.520 ;
        RECT 49.990 14.950 50.160 17.350 ;
        RECT 50.790 16.840 56.790 17.010 ;
        RECT 50.560 15.630 50.730 16.670 ;
        RECT 56.850 15.630 57.020 16.670 ;
        RECT 50.790 15.290 56.790 15.460 ;
        RECT 57.420 14.950 57.590 17.350 ;
        RECT 77.720 15.350 77.890 19.900 ;
        RECT 78.290 16.030 78.460 22.070 ;
        RECT 79.580 16.030 79.750 22.070 ;
        RECT 78.520 15.690 79.520 15.860 ;
        RECT 80.150 15.350 80.320 22.750 ;
        RECT 91.340 21.770 97.180 21.940 ;
        RECT 91.340 19.370 91.510 21.770 ;
        RECT 92.140 21.260 96.380 21.430 ;
        RECT 91.910 20.050 92.080 21.090 ;
        RECT 96.440 20.050 96.610 21.090 ;
        RECT 92.140 19.710 96.380 19.880 ;
        RECT 97.010 19.370 97.180 21.770 ;
        RECT 117.580 21.300 117.780 23.200 ;
        RECT 91.340 19.200 97.180 19.370 ;
        RECT 91.680 19.170 94.440 19.200 ;
        RECT 91.210 18.190 98.810 18.360 ;
        RECT 91.210 15.790 91.380 18.190 ;
        RECT 92.010 17.680 98.010 17.850 ;
        RECT 91.780 16.470 91.950 17.510 ;
        RECT 98.070 16.470 98.240 17.510 ;
        RECT 92.010 16.130 98.010 16.300 ;
        RECT 98.640 15.790 98.810 18.190 ;
        RECT 117.600 16.750 117.770 21.300 ;
        RECT 118.170 17.430 118.340 23.470 ;
        RECT 119.460 17.430 119.630 23.470 ;
        RECT 118.400 17.090 119.400 17.260 ;
        RECT 120.030 16.750 120.200 24.150 ;
        RECT 131.220 23.170 137.060 23.340 ;
        RECT 131.220 20.770 131.390 23.170 ;
        RECT 132.020 22.660 136.260 22.830 ;
        RECT 131.790 21.450 131.960 22.490 ;
        RECT 136.320 21.450 136.490 22.490 ;
        RECT 132.020 21.110 136.260 21.280 ;
        RECT 136.890 20.770 137.060 23.170 ;
        RECT 131.220 20.600 137.060 20.770 ;
        RECT 131.560 20.570 134.320 20.600 ;
        RECT 131.090 19.590 138.690 19.760 ;
        RECT 131.090 17.190 131.260 19.590 ;
        RECT 131.890 19.080 137.890 19.250 ;
        RECT 131.660 17.870 131.830 18.910 ;
        RECT 137.950 17.870 138.120 18.910 ;
        RECT 131.890 17.530 137.890 17.700 ;
        RECT 138.520 17.190 138.690 19.590 ;
        RECT 131.090 17.020 138.690 17.190 ;
        RECT 131.560 16.990 134.320 17.020 ;
        RECT 117.600 16.580 120.200 16.750 ;
        RECT 131.110 16.010 141.190 16.180 ;
        RECT 91.210 15.620 98.810 15.790 ;
        RECT 119.600 15.650 122.200 15.820 ;
        RECT 91.680 15.590 94.440 15.620 ;
        RECT 77.720 15.180 80.320 15.350 ;
        RECT 119.600 15.000 119.770 15.650 ;
        RECT 120.400 15.140 121.400 15.310 ;
        RECT 49.990 14.780 57.590 14.950 ;
        RECT 50.460 14.750 53.220 14.780 ;
        RECT 36.500 14.340 39.100 14.510 ;
        RECT 91.230 14.610 101.310 14.780 ;
        RECT 79.720 14.250 82.320 14.420 ;
        RECT 50.010 13.770 60.090 13.940 ;
        RECT 38.500 13.410 41.100 13.580 ;
        RECT 38.500 12.760 38.670 13.410 ;
        RECT 39.300 12.900 40.300 13.070 ;
        RECT 38.480 10.960 38.680 12.760 ;
        RECT 38.500 7.770 38.670 10.960 ;
        RECT 39.070 8.450 39.240 12.730 ;
        RECT 40.360 8.450 40.530 12.730 ;
        RECT 39.300 8.110 40.300 8.280 ;
        RECT 40.930 7.770 41.100 13.410 ;
        RECT 50.010 11.370 50.180 13.770 ;
        RECT 50.810 13.260 59.290 13.430 ;
        RECT 50.580 12.050 50.750 13.090 ;
        RECT 59.350 12.050 59.520 13.090 ;
        RECT 50.810 11.710 59.290 11.880 ;
        RECT 59.920 11.370 60.090 13.770 ;
        RECT 79.720 13.600 79.890 14.250 ;
        RECT 80.520 13.740 81.520 13.910 ;
        RECT 79.700 11.800 79.900 13.600 ;
        RECT 50.010 11.200 60.090 11.370 ;
        RECT 50.460 11.170 53.220 11.200 ;
        RECT 38.500 7.600 41.100 7.770 ;
        RECT 50.020 10.190 63.620 10.360 ;
        RECT 50.020 7.790 50.190 10.190 ;
        RECT 50.820 9.680 62.820 9.850 ;
        RECT 50.590 8.470 50.760 9.510 ;
        RECT 62.880 8.470 63.050 9.510 ;
        RECT 50.820 8.130 62.820 8.300 ;
        RECT 60.380 7.790 63.130 7.810 ;
        RECT 63.450 7.790 63.620 10.190 ;
        RECT 79.720 8.610 79.890 11.800 ;
        RECT 80.290 9.290 80.460 13.570 ;
        RECT 81.580 9.290 81.750 13.570 ;
        RECT 80.520 8.950 81.520 9.120 ;
        RECT 82.150 8.610 82.320 14.250 ;
        RECT 91.230 12.210 91.400 14.610 ;
        RECT 92.030 14.100 100.510 14.270 ;
        RECT 91.800 12.890 91.970 13.930 ;
        RECT 100.570 12.890 100.740 13.930 ;
        RECT 92.030 12.550 100.510 12.720 ;
        RECT 101.140 12.210 101.310 14.610 ;
        RECT 119.580 13.200 119.780 15.000 ;
        RECT 91.230 12.040 101.310 12.210 ;
        RECT 91.680 12.010 94.440 12.040 ;
        RECT 79.720 8.440 82.320 8.610 ;
        RECT 91.240 11.030 104.840 11.200 ;
        RECT 91.240 8.630 91.410 11.030 ;
        RECT 92.040 10.520 104.040 10.690 ;
        RECT 91.810 9.310 91.980 10.350 ;
        RECT 104.100 9.310 104.270 10.350 ;
        RECT 92.040 8.970 104.040 9.140 ;
        RECT 101.600 8.630 104.350 8.650 ;
        RECT 104.670 8.630 104.840 11.030 ;
        RECT 119.600 10.010 119.770 13.200 ;
        RECT 120.170 10.690 120.340 14.970 ;
        RECT 121.460 10.690 121.630 14.970 ;
        RECT 120.400 10.350 121.400 10.520 ;
        RECT 122.030 10.010 122.200 15.650 ;
        RECT 131.110 13.610 131.280 16.010 ;
        RECT 131.910 15.500 140.390 15.670 ;
        RECT 131.680 14.290 131.850 15.330 ;
        RECT 140.450 14.290 140.620 15.330 ;
        RECT 131.910 13.950 140.390 14.120 ;
        RECT 141.020 13.610 141.190 16.010 ;
        RECT 131.110 13.440 141.190 13.610 ;
        RECT 131.560 13.410 134.320 13.440 ;
        RECT 119.600 9.840 122.200 10.010 ;
        RECT 131.120 12.430 144.720 12.600 ;
        RECT 131.120 10.030 131.290 12.430 ;
        RECT 131.920 11.920 143.920 12.090 ;
        RECT 131.690 10.710 131.860 11.750 ;
        RECT 143.980 10.710 144.150 11.750 ;
        RECT 131.920 10.370 143.920 10.540 ;
        RECT 141.480 10.030 144.230 10.050 ;
        RECT 144.550 10.030 144.720 12.430 ;
        RECT 131.120 9.860 144.720 10.030 ;
        RECT 141.480 9.850 144.230 9.860 ;
        RECT 91.240 8.460 104.840 8.630 ;
        RECT 101.600 8.450 104.350 8.460 ;
        RECT 50.020 7.620 63.620 7.790 ;
        RECT 60.380 7.610 63.130 7.620 ;
      LAYER met1 ;
        RECT 87.160 210.160 87.480 210.220 ;
        RECT 125.340 210.160 125.660 210.220 ;
        RECT 87.160 210.020 125.660 210.160 ;
        RECT 87.160 209.960 87.480 210.020 ;
        RECT 125.340 209.960 125.660 210.020 ;
        RECT 117.060 209.820 117.380 209.880 ;
        RECT 133.620 209.820 133.940 209.880 ;
        RECT 117.060 209.680 133.940 209.820 ;
        RECT 117.060 209.620 117.380 209.680 ;
        RECT 133.620 209.620 133.940 209.680 ;
        RECT 22.690 209.000 157.810 209.480 ;
        RECT 24.615 208.800 24.905 208.845 ;
        RECT 26.900 208.800 27.220 208.860 ;
        RECT 24.615 208.660 27.220 208.800 ;
        RECT 24.615 208.615 24.905 208.660 ;
        RECT 26.900 208.600 27.220 208.660 ;
        RECT 48.980 208.600 49.300 208.860 ;
        RECT 57.260 208.600 57.580 208.860 ;
        RECT 63.700 208.600 64.020 208.860 ;
        RECT 75.290 208.660 85.550 208.800 ;
        RECT 30.120 208.165 30.440 208.180 ;
        RECT 30.120 207.935 30.525 208.165 ;
        RECT 37.480 208.120 37.800 208.180 ;
        RECT 39.335 208.120 39.625 208.165 ;
        RECT 37.480 207.980 39.625 208.120 ;
        RECT 49.070 208.120 49.210 208.600 ;
        RECT 50.375 208.120 50.665 208.165 ;
        RECT 49.070 207.980 50.665 208.120 ;
        RECT 57.350 208.120 57.490 208.600 ;
        RECT 57.735 208.120 58.025 208.165 ;
        RECT 57.350 207.980 58.025 208.120 ;
        RECT 30.120 207.920 30.440 207.935 ;
        RECT 37.480 207.920 37.800 207.980 ;
        RECT 39.335 207.935 39.625 207.980 ;
        RECT 50.375 207.935 50.665 207.980 ;
        RECT 57.735 207.935 58.025 207.980 ;
        RECT 62.795 207.935 63.085 208.165 ;
        RECT 63.790 208.120 63.930 208.600 ;
        RECT 68.775 208.460 69.065 208.505 ;
        RECT 75.290 208.460 75.430 208.660 ;
        RECT 68.775 208.320 75.430 208.460 ;
        RECT 75.750 208.320 82.790 208.460 ;
        RECT 68.775 208.275 69.065 208.320 ;
        RECT 64.175 208.120 64.465 208.165 ;
        RECT 63.790 207.980 64.465 208.120 ;
        RECT 64.175 207.935 64.465 207.980 ;
        RECT 67.395 207.935 67.685 208.165 ;
        RECT 26.925 207.780 27.215 207.825 ;
        RECT 29.445 207.780 29.735 207.825 ;
        RECT 30.635 207.780 30.925 207.825 ;
        RECT 26.925 207.640 30.925 207.780 ;
        RECT 26.925 207.595 27.215 207.640 ;
        RECT 29.445 207.595 29.735 207.640 ;
        RECT 30.635 207.595 30.925 207.640 ;
        RECT 31.500 207.580 31.820 207.840 ;
        RECT 62.870 207.780 63.010 207.935 ;
        RECT 67.470 207.780 67.610 207.935 ;
        RECT 68.300 207.920 68.620 208.180 ;
        RECT 69.220 207.920 69.540 208.180 ;
        RECT 71.520 208.120 71.840 208.180 ;
        RECT 74.755 208.120 75.045 208.165 ;
        RECT 71.520 207.980 75.045 208.120 ;
        RECT 71.520 207.920 71.840 207.980 ;
        RECT 74.755 207.935 75.045 207.980 ;
        RECT 70.615 207.780 70.905 207.825 ;
        RECT 62.870 207.640 63.930 207.780 ;
        RECT 67.470 207.640 70.905 207.780 ;
        RECT 27.360 207.440 27.650 207.485 ;
        RECT 28.930 207.440 29.220 207.485 ;
        RECT 31.030 207.440 31.320 207.485 ;
        RECT 27.360 207.300 31.320 207.440 ;
        RECT 27.360 207.255 27.650 207.300 ;
        RECT 28.930 207.255 29.220 207.300 ;
        RECT 31.030 207.255 31.320 207.300 ;
        RECT 63.790 207.160 63.930 207.640 ;
        RECT 70.615 207.595 70.905 207.640 ;
        RECT 71.060 207.780 71.380 207.840 ;
        RECT 73.375 207.780 73.665 207.825 ;
        RECT 71.060 207.640 73.665 207.780 ;
        RECT 71.060 207.580 71.380 207.640 ;
        RECT 73.375 207.595 73.665 207.640 ;
        RECT 70.155 207.440 70.445 207.485 ;
        RECT 75.200 207.440 75.520 207.500 ;
        RECT 75.750 207.485 75.890 208.320 ;
        RECT 78.420 208.120 78.740 208.180 ;
        RECT 82.650 208.165 82.790 208.320 ;
        RECT 79.815 208.120 80.105 208.165 ;
        RECT 78.420 207.980 80.105 208.120 ;
        RECT 78.420 207.920 78.740 207.980 ;
        RECT 79.815 207.935 80.105 207.980 ;
        RECT 81.655 207.935 81.945 208.165 ;
        RECT 82.575 208.120 82.865 208.165 ;
        RECT 83.480 208.120 83.800 208.180 ;
        RECT 82.575 207.980 83.800 208.120 ;
        RECT 82.575 207.935 82.865 207.980 ;
        RECT 76.120 207.580 76.440 207.840 ;
        RECT 78.880 207.580 79.200 207.840 ;
        RECT 81.730 207.780 81.870 207.935 ;
        RECT 83.480 207.920 83.800 207.980 ;
        RECT 82.100 207.780 82.420 207.840 ;
        RECT 81.730 207.640 82.420 207.780 ;
        RECT 85.410 207.780 85.550 208.660 ;
        RECT 100.500 208.600 100.820 208.860 ;
        RECT 125.340 208.800 125.660 208.860 ;
        RECT 118.070 208.660 121.890 208.800 ;
        RECT 85.780 208.120 86.100 208.180 ;
        RECT 91.315 208.120 91.605 208.165 ;
        RECT 85.780 207.980 91.605 208.120 ;
        RECT 85.780 207.920 86.100 207.980 ;
        RECT 91.315 207.935 91.605 207.980 ;
        RECT 93.140 208.120 93.460 208.180 ;
        RECT 93.615 208.120 93.905 208.165 ;
        RECT 93.140 207.980 93.905 208.120 ;
        RECT 93.140 207.920 93.460 207.980 ;
        RECT 93.615 207.935 93.905 207.980 ;
        RECT 96.360 207.920 96.680 208.180 ;
        RECT 100.590 208.120 100.730 208.600 ;
        RECT 118.070 208.520 118.210 208.660 ;
        RECT 107.860 208.460 108.180 208.520 ;
        RECT 109.255 208.460 109.545 208.505 ;
        RECT 107.860 208.320 109.545 208.460 ;
        RECT 107.860 208.260 108.180 208.320 ;
        RECT 109.255 208.275 109.545 208.320 ;
        RECT 109.790 208.320 117.750 208.460 ;
        RECT 100.975 208.120 101.265 208.165 ;
        RECT 100.590 207.980 101.265 208.120 ;
        RECT 100.975 207.935 101.265 207.980 ;
        RECT 103.720 208.120 104.040 208.180 ;
        RECT 104.655 208.120 104.945 208.165 ;
        RECT 103.720 207.980 104.945 208.120 ;
        RECT 103.720 207.920 104.040 207.980 ;
        RECT 104.655 207.935 104.945 207.980 ;
        RECT 85.410 207.640 88.310 207.780 ;
        RECT 81.960 207.580 82.420 207.640 ;
        RECT 70.155 207.300 75.520 207.440 ;
        RECT 70.155 207.255 70.445 207.300 ;
        RECT 75.200 207.240 75.520 207.300 ;
        RECT 75.675 207.255 75.965 207.485 ;
        RECT 81.960 207.440 82.100 207.580 ;
        RECT 88.170 207.500 88.310 207.640 ;
        RECT 90.380 207.580 90.700 207.840 ;
        RECT 109.790 207.780 109.930 208.320 ;
        RECT 110.160 207.920 110.480 208.180 ;
        RECT 117.060 207.920 117.380 208.180 ;
        RECT 117.610 208.165 117.750 208.320 ;
        RECT 117.980 208.260 118.300 208.520 ;
        RECT 118.440 208.260 118.760 208.520 ;
        RECT 121.215 208.460 121.505 208.505 ;
        RECT 118.990 208.320 121.505 208.460 ;
        RECT 121.750 208.460 121.890 208.660 ;
        RECT 125.340 208.660 137.070 208.800 ;
        RECT 125.340 208.600 125.660 208.660 ;
        RECT 136.930 208.505 137.070 208.660 ;
        RECT 137.300 208.600 137.620 208.860 ;
        RECT 152.020 208.600 152.340 208.860 ;
        RECT 121.750 208.320 133.390 208.460 ;
        RECT 117.535 208.120 117.825 208.165 ;
        RECT 118.530 208.120 118.670 208.260 ;
        RECT 118.990 208.165 119.130 208.320 ;
        RECT 121.215 208.275 121.505 208.320 ;
        RECT 117.535 207.980 118.670 208.120 ;
        RECT 117.535 207.935 117.825 207.980 ;
        RECT 118.915 207.935 119.205 208.165 ;
        RECT 119.835 207.935 120.125 208.165 ;
        RECT 127.655 208.120 127.945 208.165 ;
        RECT 129.940 208.120 130.260 208.180 ;
        RECT 127.655 207.980 130.260 208.120 ;
        RECT 127.655 207.935 127.945 207.980 ;
        RECT 92.310 207.640 109.930 207.780 ;
        RECT 115.220 207.780 115.540 207.840 ;
        RECT 119.910 207.780 120.050 207.935 ;
        RECT 129.940 207.920 130.260 207.980 ;
        RECT 115.220 207.640 120.050 207.780 ;
        RECT 76.210 207.300 82.100 207.440 ;
        RECT 88.080 207.440 88.400 207.500 ;
        RECT 92.310 207.485 92.450 207.640 ;
        RECT 115.220 207.580 115.540 207.640 ;
        RECT 123.960 207.580 124.280 207.840 ;
        RECT 128.560 207.580 128.880 207.840 ;
        RECT 132.240 207.580 132.560 207.840 ;
        RECT 133.250 207.780 133.390 208.320 ;
        RECT 136.855 208.275 137.145 208.505 ;
        RECT 137.390 208.460 137.530 208.600 ;
        RECT 137.390 208.320 139.370 208.460 ;
        RECT 133.620 208.120 133.940 208.180 ;
        RECT 139.230 208.165 139.370 208.320 ;
        RECT 136.395 208.120 136.685 208.165 ;
        RECT 133.620 207.980 136.685 208.120 ;
        RECT 133.620 207.920 133.940 207.980 ;
        RECT 136.395 207.935 136.685 207.980 ;
        RECT 137.315 207.935 137.605 208.165 ;
        RECT 138.235 207.935 138.525 208.165 ;
        RECT 139.155 207.935 139.445 208.165 ;
        RECT 152.110 208.120 152.250 208.600 ;
        RECT 153.415 208.120 153.705 208.165 ;
        RECT 152.110 207.980 153.705 208.120 ;
        RECT 153.415 207.935 153.705 207.980 ;
        RECT 135.920 207.780 136.240 207.840 ;
        RECT 137.390 207.780 137.530 207.935 ;
        RECT 133.250 207.640 137.530 207.780 ;
        RECT 135.920 207.580 136.240 207.640 ;
        RECT 92.235 207.440 92.525 207.485 ;
        RECT 88.080 207.300 92.525 207.440 ;
        RECT 37.940 207.100 38.260 207.160 ;
        RECT 38.415 207.100 38.705 207.145 ;
        RECT 37.940 206.960 38.705 207.100 ;
        RECT 37.940 206.900 38.260 206.960 ;
        RECT 38.415 206.915 38.705 206.960 ;
        RECT 49.440 206.900 49.760 207.160 ;
        RECT 56.800 206.900 57.120 207.160 ;
        RECT 62.320 206.900 62.640 207.160 ;
        RECT 63.700 206.900 64.020 207.160 ;
        RECT 65.095 207.100 65.385 207.145 ;
        RECT 76.210 207.100 76.350 207.300 ;
        RECT 88.080 207.240 88.400 207.300 ;
        RECT 92.235 207.255 92.525 207.300 ;
        RECT 92.680 207.440 93.000 207.500 ;
        RECT 105.575 207.440 105.865 207.485 ;
        RECT 110.620 207.440 110.940 207.500 ;
        RECT 92.680 207.300 95.670 207.440 ;
        RECT 92.680 207.240 93.000 207.300 ;
        RECT 65.095 206.960 76.350 207.100 ;
        RECT 65.095 206.915 65.385 206.960 ;
        RECT 80.720 206.900 81.040 207.160 ;
        RECT 82.115 207.100 82.405 207.145 ;
        RECT 83.020 207.100 83.340 207.160 ;
        RECT 82.115 206.960 83.340 207.100 ;
        RECT 82.115 206.915 82.405 206.960 ;
        RECT 83.020 206.900 83.340 206.960 ;
        RECT 87.620 206.900 87.940 207.160 ;
        RECT 93.140 207.100 93.460 207.160 ;
        RECT 95.530 207.145 95.670 207.300 ;
        RECT 105.575 207.300 110.940 207.440 ;
        RECT 105.575 207.255 105.865 207.300 ;
        RECT 110.620 207.240 110.940 207.300 ;
        RECT 131.335 207.440 131.625 207.485 ;
        RECT 138.310 207.440 138.450 207.935 ;
        RECT 131.335 207.300 138.450 207.440 ;
        RECT 131.335 207.255 131.625 207.300 ;
        RECT 94.535 207.100 94.825 207.145 ;
        RECT 93.140 206.960 94.825 207.100 ;
        RECT 93.140 206.900 93.460 206.960 ;
        RECT 94.535 206.915 94.825 206.960 ;
        RECT 95.455 206.915 95.745 207.145 ;
        RECT 101.880 206.900 102.200 207.160 ;
        RECT 108.780 206.900 109.100 207.160 ;
        RECT 111.080 206.900 111.400 207.160 ;
        RECT 116.155 207.100 116.445 207.145 ;
        RECT 117.520 207.100 117.840 207.160 ;
        RECT 116.155 206.960 117.840 207.100 ;
        RECT 116.155 206.915 116.445 206.960 ;
        RECT 117.520 206.900 117.840 206.960 ;
        RECT 120.280 206.900 120.600 207.160 ;
        RECT 126.720 206.900 127.040 207.160 ;
        RECT 135.000 206.900 135.320 207.160 ;
        RECT 135.460 206.900 135.780 207.160 ;
        RECT 137.760 207.100 138.080 207.160 ;
        RECT 140.075 207.100 140.365 207.145 ;
        RECT 137.760 206.960 140.365 207.100 ;
        RECT 137.760 206.900 138.080 206.960 ;
        RECT 140.075 206.915 140.365 206.960 ;
        RECT 152.480 206.900 152.800 207.160 ;
        RECT 22.690 206.280 157.010 206.760 ;
        RECT 48.535 206.080 48.825 206.125 ;
        RECT 49.440 206.080 49.760 206.140 ;
        RECT 85.795 206.080 86.085 206.125 ;
        RECT 86.240 206.080 86.560 206.140 ;
        RECT 90.380 206.080 90.700 206.140 ;
        RECT 48.535 205.940 49.760 206.080 ;
        RECT 48.535 205.895 48.825 205.940 ;
        RECT 28.320 205.740 28.610 205.785 ;
        RECT 30.420 205.740 30.710 205.785 ;
        RECT 31.990 205.740 32.280 205.785 ;
        RECT 28.320 205.600 32.280 205.740 ;
        RECT 28.320 205.555 28.610 205.600 ;
        RECT 30.420 205.555 30.710 205.600 ;
        RECT 31.990 205.555 32.280 205.600 ;
        RECT 34.260 205.740 34.580 205.800 ;
        RECT 34.735 205.740 35.025 205.785 ;
        RECT 34.260 205.600 35.025 205.740 ;
        RECT 34.260 205.540 34.580 205.600 ;
        RECT 34.735 205.555 35.025 205.600 ;
        RECT 37.060 205.740 37.350 205.785 ;
        RECT 39.160 205.740 39.450 205.785 ;
        RECT 40.730 205.740 41.020 205.785 ;
        RECT 37.060 205.600 41.020 205.740 ;
        RECT 37.060 205.555 37.350 205.600 ;
        RECT 39.160 205.555 39.450 205.600 ;
        RECT 40.730 205.555 41.020 205.600 ;
        RECT 45.775 205.740 46.065 205.785 ;
        RECT 48.610 205.740 48.750 205.895 ;
        RECT 49.440 205.880 49.760 205.940 ;
        RECT 49.990 205.940 57.030 206.080 ;
        RECT 45.775 205.600 48.750 205.740 ;
        RECT 45.775 205.555 46.065 205.600 ;
        RECT 28.715 205.400 29.005 205.445 ;
        RECT 29.905 205.400 30.195 205.445 ;
        RECT 32.425 205.400 32.715 205.445 ;
        RECT 28.715 205.260 32.715 205.400 ;
        RECT 28.715 205.215 29.005 205.260 ;
        RECT 29.905 205.215 30.195 205.260 ;
        RECT 32.425 205.215 32.715 205.260 ;
        RECT 37.455 205.400 37.745 205.445 ;
        RECT 38.645 205.400 38.935 205.445 ;
        RECT 41.165 205.400 41.455 205.445 ;
        RECT 37.455 205.260 41.455 205.400 ;
        RECT 37.455 205.215 37.745 205.260 ;
        RECT 38.645 205.215 38.935 205.260 ;
        RECT 41.165 205.215 41.455 205.260 ;
        RECT 43.935 205.400 44.225 205.445 ;
        RECT 49.990 205.400 50.130 205.940 ;
        RECT 56.890 205.800 57.030 205.940 ;
        RECT 85.795 205.940 86.560 206.080 ;
        RECT 85.795 205.895 86.085 205.940 ;
        RECT 86.240 205.880 86.560 205.940 ;
        RECT 89.090 205.940 90.700 206.080 ;
        RECT 50.375 205.555 50.665 205.785 ;
        RECT 51.320 205.740 51.610 205.785 ;
        RECT 53.420 205.740 53.710 205.785 ;
        RECT 54.990 205.740 55.280 205.785 ;
        RECT 51.320 205.600 55.280 205.740 ;
        RECT 51.320 205.555 51.610 205.600 ;
        RECT 53.420 205.555 53.710 205.600 ;
        RECT 54.990 205.555 55.280 205.600 ;
        RECT 43.935 205.260 50.130 205.400 ;
        RECT 43.935 205.215 44.225 205.260 ;
        RECT 27.835 205.060 28.125 205.105 ;
        RECT 31.500 205.060 31.820 205.120 ;
        RECT 36.575 205.060 36.865 205.105 ;
        RECT 42.540 205.060 42.860 205.120 ;
        RECT 49.070 205.105 49.210 205.260 ;
        RECT 27.835 204.920 42.860 205.060 ;
        RECT 27.835 204.875 28.125 204.920 ;
        RECT 28.830 204.440 28.970 204.920 ;
        RECT 31.500 204.860 31.820 204.920 ;
        RECT 36.575 204.875 36.865 204.920 ;
        RECT 42.540 204.860 42.860 204.920 ;
        RECT 48.995 204.875 49.285 205.105 ;
        RECT 49.440 204.860 49.760 205.120 ;
        RECT 50.450 205.060 50.590 205.555 ;
        RECT 56.800 205.540 57.120 205.800 ;
        RECT 58.655 205.740 58.945 205.785 ;
        RECT 57.810 205.600 58.945 205.740 ;
        RECT 51.715 205.400 52.005 205.445 ;
        RECT 52.905 205.400 53.195 205.445 ;
        RECT 55.425 205.400 55.715 205.445 ;
        RECT 51.715 205.260 55.715 205.400 ;
        RECT 51.715 205.215 52.005 205.260 ;
        RECT 52.905 205.215 53.195 205.260 ;
        RECT 55.425 205.215 55.715 205.260 ;
        RECT 49.990 204.920 50.590 205.060 ;
        RECT 50.835 205.060 51.125 205.105 ;
        RECT 54.040 205.060 54.360 205.120 ;
        RECT 50.835 204.920 54.360 205.060 ;
        RECT 29.200 204.765 29.520 204.780 ;
        RECT 37.940 204.765 38.260 204.780 ;
        RECT 29.170 204.535 29.520 204.765 ;
        RECT 37.910 204.720 38.260 204.765 ;
        RECT 47.140 204.720 47.460 204.780 ;
        RECT 37.745 204.580 38.260 204.720 ;
        RECT 37.910 204.535 38.260 204.580 ;
        RECT 29.200 204.520 29.520 204.535 ;
        RECT 37.940 204.520 38.260 204.535 ;
        RECT 43.550 204.580 47.460 204.720 ;
        RECT 49.990 204.720 50.130 204.920 ;
        RECT 50.835 204.875 51.125 204.920 ;
        RECT 54.040 204.860 54.360 204.920 ;
        RECT 52.060 204.720 52.350 204.765 ;
        RECT 57.260 204.720 57.580 204.780 ;
        RECT 49.990 204.580 52.350 204.720 ;
        RECT 28.740 204.180 29.060 204.440 ;
        RECT 43.550 204.425 43.690 204.580 ;
        RECT 47.140 204.520 47.460 204.580 ;
        RECT 52.060 204.535 52.350 204.580 ;
        RECT 53.210 204.580 57.580 204.720 ;
        RECT 43.475 204.195 43.765 204.425 ;
        RECT 45.760 204.380 46.080 204.440 ;
        RECT 46.235 204.380 46.525 204.425 ;
        RECT 45.760 204.240 46.525 204.380 ;
        RECT 45.760 204.180 46.080 204.240 ;
        RECT 46.235 204.195 46.525 204.240 ;
        RECT 46.695 204.380 46.985 204.425 ;
        RECT 47.600 204.380 47.920 204.440 ;
        RECT 46.695 204.240 47.920 204.380 ;
        RECT 46.695 204.195 46.985 204.240 ;
        RECT 47.600 204.180 47.920 204.240 ;
        RECT 48.980 204.380 49.300 204.440 ;
        RECT 53.210 204.380 53.350 204.580 ;
        RECT 57.260 204.520 57.580 204.580 ;
        RECT 57.810 204.720 57.950 205.600 ;
        RECT 58.655 205.555 58.945 205.600 ;
        RECT 65.540 205.740 65.830 205.785 ;
        RECT 67.110 205.740 67.400 205.785 ;
        RECT 69.210 205.740 69.500 205.785 ;
        RECT 65.540 205.600 69.500 205.740 ;
        RECT 65.540 205.555 65.830 205.600 ;
        RECT 67.110 205.555 67.400 205.600 ;
        RECT 69.210 205.555 69.500 205.600 ;
        RECT 73.360 205.740 73.650 205.785 ;
        RECT 74.930 205.740 75.220 205.785 ;
        RECT 77.030 205.740 77.320 205.785 ;
        RECT 73.360 205.600 77.320 205.740 ;
        RECT 73.360 205.555 73.650 205.600 ;
        RECT 74.930 205.555 75.220 205.600 ;
        RECT 77.030 205.555 77.320 205.600 ;
        RECT 78.460 205.740 78.750 205.785 ;
        RECT 80.560 205.740 80.850 205.785 ;
        RECT 82.130 205.740 82.420 205.785 ;
        RECT 78.460 205.600 82.420 205.740 ;
        RECT 78.460 205.555 78.750 205.600 ;
        RECT 80.560 205.555 80.850 205.600 ;
        RECT 82.130 205.555 82.420 205.600 ;
        RECT 84.860 205.740 85.180 205.800 ;
        RECT 89.090 205.740 89.230 205.940 ;
        RECT 90.380 205.880 90.700 205.940 ;
        RECT 95.915 206.080 96.205 206.125 ;
        RECT 98.200 206.080 98.520 206.140 ;
        RECT 95.915 205.940 98.520 206.080 ;
        RECT 95.915 205.895 96.205 205.940 ;
        RECT 98.200 205.880 98.520 205.940 ;
        RECT 100.975 206.080 101.265 206.125 ;
        RECT 101.880 206.080 102.200 206.140 ;
        RECT 100.975 205.940 102.200 206.080 ;
        RECT 100.975 205.895 101.265 205.940 ;
        RECT 101.880 205.880 102.200 205.940 ;
        RECT 123.515 206.080 123.805 206.125 ;
        RECT 123.960 206.080 124.280 206.140 ;
        RECT 123.515 205.940 124.280 206.080 ;
        RECT 123.515 205.895 123.805 205.940 ;
        RECT 123.960 205.880 124.280 205.940 ;
        RECT 132.240 206.080 132.560 206.140 ;
        RECT 133.160 206.080 133.480 206.140 ;
        RECT 132.240 205.940 133.480 206.080 ;
        RECT 132.240 205.880 132.560 205.940 ;
        RECT 133.160 205.880 133.480 205.940 ;
        RECT 152.480 205.880 152.800 206.140 ;
        RECT 84.860 205.600 89.230 205.740 ;
        RECT 89.500 205.740 89.790 205.785 ;
        RECT 91.600 205.740 91.890 205.785 ;
        RECT 93.170 205.740 93.460 205.785 ;
        RECT 89.500 205.600 93.460 205.740 ;
        RECT 84.860 205.540 85.180 205.600 ;
        RECT 89.500 205.555 89.790 205.600 ;
        RECT 91.600 205.555 91.890 205.600 ;
        RECT 93.170 205.555 93.460 205.600 ;
        RECT 105.100 205.540 105.420 205.800 ;
        RECT 107.860 205.740 108.150 205.785 ;
        RECT 109.430 205.740 109.720 205.785 ;
        RECT 111.530 205.740 111.820 205.785 ;
        RECT 107.860 205.600 111.820 205.740 ;
        RECT 107.860 205.555 108.150 205.600 ;
        RECT 109.430 205.555 109.720 205.600 ;
        RECT 111.530 205.555 111.820 205.600 ;
        RECT 117.100 205.740 117.390 205.785 ;
        RECT 119.200 205.740 119.490 205.785 ;
        RECT 120.770 205.740 121.060 205.785 ;
        RECT 117.100 205.600 121.060 205.740 ;
        RECT 117.100 205.555 117.390 205.600 ;
        RECT 119.200 205.555 119.490 205.600 ;
        RECT 120.770 205.555 121.060 205.600 ;
        RECT 126.760 205.740 127.050 205.785 ;
        RECT 128.860 205.740 129.150 205.785 ;
        RECT 130.430 205.740 130.720 205.785 ;
        RECT 152.570 205.740 152.710 205.880 ;
        RECT 126.760 205.600 130.720 205.740 ;
        RECT 126.760 205.555 127.050 205.600 ;
        RECT 128.860 205.555 129.150 205.600 ;
        RECT 130.430 205.555 130.720 205.600 ;
        RECT 132.790 205.600 152.710 205.740 ;
        RECT 65.105 205.400 65.395 205.445 ;
        RECT 67.625 205.400 67.915 205.445 ;
        RECT 68.815 205.400 69.105 205.445 ;
        RECT 65.105 205.260 69.105 205.400 ;
        RECT 65.105 205.215 65.395 205.260 ;
        RECT 67.625 205.215 67.915 205.260 ;
        RECT 68.815 205.215 69.105 205.260 ;
        RECT 72.925 205.400 73.215 205.445 ;
        RECT 75.445 205.400 75.735 205.445 ;
        RECT 76.635 205.400 76.925 205.445 ;
        RECT 72.925 205.260 76.925 205.400 ;
        RECT 72.925 205.215 73.215 205.260 ;
        RECT 75.445 205.215 75.735 205.260 ;
        RECT 76.635 205.215 76.925 205.260 ;
        RECT 78.855 205.400 79.145 205.445 ;
        RECT 80.045 205.400 80.335 205.445 ;
        RECT 82.565 205.400 82.855 205.445 ;
        RECT 78.855 205.260 82.855 205.400 ;
        RECT 78.855 205.215 79.145 205.260 ;
        RECT 80.045 205.215 80.335 205.260 ;
        RECT 82.565 205.215 82.855 205.260 ;
        RECT 83.020 205.200 83.340 205.460 ;
        RECT 83.940 205.400 84.260 205.460 ;
        RECT 89.015 205.400 89.305 205.445 ;
        RECT 83.940 205.260 89.305 205.400 ;
        RECT 83.940 205.200 84.260 205.260 ;
        RECT 89.015 205.215 89.305 205.260 ;
        RECT 89.895 205.400 90.185 205.445 ;
        RECT 91.085 205.400 91.375 205.445 ;
        RECT 93.605 205.400 93.895 205.445 ;
        RECT 100.055 205.400 100.345 205.445 ;
        RECT 104.640 205.400 104.960 205.460 ;
        RECT 106.480 205.400 106.800 205.460 ;
        RECT 89.895 205.260 93.895 205.400 ;
        RECT 89.895 205.215 90.185 205.260 ;
        RECT 91.085 205.215 91.375 205.260 ;
        RECT 93.605 205.215 93.895 205.260 ;
        RECT 94.150 205.260 106.800 205.400 ;
        RECT 69.695 205.060 69.985 205.105 ;
        RECT 74.740 205.060 75.060 205.120 ;
        RECT 77.515 205.060 77.805 205.105 ;
        RECT 77.975 205.060 78.265 205.105 ;
        RECT 69.695 204.920 78.265 205.060 ;
        RECT 83.110 205.060 83.250 205.200 ;
        RECT 85.320 205.060 85.640 205.120 ;
        RECT 83.110 204.920 85.640 205.060 ;
        RECT 69.695 204.875 69.985 204.920 ;
        RECT 74.740 204.860 75.060 204.920 ;
        RECT 77.515 204.875 77.805 204.920 ;
        RECT 77.975 204.875 78.265 204.920 ;
        RECT 85.320 204.860 85.640 204.920 ;
        RECT 86.255 205.060 86.545 205.105 ;
        RECT 87.620 205.060 87.940 205.120 ;
        RECT 86.255 204.920 87.940 205.060 ;
        RECT 86.255 204.875 86.545 204.920 ;
        RECT 87.620 204.860 87.940 204.920 ;
        RECT 90.350 205.060 90.640 205.105 ;
        RECT 92.680 205.060 93.000 205.120 ;
        RECT 90.350 204.920 93.000 205.060 ;
        RECT 90.350 204.875 90.640 204.920 ;
        RECT 92.680 204.860 93.000 204.920 ;
        RECT 93.140 205.060 93.460 205.120 ;
        RECT 94.150 205.060 94.290 205.260 ;
        RECT 100.055 205.215 100.345 205.260 ;
        RECT 104.640 205.200 104.960 205.260 ;
        RECT 106.480 205.200 106.800 205.260 ;
        RECT 107.425 205.400 107.715 205.445 ;
        RECT 109.945 205.400 110.235 205.445 ;
        RECT 111.135 205.400 111.425 205.445 ;
        RECT 107.425 205.260 111.425 205.400 ;
        RECT 107.425 205.215 107.715 205.260 ;
        RECT 109.945 205.215 110.235 205.260 ;
        RECT 111.135 205.215 111.425 205.260 ;
        RECT 117.495 205.400 117.785 205.445 ;
        RECT 118.685 205.400 118.975 205.445 ;
        RECT 121.205 205.400 121.495 205.445 ;
        RECT 117.495 205.260 121.495 205.400 ;
        RECT 117.495 205.215 117.785 205.260 ;
        RECT 118.685 205.215 118.975 205.260 ;
        RECT 121.205 205.215 121.495 205.260 ;
        RECT 126.260 205.200 126.580 205.460 ;
        RECT 127.155 205.400 127.445 205.445 ;
        RECT 128.345 205.400 128.635 205.445 ;
        RECT 130.865 205.400 131.155 205.445 ;
        RECT 127.155 205.260 131.155 205.400 ;
        RECT 127.155 205.215 127.445 205.260 ;
        RECT 128.345 205.215 128.635 205.260 ;
        RECT 130.865 205.215 131.155 205.260 ;
        RECT 93.140 204.920 94.290 205.060 ;
        RECT 93.140 204.860 93.460 204.920 ;
        RECT 97.295 204.875 97.585 205.105 ;
        RECT 101.435 204.875 101.725 205.105 ;
        RECT 60.020 204.720 60.340 204.780 ;
        RECT 57.810 204.580 60.340 204.720 ;
        RECT 48.980 204.240 53.350 204.380 ;
        RECT 53.580 204.380 53.900 204.440 ;
        RECT 57.810 204.425 57.950 204.580 ;
        RECT 60.020 204.520 60.340 204.580 ;
        RECT 60.495 204.720 60.785 204.765 ;
        RECT 63.240 204.720 63.560 204.780 ;
        RECT 68.360 204.720 68.650 204.765 ;
        RECT 60.495 204.580 63.010 204.720 ;
        RECT 60.495 204.535 60.785 204.580 ;
        RECT 57.735 204.380 58.025 204.425 ;
        RECT 53.580 204.240 58.025 204.380 ;
        RECT 48.980 204.180 49.300 204.240 ;
        RECT 53.580 204.180 53.900 204.240 ;
        RECT 57.735 204.195 58.025 204.240 ;
        RECT 58.180 204.180 58.500 204.440 ;
        RECT 62.870 204.425 63.010 204.580 ;
        RECT 63.240 204.580 68.650 204.720 ;
        RECT 63.240 204.520 63.560 204.580 ;
        RECT 68.360 204.535 68.650 204.580 ;
        RECT 75.200 204.720 75.520 204.780 ;
        RECT 76.180 204.720 76.470 204.765 ;
        RECT 75.200 204.580 76.470 204.720 ;
        RECT 75.200 204.520 75.520 204.580 ;
        RECT 76.180 204.535 76.470 204.580 ;
        RECT 79.310 204.720 79.600 204.765 ;
        RECT 88.540 204.720 88.860 204.780 ;
        RECT 79.310 204.580 88.860 204.720 ;
        RECT 79.310 204.535 79.600 204.580 ;
        RECT 88.540 204.520 88.860 204.580 ;
        RECT 91.300 204.720 91.620 204.780 ;
        RECT 95.440 204.720 95.760 204.780 ;
        RECT 96.835 204.720 97.125 204.765 ;
        RECT 91.300 204.580 94.750 204.720 ;
        RECT 91.300 204.520 91.620 204.580 ;
        RECT 62.795 204.380 63.085 204.425 ;
        RECT 63.700 204.380 64.020 204.440 ;
        RECT 62.795 204.240 64.020 204.380 ;
        RECT 62.795 204.195 63.085 204.240 ;
        RECT 63.700 204.180 64.020 204.240 ;
        RECT 67.840 204.380 68.160 204.440 ;
        RECT 70.615 204.380 70.905 204.425 ;
        RECT 71.060 204.380 71.380 204.440 ;
        RECT 67.840 204.240 71.380 204.380 ;
        RECT 67.840 204.180 68.160 204.240 ;
        RECT 70.615 204.195 70.905 204.240 ;
        RECT 71.060 204.180 71.380 204.240 ;
        RECT 75.660 204.380 75.980 204.440 ;
        RECT 93.140 204.380 93.460 204.440 ;
        RECT 75.660 204.240 93.460 204.380 ;
        RECT 94.610 204.380 94.750 204.580 ;
        RECT 95.440 204.580 97.125 204.720 ;
        RECT 97.370 204.720 97.510 204.875 ;
        RECT 97.740 204.720 98.060 204.780 ;
        RECT 97.370 204.580 100.730 204.720 ;
        RECT 95.440 204.520 95.760 204.580 ;
        RECT 96.835 204.535 97.125 204.580 ;
        RECT 97.740 204.520 98.060 204.580 ;
        RECT 100.590 204.440 100.730 204.580 ;
        RECT 98.675 204.380 98.965 204.425 ;
        RECT 94.610 204.240 98.965 204.380 ;
        RECT 75.660 204.180 75.980 204.240 ;
        RECT 93.140 204.180 93.460 204.240 ;
        RECT 98.675 204.195 98.965 204.240 ;
        RECT 100.500 204.180 100.820 204.440 ;
        RECT 101.510 204.380 101.650 204.875 ;
        RECT 101.880 204.860 102.200 205.120 ;
        RECT 110.620 205.105 110.940 205.120 ;
        RECT 110.620 205.060 110.970 205.105 ;
        RECT 112.015 205.060 112.305 205.105 ;
        RECT 116.615 205.060 116.905 205.105 ;
        RECT 117.060 205.060 117.380 205.120 ;
        RECT 110.620 204.920 111.135 205.060 ;
        RECT 112.015 204.920 117.380 205.060 ;
        RECT 110.620 204.875 110.970 204.920 ;
        RECT 112.015 204.875 112.305 204.920 ;
        RECT 116.615 204.875 116.905 204.920 ;
        RECT 110.620 204.860 110.940 204.875 ;
        RECT 117.060 204.860 117.380 204.920 ;
        RECT 117.950 204.875 118.240 205.105 ;
        RECT 122.120 205.060 122.440 205.120 ;
        RECT 123.975 205.060 124.265 205.105 ;
        RECT 132.790 205.060 132.930 205.600 ;
        RECT 133.620 205.400 133.940 205.460 ;
        RECT 135.000 205.400 135.320 205.460 ;
        RECT 142.835 205.400 143.125 205.445 ;
        RECT 133.620 205.260 134.770 205.400 ;
        RECT 133.620 205.200 133.940 205.260 ;
        RECT 122.120 204.920 124.265 205.060 ;
        RECT 102.800 204.720 103.120 204.780 ;
        RECT 103.275 204.720 103.565 204.765 ;
        RECT 117.520 204.720 117.840 204.780 ;
        RECT 118.070 204.720 118.210 204.875 ;
        RECT 122.120 204.860 122.440 204.920 ;
        RECT 123.975 204.875 124.265 204.920 ;
        RECT 124.510 204.920 132.930 205.060 ;
        RECT 133.160 205.060 133.480 205.120 ;
        RECT 134.630 205.105 134.770 205.260 ;
        RECT 135.000 205.260 136.610 205.400 ;
        RECT 135.000 205.200 135.320 205.260 ;
        RECT 136.470 205.105 136.610 205.260 ;
        RECT 140.150 205.260 143.125 205.400 ;
        RECT 140.150 205.105 140.290 205.260 ;
        RECT 142.835 205.215 143.125 205.260 ;
        RECT 133.160 204.920 134.310 205.060 ;
        RECT 124.510 204.720 124.650 204.920 ;
        RECT 133.160 204.860 133.480 204.920 ;
        RECT 102.800 204.580 103.565 204.720 ;
        RECT 102.800 204.520 103.120 204.580 ;
        RECT 103.275 204.535 103.565 204.580 ;
        RECT 105.190 204.580 117.290 204.720 ;
        RECT 105.190 204.380 105.330 204.580 ;
        RECT 101.510 204.240 105.330 204.380 ;
        RECT 117.150 204.380 117.290 204.580 ;
        RECT 117.520 204.580 118.210 204.720 ;
        RECT 123.130 204.580 124.650 204.720 ;
        RECT 127.610 204.720 127.900 204.765 ;
        RECT 127.610 204.580 133.850 204.720 ;
        RECT 117.520 204.520 117.840 204.580 ;
        RECT 123.130 204.380 123.270 204.580 ;
        RECT 127.610 204.535 127.900 204.580 ;
        RECT 117.150 204.240 123.270 204.380 ;
        RECT 124.880 204.180 125.200 204.440 ;
        RECT 133.710 204.425 133.850 204.580 ;
        RECT 133.635 204.195 133.925 204.425 ;
        RECT 134.170 204.380 134.310 204.920 ;
        RECT 134.555 204.875 134.845 205.105 ;
        RECT 136.395 204.875 136.685 205.105 ;
        RECT 136.855 204.875 137.145 205.105 ;
        RECT 140.075 204.875 140.365 205.105 ;
        RECT 142.375 205.060 142.665 205.105 ;
        RECT 140.610 204.920 142.665 205.060 ;
        RECT 135.000 204.520 135.320 204.780 ;
        RECT 135.475 204.720 135.765 204.765 ;
        RECT 135.920 204.720 136.240 204.780 ;
        RECT 135.475 204.580 136.240 204.720 ;
        RECT 135.475 204.535 135.765 204.580 ;
        RECT 135.920 204.520 136.240 204.580 ;
        RECT 136.930 204.380 137.070 204.875 ;
        RECT 137.300 204.720 137.620 204.780 ;
        RECT 140.610 204.720 140.750 204.920 ;
        RECT 142.375 204.875 142.665 204.920 ;
        RECT 143.295 204.875 143.585 205.105 ;
        RECT 144.675 205.060 144.965 205.105 ;
        RECT 144.675 204.920 146.270 205.060 ;
        RECT 144.675 204.875 144.965 204.920 ;
        RECT 137.300 204.580 140.750 204.720 ;
        RECT 137.300 204.520 137.620 204.580 ;
        RECT 141.900 204.520 142.220 204.780 ;
        RECT 143.370 204.720 143.510 204.875 ;
        RECT 142.450 204.580 143.510 204.720 ;
        RECT 142.450 204.440 142.590 204.580 ;
        RECT 146.130 204.440 146.270 204.920 ;
        RECT 134.170 204.240 137.070 204.380 ;
        RECT 138.220 204.380 138.540 204.440 ;
        RECT 139.155 204.380 139.445 204.425 ;
        RECT 138.220 204.240 139.445 204.380 ;
        RECT 138.220 204.180 138.540 204.240 ;
        RECT 139.155 204.195 139.445 204.240 ;
        RECT 139.600 204.380 139.920 204.440 ;
        RECT 140.535 204.380 140.825 204.425 ;
        RECT 139.600 204.240 140.825 204.380 ;
        RECT 139.600 204.180 139.920 204.240 ;
        RECT 140.535 204.195 140.825 204.240 ;
        RECT 140.980 204.180 141.300 204.440 ;
        RECT 142.360 204.180 142.680 204.440 ;
        RECT 144.200 204.180 144.520 204.440 ;
        RECT 146.040 204.180 146.360 204.440 ;
        RECT 22.690 203.560 157.810 204.040 ;
        RECT 37.480 203.360 37.800 203.420 ;
        RECT 40.255 203.360 40.545 203.405 ;
        RECT 48.980 203.360 49.300 203.420 ;
        RECT 37.480 203.220 40.545 203.360 ;
        RECT 37.480 203.160 37.800 203.220 ;
        RECT 40.255 203.175 40.545 203.220 ;
        RECT 43.550 203.220 49.300 203.360 ;
        RECT 39.335 203.020 39.625 203.065 ;
        RECT 40.700 203.020 41.020 203.080 ;
        RECT 42.555 203.020 42.845 203.065 ;
        RECT 39.335 202.880 41.020 203.020 ;
        RECT 39.335 202.835 39.625 202.880 ;
        RECT 40.700 202.820 41.020 202.880 ;
        RECT 41.250 202.880 42.845 203.020 ;
        RECT 29.675 202.680 29.965 202.725 ;
        RECT 29.290 202.540 29.965 202.680 ;
        RECT 29.290 202.400 29.430 202.540 ;
        RECT 29.675 202.495 29.965 202.540 ;
        RECT 30.120 202.680 30.440 202.740 ;
        RECT 30.955 202.680 31.245 202.725 ;
        RECT 30.120 202.540 31.245 202.680 ;
        RECT 30.120 202.480 30.440 202.540 ;
        RECT 30.955 202.495 31.245 202.540 ;
        RECT 37.495 202.680 37.785 202.725 ;
        RECT 37.940 202.680 38.260 202.740 ;
        RECT 41.250 202.725 41.390 202.880 ;
        RECT 42.555 202.835 42.845 202.880 ;
        RECT 43.550 202.725 43.690 203.220 ;
        RECT 48.980 203.160 49.300 203.220 ;
        RECT 49.440 203.360 49.760 203.420 ;
        RECT 50.835 203.360 51.125 203.405 ;
        RECT 49.440 203.220 51.125 203.360 ;
        RECT 49.440 203.160 49.760 203.220 ;
        RECT 50.835 203.175 51.125 203.220 ;
        RECT 54.975 203.360 55.265 203.405 ;
        RECT 54.975 203.220 55.650 203.360 ;
        RECT 54.975 203.175 55.265 203.220 ;
        RECT 53.580 203.020 53.900 203.080 ;
        RECT 45.850 202.880 53.900 203.020 ;
        RECT 45.850 202.725 45.990 202.880 ;
        RECT 53.580 202.820 53.900 202.880 ;
        RECT 55.510 202.740 55.650 203.220 ;
        RECT 55.895 203.175 56.185 203.405 ;
        RECT 57.260 203.360 57.580 203.420 ;
        RECT 59.560 203.360 59.880 203.420 ;
        RECT 78.880 203.360 79.200 203.420 ;
        RECT 81.655 203.360 81.945 203.405 ;
        RECT 57.260 203.220 60.710 203.360 ;
        RECT 55.970 203.020 56.110 203.175 ;
        RECT 57.260 203.160 57.580 203.220 ;
        RECT 59.560 203.160 59.880 203.220 ;
        RECT 59.100 203.020 59.420 203.080 ;
        RECT 55.970 202.880 59.420 203.020 ;
        RECT 59.100 202.820 59.420 202.880 ;
        RECT 41.175 202.680 41.465 202.725 ;
        RECT 37.495 202.540 41.465 202.680 ;
        RECT 37.495 202.495 37.785 202.540 ;
        RECT 37.940 202.480 38.260 202.540 ;
        RECT 41.175 202.495 41.465 202.540 ;
        RECT 42.095 202.680 42.385 202.725 ;
        RECT 43.475 202.680 43.765 202.725 ;
        RECT 42.095 202.540 43.765 202.680 ;
        RECT 42.095 202.495 42.385 202.540 ;
        RECT 43.475 202.495 43.765 202.540 ;
        RECT 45.775 202.495 46.065 202.725 ;
        RECT 49.915 202.680 50.205 202.725 ;
        RECT 47.690 202.540 50.205 202.680 ;
        RECT 29.200 202.140 29.520 202.400 ;
        RECT 30.555 202.340 30.845 202.385 ;
        RECT 31.745 202.340 32.035 202.385 ;
        RECT 34.265 202.340 34.555 202.385 ;
        RECT 30.555 202.200 34.555 202.340 ;
        RECT 30.555 202.155 30.845 202.200 ;
        RECT 31.745 202.155 32.035 202.200 ;
        RECT 34.265 202.155 34.555 202.200 ;
        RECT 41.635 202.340 41.925 202.385 ;
        RECT 45.300 202.340 45.620 202.400 ;
        RECT 41.635 202.200 45.620 202.340 ;
        RECT 41.635 202.155 41.925 202.200 ;
        RECT 45.300 202.140 45.620 202.200 ;
        RECT 47.690 202.045 47.830 202.540 ;
        RECT 49.915 202.495 50.205 202.540 ;
        RECT 54.055 202.495 54.345 202.725 ;
        RECT 48.995 202.340 49.285 202.385 ;
        RECT 48.150 202.200 49.285 202.340 ;
        RECT 30.160 202.000 30.450 202.045 ;
        RECT 32.260 202.000 32.550 202.045 ;
        RECT 33.830 202.000 34.120 202.045 ;
        RECT 30.160 201.860 34.120 202.000 ;
        RECT 30.160 201.815 30.450 201.860 ;
        RECT 32.260 201.815 32.550 201.860 ;
        RECT 33.830 201.815 34.120 201.860 ;
        RECT 38.950 201.860 41.850 202.000 ;
        RECT 36.575 201.660 36.865 201.705 ;
        RECT 38.950 201.660 39.090 201.860 ;
        RECT 41.710 201.720 41.850 201.860 ;
        RECT 44.010 201.860 47.370 202.000 ;
        RECT 44.010 201.720 44.150 201.860 ;
        RECT 36.575 201.520 39.090 201.660 ;
        RECT 39.335 201.660 39.625 201.705 ;
        RECT 41.160 201.660 41.480 201.720 ;
        RECT 39.335 201.520 41.480 201.660 ;
        RECT 36.575 201.475 36.865 201.520 ;
        RECT 39.335 201.475 39.625 201.520 ;
        RECT 41.160 201.460 41.480 201.520 ;
        RECT 41.620 201.460 41.940 201.720 ;
        RECT 43.920 201.460 44.240 201.720 ;
        RECT 44.380 201.460 44.700 201.720 ;
        RECT 47.230 201.660 47.370 201.860 ;
        RECT 47.615 201.815 47.905 202.045 ;
        RECT 48.150 201.660 48.290 202.200 ;
        RECT 48.995 202.155 49.285 202.200 ;
        RECT 51.740 202.140 52.060 202.400 ;
        RECT 54.130 202.340 54.270 202.495 ;
        RECT 54.500 202.480 54.820 202.740 ;
        RECT 55.420 202.480 55.740 202.740 ;
        RECT 58.640 202.725 58.960 202.740 ;
        RECT 60.570 202.725 60.710 203.220 ;
        RECT 68.390 203.220 81.945 203.360 ;
        RECT 67.840 203.020 68.160 203.080 ;
        RECT 63.330 202.880 68.160 203.020 ;
        RECT 56.355 202.680 56.645 202.725 ;
        RECT 58.610 202.680 58.960 202.725 ;
        RECT 56.355 202.540 58.410 202.680 ;
        RECT 56.355 202.495 56.645 202.540 ;
        RECT 58.270 202.400 58.410 202.540 ;
        RECT 58.610 202.540 59.110 202.680 ;
        RECT 58.610 202.495 58.960 202.540 ;
        RECT 60.495 202.495 60.785 202.725 ;
        RECT 61.400 202.680 61.720 202.740 ;
        RECT 63.330 202.725 63.470 202.880 ;
        RECT 67.840 202.820 68.160 202.880 ;
        RECT 62.795 202.680 63.085 202.725 ;
        RECT 61.400 202.540 63.085 202.680 ;
        RECT 58.640 202.480 58.960 202.495 ;
        RECT 61.400 202.480 61.720 202.540 ;
        RECT 62.795 202.495 63.085 202.540 ;
        RECT 63.255 202.495 63.545 202.725 ;
        RECT 63.700 202.480 64.020 202.740 ;
        RECT 68.390 202.725 68.530 203.220 ;
        RECT 78.880 203.160 79.200 203.220 ;
        RECT 81.655 203.175 81.945 203.220 ;
        RECT 83.480 203.160 83.800 203.420 ;
        RECT 84.860 203.360 85.180 203.420 ;
        RECT 91.300 203.360 91.620 203.420 ;
        RECT 84.490 203.220 85.180 203.360 ;
        RECT 69.220 203.020 69.540 203.080 ;
        RECT 75.980 203.020 76.270 203.065 ;
        RECT 68.850 202.880 72.210 203.020 ;
        RECT 68.315 202.495 68.605 202.725 ;
        RECT 54.960 202.340 55.280 202.400 ;
        RECT 54.130 202.200 55.280 202.340 ;
        RECT 54.960 202.140 55.280 202.200 ;
        RECT 55.880 202.140 56.200 202.400 ;
        RECT 57.735 202.340 58.025 202.385 ;
        RECT 56.430 202.200 58.025 202.340 ;
        RECT 51.830 202.000 51.970 202.140 ;
        RECT 56.430 202.000 56.570 202.200 ;
        RECT 57.735 202.155 58.025 202.200 ;
        RECT 58.180 202.140 58.500 202.400 ;
        RECT 67.855 202.340 68.145 202.385 ;
        RECT 59.190 202.200 68.145 202.340 ;
        RECT 51.830 201.860 56.570 202.000 ;
        RECT 56.815 201.815 57.105 202.045 ;
        RECT 58.640 202.000 58.960 202.060 ;
        RECT 59.190 202.000 59.330 202.200 ;
        RECT 67.855 202.155 68.145 202.200 ;
        RECT 68.850 202.000 68.990 202.880 ;
        RECT 69.220 202.820 69.540 202.880 ;
        RECT 70.155 202.495 70.445 202.725 ;
        RECT 58.640 201.860 59.330 202.000 ;
        RECT 63.790 201.860 68.990 202.000 ;
        RECT 47.230 201.520 48.290 201.660 ;
        RECT 55.420 201.660 55.740 201.720 ;
        RECT 56.890 201.660 57.030 201.815 ;
        RECT 58.640 201.800 58.960 201.860 ;
        RECT 63.790 201.720 63.930 201.860 ;
        RECT 57.720 201.660 58.040 201.720 ;
        RECT 55.420 201.520 58.040 201.660 ;
        RECT 55.420 201.460 55.740 201.520 ;
        RECT 57.720 201.460 58.040 201.520 ;
        RECT 63.700 201.460 64.020 201.720 ;
        RECT 66.920 201.460 67.240 201.720 ;
        RECT 70.230 201.660 70.370 202.495 ;
        RECT 71.060 202.480 71.380 202.740 ;
        RECT 71.520 202.480 71.840 202.740 ;
        RECT 72.070 202.725 72.210 202.880 ;
        RECT 72.990 202.880 76.270 203.020 ;
        RECT 71.995 202.495 72.285 202.725 ;
        RECT 72.990 202.045 73.130 202.880 ;
        RECT 75.980 202.835 76.270 202.880 ;
        RECT 82.100 202.820 82.420 203.080 ;
        RECT 84.490 203.065 84.630 203.220 ;
        RECT 84.860 203.160 85.180 203.220 ;
        RECT 90.010 203.220 91.620 203.360 ;
        RECT 90.010 203.065 90.150 203.220 ;
        RECT 91.300 203.160 91.620 203.220 ;
        RECT 91.775 203.360 92.065 203.405 ;
        RECT 94.980 203.360 95.300 203.420 ;
        RECT 95.535 203.360 95.825 203.405 ;
        RECT 91.775 203.220 95.825 203.360 ;
        RECT 91.775 203.175 92.065 203.220 ;
        RECT 94.980 203.160 95.300 203.220 ;
        RECT 95.535 203.175 95.825 203.220 ;
        RECT 96.360 203.160 96.680 203.420 ;
        RECT 100.500 203.360 100.820 203.420 ;
        RECT 101.435 203.360 101.725 203.405 ;
        RECT 100.500 203.220 103.030 203.360 ;
        RECT 100.500 203.160 100.820 203.220 ;
        RECT 101.435 203.175 101.725 203.220 ;
        RECT 92.220 203.065 92.540 203.080 ;
        RECT 84.415 202.835 84.705 203.065 ;
        RECT 89.935 202.835 90.225 203.065 ;
        RECT 92.220 202.835 92.615 203.065 ;
        RECT 94.535 203.020 94.825 203.065 ;
        RECT 96.820 203.020 97.140 203.080 ;
        RECT 94.535 202.880 97.140 203.020 ;
        RECT 94.535 202.835 94.825 202.880 ;
        RECT 92.220 202.820 92.540 202.835 ;
        RECT 96.820 202.820 97.140 202.880 ;
        RECT 97.740 203.065 98.060 203.080 ;
        RECT 97.740 202.835 98.275 203.065 ;
        RECT 98.835 203.020 99.125 203.065 ;
        RECT 100.960 203.020 101.280 203.080 ;
        RECT 98.750 202.880 101.280 203.020 ;
        RECT 98.750 202.835 99.125 202.880 ;
        RECT 97.740 202.820 98.060 202.835 ;
        RECT 85.320 202.680 85.640 202.740 ;
        RECT 89.200 202.680 89.490 202.725 ;
        RECT 85.320 202.540 89.490 202.680 ;
        RECT 85.320 202.480 85.640 202.540 ;
        RECT 89.200 202.495 89.490 202.540 ;
        RECT 90.855 202.495 91.145 202.725 ;
        RECT 91.775 202.670 92.065 202.725 ;
        RECT 93.155 202.680 93.445 202.725 ;
        RECT 92.770 202.670 93.445 202.680 ;
        RECT 91.775 202.540 93.445 202.670 ;
        RECT 91.775 202.530 92.910 202.540 ;
        RECT 91.775 202.495 92.065 202.530 ;
        RECT 93.155 202.495 93.445 202.540 ;
        RECT 74.740 202.140 75.060 202.400 ;
        RECT 75.635 202.340 75.925 202.385 ;
        RECT 76.825 202.340 77.115 202.385 ;
        RECT 79.345 202.340 79.635 202.385 ;
        RECT 75.635 202.200 79.635 202.340 ;
        RECT 75.635 202.155 75.925 202.200 ;
        RECT 76.825 202.155 77.115 202.200 ;
        RECT 79.345 202.155 79.635 202.200 ;
        RECT 80.720 202.340 81.040 202.400 ;
        RECT 82.100 202.340 82.420 202.400 ;
        RECT 80.720 202.200 82.420 202.340 ;
        RECT 80.720 202.140 81.040 202.200 ;
        RECT 82.100 202.140 82.420 202.200 ;
        RECT 83.955 202.340 84.245 202.385 ;
        RECT 87.620 202.340 87.940 202.400 ;
        RECT 83.955 202.200 87.940 202.340 ;
        RECT 83.955 202.155 84.245 202.200 ;
        RECT 87.620 202.140 87.940 202.200 ;
        RECT 88.095 202.155 88.385 202.385 ;
        RECT 72.915 201.815 73.205 202.045 ;
        RECT 75.240 202.000 75.530 202.045 ;
        RECT 77.340 202.000 77.630 202.045 ;
        RECT 78.910 202.000 79.200 202.045 ;
        RECT 86.700 202.000 87.020 202.060 ;
        RECT 75.240 201.860 79.200 202.000 ;
        RECT 75.240 201.815 75.530 201.860 ;
        RECT 77.340 201.815 77.630 201.860 ;
        RECT 78.910 201.815 79.200 201.860 ;
        RECT 84.950 201.860 87.020 202.000 ;
        RECT 84.950 201.720 85.090 201.860 ;
        RECT 86.700 201.800 87.020 201.860 ;
        RECT 87.160 202.000 87.480 202.060 ;
        RECT 88.170 202.000 88.310 202.155 ;
        RECT 87.160 201.860 88.310 202.000 ;
        RECT 90.930 202.000 91.070 202.495 ;
        RECT 93.230 202.340 93.370 202.495 ;
        RECT 97.740 202.340 98.060 202.400 ;
        RECT 98.750 202.340 98.890 202.835 ;
        RECT 100.960 202.820 101.280 202.880 ;
        RECT 102.340 202.820 102.660 203.080 ;
        RECT 102.890 203.020 103.030 203.220 ;
        RECT 103.720 203.160 104.040 203.420 ;
        RECT 105.100 203.360 105.420 203.420 ;
        RECT 104.270 203.220 105.420 203.360 ;
        RECT 104.270 203.020 104.410 203.220 ;
        RECT 105.100 203.160 105.420 203.220 ;
        RECT 123.040 203.360 123.360 203.420 ;
        RECT 134.555 203.360 134.845 203.405 ;
        RECT 139.140 203.360 139.460 203.420 ;
        RECT 141.455 203.360 141.745 203.405 ;
        RECT 141.900 203.360 142.220 203.420 ;
        RECT 123.040 203.220 137.070 203.360 ;
        RECT 123.040 203.160 123.360 203.220 ;
        RECT 134.555 203.175 134.845 203.220 ;
        RECT 102.890 202.880 104.410 203.020 ;
        RECT 104.640 202.820 104.960 203.080 ;
        RECT 111.080 203.020 111.400 203.080 ;
        RECT 112.980 203.020 113.270 203.065 ;
        RECT 111.080 202.880 113.270 203.020 ;
        RECT 111.080 202.820 111.400 202.880 ;
        RECT 112.980 202.835 113.270 202.880 ;
        RECT 114.760 203.020 115.080 203.080 ;
        RECT 127.640 203.020 127.960 203.080 ;
        RECT 114.760 202.880 127.960 203.020 ;
        RECT 136.930 203.020 137.070 203.220 ;
        RECT 139.140 203.220 141.210 203.360 ;
        RECT 139.140 203.160 139.460 203.220 ;
        RECT 136.930 202.880 138.450 203.020 ;
        RECT 114.760 202.820 115.080 202.880 ;
        RECT 127.640 202.820 127.960 202.880 ;
        RECT 101.895 202.680 102.185 202.725 ;
        RECT 93.230 202.200 98.060 202.340 ;
        RECT 97.740 202.140 98.060 202.200 ;
        RECT 98.290 202.200 98.890 202.340 ;
        RECT 99.210 202.540 102.185 202.680 ;
        RECT 92.220 202.000 92.540 202.060 ;
        RECT 93.140 202.000 93.460 202.060 ;
        RECT 98.290 202.000 98.430 202.200 ;
        RECT 90.930 201.860 98.430 202.000 ;
        RECT 87.160 201.800 87.480 201.860 ;
        RECT 92.220 201.800 92.540 201.860 ;
        RECT 93.140 201.800 93.460 201.860 ;
        RECT 76.120 201.660 76.440 201.720 ;
        RECT 70.230 201.520 76.440 201.660 ;
        RECT 76.120 201.460 76.440 201.520 ;
        RECT 84.860 201.460 85.180 201.720 ;
        RECT 85.320 201.460 85.640 201.720 ;
        RECT 88.080 201.660 88.400 201.720 ;
        RECT 88.555 201.660 88.845 201.705 ;
        RECT 88.080 201.520 88.845 201.660 ;
        RECT 88.080 201.460 88.400 201.520 ;
        RECT 88.555 201.475 88.845 201.520 ;
        RECT 94.075 201.660 94.365 201.705 ;
        RECT 95.455 201.660 95.745 201.705 ;
        RECT 94.075 201.520 95.745 201.660 ;
        RECT 94.075 201.475 94.365 201.520 ;
        RECT 95.455 201.475 95.745 201.520 ;
        RECT 98.200 201.660 98.520 201.720 ;
        RECT 98.675 201.660 98.965 201.705 ;
        RECT 99.210 201.660 99.350 202.540 ;
        RECT 101.895 202.495 102.185 202.540 ;
        RECT 106.480 202.680 106.800 202.740 ;
        RECT 114.315 202.680 114.605 202.725 ;
        RECT 117.075 202.680 117.365 202.725 ;
        RECT 117.520 202.680 117.840 202.740 ;
        RECT 118.440 202.725 118.760 202.740 ;
        RECT 106.480 202.540 114.070 202.680 ;
        RECT 106.480 202.480 106.800 202.540 ;
        RECT 109.725 202.340 110.015 202.385 ;
        RECT 112.245 202.340 112.535 202.385 ;
        RECT 113.435 202.340 113.725 202.385 ;
        RECT 100.590 202.200 107.630 202.340 ;
        RECT 100.590 202.060 100.730 202.200 ;
        RECT 100.500 201.800 100.820 202.060 ;
        RECT 105.100 202.000 105.420 202.060 ;
        RECT 106.495 202.000 106.785 202.045 ;
        RECT 105.100 201.860 106.785 202.000 ;
        RECT 105.100 201.800 105.420 201.860 ;
        RECT 106.495 201.815 106.785 201.860 ;
        RECT 98.200 201.520 99.350 201.660 ;
        RECT 98.200 201.460 98.520 201.520 ;
        RECT 98.675 201.475 98.965 201.520 ;
        RECT 99.580 201.460 99.900 201.720 ;
        RECT 103.260 201.460 103.580 201.720 ;
        RECT 103.720 201.660 104.040 201.720 ;
        RECT 107.490 201.705 107.630 202.200 ;
        RECT 109.725 202.200 113.725 202.340 ;
        RECT 113.930 202.340 114.070 202.540 ;
        RECT 114.315 202.540 117.840 202.680 ;
        RECT 114.315 202.495 114.605 202.540 ;
        RECT 117.075 202.495 117.365 202.540 ;
        RECT 117.520 202.480 117.840 202.540 ;
        RECT 118.410 202.495 118.760 202.725 ;
        RECT 131.895 202.680 132.185 202.725 ;
        RECT 134.540 202.680 134.860 202.740 ;
        RECT 131.895 202.540 133.850 202.680 ;
        RECT 134.345 202.540 134.860 202.680 ;
        RECT 131.895 202.495 132.185 202.540 ;
        RECT 118.440 202.480 118.760 202.495 ;
        RECT 116.140 202.340 116.460 202.400 ;
        RECT 113.930 202.200 116.460 202.340 ;
        RECT 109.725 202.155 110.015 202.200 ;
        RECT 112.245 202.155 112.535 202.200 ;
        RECT 113.435 202.155 113.725 202.200 ;
        RECT 116.140 202.140 116.460 202.200 ;
        RECT 117.955 202.340 118.245 202.385 ;
        RECT 119.145 202.340 119.435 202.385 ;
        RECT 121.665 202.340 121.955 202.385 ;
        RECT 117.955 202.200 121.955 202.340 ;
        RECT 117.955 202.155 118.245 202.200 ;
        RECT 119.145 202.155 119.435 202.200 ;
        RECT 121.665 202.155 121.955 202.200 ;
        RECT 128.585 202.340 128.875 202.385 ;
        RECT 131.105 202.340 131.395 202.385 ;
        RECT 132.295 202.340 132.585 202.385 ;
        RECT 128.585 202.200 132.585 202.340 ;
        RECT 128.585 202.155 128.875 202.200 ;
        RECT 131.105 202.155 131.395 202.200 ;
        RECT 132.295 202.155 132.585 202.200 ;
        RECT 133.160 202.140 133.480 202.400 ;
        RECT 133.710 202.340 133.850 202.540 ;
        RECT 134.540 202.480 134.860 202.540 ;
        RECT 136.840 202.480 137.160 202.740 ;
        RECT 138.310 202.725 138.450 202.880 ;
        RECT 139.230 202.725 139.370 203.160 ;
        RECT 137.315 202.495 137.605 202.725 ;
        RECT 138.235 202.495 138.525 202.725 ;
        RECT 139.155 202.495 139.445 202.725 ;
        RECT 139.990 202.680 140.280 202.725 ;
        RECT 141.070 202.680 141.210 203.220 ;
        RECT 141.455 203.220 142.220 203.360 ;
        RECT 141.455 203.175 141.745 203.220 ;
        RECT 141.900 203.160 142.220 203.220 ;
        RECT 142.375 203.360 142.665 203.405 ;
        RECT 142.375 203.220 143.510 203.360 ;
        RECT 142.375 203.175 142.665 203.220 ;
        RECT 143.370 203.080 143.510 203.220 ;
        RECT 144.200 203.160 144.520 203.420 ;
        RECT 143.280 202.820 143.600 203.080 ;
        RECT 142.080 202.680 142.370 202.725 ;
        RECT 139.990 202.670 140.290 202.680 ;
        RECT 139.990 202.530 140.750 202.670 ;
        RECT 141.070 202.540 142.370 202.680 ;
        RECT 139.990 202.495 140.280 202.530 ;
        RECT 135.460 202.340 135.780 202.400 ;
        RECT 133.710 202.200 135.780 202.340 ;
        RECT 135.460 202.140 135.780 202.200 ;
        RECT 110.160 202.000 110.450 202.045 ;
        RECT 111.730 202.000 112.020 202.045 ;
        RECT 113.830 202.000 114.120 202.045 ;
        RECT 110.160 201.860 114.120 202.000 ;
        RECT 110.160 201.815 110.450 201.860 ;
        RECT 111.730 201.815 112.020 201.860 ;
        RECT 113.830 201.815 114.120 201.860 ;
        RECT 117.560 202.000 117.850 202.045 ;
        RECT 119.660 202.000 119.950 202.045 ;
        RECT 121.230 202.000 121.520 202.045 ;
        RECT 117.560 201.860 121.520 202.000 ;
        RECT 117.560 201.815 117.850 201.860 ;
        RECT 119.660 201.815 119.950 201.860 ;
        RECT 121.230 201.815 121.520 201.860 ;
        RECT 129.020 202.000 129.310 202.045 ;
        RECT 130.590 202.000 130.880 202.045 ;
        RECT 132.690 202.000 132.980 202.045 ;
        RECT 129.020 201.860 132.980 202.000 ;
        RECT 129.020 201.815 129.310 201.860 ;
        RECT 130.590 201.815 130.880 201.860 ;
        RECT 132.690 201.815 132.980 201.860 ;
        RECT 133.635 202.000 133.925 202.045 ;
        RECT 137.390 202.000 137.530 202.495 ;
        RECT 138.680 202.140 139.000 202.400 ;
        RECT 140.610 202.340 140.750 202.530 ;
        RECT 142.080 202.495 142.370 202.540 ;
        RECT 143.370 202.340 143.510 202.820 ;
        RECT 144.290 202.725 144.430 203.160 ;
        RECT 144.215 202.495 144.505 202.725 ;
        RECT 144.675 202.680 144.965 202.725 ;
        RECT 147.435 202.680 147.725 202.725 ;
        RECT 149.720 202.680 150.040 202.740 ;
        RECT 144.675 202.540 150.040 202.680 ;
        RECT 144.675 202.495 144.965 202.540 ;
        RECT 147.435 202.495 147.725 202.540 ;
        RECT 149.720 202.480 150.040 202.540 ;
        RECT 140.610 202.200 143.510 202.340 ;
        RECT 142.820 202.000 143.140 202.060 ;
        RECT 145.135 202.000 145.425 202.045 ;
        RECT 133.635 201.860 137.070 202.000 ;
        RECT 137.390 201.860 145.425 202.000 ;
        RECT 133.635 201.815 133.925 201.860 ;
        RECT 104.655 201.660 104.945 201.705 ;
        RECT 103.720 201.520 104.945 201.660 ;
        RECT 103.720 201.460 104.040 201.520 ;
        RECT 104.655 201.475 104.945 201.520 ;
        RECT 107.415 201.660 107.705 201.705 ;
        RECT 107.860 201.660 108.180 201.720 ;
        RECT 107.415 201.520 108.180 201.660 ;
        RECT 107.415 201.475 107.705 201.520 ;
        RECT 107.860 201.460 108.180 201.520 ;
        RECT 110.620 201.660 110.940 201.720 ;
        RECT 115.680 201.660 116.000 201.720 ;
        RECT 117.980 201.660 118.300 201.720 ;
        RECT 120.280 201.660 120.600 201.720 ;
        RECT 110.620 201.520 120.600 201.660 ;
        RECT 110.620 201.460 110.940 201.520 ;
        RECT 115.680 201.460 116.000 201.520 ;
        RECT 117.980 201.460 118.300 201.520 ;
        RECT 120.280 201.460 120.600 201.520 ;
        RECT 123.040 201.660 123.360 201.720 ;
        RECT 123.975 201.660 124.265 201.705 ;
        RECT 123.040 201.520 124.265 201.660 ;
        RECT 123.040 201.460 123.360 201.520 ;
        RECT 123.975 201.475 124.265 201.520 ;
        RECT 126.275 201.660 126.565 201.705 ;
        RECT 128.560 201.660 128.880 201.720 ;
        RECT 134.080 201.660 134.400 201.720 ;
        RECT 126.275 201.520 134.400 201.660 ;
        RECT 126.275 201.475 126.565 201.520 ;
        RECT 128.560 201.460 128.880 201.520 ;
        RECT 134.080 201.460 134.400 201.520 ;
        RECT 136.380 201.460 136.700 201.720 ;
        RECT 136.930 201.660 137.070 201.860 ;
        RECT 142.820 201.800 143.140 201.860 ;
        RECT 145.135 201.815 145.425 201.860 ;
        RECT 138.680 201.660 139.000 201.720 ;
        RECT 136.930 201.520 139.000 201.660 ;
        RECT 138.680 201.460 139.000 201.520 ;
        RECT 140.980 201.460 141.300 201.720 ;
        RECT 146.040 201.460 146.360 201.720 ;
        RECT 22.690 200.840 157.010 201.320 ;
        RECT 37.940 200.640 38.260 200.700 ;
        RECT 38.415 200.640 38.705 200.685 ;
        RECT 37.940 200.500 38.705 200.640 ;
        RECT 37.940 200.440 38.260 200.500 ;
        RECT 38.415 200.455 38.705 200.500 ;
        RECT 40.700 200.640 41.020 200.700 ;
        RECT 42.555 200.640 42.845 200.685 ;
        RECT 40.700 200.500 42.845 200.640 ;
        RECT 40.700 200.440 41.020 200.500 ;
        RECT 42.555 200.455 42.845 200.500 ;
        RECT 44.380 200.640 44.700 200.700 ;
        RECT 44.855 200.640 45.145 200.685 ;
        RECT 44.380 200.500 45.145 200.640 ;
        RECT 44.380 200.440 44.700 200.500 ;
        RECT 44.855 200.455 45.145 200.500 ;
        RECT 45.300 200.440 45.620 200.700 ;
        RECT 52.200 200.440 52.520 200.700 ;
        RECT 54.500 200.440 54.820 200.700 ;
        RECT 55.880 200.440 56.200 200.700 ;
        RECT 57.275 200.640 57.565 200.685 ;
        RECT 58.180 200.640 58.500 200.700 ;
        RECT 57.275 200.500 58.500 200.640 ;
        RECT 57.275 200.455 57.565 200.500 ;
        RECT 58.180 200.440 58.500 200.500 ;
        RECT 60.495 200.640 60.785 200.685 ;
        RECT 62.320 200.640 62.640 200.700 ;
        RECT 60.495 200.500 62.640 200.640 ;
        RECT 60.495 200.455 60.785 200.500 ;
        RECT 62.320 200.440 62.640 200.500 ;
        RECT 63.240 200.440 63.560 200.700 ;
        RECT 66.920 200.440 67.240 200.700 ;
        RECT 67.380 200.640 67.700 200.700 ;
        RECT 68.300 200.640 68.620 200.700 ;
        RECT 71.060 200.640 71.380 200.700 ;
        RECT 67.380 200.500 71.380 200.640 ;
        RECT 67.380 200.440 67.700 200.500 ;
        RECT 68.300 200.440 68.620 200.500 ;
        RECT 71.060 200.440 71.380 200.500 ;
        RECT 71.520 200.640 71.840 200.700 ;
        RECT 75.660 200.640 75.980 200.700 ;
        RECT 71.520 200.500 75.980 200.640 ;
        RECT 71.520 200.440 71.840 200.500 ;
        RECT 75.660 200.440 75.980 200.500 ;
        RECT 86.240 200.440 86.560 200.700 ;
        RECT 87.620 200.440 87.940 200.700 ;
        RECT 88.540 200.640 88.860 200.700 ;
        RECT 89.015 200.640 89.305 200.685 ;
        RECT 102.800 200.640 103.120 200.700 ;
        RECT 88.540 200.500 89.305 200.640 ;
        RECT 88.540 200.440 88.860 200.500 ;
        RECT 89.015 200.455 89.305 200.500 ;
        RECT 97.830 200.500 103.120 200.640 ;
        RECT 41.175 200.300 41.465 200.345 ;
        RECT 39.410 200.160 42.310 200.300 ;
        RECT 35.180 199.620 35.500 199.680 ;
        RECT 39.410 199.665 39.550 200.160 ;
        RECT 41.175 200.115 41.465 200.160 ;
        RECT 38.415 199.620 38.705 199.665 ;
        RECT 35.180 199.480 38.705 199.620 ;
        RECT 35.180 199.420 35.500 199.480 ;
        RECT 38.415 199.435 38.705 199.480 ;
        RECT 39.335 199.435 39.625 199.665 ;
        RECT 41.595 199.630 41.885 199.675 ;
        RECT 42.170 199.665 42.310 200.160 ;
        RECT 41.090 199.490 41.885 199.630 ;
        RECT 38.490 199.280 38.630 199.435 ;
        RECT 39.780 199.280 40.100 199.340 ;
        RECT 38.490 199.140 40.100 199.280 ;
        RECT 41.090 199.280 41.230 199.490 ;
        RECT 41.595 199.445 41.885 199.490 ;
        RECT 42.095 199.435 42.385 199.665 ;
        RECT 43.000 199.420 43.320 199.680 ;
        RECT 41.090 199.170 41.390 199.280 ;
        RECT 41.090 199.140 41.850 199.170 ;
        RECT 39.780 199.080 40.100 199.140 ;
        RECT 41.250 199.030 41.850 199.140 ;
        RECT 43.920 199.080 44.240 199.340 ;
        RECT 44.960 199.280 45.250 199.325 ;
        RECT 45.390 199.280 45.530 200.440 ;
        RECT 45.775 200.115 46.065 200.345 ;
        RECT 47.155 200.300 47.445 200.345 ;
        RECT 49.440 200.300 49.760 200.360 ;
        RECT 47.155 200.160 49.760 200.300 ;
        RECT 47.155 200.115 47.445 200.160 ;
        RECT 45.850 199.620 45.990 200.115 ;
        RECT 49.440 200.100 49.760 200.160 ;
        RECT 54.590 199.960 54.730 200.440 ;
        RECT 55.970 200.300 56.110 200.440 ;
        RECT 55.970 200.160 57.950 200.300 ;
        RECT 54.590 199.820 56.570 199.960 ;
        RECT 46.235 199.620 46.525 199.665 ;
        RECT 45.850 199.480 46.525 199.620 ;
        RECT 46.235 199.435 46.525 199.480 ;
        RECT 47.140 199.620 47.460 199.680 ;
        RECT 51.740 199.620 52.060 199.680 ;
        RECT 47.140 199.480 52.060 199.620 ;
        RECT 47.140 199.420 47.460 199.480 ;
        RECT 51.740 199.420 52.060 199.480 ;
        RECT 53.120 199.420 53.440 199.680 ;
        RECT 56.430 199.665 56.570 199.820 ;
        RECT 57.810 199.665 57.950 200.160 ;
        RECT 61.400 200.100 61.720 200.360 ;
        RECT 61.490 199.960 61.630 200.100 ;
        RECT 59.190 199.820 61.630 199.960 ;
        RECT 59.190 199.665 59.330 199.820 ;
        RECT 53.595 199.435 53.885 199.665 ;
        RECT 55.895 199.435 56.185 199.665 ;
        RECT 56.355 199.435 56.645 199.665 ;
        RECT 57.735 199.435 58.025 199.665 ;
        RECT 59.115 199.435 59.405 199.665 ;
        RECT 47.230 199.280 47.370 199.420 ;
        RECT 44.960 199.140 45.530 199.280 ;
        RECT 45.850 199.140 47.370 199.280 ;
        RECT 53.670 199.280 53.810 199.435 ;
        RECT 55.970 199.280 56.110 199.435 ;
        RECT 57.260 199.280 57.580 199.340 ;
        RECT 53.670 199.140 55.650 199.280 ;
        RECT 55.970 199.140 57.580 199.280 ;
        RECT 57.810 199.280 57.950 199.435 ;
        RECT 59.560 199.420 59.880 199.680 ;
        RECT 60.020 199.620 60.340 199.680 ;
        RECT 60.955 199.620 61.245 199.665 ;
        RECT 60.020 199.480 61.245 199.620 ;
        RECT 60.020 199.420 60.340 199.480 ;
        RECT 60.955 199.435 61.245 199.480 ;
        RECT 63.700 199.620 64.020 199.680 ;
        RECT 64.175 199.620 64.465 199.665 ;
        RECT 66.015 199.620 66.305 199.665 ;
        RECT 67.010 199.620 67.150 200.440 ;
        RECT 82.100 200.300 82.420 200.360 ;
        RECT 63.700 199.480 64.465 199.620 ;
        RECT 63.700 199.420 64.020 199.480 ;
        RECT 64.175 199.435 64.465 199.480 ;
        RECT 64.710 199.480 65.770 199.620 ;
        RECT 64.710 199.340 64.850 199.480 ;
        RECT 58.180 199.280 58.500 199.340 ;
        RECT 57.810 199.140 58.500 199.280 ;
        RECT 44.960 199.095 45.250 199.140 ;
        RECT 41.710 198.940 41.850 199.030 ;
        RECT 45.850 198.940 45.990 199.140 ;
        RECT 41.710 198.800 45.990 198.940 ;
        RECT 54.960 198.740 55.280 199.000 ;
        RECT 55.510 198.940 55.650 199.140 ;
        RECT 57.260 199.080 57.580 199.140 ;
        RECT 58.180 199.080 58.500 199.140 ;
        RECT 61.860 199.080 62.180 199.340 ;
        RECT 64.620 199.080 64.940 199.340 ;
        RECT 65.095 199.095 65.385 199.325 ;
        RECT 65.630 199.280 65.770 199.480 ;
        RECT 66.015 199.480 67.150 199.620 ;
        RECT 70.690 200.160 84.630 200.300 ;
        RECT 66.015 199.435 66.305 199.480 ;
        RECT 70.690 199.280 70.830 200.160 ;
        RECT 82.100 200.100 82.420 200.160 ;
        RECT 79.355 199.620 79.645 199.665 ;
        RECT 81.195 199.620 81.485 199.665 ;
        RECT 81.655 199.620 81.945 199.665 ;
        RECT 79.355 199.480 80.950 199.620 ;
        RECT 79.355 199.435 79.645 199.480 ;
        RECT 65.630 199.140 70.830 199.280 ;
        RECT 75.215 199.280 75.505 199.325 ;
        RECT 77.960 199.280 78.280 199.340 ;
        RECT 75.215 199.140 78.280 199.280 ;
        RECT 75.215 199.095 75.505 199.140 ;
        RECT 58.640 198.940 58.960 199.000 ;
        RECT 55.510 198.800 58.960 198.940 ;
        RECT 61.950 198.940 62.090 199.080 ;
        RECT 65.170 198.940 65.310 199.095 ;
        RECT 77.960 199.080 78.280 199.140 ;
        RECT 79.800 199.080 80.120 199.340 ;
        RECT 80.260 199.080 80.580 199.340 ;
        RECT 80.810 199.280 80.950 199.480 ;
        RECT 81.195 199.480 81.945 199.620 ;
        RECT 81.195 199.435 81.485 199.480 ;
        RECT 81.655 199.435 81.945 199.480 ;
        RECT 80.810 199.140 82.100 199.280 ;
        RECT 67.380 198.940 67.700 199.000 ;
        RECT 61.950 198.800 67.700 198.940 ;
        RECT 58.640 198.740 58.960 198.800 ;
        RECT 67.380 198.740 67.700 198.800 ;
        RECT 67.855 198.940 68.145 198.985 ;
        RECT 68.300 198.940 68.620 199.000 ;
        RECT 67.855 198.800 68.620 198.940 ;
        RECT 67.855 198.755 68.145 198.800 ;
        RECT 68.300 198.740 68.620 198.800 ;
        RECT 78.420 198.740 78.740 199.000 ;
        RECT 81.960 198.940 82.100 199.140 ;
        RECT 83.020 198.940 83.340 199.000 ;
        RECT 81.960 198.800 83.340 198.940 ;
        RECT 84.490 198.940 84.630 200.160 ;
        RECT 84.875 199.435 85.165 199.665 ;
        RECT 86.330 199.620 86.470 200.440 ;
        RECT 87.710 200.300 87.850 200.440 ;
        RECT 97.830 200.300 97.970 200.500 ;
        RECT 102.800 200.440 103.120 200.500 ;
        RECT 104.640 200.440 104.960 200.700 ;
        RECT 105.560 200.440 105.880 200.700 ;
        RECT 106.495 200.640 106.785 200.685 ;
        RECT 110.160 200.640 110.480 200.700 ;
        RECT 116.600 200.640 116.920 200.700 ;
        RECT 106.495 200.500 110.480 200.640 ;
        RECT 106.495 200.455 106.785 200.500 ;
        RECT 110.160 200.440 110.480 200.500 ;
        RECT 111.630 200.500 116.920 200.640 ;
        RECT 100.500 200.300 100.820 200.360 ;
        RECT 87.710 200.160 97.970 200.300 ;
        RECT 98.290 200.160 100.820 200.300 ;
        RECT 86.700 199.960 87.020 200.020 ;
        RECT 94.980 199.960 95.300 200.020 ;
        RECT 86.700 199.820 88.310 199.960 ;
        RECT 86.700 199.760 87.020 199.820 ;
        RECT 88.170 199.665 88.310 199.820 ;
        RECT 94.610 199.820 95.300 199.960 ;
        RECT 87.635 199.620 87.925 199.665 ;
        RECT 86.330 199.480 87.925 199.620 ;
        RECT 87.635 199.435 87.925 199.480 ;
        RECT 88.095 199.435 88.385 199.665 ;
        RECT 89.935 199.620 90.225 199.665 ;
        RECT 92.220 199.620 92.540 199.680 ;
        RECT 94.610 199.665 94.750 199.820 ;
        RECT 94.980 199.760 95.300 199.820 ;
        RECT 89.935 199.480 92.540 199.620 ;
        RECT 89.935 199.435 90.225 199.480 ;
        RECT 84.950 199.280 85.090 199.435 ;
        RECT 92.220 199.420 92.540 199.480 ;
        RECT 94.535 199.435 94.825 199.665 ;
        RECT 95.440 199.420 95.760 199.680 ;
        RECT 98.290 199.665 98.430 200.160 ;
        RECT 100.500 200.100 100.820 200.160 ;
        RECT 103.260 200.300 103.580 200.360 ;
        RECT 103.735 200.300 104.025 200.345 ;
        RECT 103.260 200.160 104.025 200.300 ;
        RECT 103.260 200.100 103.580 200.160 ;
        RECT 103.735 200.115 104.025 200.160 ;
        RECT 104.730 199.960 104.870 200.440 ;
        RECT 99.210 199.820 104.870 199.960 ;
        RECT 98.215 199.435 98.505 199.665 ;
        RECT 98.660 199.420 98.980 199.680 ;
        RECT 94.995 199.280 95.285 199.325 ;
        RECT 99.210 199.280 99.350 199.820 ;
        RECT 105.100 199.420 105.420 199.680 ;
        RECT 108.795 199.620 109.085 199.665 ;
        RECT 105.650 199.480 109.085 199.620 ;
        RECT 84.950 199.140 87.850 199.280 ;
        RECT 87.710 199.000 87.850 199.140 ;
        RECT 94.995 199.140 99.350 199.280 ;
        RECT 99.580 199.280 99.900 199.340 ;
        RECT 105.190 199.280 105.330 199.420 ;
        RECT 105.650 199.325 105.790 199.480 ;
        RECT 108.795 199.435 109.085 199.480 ;
        RECT 109.715 199.435 110.005 199.665 ;
        RECT 99.580 199.140 105.330 199.280 ;
        RECT 94.995 199.095 95.285 199.140 ;
        RECT 99.580 199.080 99.900 199.140 ;
        RECT 87.160 198.940 87.480 199.000 ;
        RECT 84.490 198.800 87.480 198.940 ;
        RECT 83.020 198.740 83.340 198.800 ;
        RECT 87.160 198.740 87.480 198.800 ;
        RECT 87.620 198.740 87.940 199.000 ;
        RECT 97.740 198.740 98.060 199.000 ;
        RECT 99.120 198.740 99.440 199.000 ;
        RECT 101.880 198.940 102.200 199.000 ;
        RECT 103.720 198.940 104.040 199.000 ;
        RECT 101.880 198.800 104.040 198.940 ;
        RECT 105.190 198.940 105.330 199.140 ;
        RECT 105.575 199.095 105.865 199.325 ;
        RECT 106.955 199.280 107.245 199.325 ;
        RECT 106.110 199.140 107.245 199.280 ;
        RECT 106.110 198.940 106.250 199.140 ;
        RECT 106.955 199.095 107.245 199.140 ;
        RECT 107.860 199.080 108.180 199.340 ;
        RECT 109.790 199.280 109.930 199.435 ;
        RECT 110.620 199.420 110.940 199.680 ;
        RECT 111.630 199.665 111.770 200.500 ;
        RECT 116.600 200.440 116.920 200.500 ;
        RECT 117.535 200.640 117.825 200.685 ;
        RECT 118.440 200.640 118.760 200.700 ;
        RECT 135.000 200.640 135.320 200.700 ;
        RECT 117.535 200.500 118.760 200.640 ;
        RECT 117.535 200.455 117.825 200.500 ;
        RECT 118.440 200.440 118.760 200.500 ;
        RECT 130.260 200.500 135.320 200.640 ;
        RECT 112.475 200.300 112.765 200.345 ;
        RECT 117.980 200.300 118.300 200.360 ;
        RECT 112.475 200.160 118.300 200.300 ;
        RECT 112.475 200.115 112.765 200.160 ;
        RECT 117.980 200.100 118.300 200.160 ;
        RECT 127.640 200.300 127.960 200.360 ;
        RECT 130.260 200.300 130.400 200.500 ;
        RECT 135.000 200.440 135.320 200.500 ;
        RECT 138.680 200.440 139.000 200.700 ;
        RECT 140.995 200.640 141.285 200.685 ;
        RECT 141.440 200.640 141.760 200.700 ;
        RECT 140.995 200.500 141.760 200.640 ;
        RECT 140.995 200.455 141.285 200.500 ;
        RECT 141.440 200.440 141.760 200.500 ;
        RECT 141.900 200.440 142.220 200.700 ;
        RECT 127.640 200.160 130.400 200.300 ;
        RECT 138.770 200.300 138.910 200.440 ;
        RECT 139.155 200.300 139.445 200.345 ;
        RECT 138.770 200.160 139.445 200.300 ;
        RECT 127.640 200.100 127.960 200.160 ;
        RECT 139.155 200.115 139.445 200.160 ;
        RECT 119.835 199.960 120.125 200.005 ;
        RECT 114.850 199.820 120.125 199.960 ;
        RECT 111.555 199.435 111.845 199.665 ;
        RECT 113.380 199.420 113.700 199.680 ;
        RECT 114.850 199.665 114.990 199.820 ;
        RECT 119.835 199.775 120.125 199.820 ;
        RECT 123.040 199.760 123.360 200.020 ;
        RECT 141.440 199.960 141.760 200.020 ;
        RECT 140.610 199.820 141.760 199.960 ;
        RECT 114.775 199.435 115.065 199.665 ;
        RECT 115.680 199.420 116.000 199.680 ;
        RECT 116.140 199.420 116.460 199.680 ;
        RECT 116.600 199.620 116.920 199.680 ;
        RECT 118.900 199.620 119.220 199.680 ;
        RECT 116.600 199.480 119.220 199.620 ;
        RECT 116.600 199.420 116.920 199.480 ;
        RECT 118.900 199.420 119.220 199.480 ;
        RECT 125.800 199.620 126.120 199.680 ;
        RECT 126.275 199.620 126.565 199.665 ;
        RECT 125.800 199.480 126.565 199.620 ;
        RECT 125.800 199.420 126.120 199.480 ;
        RECT 126.275 199.435 126.565 199.480 ;
        RECT 128.100 199.420 128.420 199.680 ;
        RECT 136.380 199.620 136.700 199.680 ;
        RECT 140.610 199.620 140.750 199.820 ;
        RECT 141.440 199.760 141.760 199.820 ;
        RECT 141.990 199.960 142.130 200.440 ;
        RECT 142.820 200.100 143.140 200.360 ;
        RECT 146.515 200.115 146.805 200.345 ;
        RECT 149.260 200.300 149.550 200.345 ;
        RECT 150.830 200.300 151.120 200.345 ;
        RECT 152.930 200.300 153.220 200.345 ;
        RECT 149.260 200.160 153.220 200.300 ;
        RECT 149.260 200.115 149.550 200.160 ;
        RECT 150.830 200.115 151.120 200.160 ;
        RECT 152.930 200.115 153.220 200.160 ;
        RECT 144.675 199.960 144.965 200.005 ;
        RECT 141.990 199.820 144.965 199.960 ;
        RECT 136.380 199.480 140.750 199.620 ;
        RECT 136.380 199.420 136.700 199.480 ;
        RECT 109.790 199.140 110.850 199.280 ;
        RECT 105.190 198.800 106.250 198.940 ;
        RECT 110.710 198.940 110.850 199.140 ;
        RECT 111.080 199.080 111.400 199.340 ;
        RECT 123.515 199.280 123.805 199.325 ;
        RECT 111.630 199.140 123.805 199.280 ;
        RECT 111.630 198.940 111.770 199.140 ;
        RECT 123.515 199.095 123.805 199.140 ;
        RECT 140.995 199.280 141.285 199.325 ;
        RECT 141.990 199.280 142.130 199.820 ;
        RECT 144.675 199.775 144.965 199.820 ;
        RECT 146.590 199.680 146.730 200.115 ;
        RECT 148.825 199.960 149.115 200.005 ;
        RECT 151.345 199.960 151.635 200.005 ;
        RECT 152.535 199.960 152.825 200.005 ;
        RECT 148.825 199.820 152.825 199.960 ;
        RECT 148.825 199.775 149.115 199.820 ;
        RECT 151.345 199.775 151.635 199.820 ;
        RECT 152.535 199.775 152.825 199.820 ;
        RECT 142.360 199.620 142.680 199.680 ;
        RECT 143.740 199.620 144.060 199.680 ;
        RECT 146.500 199.620 146.820 199.680 ;
        RECT 153.415 199.620 153.705 199.665 ;
        RECT 142.360 199.480 146.820 199.620 ;
        RECT 142.360 199.420 142.680 199.480 ;
        RECT 143.740 199.420 144.060 199.480 ;
        RECT 146.500 199.420 146.820 199.480 ;
        RECT 151.190 199.480 153.705 199.620 ;
        RECT 140.995 199.140 142.130 199.280 ;
        RECT 140.995 199.095 141.285 199.140 ;
        RECT 151.190 199.000 151.330 199.480 ;
        RECT 153.415 199.435 153.705 199.480 ;
        RECT 152.020 199.325 152.340 199.340 ;
        RECT 152.020 199.095 152.370 199.325 ;
        RECT 152.020 199.080 152.340 199.095 ;
        RECT 110.710 198.800 111.770 198.940 ;
        RECT 101.880 198.740 102.200 198.800 ;
        RECT 103.720 198.740 104.040 198.800 ;
        RECT 114.300 198.740 114.620 199.000 ;
        RECT 127.195 198.940 127.485 198.985 ;
        RECT 128.560 198.940 128.880 199.000 ;
        RECT 127.195 198.800 128.880 198.940 ;
        RECT 127.195 198.755 127.485 198.800 ;
        RECT 128.560 198.740 128.880 198.800 ;
        RECT 141.900 198.740 142.220 199.000 ;
        RECT 142.360 198.740 142.680 199.000 ;
        RECT 151.100 198.740 151.420 199.000 ;
        RECT 22.690 198.120 157.810 198.600 ;
        RECT 36.100 197.920 36.420 197.980 ;
        RECT 53.120 197.920 53.440 197.980 ;
        RECT 56.340 197.920 56.660 197.980 ;
        RECT 36.100 197.780 39.090 197.920 ;
        RECT 36.100 197.720 36.420 197.780 ;
        RECT 30.580 197.285 30.900 197.300 ;
        RECT 30.550 197.055 30.900 197.285 ;
        RECT 37.495 197.055 37.785 197.285 ;
        RECT 30.580 197.040 30.900 197.055 ;
        RECT 29.200 196.700 29.520 196.960 ;
        RECT 30.095 196.900 30.385 196.945 ;
        RECT 31.285 196.900 31.575 196.945 ;
        RECT 33.805 196.900 34.095 196.945 ;
        RECT 30.095 196.760 34.095 196.900 ;
        RECT 30.095 196.715 30.385 196.760 ;
        RECT 31.285 196.715 31.575 196.760 ;
        RECT 33.805 196.715 34.095 196.760 ;
        RECT 37.570 196.900 37.710 197.055 ;
        RECT 37.940 197.040 38.260 197.300 ;
        RECT 38.950 197.285 39.090 197.780 ;
        RECT 44.470 197.780 56.660 197.920 ;
        RECT 41.160 197.625 41.480 197.640 ;
        RECT 41.015 197.395 41.480 197.625 ;
        RECT 41.160 197.380 41.480 197.395 ;
        RECT 42.080 197.580 42.400 197.640 ;
        RECT 43.920 197.580 44.240 197.640 ;
        RECT 42.080 197.440 44.240 197.580 ;
        RECT 42.080 197.380 42.400 197.440 ;
        RECT 43.920 197.380 44.240 197.440 ;
        RECT 38.875 197.240 39.165 197.285 ;
        RECT 44.470 197.240 44.610 197.780 ;
        RECT 53.120 197.720 53.440 197.780 ;
        RECT 56.340 197.720 56.660 197.780 ;
        RECT 56.815 197.920 57.105 197.965 ;
        RECT 57.260 197.920 57.580 197.980 ;
        RECT 56.815 197.780 57.580 197.920 ;
        RECT 56.815 197.735 57.105 197.780 ;
        RECT 57.260 197.720 57.580 197.780 ;
        RECT 57.720 197.720 58.040 197.980 ;
        RECT 70.155 197.920 70.445 197.965 ;
        RECT 62.870 197.780 70.445 197.920 ;
        RECT 57.810 197.580 57.950 197.720 ;
        RECT 49.070 197.440 54.270 197.580 ;
        RECT 49.070 197.285 49.210 197.440 ;
        RECT 38.875 197.100 44.610 197.240 ;
        RECT 38.875 197.055 39.165 197.100 ;
        RECT 48.995 197.055 49.285 197.285 ;
        RECT 49.440 197.240 49.760 197.300 ;
        RECT 50.275 197.240 50.565 197.285 ;
        RECT 49.440 197.100 50.565 197.240 ;
        RECT 49.440 197.040 49.760 197.100 ;
        RECT 50.275 197.055 50.565 197.100 ;
        RECT 54.130 196.960 54.270 197.440 ;
        RECT 57.350 197.440 57.950 197.580 ;
        RECT 55.880 197.230 56.200 197.300 ;
        RECT 57.350 197.285 57.490 197.440 ;
        RECT 56.355 197.230 56.645 197.285 ;
        RECT 55.880 197.090 56.645 197.230 ;
        RECT 55.880 197.040 56.200 197.090 ;
        RECT 56.355 197.055 56.645 197.090 ;
        RECT 57.275 197.055 57.565 197.285 ;
        RECT 57.720 197.040 58.040 197.300 ;
        RECT 58.640 197.240 58.960 197.300 ;
        RECT 62.870 197.285 63.010 197.780 ;
        RECT 70.155 197.735 70.445 197.780 ;
        RECT 96.820 197.920 97.140 197.980 ;
        RECT 99.580 197.920 99.900 197.980 ;
        RECT 102.435 197.920 102.725 197.965 ;
        RECT 96.820 197.780 98.430 197.920 ;
        RECT 64.620 197.285 64.940 197.300 ;
        RECT 62.335 197.240 62.625 197.285 ;
        RECT 58.640 197.100 62.625 197.240 ;
        RECT 58.640 197.040 58.960 197.100 ;
        RECT 62.335 197.055 62.625 197.100 ;
        RECT 62.795 197.055 63.085 197.285 ;
        RECT 64.590 197.055 64.940 197.285 ;
        RECT 70.230 197.240 70.370 197.735 ;
        RECT 96.820 197.720 97.140 197.780 ;
        RECT 76.090 197.580 76.380 197.625 ;
        RECT 78.420 197.580 78.740 197.640 ;
        RECT 76.090 197.440 78.740 197.580 ;
        RECT 76.090 197.395 76.380 197.440 ;
        RECT 78.420 197.380 78.740 197.440 ;
        RECT 92.680 197.580 93.000 197.640 ;
        RECT 98.290 197.580 98.430 197.780 ;
        RECT 99.580 197.780 102.725 197.920 ;
        RECT 99.580 197.720 99.900 197.780 ;
        RECT 102.435 197.735 102.725 197.780 ;
        RECT 106.955 197.920 107.245 197.965 ;
        RECT 113.380 197.920 113.700 197.980 ;
        RECT 106.955 197.780 113.700 197.920 ;
        RECT 106.955 197.735 107.245 197.780 ;
        RECT 113.380 197.720 113.700 197.780 ;
        RECT 144.215 197.735 144.505 197.965 ;
        RECT 101.435 197.580 101.725 197.625 ;
        RECT 92.680 197.440 97.970 197.580 ;
        RECT 98.290 197.440 100.270 197.580 ;
        RECT 92.680 197.380 93.000 197.440 ;
        RECT 73.375 197.240 73.665 197.285 ;
        RECT 70.230 197.100 73.665 197.240 ;
        RECT 73.375 197.055 73.665 197.100 ;
        RECT 83.480 197.240 83.800 197.300 ;
        RECT 97.830 197.285 97.970 197.440 ;
        RECT 85.235 197.240 85.525 197.285 ;
        RECT 83.480 197.100 85.525 197.240 ;
        RECT 64.620 197.040 64.940 197.055 ;
        RECT 83.480 197.040 83.800 197.100 ;
        RECT 85.235 197.055 85.525 197.100 ;
        RECT 97.295 197.055 97.585 197.285 ;
        RECT 97.755 197.055 98.045 197.285 ;
        RECT 98.200 197.240 98.520 197.300 ;
        RECT 98.675 197.240 98.965 197.285 ;
        RECT 99.580 197.240 99.900 197.300 ;
        RECT 98.200 197.100 99.900 197.240 ;
        RECT 100.130 197.240 100.270 197.440 ;
        RECT 101.435 197.440 103.030 197.580 ;
        RECT 101.435 197.395 101.725 197.440 ;
        RECT 101.880 197.240 102.200 197.300 ;
        RECT 100.130 197.100 102.200 197.240 ;
        RECT 41.160 196.900 41.480 196.960 ;
        RECT 37.570 196.760 41.480 196.900 ;
        RECT 29.290 196.220 29.430 196.700 ;
        RECT 29.700 196.560 29.990 196.605 ;
        RECT 31.800 196.560 32.090 196.605 ;
        RECT 33.370 196.560 33.660 196.605 ;
        RECT 37.570 196.560 37.710 196.760 ;
        RECT 41.160 196.700 41.480 196.760 ;
        RECT 49.875 196.900 50.165 196.945 ;
        RECT 51.065 196.900 51.355 196.945 ;
        RECT 53.585 196.900 53.875 196.945 ;
        RECT 49.875 196.760 53.875 196.900 ;
        RECT 49.875 196.715 50.165 196.760 ;
        RECT 51.065 196.715 51.355 196.760 ;
        RECT 53.585 196.715 53.875 196.760 ;
        RECT 54.040 196.900 54.360 196.960 ;
        RECT 63.255 196.900 63.545 196.945 ;
        RECT 54.040 196.760 63.545 196.900 ;
        RECT 54.040 196.700 54.360 196.760 ;
        RECT 63.255 196.715 63.545 196.760 ;
        RECT 64.135 196.900 64.425 196.945 ;
        RECT 65.325 196.900 65.615 196.945 ;
        RECT 67.845 196.900 68.135 196.945 ;
        RECT 64.135 196.760 68.135 196.900 ;
        RECT 64.135 196.715 64.425 196.760 ;
        RECT 65.325 196.715 65.615 196.760 ;
        RECT 67.845 196.715 68.135 196.760 ;
        RECT 29.700 196.420 33.660 196.560 ;
        RECT 29.700 196.375 29.990 196.420 ;
        RECT 31.800 196.375 32.090 196.420 ;
        RECT 33.370 196.375 33.660 196.420 ;
        RECT 33.890 196.420 37.710 196.560 ;
        RECT 39.795 196.560 40.085 196.605 ;
        RECT 49.480 196.560 49.770 196.605 ;
        RECT 51.580 196.560 51.870 196.605 ;
        RECT 53.150 196.560 53.440 196.605 ;
        RECT 39.795 196.420 41.390 196.560 ;
        RECT 33.890 196.280 34.030 196.420 ;
        RECT 39.795 196.375 40.085 196.420 ;
        RECT 31.040 196.220 31.360 196.280 ;
        RECT 29.290 196.080 31.360 196.220 ;
        RECT 31.040 196.020 31.360 196.080 ;
        RECT 33.800 196.020 34.120 196.280 ;
        RECT 37.020 196.220 37.340 196.280 ;
        RECT 41.250 196.265 41.390 196.420 ;
        RECT 49.480 196.420 53.440 196.560 ;
        RECT 49.480 196.375 49.770 196.420 ;
        RECT 51.580 196.375 51.870 196.420 ;
        RECT 53.150 196.375 53.440 196.420 ;
        RECT 54.500 196.560 54.820 196.620 ;
        RECT 58.195 196.560 58.485 196.605 ;
        RECT 54.500 196.420 58.485 196.560 ;
        RECT 54.500 196.360 54.820 196.420 ;
        RECT 58.195 196.375 58.485 196.420 ;
        RECT 59.560 196.360 59.880 196.620 ;
        RECT 40.255 196.220 40.545 196.265 ;
        RECT 37.020 196.080 40.545 196.220 ;
        RECT 37.020 196.020 37.340 196.080 ;
        RECT 40.255 196.035 40.545 196.080 ;
        RECT 41.175 196.035 41.465 196.265 ;
        RECT 55.895 196.220 56.185 196.265 ;
        RECT 59.650 196.220 59.790 196.360 ;
        RECT 55.895 196.080 59.790 196.220 ;
        RECT 63.330 196.220 63.470 196.715 ;
        RECT 74.740 196.700 75.060 196.960 ;
        RECT 75.635 196.900 75.925 196.945 ;
        RECT 76.825 196.900 77.115 196.945 ;
        RECT 79.345 196.900 79.635 196.945 ;
        RECT 75.635 196.760 79.635 196.900 ;
        RECT 75.635 196.715 75.925 196.760 ;
        RECT 76.825 196.715 77.115 196.760 ;
        RECT 79.345 196.715 79.635 196.760 ;
        RECT 83.940 196.700 84.260 196.960 ;
        RECT 84.835 196.900 85.125 196.945 ;
        RECT 86.025 196.900 86.315 196.945 ;
        RECT 88.545 196.900 88.835 196.945 ;
        RECT 84.835 196.760 88.835 196.900 ;
        RECT 84.835 196.715 85.125 196.760 ;
        RECT 86.025 196.715 86.315 196.760 ;
        RECT 88.545 196.715 88.835 196.760 ;
        RECT 94.535 196.715 94.825 196.945 ;
        RECT 97.370 196.900 97.510 197.055 ;
        RECT 98.200 197.040 98.520 197.100 ;
        RECT 98.675 197.055 98.965 197.100 ;
        RECT 99.580 197.040 99.900 197.100 ;
        RECT 101.880 197.040 102.200 197.100 ;
        RECT 102.890 196.960 103.030 197.440 ;
        RECT 103.260 197.380 103.580 197.640 ;
        RECT 106.035 197.580 106.325 197.625 ;
        RECT 109.255 197.580 109.545 197.625 ;
        RECT 106.035 197.440 109.545 197.580 ;
        RECT 106.035 197.395 106.325 197.440 ;
        RECT 109.255 197.395 109.545 197.440 ;
        RECT 114.300 197.580 114.620 197.640 ;
        RECT 115.280 197.580 115.570 197.625 ;
        RECT 127.610 197.580 127.900 197.625 ;
        RECT 128.560 197.580 128.880 197.640 ;
        RECT 114.300 197.440 115.570 197.580 ;
        RECT 114.300 197.380 114.620 197.440 ;
        RECT 115.280 197.395 115.570 197.440 ;
        RECT 117.610 197.440 126.490 197.580 ;
        RECT 103.350 197.240 103.490 197.380 ;
        RECT 107.415 197.240 107.705 197.285 ;
        RECT 107.860 197.240 108.180 197.300 ;
        RECT 103.350 197.100 108.180 197.240 ;
        RECT 107.415 197.055 107.705 197.100 ;
        RECT 107.860 197.040 108.180 197.100 ;
        RECT 108.335 197.240 108.625 197.285 ;
        RECT 108.335 197.100 109.930 197.240 ;
        RECT 108.335 197.055 108.625 197.100 ;
        RECT 102.800 196.900 103.120 196.960 ;
        RECT 108.410 196.900 108.550 197.055 ;
        RECT 97.370 196.760 108.550 196.900 ;
        RECT 63.740 196.560 64.030 196.605 ;
        RECT 65.840 196.560 66.130 196.605 ;
        RECT 67.410 196.560 67.700 196.605 ;
        RECT 74.830 196.560 74.970 196.700 ;
        RECT 63.740 196.420 67.700 196.560 ;
        RECT 63.740 196.375 64.030 196.420 ;
        RECT 65.840 196.375 66.130 196.420 ;
        RECT 67.410 196.375 67.700 196.420 ;
        RECT 68.390 196.420 74.970 196.560 ;
        RECT 75.240 196.560 75.530 196.605 ;
        RECT 77.340 196.560 77.630 196.605 ;
        RECT 78.910 196.560 79.200 196.605 ;
        RECT 75.240 196.420 79.200 196.560 ;
        RECT 68.390 196.280 68.530 196.420 ;
        RECT 75.240 196.375 75.530 196.420 ;
        RECT 77.340 196.375 77.630 196.420 ;
        RECT 78.910 196.375 79.200 196.420 ;
        RECT 84.440 196.560 84.730 196.605 ;
        RECT 86.540 196.560 86.830 196.605 ;
        RECT 88.110 196.560 88.400 196.605 ;
        RECT 84.440 196.420 88.400 196.560 ;
        RECT 84.440 196.375 84.730 196.420 ;
        RECT 86.540 196.375 86.830 196.420 ;
        RECT 88.110 196.375 88.400 196.420 ;
        RECT 90.855 196.560 91.145 196.605 ;
        RECT 94.610 196.560 94.750 196.715 ;
        RECT 102.800 196.700 103.120 196.760 ;
        RECT 103.260 196.560 103.580 196.620 ;
        RECT 109.790 196.605 109.930 197.100 ;
        RECT 117.610 196.960 117.750 197.440 ;
        RECT 126.350 197.300 126.490 197.440 ;
        RECT 127.610 197.440 128.880 197.580 ;
        RECT 127.610 197.395 127.900 197.440 ;
        RECT 128.560 197.380 128.880 197.440 ;
        RECT 117.980 197.240 118.300 197.300 ;
        RECT 118.815 197.240 119.105 197.285 ;
        RECT 117.980 197.100 119.105 197.240 ;
        RECT 117.980 197.040 118.300 197.100 ;
        RECT 118.815 197.055 119.105 197.100 ;
        RECT 126.260 197.040 126.580 197.300 ;
        RECT 135.460 197.040 135.780 197.300 ;
        RECT 142.835 197.240 143.125 197.285 ;
        RECT 144.290 197.240 144.430 197.735 ;
        RECT 146.500 197.720 146.820 197.980 ;
        RECT 148.340 197.720 148.660 197.980 ;
        RECT 145.120 197.625 145.440 197.640 ;
        RECT 145.055 197.395 145.440 197.625 ;
        RECT 145.120 197.380 145.440 197.395 ;
        RECT 146.040 197.380 146.360 197.640 ;
        RECT 146.590 197.580 146.730 197.720 ;
        RECT 146.590 197.440 147.190 197.580 ;
        RECT 142.835 197.100 144.430 197.240 ;
        RECT 142.835 197.055 143.125 197.100 ;
        RECT 146.515 197.055 146.805 197.285 ;
        RECT 147.050 197.240 147.190 197.440 ;
        RECT 147.390 197.240 147.680 197.285 ;
        RECT 147.050 197.100 147.680 197.240 ;
        RECT 147.390 197.055 147.680 197.100 ;
        RECT 112.025 196.900 112.315 196.945 ;
        RECT 114.545 196.900 114.835 196.945 ;
        RECT 115.735 196.900 116.025 196.945 ;
        RECT 112.025 196.760 116.025 196.900 ;
        RECT 112.025 196.715 112.315 196.760 ;
        RECT 114.545 196.715 114.835 196.760 ;
        RECT 115.735 196.715 116.025 196.760 ;
        RECT 116.615 196.900 116.905 196.945 ;
        RECT 117.520 196.900 117.840 196.960 ;
        RECT 116.615 196.760 117.840 196.900 ;
        RECT 116.615 196.715 116.905 196.760 ;
        RECT 117.520 196.700 117.840 196.760 ;
        RECT 118.415 196.900 118.705 196.945 ;
        RECT 119.605 196.900 119.895 196.945 ;
        RECT 122.125 196.900 122.415 196.945 ;
        RECT 118.415 196.760 122.415 196.900 ;
        RECT 118.415 196.715 118.705 196.760 ;
        RECT 119.605 196.715 119.895 196.760 ;
        RECT 122.125 196.715 122.415 196.760 ;
        RECT 127.155 196.900 127.445 196.945 ;
        RECT 128.345 196.900 128.635 196.945 ;
        RECT 130.865 196.900 131.155 196.945 ;
        RECT 146.590 196.900 146.730 197.055 ;
        RECT 147.880 197.040 148.200 197.300 ;
        RECT 149.260 197.040 149.580 197.300 ;
        RECT 152.020 197.040 152.340 197.300 ;
        RECT 127.155 196.760 131.155 196.900 ;
        RECT 127.155 196.715 127.445 196.760 ;
        RECT 128.345 196.715 128.635 196.760 ;
        RECT 130.865 196.715 131.155 196.760 ;
        RECT 142.910 196.760 146.730 196.900 ;
        RECT 104.195 196.560 104.485 196.605 ;
        RECT 90.855 196.420 98.890 196.560 ;
        RECT 90.855 196.375 91.145 196.420 ;
        RECT 68.300 196.220 68.620 196.280 ;
        RECT 63.330 196.080 68.620 196.220 ;
        RECT 55.895 196.035 56.185 196.080 ;
        RECT 68.300 196.020 68.620 196.080 ;
        RECT 70.600 196.020 70.920 196.280 ;
        RECT 81.655 196.220 81.945 196.265 ;
        RECT 87.620 196.220 87.940 196.280 ;
        RECT 81.655 196.080 87.940 196.220 ;
        RECT 81.655 196.035 81.945 196.080 ;
        RECT 87.620 196.020 87.940 196.080 ;
        RECT 91.300 196.020 91.620 196.280 ;
        RECT 94.995 196.220 95.285 196.265 ;
        RECT 96.360 196.220 96.680 196.280 ;
        RECT 96.910 196.265 97.050 196.420 ;
        RECT 98.750 196.280 98.890 196.420 ;
        RECT 103.260 196.420 104.485 196.560 ;
        RECT 103.260 196.360 103.580 196.420 ;
        RECT 104.195 196.375 104.485 196.420 ;
        RECT 109.715 196.375 110.005 196.605 ;
        RECT 112.460 196.560 112.750 196.605 ;
        RECT 114.030 196.560 114.320 196.605 ;
        RECT 116.130 196.560 116.420 196.605 ;
        RECT 112.460 196.420 116.420 196.560 ;
        RECT 112.460 196.375 112.750 196.420 ;
        RECT 114.030 196.375 114.320 196.420 ;
        RECT 116.130 196.375 116.420 196.420 ;
        RECT 118.020 196.560 118.310 196.605 ;
        RECT 120.120 196.560 120.410 196.605 ;
        RECT 121.690 196.560 121.980 196.605 ;
        RECT 118.020 196.420 121.980 196.560 ;
        RECT 118.020 196.375 118.310 196.420 ;
        RECT 120.120 196.375 120.410 196.420 ;
        RECT 121.690 196.375 121.980 196.420 ;
        RECT 126.760 196.560 127.050 196.605 ;
        RECT 128.860 196.560 129.150 196.605 ;
        RECT 130.430 196.560 130.720 196.605 ;
        RECT 126.760 196.420 130.720 196.560 ;
        RECT 126.760 196.375 127.050 196.420 ;
        RECT 128.860 196.375 129.150 196.420 ;
        RECT 130.430 196.375 130.720 196.420 ;
        RECT 142.910 196.280 143.050 196.760 ;
        RECT 143.755 196.560 144.045 196.605 ;
        RECT 152.110 196.560 152.250 197.040 ;
        RECT 143.755 196.420 152.250 196.560 ;
        RECT 143.755 196.375 144.045 196.420 ;
        RECT 94.995 196.080 96.680 196.220 ;
        RECT 94.995 196.035 95.285 196.080 ;
        RECT 96.360 196.020 96.680 196.080 ;
        RECT 96.835 196.035 97.125 196.265 ;
        RECT 98.200 196.020 98.520 196.280 ;
        RECT 98.660 196.020 98.980 196.280 ;
        RECT 100.500 196.220 100.820 196.280 ;
        RECT 102.355 196.220 102.645 196.265 ;
        RECT 100.500 196.080 102.645 196.220 ;
        RECT 100.500 196.020 100.820 196.080 ;
        RECT 102.355 196.035 102.645 196.080 ;
        RECT 103.720 196.220 104.040 196.280 ;
        RECT 105.560 196.220 105.880 196.280 ;
        RECT 106.035 196.220 106.325 196.265 ;
        RECT 103.720 196.080 106.325 196.220 ;
        RECT 103.720 196.020 104.040 196.080 ;
        RECT 105.560 196.020 105.880 196.080 ;
        RECT 106.035 196.035 106.325 196.080 ;
        RECT 124.435 196.220 124.725 196.265 ;
        RECT 125.800 196.220 126.120 196.280 ;
        RECT 129.940 196.220 130.260 196.280 ;
        RECT 124.435 196.080 130.260 196.220 ;
        RECT 124.435 196.035 124.725 196.080 ;
        RECT 125.800 196.020 126.120 196.080 ;
        RECT 129.940 196.020 130.260 196.080 ;
        RECT 133.175 196.220 133.465 196.265 ;
        RECT 134.080 196.220 134.400 196.280 ;
        RECT 133.175 196.080 134.400 196.220 ;
        RECT 133.175 196.035 133.465 196.080 ;
        RECT 134.080 196.020 134.400 196.080 ;
        RECT 134.540 196.020 134.860 196.280 ;
        RECT 142.820 196.020 143.140 196.280 ;
        RECT 145.120 196.020 145.440 196.280 ;
        RECT 145.580 196.220 145.900 196.280 ;
        RECT 146.975 196.220 147.265 196.265 ;
        RECT 148.800 196.220 149.120 196.280 ;
        RECT 145.580 196.080 149.120 196.220 ;
        RECT 145.580 196.020 145.900 196.080 ;
        RECT 146.975 196.035 147.265 196.080 ;
        RECT 148.800 196.020 149.120 196.080 ;
        RECT 150.180 196.020 150.500 196.280 ;
        RECT 22.690 195.400 157.010 195.880 ;
        RECT 30.580 195.200 30.900 195.260 ;
        RECT 31.055 195.200 31.345 195.245 ;
        RECT 37.020 195.200 37.340 195.260 ;
        RECT 30.580 195.060 31.345 195.200 ;
        RECT 30.580 195.000 30.900 195.060 ;
        RECT 31.055 195.015 31.345 195.060 ;
        RECT 33.660 195.060 37.340 195.200 ;
        RECT 33.660 194.520 33.800 195.060 ;
        RECT 37.020 195.000 37.340 195.060 ;
        RECT 42.540 195.000 42.860 195.260 ;
        RECT 54.960 195.000 55.280 195.260 ;
        RECT 68.300 195.200 68.620 195.260 ;
        RECT 67.470 195.060 68.620 195.200 ;
        RECT 35.180 194.660 35.500 194.920 ;
        RECT 36.100 194.660 36.420 194.920 ;
        RECT 52.660 194.860 52.980 194.920 ;
        RECT 54.055 194.860 54.345 194.905 ;
        RECT 52.660 194.720 54.345 194.860 ;
        RECT 52.660 194.660 52.980 194.720 ;
        RECT 54.055 194.675 54.345 194.720 ;
        RECT 32.050 194.380 33.800 194.520 ;
        RECT 32.050 194.225 32.190 194.380 ;
        RECT 31.975 193.995 32.265 194.225 ;
        RECT 33.355 194.180 33.645 194.225 ;
        RECT 34.260 194.180 34.580 194.240 ;
        RECT 33.355 194.040 34.580 194.180 ;
        RECT 33.355 193.995 33.645 194.040 ;
        RECT 34.260 193.980 34.580 194.040 ;
        RECT 35.195 194.180 35.485 194.225 ;
        RECT 36.190 194.180 36.330 194.660 ;
        RECT 54.515 194.520 54.805 194.565 ;
        RECT 55.050 194.520 55.190 195.000 ;
        RECT 54.515 194.380 55.190 194.520 ;
        RECT 63.700 194.520 64.020 194.580 ;
        RECT 66.000 194.520 66.320 194.580 ;
        RECT 67.470 194.565 67.610 195.060 ;
        RECT 68.300 195.000 68.620 195.060 ;
        RECT 83.480 195.000 83.800 195.260 ;
        RECT 87.160 195.000 87.480 195.260 ;
        RECT 91.300 195.000 91.620 195.260 ;
        RECT 99.120 195.200 99.440 195.260 ;
        RECT 100.055 195.200 100.345 195.245 ;
        RECT 99.120 195.060 100.345 195.200 ;
        RECT 99.120 195.000 99.440 195.060 ;
        RECT 100.055 195.015 100.345 195.060 ;
        RECT 102.800 195.000 103.120 195.260 ;
        RECT 103.260 195.000 103.580 195.260 ;
        RECT 128.100 195.000 128.420 195.260 ;
        RECT 129.035 195.200 129.325 195.245 ;
        RECT 130.860 195.200 131.180 195.260 ;
        RECT 133.160 195.200 133.480 195.260 ;
        RECT 129.035 195.060 131.180 195.200 ;
        RECT 129.035 195.015 129.325 195.060 ;
        RECT 130.860 195.000 131.180 195.060 ;
        RECT 131.410 195.060 133.480 195.200 ;
        RECT 67.880 194.860 68.170 194.905 ;
        RECT 69.980 194.860 70.270 194.905 ;
        RECT 71.550 194.860 71.840 194.905 ;
        RECT 67.880 194.720 71.840 194.860 ;
        RECT 67.880 194.675 68.170 194.720 ;
        RECT 69.980 194.675 70.270 194.720 ;
        RECT 71.550 194.675 71.840 194.720 ;
        RECT 74.280 194.860 74.600 194.920 ;
        RECT 87.250 194.860 87.390 195.000 ;
        RECT 74.280 194.720 77.730 194.860 ;
        RECT 74.280 194.660 74.600 194.720 ;
        RECT 77.590 194.565 77.730 194.720 ;
        RECT 84.950 194.720 87.390 194.860 ;
        RECT 63.700 194.380 65.310 194.520 ;
        RECT 54.515 194.335 54.805 194.380 ;
        RECT 63.700 194.320 64.020 194.380 ;
        RECT 35.195 194.040 36.330 194.180 ;
        RECT 35.195 193.995 35.485 194.040 ;
        RECT 53.135 193.995 53.425 194.225 ;
        RECT 33.800 193.640 34.120 193.900 ;
        RECT 34.735 193.655 35.025 193.885 ;
        RECT 32.420 193.300 32.740 193.560 ;
        RECT 34.810 193.500 34.950 193.655 ;
        RECT 36.100 193.640 36.420 193.900 ;
        RECT 37.940 193.640 38.260 193.900 ;
        RECT 53.210 193.840 53.350 193.995 ;
        RECT 53.580 193.980 53.900 194.240 ;
        RECT 59.575 193.995 59.865 194.225 ;
        RECT 57.720 193.840 58.040 193.900 ;
        RECT 59.100 193.840 59.420 193.900 ;
        RECT 53.210 193.700 59.420 193.840 ;
        RECT 57.720 193.640 58.040 193.700 ;
        RECT 59.100 193.640 59.420 193.700 ;
        RECT 38.030 193.500 38.170 193.640 ;
        RECT 59.650 193.560 59.790 193.995 ;
        RECT 60.020 193.980 60.340 194.240 ;
        RECT 63.255 194.180 63.545 194.225 ;
        RECT 64.160 194.180 64.480 194.240 ;
        RECT 65.170 194.225 65.310 194.380 ;
        RECT 65.630 194.380 66.320 194.520 ;
        RECT 65.630 194.225 65.770 194.380 ;
        RECT 66.000 194.320 66.320 194.380 ;
        RECT 67.395 194.335 67.685 194.565 ;
        RECT 68.275 194.520 68.565 194.565 ;
        RECT 69.465 194.520 69.755 194.565 ;
        RECT 71.985 194.520 72.275 194.565 ;
        RECT 68.275 194.380 72.275 194.520 ;
        RECT 68.275 194.335 68.565 194.380 ;
        RECT 69.465 194.335 69.755 194.380 ;
        RECT 71.985 194.335 72.275 194.380 ;
        RECT 77.515 194.335 77.805 194.565 ;
        RECT 63.255 194.040 64.480 194.180 ;
        RECT 63.255 193.995 63.545 194.040 ;
        RECT 64.160 193.980 64.480 194.040 ;
        RECT 65.095 193.995 65.385 194.225 ;
        RECT 65.555 194.180 65.845 194.225 ;
        RECT 65.555 194.040 66.690 194.180 ;
        RECT 65.555 193.995 65.845 194.040 ;
        RECT 61.860 193.840 62.180 193.900 ;
        RECT 66.015 193.840 66.305 193.885 ;
        RECT 61.860 193.700 66.305 193.840 ;
        RECT 66.550 193.840 66.690 194.040 ;
        RECT 66.920 193.980 67.240 194.240 ;
        RECT 78.420 194.180 78.740 194.240 ;
        RECT 68.390 194.040 78.740 194.180 ;
        RECT 68.390 193.840 68.530 194.040 ;
        RECT 78.420 193.980 78.740 194.040 ;
        RECT 82.560 193.980 82.880 194.240 ;
        RECT 83.020 194.180 83.340 194.240 ;
        RECT 84.950 194.225 85.090 194.720 ;
        RECT 91.390 194.520 91.530 195.000 ;
        RECT 96.360 194.860 96.680 194.920 ;
        RECT 86.330 194.380 91.530 194.520 ;
        RECT 93.230 194.720 96.680 194.860 ;
        RECT 86.330 194.225 86.470 194.380 ;
        RECT 84.415 194.180 84.705 194.225 ;
        RECT 83.020 194.040 84.705 194.180 ;
        RECT 83.020 193.980 83.340 194.040 ;
        RECT 84.415 193.995 84.705 194.040 ;
        RECT 84.875 193.995 85.165 194.225 ;
        RECT 86.255 193.995 86.545 194.225 ;
        RECT 87.620 193.980 87.940 194.240 ;
        RECT 88.095 194.180 88.385 194.225 ;
        RECT 92.680 194.180 93.000 194.240 ;
        RECT 93.230 194.225 93.370 194.720 ;
        RECT 96.360 194.660 96.680 194.720 ;
        RECT 100.515 194.520 100.805 194.565 ;
        RECT 102.890 194.520 103.030 195.000 ;
        RECT 95.570 194.380 98.135 194.520 ;
        RECT 88.095 194.040 93.000 194.180 ;
        RECT 88.095 193.995 88.385 194.040 ;
        RECT 92.680 193.980 93.000 194.040 ;
        RECT 93.155 193.995 93.445 194.225 ;
        RECT 94.075 193.995 94.365 194.225 ;
        RECT 94.535 193.995 94.825 194.225 ;
        RECT 94.980 194.180 95.300 194.240 ;
        RECT 95.570 194.180 95.710 194.380 ;
        RECT 97.995 194.225 98.135 194.380 ;
        RECT 100.515 194.380 103.030 194.520 ;
        RECT 100.515 194.335 100.805 194.380 ;
        RECT 103.350 194.225 103.490 195.000 ;
        RECT 106.060 194.860 106.350 194.905 ;
        RECT 108.160 194.860 108.450 194.905 ;
        RECT 109.730 194.860 110.020 194.905 ;
        RECT 106.060 194.720 110.020 194.860 ;
        RECT 106.060 194.675 106.350 194.720 ;
        RECT 108.160 194.675 108.450 194.720 ;
        RECT 109.730 194.675 110.020 194.720 ;
        RECT 104.640 194.520 104.960 194.580 ;
        RECT 103.810 194.380 104.960 194.520 ;
        RECT 103.810 194.225 103.950 194.380 ;
        RECT 104.640 194.320 104.960 194.380 ;
        RECT 106.455 194.520 106.745 194.565 ;
        RECT 107.645 194.520 107.935 194.565 ;
        RECT 110.165 194.520 110.455 194.565 ;
        RECT 106.455 194.380 110.455 194.520 ;
        RECT 106.455 194.335 106.745 194.380 ;
        RECT 107.645 194.335 107.935 194.380 ;
        RECT 110.165 194.335 110.455 194.380 ;
        RECT 126.260 194.520 126.580 194.580 ;
        RECT 131.410 194.565 131.550 195.060 ;
        RECT 133.160 195.000 133.480 195.060 ;
        RECT 136.380 195.000 136.700 195.260 ;
        RECT 144.675 195.200 144.965 195.245 ;
        RECT 145.120 195.200 145.440 195.260 ;
        RECT 144.675 195.060 145.440 195.200 ;
        RECT 144.675 195.015 144.965 195.060 ;
        RECT 145.120 195.000 145.440 195.060 ;
        RECT 146.975 195.015 147.265 195.245 ;
        RECT 147.895 195.200 148.185 195.245 ;
        RECT 149.260 195.200 149.580 195.260 ;
        RECT 147.895 195.060 149.580 195.200 ;
        RECT 147.895 195.015 148.185 195.060 ;
        RECT 131.820 194.860 132.110 194.905 ;
        RECT 133.920 194.860 134.210 194.905 ;
        RECT 135.490 194.860 135.780 194.905 ;
        RECT 131.820 194.720 135.780 194.860 ;
        RECT 136.470 194.860 136.610 195.000 ;
        RECT 146.040 194.860 146.360 194.920 ;
        RECT 147.050 194.860 147.190 195.015 ;
        RECT 149.260 195.000 149.580 195.060 ;
        RECT 150.180 195.000 150.500 195.260 ;
        RECT 136.470 194.720 147.190 194.860 ;
        RECT 131.820 194.675 132.110 194.720 ;
        RECT 133.920 194.675 134.210 194.720 ;
        RECT 135.490 194.675 135.780 194.720 ;
        RECT 146.040 194.660 146.360 194.720 ;
        RECT 131.335 194.520 131.625 194.565 ;
        RECT 126.260 194.380 131.625 194.520 ;
        RECT 126.260 194.320 126.580 194.380 ;
        RECT 131.335 194.335 131.625 194.380 ;
        RECT 132.215 194.520 132.505 194.565 ;
        RECT 133.405 194.520 133.695 194.565 ;
        RECT 135.925 194.520 136.215 194.565 ;
        RECT 132.215 194.380 136.215 194.520 ;
        RECT 132.215 194.335 132.505 194.380 ;
        RECT 133.405 194.335 133.695 194.380 ;
        RECT 135.925 194.335 136.215 194.380 ;
        RECT 136.470 194.380 146.730 194.520 ;
        RECT 94.980 194.040 95.710 194.180 ;
        RECT 68.760 193.885 69.080 193.900 ;
        RECT 66.550 193.700 68.530 193.840 ;
        RECT 61.860 193.640 62.180 193.700 ;
        RECT 66.015 193.655 66.305 193.700 ;
        RECT 68.730 193.655 69.080 193.885 ;
        RECT 68.760 193.640 69.080 193.655 ;
        RECT 34.810 193.360 38.170 193.500 ;
        RECT 58.640 193.300 58.960 193.560 ;
        RECT 59.560 193.300 59.880 193.560 ;
        RECT 62.780 193.300 63.100 193.560 ;
        RECT 64.175 193.500 64.465 193.545 ;
        RECT 69.220 193.500 69.540 193.560 ;
        RECT 64.175 193.360 69.540 193.500 ;
        RECT 64.175 193.315 64.465 193.360 ;
        RECT 69.220 193.300 69.540 193.360 ;
        RECT 74.740 193.300 75.060 193.560 ;
        RECT 77.500 193.500 77.820 193.560 ;
        RECT 79.815 193.500 80.105 193.545 ;
        RECT 77.500 193.360 80.105 193.500 ;
        RECT 82.650 193.500 82.790 193.980 ;
        RECT 85.320 193.640 85.640 193.900 ;
        RECT 94.150 193.560 94.290 193.995 ;
        RECT 94.610 193.840 94.750 193.995 ;
        RECT 94.980 193.980 95.300 194.040 ;
        RECT 95.915 193.995 96.205 194.225 ;
        RECT 97.920 193.995 98.210 194.225 ;
        RECT 101.895 193.995 102.185 194.225 ;
        RECT 102.815 193.995 103.105 194.225 ;
        RECT 103.275 193.995 103.565 194.225 ;
        RECT 103.735 193.995 104.025 194.225 ;
        RECT 105.560 194.180 105.880 194.240 ;
        RECT 108.780 194.180 109.100 194.240 ;
        RECT 105.560 194.040 109.100 194.180 ;
        RECT 95.440 193.840 95.760 193.900 ;
        RECT 94.610 193.700 95.760 193.840 ;
        RECT 95.990 193.840 96.130 193.995 ;
        RECT 95.990 193.700 97.970 193.840 ;
        RECT 95.440 193.640 95.760 193.700 ;
        RECT 97.830 193.560 97.970 193.700 ;
        RECT 101.970 193.560 102.110 193.995 ;
        RECT 94.060 193.500 94.380 193.560 ;
        RECT 82.650 193.360 94.380 193.500 ;
        RECT 77.500 193.300 77.820 193.360 ;
        RECT 79.815 193.315 80.105 193.360 ;
        RECT 94.060 193.300 94.380 193.360 ;
        RECT 96.820 193.300 97.140 193.560 ;
        RECT 97.280 193.300 97.600 193.560 ;
        RECT 97.740 193.500 98.060 193.560 ;
        RECT 98.215 193.500 98.505 193.545 ;
        RECT 97.740 193.360 98.505 193.500 ;
        RECT 97.740 193.300 98.060 193.360 ;
        RECT 98.215 193.315 98.505 193.360 ;
        RECT 101.880 193.300 102.200 193.560 ;
        RECT 102.890 193.500 103.030 193.995 ;
        RECT 105.560 193.980 105.880 194.040 ;
        RECT 108.780 193.980 109.100 194.040 ;
        RECT 130.875 194.180 131.165 194.225 ;
        RECT 131.780 194.180 132.100 194.240 ;
        RECT 136.470 194.180 136.610 194.380 ;
        RECT 130.875 194.040 132.100 194.180 ;
        RECT 130.875 193.995 131.165 194.040 ;
        RECT 131.780 193.980 132.100 194.040 ;
        RECT 132.330 194.040 136.610 194.180 ;
        RECT 138.220 194.180 138.540 194.240 ;
        RECT 139.155 194.180 139.445 194.225 ;
        RECT 138.220 194.040 139.445 194.180 ;
        RECT 105.115 193.840 105.405 193.885 ;
        RECT 106.800 193.840 107.090 193.885 ;
        RECT 105.115 193.700 107.090 193.840 ;
        RECT 105.115 193.655 105.405 193.700 ;
        RECT 106.800 193.655 107.090 193.700 ;
        RECT 118.915 193.655 119.205 193.885 ;
        RECT 127.655 193.840 127.945 193.885 ;
        RECT 132.330 193.840 132.470 194.040 ;
        RECT 138.220 193.980 138.540 194.040 ;
        RECT 139.155 193.995 139.445 194.040 ;
        RECT 140.075 193.995 140.365 194.225 ;
        RECT 140.535 194.180 140.825 194.225 ;
        RECT 140.980 194.180 141.300 194.240 ;
        RECT 140.535 194.040 141.300 194.180 ;
        RECT 140.535 193.995 140.825 194.040 ;
        RECT 127.655 193.700 132.470 193.840 ;
        RECT 132.670 193.840 132.960 193.885 ;
        RECT 134.540 193.840 134.860 193.900 ;
        RECT 132.670 193.700 134.860 193.840 ;
        RECT 127.655 193.655 127.945 193.700 ;
        RECT 132.670 193.655 132.960 193.700 ;
        RECT 103.260 193.500 103.580 193.560 ;
        RECT 102.890 193.360 103.580 193.500 ;
        RECT 103.260 193.300 103.580 193.360 ;
        RECT 106.020 193.500 106.340 193.560 ;
        RECT 111.540 193.500 111.860 193.560 ;
        RECT 106.020 193.360 111.860 193.500 ;
        RECT 106.020 193.300 106.340 193.360 ;
        RECT 111.540 193.300 111.860 193.360 ;
        RECT 112.460 193.300 112.780 193.560 ;
        RECT 117.520 193.500 117.840 193.560 ;
        RECT 118.990 193.500 119.130 193.655 ;
        RECT 134.540 193.640 134.860 193.700 ;
        RECT 137.760 193.840 138.080 193.900 ;
        RECT 140.150 193.840 140.290 193.995 ;
        RECT 140.980 193.980 141.300 194.040 ;
        RECT 141.455 193.995 141.745 194.225 ;
        RECT 137.760 193.700 140.290 193.840 ;
        RECT 141.530 193.840 141.670 193.995 ;
        RECT 141.900 193.980 142.220 194.240 ;
        RECT 142.360 193.980 142.680 194.240 ;
        RECT 145.135 194.180 145.425 194.225 ;
        RECT 146.040 194.180 146.360 194.240 ;
        RECT 145.135 194.040 146.360 194.180 ;
        RECT 145.135 193.995 145.425 194.040 ;
        RECT 146.040 193.980 146.360 194.040 ;
        RECT 142.450 193.840 142.590 193.980 ;
        RECT 146.590 193.900 146.730 194.380 ;
        RECT 141.530 193.700 142.590 193.840 ;
        RECT 137.760 193.640 138.080 193.700 ;
        RECT 117.520 193.360 119.130 193.500 ;
        RECT 117.520 193.300 117.840 193.360 ;
        RECT 129.020 193.300 129.340 193.560 ;
        RECT 130.860 193.500 131.180 193.560 ;
        RECT 133.160 193.500 133.480 193.560 ;
        RECT 136.380 193.500 136.700 193.560 ;
        RECT 130.860 193.360 136.700 193.500 ;
        RECT 130.860 193.300 131.180 193.360 ;
        RECT 133.160 193.300 133.480 193.360 ;
        RECT 136.380 193.300 136.700 193.360 ;
        RECT 136.840 193.500 137.160 193.560 ;
        RECT 138.235 193.500 138.525 193.545 ;
        RECT 136.840 193.360 138.525 193.500 ;
        RECT 140.150 193.500 140.290 193.700 ;
        RECT 142.820 193.640 143.140 193.900 ;
        RECT 143.740 193.640 144.060 193.900 ;
        RECT 146.500 193.640 146.820 193.900 ;
        RECT 150.270 193.840 150.410 195.000 ;
        RECT 151.100 194.860 151.390 194.905 ;
        RECT 152.670 194.860 152.960 194.905 ;
        RECT 154.770 194.860 155.060 194.905 ;
        RECT 151.100 194.720 155.060 194.860 ;
        RECT 151.100 194.675 151.390 194.720 ;
        RECT 152.670 194.675 152.960 194.720 ;
        RECT 154.770 194.675 155.060 194.720 ;
        RECT 150.665 194.520 150.955 194.565 ;
        RECT 153.185 194.520 153.475 194.565 ;
        RECT 154.375 194.520 154.665 194.565 ;
        RECT 150.665 194.380 154.665 194.520 ;
        RECT 150.665 194.335 150.955 194.380 ;
        RECT 153.185 194.335 153.475 194.380 ;
        RECT 154.375 194.335 154.665 194.380 ;
        RECT 151.100 194.180 151.420 194.240 ;
        RECT 155.255 194.180 155.545 194.225 ;
        RECT 151.100 194.040 155.545 194.180 ;
        RECT 151.100 193.980 151.420 194.040 ;
        RECT 155.255 193.995 155.545 194.040 ;
        RECT 153.920 193.840 154.210 193.885 ;
        RECT 150.270 193.700 154.210 193.840 ;
        RECT 153.920 193.655 154.210 193.700 ;
        RECT 142.360 193.500 142.680 193.560 ;
        RECT 140.150 193.360 142.680 193.500 ;
        RECT 136.840 193.300 137.160 193.360 ;
        RECT 138.235 193.315 138.525 193.360 ;
        RECT 142.360 193.300 142.680 193.360 ;
        RECT 146.975 193.500 147.265 193.545 ;
        RECT 147.420 193.500 147.740 193.560 ;
        RECT 146.975 193.360 147.740 193.500 ;
        RECT 146.975 193.315 147.265 193.360 ;
        RECT 147.420 193.300 147.740 193.360 ;
        RECT 147.880 193.500 148.200 193.560 ;
        RECT 148.355 193.500 148.645 193.545 ;
        RECT 147.880 193.360 148.645 193.500 ;
        RECT 147.880 193.300 148.200 193.360 ;
        RECT 148.355 193.315 148.645 193.360 ;
        RECT 22.690 192.680 157.810 193.160 ;
        RECT 34.260 192.480 34.580 192.540 ;
        RECT 38.415 192.480 38.705 192.525 ;
        RECT 42.080 192.480 42.400 192.540 ;
        RECT 34.260 192.340 38.705 192.480 ;
        RECT 34.260 192.280 34.580 192.340 ;
        RECT 38.415 192.295 38.705 192.340 ;
        RECT 40.330 192.340 42.400 192.480 ;
        RECT 32.420 192.185 32.740 192.200 ;
        RECT 40.330 192.185 40.470 192.340 ;
        RECT 42.080 192.280 42.400 192.340 ;
        RECT 55.895 192.295 56.185 192.525 ;
        RECT 64.175 192.480 64.465 192.525 ;
        RECT 64.620 192.480 64.940 192.540 ;
        RECT 64.175 192.340 64.940 192.480 ;
        RECT 64.175 192.295 64.465 192.340 ;
        RECT 32.390 192.140 32.740 192.185 ;
        RECT 32.225 192.000 32.740 192.140 ;
        RECT 32.390 191.955 32.740 192.000 ;
        RECT 39.255 192.140 39.545 192.185 ;
        RECT 39.255 192.000 40.010 192.140 ;
        RECT 39.255 191.955 39.545 192.000 ;
        RECT 32.420 191.940 32.740 191.955 ;
        RECT 31.040 191.260 31.360 191.520 ;
        RECT 31.935 191.460 32.225 191.505 ;
        RECT 33.125 191.460 33.415 191.505 ;
        RECT 35.645 191.460 35.935 191.505 ;
        RECT 31.935 191.320 35.935 191.460 ;
        RECT 39.870 191.460 40.010 192.000 ;
        RECT 40.255 191.955 40.545 192.185 ;
        RECT 41.160 192.140 41.480 192.200 ;
        RECT 42.555 192.140 42.845 192.185 ;
        RECT 55.970 192.140 56.110 192.295 ;
        RECT 64.620 192.280 64.940 192.340 ;
        RECT 66.920 192.480 67.240 192.540 ;
        RECT 67.855 192.480 68.145 192.525 ;
        RECT 66.920 192.340 68.145 192.480 ;
        RECT 66.920 192.280 67.240 192.340 ;
        RECT 67.855 192.295 68.145 192.340 ;
        RECT 68.315 192.480 68.605 192.525 ;
        RECT 68.760 192.480 69.080 192.540 ;
        RECT 74.740 192.480 75.060 192.540 ;
        RECT 68.315 192.340 69.080 192.480 ;
        RECT 68.315 192.295 68.605 192.340 ;
        RECT 68.760 192.280 69.080 192.340 ;
        RECT 71.150 192.340 75.060 192.480 ;
        RECT 41.160 192.000 44.610 192.140 ;
        RECT 41.160 191.940 41.480 192.000 ;
        RECT 42.555 191.955 42.845 192.000 ;
        RECT 41.635 191.800 41.925 191.845 ;
        RECT 43.000 191.800 43.320 191.860 ;
        RECT 41.635 191.660 43.320 191.800 ;
        RECT 41.635 191.615 41.925 191.660 ;
        RECT 43.000 191.600 43.320 191.660 ;
        RECT 43.935 191.800 44.225 191.845 ;
        RECT 44.470 191.800 44.610 192.000 ;
        RECT 49.070 192.000 54.270 192.140 ;
        RECT 55.970 192.000 58.870 192.140 ;
        RECT 43.935 191.660 44.610 191.800 ;
        RECT 43.935 191.615 44.225 191.660 ;
        RECT 46.220 191.600 46.540 191.860 ;
        RECT 49.070 191.845 49.210 192.000 ;
        RECT 54.130 191.860 54.270 192.000 ;
        RECT 48.995 191.615 49.285 191.845 ;
        RECT 50.275 191.800 50.565 191.845 ;
        RECT 49.530 191.660 50.565 191.800 ;
        RECT 43.475 191.460 43.765 191.505 ;
        RECT 49.530 191.460 49.670 191.660 ;
        RECT 50.275 191.615 50.565 191.660 ;
        RECT 54.040 191.600 54.360 191.860 ;
        RECT 58.730 191.845 58.870 192.000 ;
        RECT 61.490 192.000 70.830 192.140 ;
        RECT 58.195 191.615 58.485 191.845 ;
        RECT 58.655 191.800 58.945 191.845 ;
        RECT 59.100 191.800 59.420 191.860 ;
        RECT 58.655 191.660 59.420 191.800 ;
        RECT 58.655 191.615 58.945 191.660 ;
        RECT 39.870 191.320 43.765 191.460 ;
        RECT 31.935 191.275 32.225 191.320 ;
        RECT 33.125 191.275 33.415 191.320 ;
        RECT 35.645 191.275 35.935 191.320 ;
        RECT 43.475 191.275 43.765 191.320 ;
        RECT 47.230 191.320 49.670 191.460 ;
        RECT 49.875 191.460 50.165 191.505 ;
        RECT 51.065 191.460 51.355 191.505 ;
        RECT 53.585 191.460 53.875 191.505 ;
        RECT 49.875 191.320 53.875 191.460 ;
        RECT 58.270 191.460 58.410 191.615 ;
        RECT 59.100 191.600 59.420 191.660 ;
        RECT 60.020 191.600 60.340 191.860 ;
        RECT 61.490 191.845 61.630 192.000 ;
        RECT 70.690 191.860 70.830 192.000 ;
        RECT 61.415 191.615 61.705 191.845 ;
        RECT 61.860 191.800 62.180 191.860 ;
        RECT 62.335 191.800 62.625 191.845 ;
        RECT 61.860 191.660 62.625 191.800 ;
        RECT 61.860 191.600 62.180 191.660 ;
        RECT 62.335 191.615 62.625 191.660 ;
        RECT 62.795 191.615 63.085 191.845 ;
        RECT 63.255 191.820 63.545 191.845 ;
        RECT 63.700 191.820 64.020 191.860 ;
        RECT 63.255 191.800 64.020 191.820 ;
        RECT 67.840 191.800 68.160 191.860 ;
        RECT 69.235 191.820 69.525 191.845 ;
        RECT 68.390 191.800 69.525 191.820 ;
        RECT 63.255 191.680 69.525 191.800 ;
        RECT 63.255 191.615 63.545 191.680 ;
        RECT 63.700 191.660 68.530 191.680 ;
        RECT 62.870 191.460 63.010 191.615 ;
        RECT 63.700 191.600 64.020 191.660 ;
        RECT 67.840 191.600 68.160 191.660 ;
        RECT 69.235 191.615 69.525 191.680 ;
        RECT 69.680 191.600 70.000 191.860 ;
        RECT 70.155 191.615 70.445 191.845 ;
        RECT 64.160 191.460 64.480 191.520 ;
        RECT 64.635 191.460 64.925 191.505 ;
        RECT 58.270 191.320 60.710 191.460 ;
        RECT 62.870 191.320 63.470 191.460 ;
        RECT 31.540 191.120 31.830 191.165 ;
        RECT 33.640 191.120 33.930 191.165 ;
        RECT 35.210 191.120 35.500 191.165 ;
        RECT 31.540 190.980 35.500 191.120 ;
        RECT 31.540 190.935 31.830 190.980 ;
        RECT 33.640 190.935 33.930 190.980 ;
        RECT 35.210 190.935 35.500 190.980 ;
        RECT 37.940 191.120 38.260 191.180 ;
        RECT 47.230 191.165 47.370 191.320 ;
        RECT 49.875 191.275 50.165 191.320 ;
        RECT 51.065 191.275 51.355 191.320 ;
        RECT 53.585 191.275 53.875 191.320 ;
        RECT 37.940 190.980 43.230 191.120 ;
        RECT 37.940 190.920 38.260 190.980 ;
        RECT 43.090 190.840 43.230 190.980 ;
        RECT 47.155 190.935 47.445 191.165 ;
        RECT 49.480 191.120 49.770 191.165 ;
        RECT 51.580 191.120 51.870 191.165 ;
        RECT 53.150 191.120 53.440 191.165 ;
        RECT 60.020 191.120 60.340 191.180 ;
        RECT 49.480 190.980 53.440 191.120 ;
        RECT 49.480 190.935 49.770 190.980 ;
        RECT 51.580 190.935 51.870 190.980 ;
        RECT 53.150 190.935 53.440 190.980 ;
        RECT 53.670 190.980 60.340 191.120 ;
        RECT 60.570 191.120 60.710 191.320 ;
        RECT 62.780 191.120 63.100 191.180 ;
        RECT 60.570 190.980 63.100 191.120 ;
        RECT 63.330 191.120 63.470 191.320 ;
        RECT 64.160 191.320 64.925 191.460 ;
        RECT 64.160 191.260 64.480 191.320 ;
        RECT 64.635 191.275 64.925 191.320 ;
        RECT 70.230 191.180 70.370 191.615 ;
        RECT 70.600 191.600 70.920 191.860 ;
        RECT 71.150 191.845 71.290 192.340 ;
        RECT 74.740 192.280 75.060 192.340 ;
        RECT 94.060 192.480 94.380 192.540 ;
        RECT 94.535 192.480 94.825 192.525 ;
        RECT 94.060 192.340 94.825 192.480 ;
        RECT 94.060 192.280 94.380 192.340 ;
        RECT 94.535 192.295 94.825 192.340 ;
        RECT 101.880 192.480 102.200 192.540 ;
        RECT 103.260 192.480 103.580 192.540 ;
        RECT 106.020 192.480 106.340 192.540 ;
        RECT 101.880 192.340 103.580 192.480 ;
        RECT 101.880 192.280 102.200 192.340 ;
        RECT 103.260 192.280 103.580 192.340 ;
        RECT 103.890 192.340 106.340 192.480 ;
        RECT 103.890 192.270 104.030 192.340 ;
        RECT 106.020 192.280 106.340 192.340 ;
        RECT 108.780 192.480 109.100 192.540 ;
        RECT 127.640 192.480 127.960 192.540 ;
        RECT 134.555 192.480 134.845 192.525 ;
        RECT 135.460 192.480 135.780 192.540 ;
        RECT 142.820 192.480 143.140 192.540 ;
        RECT 144.675 192.480 144.965 192.525 ;
        RECT 146.845 192.480 147.135 192.525 ;
        RECT 108.780 192.340 118.210 192.480 ;
        RECT 108.780 192.280 109.100 192.340 ;
        RECT 74.280 192.140 74.600 192.200 ;
        RECT 72.530 192.000 74.600 192.140 ;
        RECT 72.530 191.845 72.670 192.000 ;
        RECT 74.280 191.940 74.600 192.000 ;
        RECT 74.830 192.000 82.100 192.140 ;
        RECT 74.830 191.860 74.970 192.000 ;
        RECT 71.075 191.615 71.365 191.845 ;
        RECT 72.455 191.615 72.745 191.845 ;
        RECT 74.740 191.600 75.060 191.860 ;
        RECT 75.200 191.800 75.520 191.860 ;
        RECT 76.035 191.800 76.325 191.845 ;
        RECT 75.200 191.660 76.325 191.800 ;
        RECT 81.960 191.800 82.100 192.000 ;
        RECT 97.740 191.940 98.060 192.200 ;
        RECT 103.810 192.185 104.030 192.270 ;
        RECT 102.815 192.140 103.105 192.185 ;
        RECT 102.815 192.000 103.490 192.140 ;
        RECT 103.810 192.000 104.105 192.185 ;
        RECT 102.815 191.955 103.105 192.000 ;
        RECT 83.940 191.800 84.260 191.860 ;
        RECT 81.960 191.660 84.260 191.800 ;
        RECT 75.200 191.600 75.520 191.660 ;
        RECT 76.035 191.615 76.325 191.660 ;
        RECT 83.940 191.600 84.260 191.660 ;
        RECT 84.400 191.800 84.720 191.860 ;
        RECT 85.235 191.800 85.525 191.845 ;
        RECT 84.400 191.660 85.525 191.800 ;
        RECT 84.400 191.600 84.720 191.660 ;
        RECT 85.235 191.615 85.525 191.660 ;
        RECT 92.235 191.800 92.525 191.845 ;
        RECT 92.680 191.800 93.000 191.860 ;
        RECT 92.235 191.660 93.000 191.800 ;
        RECT 92.235 191.615 92.525 191.660 ;
        RECT 92.680 191.600 93.000 191.660 ;
        RECT 94.830 191.800 95.120 191.845 ;
        RECT 95.440 191.800 95.760 191.860 ;
        RECT 94.830 191.660 95.760 191.800 ;
        RECT 94.830 191.615 95.120 191.660 ;
        RECT 95.440 191.600 95.760 191.660 ;
        RECT 75.635 191.460 75.925 191.505 ;
        RECT 76.825 191.460 77.115 191.505 ;
        RECT 79.345 191.460 79.635 191.505 ;
        RECT 75.635 191.320 79.635 191.460 ;
        RECT 75.635 191.275 75.925 191.320 ;
        RECT 76.825 191.275 77.115 191.320 ;
        RECT 79.345 191.275 79.635 191.320 ;
        RECT 84.835 191.460 85.125 191.505 ;
        RECT 86.025 191.460 86.315 191.505 ;
        RECT 88.545 191.460 88.835 191.505 ;
        RECT 84.835 191.320 88.835 191.460 ;
        RECT 103.350 191.460 103.490 192.000 ;
        RECT 103.815 191.955 104.105 192.000 ;
        RECT 112.460 191.940 112.780 192.200 ;
        RECT 104.640 191.800 104.960 191.860 ;
        RECT 105.115 191.800 105.405 191.845 ;
        RECT 104.640 191.660 105.405 191.800 ;
        RECT 104.640 191.600 104.960 191.660 ;
        RECT 105.115 191.615 105.405 191.660 ;
        RECT 108.335 191.800 108.625 191.845 ;
        RECT 109.715 191.800 110.005 191.845 ;
        RECT 112.550 191.800 112.690 191.940 ;
        RECT 108.335 191.660 112.690 191.800 ;
        RECT 116.600 191.845 116.920 191.860 ;
        RECT 108.335 191.615 108.625 191.660 ;
        RECT 109.715 191.615 110.005 191.660 ;
        RECT 116.600 191.615 116.950 191.845 ;
        RECT 117.520 191.800 117.840 191.860 ;
        RECT 118.070 191.845 118.210 192.340 ;
        RECT 127.640 192.340 131.090 192.480 ;
        RECT 127.640 192.280 127.960 192.340 ;
        RECT 120.280 191.940 120.600 192.200 ;
        RECT 129.020 192.140 129.340 192.200 ;
        RECT 130.415 192.140 130.705 192.185 ;
        RECT 129.020 192.000 130.705 192.140 ;
        RECT 129.020 191.940 129.340 192.000 ;
        RECT 130.415 191.955 130.705 192.000 ;
        RECT 117.995 191.800 118.285 191.845 ;
        RECT 117.520 191.660 118.285 191.800 ;
        RECT 108.410 191.460 108.550 191.615 ;
        RECT 116.600 191.600 116.920 191.615 ;
        RECT 117.520 191.600 117.840 191.660 ;
        RECT 117.995 191.615 118.285 191.660 ;
        RECT 118.900 191.800 119.220 191.860 ;
        RECT 119.375 191.800 119.665 191.845 ;
        RECT 118.900 191.660 119.665 191.800 ;
        RECT 118.900 191.600 119.220 191.660 ;
        RECT 119.375 191.615 119.665 191.660 ;
        RECT 119.820 191.600 120.140 191.860 ;
        RECT 121.215 191.800 121.505 191.845 ;
        RECT 126.275 191.800 126.565 191.845 ;
        RECT 121.215 191.660 126.565 191.800 ;
        RECT 121.215 191.615 121.505 191.660 ;
        RECT 126.275 191.615 126.565 191.660 ;
        RECT 128.560 191.800 128.880 191.860 ;
        RECT 130.950 191.845 131.090 192.340 ;
        RECT 134.555 192.340 135.780 192.480 ;
        RECT 134.555 192.295 134.845 192.340 ;
        RECT 135.460 192.280 135.780 192.340 ;
        RECT 140.150 192.340 147.135 192.480 ;
        RECT 133.620 191.940 133.940 192.200 ;
        RECT 134.080 192.140 134.400 192.200 ;
        RECT 134.080 192.000 135.230 192.140 ;
        RECT 134.080 191.940 134.400 192.000 ;
        RECT 129.955 191.800 130.245 191.845 ;
        RECT 130.830 191.830 131.120 191.845 ;
        RECT 128.560 191.660 130.245 191.800 ;
        RECT 128.560 191.600 128.880 191.660 ;
        RECT 129.955 191.615 130.245 191.660 ;
        RECT 130.795 191.615 131.120 191.830 ;
        RECT 131.320 191.800 131.640 191.860 ;
        RECT 134.540 191.800 134.860 191.860 ;
        RECT 135.090 191.845 135.230 192.000 ;
        RECT 131.320 191.660 134.860 191.800 ;
        RECT 103.350 191.320 108.550 191.460 ;
        RECT 113.405 191.460 113.695 191.505 ;
        RECT 115.925 191.460 116.215 191.505 ;
        RECT 117.115 191.460 117.405 191.505 ;
        RECT 113.405 191.320 117.405 191.460 ;
        RECT 84.835 191.275 85.125 191.320 ;
        RECT 86.025 191.275 86.315 191.320 ;
        RECT 88.545 191.275 88.835 191.320 ;
        RECT 113.405 191.275 113.695 191.320 ;
        RECT 115.925 191.275 116.215 191.320 ;
        RECT 117.115 191.275 117.405 191.320 ;
        RECT 129.035 191.460 129.325 191.505 ;
        RECT 130.795 191.460 130.935 191.615 ;
        RECT 131.320 191.600 131.640 191.660 ;
        RECT 134.540 191.600 134.860 191.660 ;
        RECT 135.015 191.615 135.305 191.845 ;
        RECT 135.475 191.460 135.765 191.505 ;
        RECT 129.035 191.320 129.435 191.460 ;
        RECT 130.795 191.320 135.765 191.460 ;
        RECT 129.035 191.275 129.325 191.320 ;
        RECT 135.475 191.275 135.765 191.320 ;
        RECT 66.460 191.120 66.780 191.180 ;
        RECT 63.330 190.980 66.780 191.120 ;
        RECT 39.335 190.780 39.625 190.825 ;
        RECT 40.715 190.780 41.005 190.825 ;
        RECT 39.335 190.640 41.005 190.780 ;
        RECT 39.335 190.595 39.625 190.640 ;
        RECT 40.715 190.595 41.005 190.640 ;
        RECT 43.000 190.780 43.320 190.840 ;
        RECT 53.670 190.780 53.810 190.980 ;
        RECT 60.020 190.920 60.340 190.980 ;
        RECT 62.780 190.920 63.100 190.980 ;
        RECT 66.460 190.920 66.780 190.980 ;
        RECT 70.140 190.920 70.460 191.180 ;
        RECT 75.240 191.120 75.530 191.165 ;
        RECT 77.340 191.120 77.630 191.165 ;
        RECT 78.910 191.120 79.200 191.165 ;
        RECT 75.240 190.980 79.200 191.120 ;
        RECT 75.240 190.935 75.530 190.980 ;
        RECT 77.340 190.935 77.630 190.980 ;
        RECT 78.910 190.935 79.200 190.980 ;
        RECT 81.655 191.120 81.945 191.165 ;
        RECT 82.560 191.120 82.880 191.180 ;
        RECT 81.655 190.980 82.880 191.120 ;
        RECT 81.655 190.935 81.945 190.980 ;
        RECT 82.560 190.920 82.880 190.980 ;
        RECT 84.440 191.120 84.730 191.165 ;
        RECT 86.540 191.120 86.830 191.165 ;
        RECT 88.110 191.120 88.400 191.165 ;
        RECT 84.440 190.980 88.400 191.120 ;
        RECT 84.440 190.935 84.730 190.980 ;
        RECT 86.540 190.935 86.830 190.980 ;
        RECT 88.110 190.935 88.400 190.980 ;
        RECT 90.840 191.120 91.160 191.180 ;
        RECT 94.980 191.120 95.300 191.180 ;
        RECT 90.840 190.980 95.300 191.120 ;
        RECT 90.840 190.920 91.160 190.980 ;
        RECT 94.980 190.920 95.300 190.980 ;
        RECT 95.455 191.120 95.745 191.165 ;
        RECT 95.900 191.120 96.220 191.180 ;
        RECT 99.580 191.120 99.900 191.180 ;
        RECT 112.000 191.120 112.320 191.180 ;
        RECT 95.455 190.980 96.220 191.120 ;
        RECT 95.455 190.935 95.745 190.980 ;
        RECT 95.900 190.920 96.220 190.980 ;
        RECT 96.450 190.980 99.900 191.120 ;
        RECT 43.000 190.640 53.810 190.780 ;
        RECT 56.340 190.780 56.660 190.840 ;
        RECT 57.275 190.780 57.565 190.825 ;
        RECT 56.340 190.640 57.565 190.780 ;
        RECT 43.000 190.580 43.320 190.640 ;
        RECT 56.340 190.580 56.660 190.640 ;
        RECT 57.275 190.595 57.565 190.640 ;
        RECT 59.560 190.780 59.880 190.840 ;
        RECT 71.995 190.780 72.285 190.825 ;
        RECT 59.560 190.640 72.285 190.780 ;
        RECT 59.560 190.580 59.880 190.640 ;
        RECT 71.995 190.595 72.285 190.640 ;
        RECT 92.695 190.780 92.985 190.825 ;
        RECT 96.450 190.780 96.590 190.980 ;
        RECT 99.580 190.920 99.900 190.980 ;
        RECT 102.430 190.980 112.320 191.120 ;
        RECT 102.430 190.840 102.570 190.980 ;
        RECT 112.000 190.920 112.320 190.980 ;
        RECT 113.840 191.120 114.130 191.165 ;
        RECT 115.410 191.120 115.700 191.165 ;
        RECT 117.510 191.120 117.800 191.165 ;
        RECT 129.110 191.120 129.250 191.275 ;
        RECT 131.320 191.120 131.640 191.180 ;
        RECT 113.840 190.980 117.800 191.120 ;
        RECT 113.840 190.935 114.130 190.980 ;
        RECT 115.410 190.935 115.700 190.980 ;
        RECT 117.510 190.935 117.800 190.980 ;
        RECT 128.650 190.980 131.640 191.120 ;
        RECT 92.695 190.640 96.590 190.780 ;
        RECT 96.820 190.780 97.140 190.840 ;
        RECT 97.755 190.780 98.045 190.825 ;
        RECT 96.820 190.640 98.045 190.780 ;
        RECT 92.695 190.595 92.985 190.640 ;
        RECT 96.820 190.580 97.140 190.640 ;
        RECT 97.755 190.595 98.045 190.640 ;
        RECT 98.675 190.780 98.965 190.825 ;
        RECT 99.120 190.780 99.440 190.840 ;
        RECT 98.675 190.640 99.440 190.780 ;
        RECT 98.675 190.595 98.965 190.640 ;
        RECT 99.120 190.580 99.440 190.640 ;
        RECT 102.340 190.580 102.660 190.840 ;
        RECT 102.800 190.780 103.120 190.840 ;
        RECT 103.735 190.780 104.025 190.825 ;
        RECT 102.800 190.640 104.025 190.780 ;
        RECT 102.800 190.580 103.120 190.640 ;
        RECT 103.735 190.595 104.025 190.640 ;
        RECT 104.640 190.580 104.960 190.840 ;
        RECT 108.780 190.780 109.100 190.840 ;
        RECT 109.255 190.780 109.545 190.825 ;
        RECT 108.780 190.640 109.545 190.780 ;
        RECT 108.780 190.580 109.100 190.640 ;
        RECT 109.255 190.595 109.545 190.640 ;
        RECT 110.160 190.780 110.480 190.840 ;
        RECT 111.095 190.780 111.385 190.825 ;
        RECT 110.160 190.640 111.385 190.780 ;
        RECT 110.160 190.580 110.480 190.640 ;
        RECT 111.095 190.595 111.385 190.640 ;
        RECT 118.455 190.780 118.745 190.825 ;
        RECT 118.900 190.780 119.220 190.840 ;
        RECT 118.455 190.640 119.220 190.780 ;
        RECT 118.455 190.595 118.745 190.640 ;
        RECT 118.900 190.580 119.220 190.640 ;
        RECT 124.420 190.780 124.740 190.840 ;
        RECT 128.650 190.780 128.790 190.980 ;
        RECT 131.320 190.920 131.640 190.980 ;
        RECT 131.795 191.120 132.085 191.165 ;
        RECT 140.150 191.120 140.290 192.340 ;
        RECT 142.820 192.280 143.140 192.340 ;
        RECT 144.675 192.295 144.965 192.340 ;
        RECT 146.845 192.295 147.135 192.340 ;
        RECT 147.420 192.480 147.740 192.540 ;
        RECT 148.355 192.480 148.645 192.525 ;
        RECT 147.420 192.340 148.645 192.480 ;
        RECT 147.420 192.280 147.740 192.340 ;
        RECT 148.355 192.295 148.645 192.340 ;
        RECT 141.915 192.140 142.205 192.185 ;
        RECT 143.280 192.140 143.600 192.200 ;
        RECT 141.915 192.000 143.600 192.140 ;
        RECT 141.915 191.955 142.205 192.000 ;
        RECT 143.280 191.940 143.600 192.000 ;
        RECT 143.755 192.140 144.045 192.185 ;
        RECT 147.880 192.140 148.200 192.200 ;
        RECT 143.755 192.000 148.200 192.140 ;
        RECT 143.755 191.955 144.045 192.000 ;
        RECT 147.880 191.940 148.200 192.000 ;
        RECT 142.375 191.800 142.665 191.845 ;
        RECT 142.820 191.800 143.140 191.860 ;
        RECT 142.375 191.660 143.140 191.800 ;
        RECT 142.375 191.615 142.665 191.660 ;
        RECT 142.820 191.600 143.140 191.660 ;
        RECT 144.200 191.600 144.520 191.860 ;
        RECT 148.340 191.600 148.660 191.860 ;
        RECT 148.800 191.800 149.120 191.860 ;
        RECT 149.275 191.800 149.565 191.845 ;
        RECT 148.800 191.660 149.565 191.800 ;
        RECT 148.800 191.600 149.120 191.660 ;
        RECT 149.275 191.615 149.565 191.660 ;
        RECT 144.290 191.460 144.430 191.600 ;
        RECT 144.290 191.320 147.190 191.460 ;
        RECT 131.795 190.980 140.290 191.120 ;
        RECT 131.795 190.935 132.085 190.980 ;
        RECT 124.420 190.640 128.790 190.780 ;
        RECT 130.860 190.780 131.180 190.840 ;
        RECT 131.870 190.780 132.010 190.935 ;
        RECT 130.860 190.640 132.010 190.780 ;
        RECT 133.160 190.780 133.480 190.840 ;
        RECT 133.635 190.780 133.925 190.825 ;
        RECT 133.160 190.640 133.925 190.780 ;
        RECT 124.420 190.580 124.740 190.640 ;
        RECT 130.860 190.580 131.180 190.640 ;
        RECT 133.160 190.580 133.480 190.640 ;
        RECT 133.635 190.595 133.925 190.640 ;
        RECT 145.580 190.580 145.900 190.840 ;
        RECT 146.040 190.580 146.360 190.840 ;
        RECT 147.050 190.825 147.190 191.320 ;
        RECT 146.975 190.595 147.265 190.825 ;
        RECT 22.690 189.960 157.010 190.440 ;
        RECT 41.160 189.560 41.480 189.820 ;
        RECT 45.315 189.575 45.605 189.805 ;
        RECT 41.250 189.420 41.390 189.560 ;
        RECT 43.475 189.420 43.765 189.465 ;
        RECT 41.250 189.280 43.765 189.420 ;
        RECT 45.390 189.420 45.530 189.575 ;
        RECT 46.220 189.560 46.540 189.820 ;
        RECT 46.680 189.560 47.000 189.820 ;
        RECT 47.615 189.760 47.905 189.805 ;
        RECT 50.360 189.760 50.680 189.820 ;
        RECT 47.615 189.620 50.680 189.760 ;
        RECT 47.615 189.575 47.905 189.620 ;
        RECT 50.360 189.560 50.680 189.620 ;
        RECT 53.580 189.560 53.900 189.820 ;
        RECT 59.575 189.760 59.865 189.805 ;
        RECT 61.875 189.760 62.165 189.805 ;
        RECT 54.130 189.620 59.330 189.760 ;
        RECT 50.835 189.420 51.125 189.465 ;
        RECT 45.390 189.280 46.910 189.420 ;
        RECT 43.475 189.235 43.765 189.280 ;
        RECT 43.550 189.080 43.690 189.235 ;
        RECT 46.220 189.080 46.540 189.140 ;
        RECT 43.550 188.940 46.540 189.080 ;
        RECT 46.220 188.880 46.540 188.940 ;
        RECT 31.055 188.740 31.345 188.785 ;
        RECT 32.420 188.740 32.740 188.800 ;
        RECT 31.055 188.600 32.740 188.740 ;
        RECT 31.055 188.555 31.345 188.600 ;
        RECT 32.420 188.540 32.740 188.600 ;
        RECT 45.300 188.540 45.620 188.800 ;
        RECT 46.770 188.740 46.910 189.280 ;
        RECT 48.150 189.280 51.125 189.420 ;
        RECT 48.150 188.740 48.290 189.280 ;
        RECT 50.835 189.235 51.125 189.280 ;
        RECT 49.915 188.740 50.205 188.785 ;
        RECT 54.130 188.740 54.270 189.620 ;
        RECT 54.975 189.420 55.265 189.465 ;
        RECT 57.260 189.420 57.580 189.480 ;
        RECT 54.975 189.280 57.580 189.420 ;
        RECT 54.975 189.235 55.265 189.280 ;
        RECT 57.260 189.220 57.580 189.280 ;
        RECT 59.190 189.140 59.330 189.620 ;
        RECT 59.575 189.620 62.165 189.760 ;
        RECT 59.575 189.575 59.865 189.620 ;
        RECT 61.875 189.575 62.165 189.620 ;
        RECT 64.160 189.760 64.480 189.820 ;
        RECT 64.635 189.760 64.925 189.805 ;
        RECT 64.160 189.620 64.925 189.760 ;
        RECT 64.160 189.560 64.480 189.620 ;
        RECT 64.635 189.575 64.925 189.620 ;
        RECT 65.080 189.760 65.400 189.820 ;
        RECT 70.140 189.760 70.460 189.820 ;
        RECT 65.080 189.620 70.460 189.760 ;
        RECT 65.080 189.560 65.400 189.620 ;
        RECT 70.140 189.560 70.460 189.620 ;
        RECT 74.755 189.760 75.045 189.805 ;
        RECT 75.200 189.760 75.520 189.820 ;
        RECT 74.755 189.620 75.520 189.760 ;
        RECT 74.755 189.575 75.045 189.620 ;
        RECT 75.200 189.560 75.520 189.620 ;
        RECT 83.940 189.760 84.260 189.820 ;
        RECT 84.415 189.760 84.705 189.805 ;
        RECT 83.940 189.620 84.705 189.760 ;
        RECT 83.940 189.560 84.260 189.620 ;
        RECT 84.415 189.575 84.705 189.620 ;
        RECT 95.900 189.560 96.220 189.820 ;
        RECT 104.640 189.560 104.960 189.820 ;
        RECT 108.335 189.760 108.625 189.805 ;
        RECT 109.715 189.760 110.005 189.805 ;
        RECT 108.335 189.620 110.005 189.760 ;
        RECT 108.335 189.575 108.625 189.620 ;
        RECT 109.715 189.575 110.005 189.620 ;
        RECT 110.160 189.560 110.480 189.820 ;
        RECT 111.540 189.560 111.860 189.820 ;
        RECT 112.000 189.560 112.320 189.820 ;
        RECT 115.695 189.760 115.985 189.805 ;
        RECT 116.600 189.760 116.920 189.820 ;
        RECT 115.695 189.620 116.920 189.760 ;
        RECT 115.695 189.575 115.985 189.620 ;
        RECT 116.600 189.560 116.920 189.620 ;
        RECT 117.655 189.620 122.305 189.760 ;
        RECT 67.380 189.420 67.670 189.465 ;
        RECT 68.950 189.420 69.240 189.465 ;
        RECT 71.050 189.420 71.340 189.465 ;
        RECT 67.380 189.280 71.340 189.420 ;
        RECT 67.380 189.235 67.670 189.280 ;
        RECT 68.950 189.235 69.240 189.280 ;
        RECT 71.050 189.235 71.340 189.280 ;
        RECT 55.895 189.080 56.185 189.125 ;
        RECT 56.340 189.080 56.660 189.140 ;
        RECT 55.895 188.940 56.660 189.080 ;
        RECT 55.895 188.895 56.185 188.940 ;
        RECT 56.340 188.880 56.660 188.940 ;
        RECT 58.640 188.880 58.960 189.140 ;
        RECT 59.100 189.080 59.420 189.140 ;
        RECT 63.715 189.080 64.005 189.125 ;
        RECT 59.100 188.940 64.005 189.080 ;
        RECT 59.100 188.880 59.420 188.940 ;
        RECT 63.715 188.895 64.005 188.940 ;
        RECT 66.945 189.080 67.235 189.125 ;
        RECT 69.465 189.080 69.755 189.125 ;
        RECT 70.655 189.080 70.945 189.125 ;
        RECT 66.945 188.940 70.945 189.080 ;
        RECT 66.945 188.895 67.235 188.940 ;
        RECT 69.465 188.895 69.755 188.940 ;
        RECT 70.655 188.895 70.945 188.940 ;
        RECT 90.840 188.880 91.160 189.140 ;
        RECT 46.770 188.600 48.290 188.740 ;
        RECT 48.610 188.600 54.270 188.740 ;
        RECT 31.500 188.400 31.820 188.460 ;
        RECT 31.975 188.400 32.265 188.445 ;
        RECT 31.500 188.260 32.265 188.400 ;
        RECT 45.390 188.400 45.530 188.540 ;
        RECT 48.610 188.445 48.750 188.600 ;
        RECT 49.915 188.555 50.205 188.600 ;
        RECT 54.515 188.555 54.805 188.785 ;
        RECT 55.435 188.555 55.725 188.785 ;
        RECT 47.455 188.400 47.745 188.445 ;
        RECT 45.390 188.260 47.745 188.400 ;
        RECT 31.500 188.200 31.820 188.260 ;
        RECT 31.975 188.215 32.265 188.260 ;
        RECT 47.455 188.215 47.745 188.260 ;
        RECT 48.535 188.215 48.825 188.445 ;
        RECT 48.980 188.200 49.300 188.460 ;
        RECT 54.590 188.120 54.730 188.555 ;
        RECT 32.880 187.860 33.200 188.120 ;
        RECT 33.340 188.060 33.660 188.120 ;
        RECT 45.315 188.060 45.605 188.105 ;
        RECT 33.340 187.920 45.605 188.060 ;
        RECT 33.340 187.860 33.660 187.920 ;
        RECT 45.315 187.875 45.605 187.920 ;
        RECT 54.500 187.860 54.820 188.120 ;
        RECT 54.960 188.060 55.280 188.120 ;
        RECT 55.510 188.060 55.650 188.555 ;
        RECT 56.430 188.400 56.570 188.880 ;
        RECT 56.815 188.740 57.105 188.785 ;
        RECT 58.730 188.740 58.870 188.880 ;
        RECT 56.815 188.600 58.870 188.740 ;
        RECT 56.815 188.555 57.105 188.600 ;
        RECT 60.035 188.555 60.325 188.785 ;
        RECT 60.110 188.400 60.250 188.555 ;
        RECT 62.780 188.540 63.100 188.800 ;
        RECT 68.300 188.740 68.620 188.800 ;
        RECT 71.535 188.740 71.825 188.785 ;
        RECT 68.300 188.600 71.825 188.740 ;
        RECT 68.300 188.540 68.620 188.600 ;
        RECT 71.535 188.555 71.825 188.600 ;
        RECT 75.675 188.740 75.965 188.785 ;
        RECT 77.040 188.740 77.360 188.800 ;
        RECT 75.675 188.600 77.360 188.740 ;
        RECT 75.675 188.555 75.965 188.600 ;
        RECT 77.040 188.540 77.360 188.600 ;
        RECT 77.500 188.540 77.820 188.800 ;
        RECT 77.960 188.540 78.280 188.800 ;
        RECT 83.940 188.740 84.260 188.800 ;
        RECT 88.080 188.740 88.400 188.800 ;
        RECT 83.940 188.600 88.400 188.740 ;
        RECT 95.990 188.740 96.130 189.560 ;
        RECT 96.360 189.420 96.680 189.480 ;
        RECT 99.135 189.420 99.425 189.465 ;
        RECT 96.360 189.280 99.425 189.420 ;
        RECT 96.360 189.220 96.680 189.280 ;
        RECT 99.135 189.235 99.425 189.280 ;
        RECT 96.835 188.740 97.125 188.785 ;
        RECT 95.990 188.600 97.125 188.740 ;
        RECT 83.940 188.540 84.260 188.600 ;
        RECT 88.080 188.540 88.400 188.600 ;
        RECT 96.835 188.555 97.125 188.600 ;
        RECT 97.295 188.740 97.585 188.785 ;
        RECT 98.200 188.740 98.520 188.800 ;
        RECT 97.295 188.600 98.520 188.740 ;
        RECT 104.730 188.740 104.870 189.560 ;
        RECT 105.575 189.420 105.865 189.465 ;
        RECT 109.240 189.420 109.560 189.480 ;
        RECT 105.575 189.280 109.560 189.420 ;
        RECT 105.575 189.235 105.865 189.280 ;
        RECT 109.240 189.220 109.560 189.280 ;
        RECT 110.250 189.080 110.390 189.560 ;
        RECT 110.635 189.235 110.925 189.465 ;
        RECT 112.090 189.420 112.230 189.560 ;
        RECT 117.655 189.420 117.795 189.620 ;
        RECT 112.090 189.280 117.795 189.420 ;
        RECT 118.020 189.420 118.310 189.465 ;
        RECT 120.120 189.420 120.410 189.465 ;
        RECT 121.690 189.420 121.980 189.465 ;
        RECT 118.020 189.280 121.980 189.420 ;
        RECT 122.165 189.420 122.305 189.620 ;
        RECT 124.420 189.560 124.740 189.820 ;
        RECT 127.180 189.760 127.500 189.820 ;
        RECT 128.115 189.760 128.405 189.805 ;
        RECT 127.180 189.620 128.405 189.760 ;
        RECT 127.180 189.560 127.500 189.620 ;
        RECT 128.115 189.575 128.405 189.620 ;
        RECT 129.480 189.560 129.800 189.820 ;
        RECT 130.415 189.760 130.705 189.805 ;
        RECT 132.240 189.760 132.560 189.820 ;
        RECT 130.415 189.620 132.930 189.760 ;
        RECT 130.415 189.575 130.705 189.620 ;
        RECT 132.240 189.560 132.560 189.620 ;
        RECT 126.260 189.420 126.580 189.480 ;
        RECT 122.165 189.280 126.580 189.420 ;
        RECT 118.020 189.235 118.310 189.280 ;
        RECT 120.120 189.235 120.410 189.280 ;
        RECT 121.690 189.235 121.980 189.280 ;
        RECT 106.110 188.940 110.390 189.080 ;
        RECT 110.710 189.080 110.850 189.235 ;
        RECT 126.260 189.220 126.580 189.280 ;
        RECT 129.035 189.420 129.325 189.465 ;
        RECT 132.790 189.420 132.930 189.620 ;
        RECT 133.620 189.560 133.940 189.820 ;
        RECT 134.080 189.560 134.400 189.820 ;
        RECT 136.840 189.560 137.160 189.820 ;
        RECT 134.170 189.420 134.310 189.560 ;
        RECT 129.035 189.280 129.710 189.420 ;
        RECT 132.790 189.280 134.310 189.420 ;
        RECT 129.035 189.235 129.325 189.280 ;
        RECT 110.710 188.940 114.990 189.080 ;
        RECT 106.110 188.785 106.250 188.940 ;
        RECT 105.115 188.740 105.405 188.785 ;
        RECT 104.730 188.600 105.405 188.740 ;
        RECT 97.295 188.555 97.585 188.600 ;
        RECT 98.200 188.540 98.520 188.600 ;
        RECT 105.115 188.555 105.405 188.600 ;
        RECT 106.035 188.740 106.325 188.785 ;
        RECT 107.400 188.750 107.720 188.800 ;
        RECT 107.030 188.740 107.720 188.750 ;
        RECT 111.095 188.740 111.385 188.785 ;
        RECT 106.035 188.610 107.720 188.740 ;
        RECT 106.035 188.600 107.170 188.610 ;
        RECT 106.035 188.555 106.325 188.600 ;
        RECT 56.430 188.260 60.250 188.400 ;
        RECT 69.220 188.400 69.540 188.460 ;
        RECT 70.200 188.400 70.490 188.445 ;
        RECT 69.220 188.260 70.490 188.400 ;
        RECT 69.220 188.200 69.540 188.260 ;
        RECT 70.200 188.215 70.490 188.260 ;
        RECT 75.200 188.400 75.520 188.460 ;
        RECT 76.135 188.400 76.425 188.445 ;
        RECT 75.200 188.260 76.425 188.400 ;
        RECT 75.200 188.200 75.520 188.260 ;
        RECT 76.135 188.215 76.425 188.260 ;
        RECT 76.580 188.200 76.900 188.460 ;
        RECT 95.455 188.400 95.745 188.445 ;
        RECT 97.740 188.400 98.060 188.460 ;
        RECT 100.975 188.400 101.265 188.445 ;
        RECT 95.455 188.260 101.265 188.400 ;
        RECT 105.190 188.400 105.330 188.555 ;
        RECT 107.400 188.540 107.720 188.610 ;
        RECT 109.330 188.600 111.385 188.740 ;
        RECT 106.495 188.400 106.785 188.445 ;
        RECT 105.190 188.260 106.785 188.400 ;
        RECT 95.455 188.215 95.745 188.260 ;
        RECT 97.740 188.200 98.060 188.260 ;
        RECT 100.975 188.215 101.265 188.260 ;
        RECT 106.495 188.215 106.785 188.260 ;
        RECT 106.940 188.400 107.260 188.460 ;
        RECT 108.795 188.400 109.085 188.445 ;
        RECT 106.940 188.260 109.085 188.400 ;
        RECT 58.180 188.060 58.500 188.120 ;
        RECT 54.960 187.920 58.500 188.060 ;
        RECT 54.960 187.860 55.280 187.920 ;
        RECT 58.180 187.860 58.500 187.920 ;
        RECT 87.620 187.860 87.940 188.120 ;
        RECT 96.375 188.060 96.665 188.105 ;
        RECT 96.820 188.060 97.140 188.120 ;
        RECT 96.375 187.920 97.140 188.060 ;
        RECT 96.375 187.875 96.665 187.920 ;
        RECT 96.820 187.860 97.140 187.920 ;
        RECT 98.200 187.860 98.520 188.120 ;
        RECT 98.660 187.860 98.980 188.120 ;
        RECT 106.570 188.060 106.710 188.215 ;
        RECT 106.940 188.200 107.260 188.260 ;
        RECT 108.795 188.215 109.085 188.260 ;
        RECT 109.330 188.060 109.470 188.600 ;
        RECT 111.095 188.555 111.385 188.600 ;
        RECT 112.460 188.740 112.780 188.800 ;
        RECT 114.850 188.785 114.990 188.940 ;
        RECT 117.520 188.880 117.840 189.140 ;
        RECT 118.415 189.080 118.705 189.125 ;
        RECT 119.605 189.080 119.895 189.125 ;
        RECT 122.125 189.080 122.415 189.125 ;
        RECT 127.640 189.080 127.960 189.140 ;
        RECT 118.415 188.940 122.415 189.080 ;
        RECT 118.415 188.895 118.705 188.940 ;
        RECT 119.605 188.895 119.895 188.940 ;
        RECT 122.125 188.895 122.415 188.940 ;
        RECT 125.890 188.940 127.960 189.080 ;
        RECT 129.570 189.080 129.710 189.280 ;
        RECT 130.860 189.080 131.180 189.140 ;
        RECT 129.570 188.940 131.180 189.080 ;
        RECT 118.900 188.785 119.220 188.800 ;
        RECT 125.890 188.785 126.030 188.940 ;
        RECT 127.640 188.880 127.960 188.940 ;
        RECT 130.860 188.880 131.180 188.940 ;
        RECT 113.395 188.740 113.685 188.785 ;
        RECT 112.460 188.600 113.685 188.740 ;
        RECT 112.460 188.540 112.780 188.600 ;
        RECT 113.395 188.555 113.685 188.600 ;
        RECT 114.315 188.555 114.605 188.785 ;
        RECT 114.775 188.555 115.065 188.785 ;
        RECT 118.870 188.740 119.220 188.785 ;
        RECT 118.705 188.600 119.220 188.740 ;
        RECT 118.870 188.555 119.220 188.600 ;
        RECT 125.815 188.555 126.105 188.785 ;
        RECT 126.260 188.740 126.580 188.800 ;
        RECT 126.735 188.740 127.025 188.785 ;
        RECT 131.780 188.740 132.100 188.800 ;
        RECT 126.260 188.600 127.025 188.740 ;
        RECT 114.390 188.400 114.530 188.555 ;
        RECT 118.900 188.540 119.220 188.555 ;
        RECT 126.260 188.540 126.580 188.600 ;
        RECT 126.735 188.555 127.025 188.600 ;
        RECT 130.075 188.600 132.100 188.740 ;
        RECT 111.170 188.260 114.530 188.400 ;
        RECT 127.195 188.400 127.485 188.445 ;
        RECT 127.640 188.400 127.960 188.460 ;
        RECT 127.195 188.260 127.960 188.400 ;
        RECT 106.570 187.920 109.470 188.060 ;
        RECT 109.700 188.105 110.020 188.120 ;
        RECT 109.700 188.060 110.085 188.105 ;
        RECT 111.170 188.060 111.310 188.260 ;
        RECT 127.195 188.215 127.485 188.260 ;
        RECT 127.640 188.200 127.960 188.260 ;
        RECT 128.275 188.400 128.565 188.445 ;
        RECT 129.020 188.400 129.340 188.460 ;
        RECT 130.075 188.400 130.215 188.600 ;
        RECT 131.780 188.540 132.100 188.600 ;
        RECT 134.540 188.740 134.860 188.800 ;
        RECT 135.935 188.740 136.225 188.785 ;
        RECT 134.540 188.600 136.225 188.740 ;
        RECT 134.540 188.540 134.860 188.600 ;
        RECT 135.935 188.555 136.225 188.600 ;
        RECT 137.300 188.740 137.620 188.800 ;
        RECT 143.280 188.740 143.600 188.800 ;
        RECT 137.300 188.600 143.600 188.740 ;
        RECT 137.300 188.540 137.620 188.600 ;
        RECT 143.280 188.540 143.600 188.600 ;
        RECT 128.275 188.260 129.340 188.400 ;
        RECT 128.275 188.215 128.565 188.260 ;
        RECT 129.020 188.200 129.340 188.260 ;
        RECT 129.570 188.260 130.215 188.400 ;
        RECT 131.335 188.400 131.625 188.445 ;
        RECT 132.660 188.400 132.950 188.445 ;
        RECT 131.335 188.260 132.950 188.400 ;
        RECT 109.700 187.920 111.310 188.060 ;
        RECT 109.700 187.875 110.085 187.920 ;
        RECT 109.700 187.860 110.020 187.875 ;
        RECT 113.380 187.860 113.700 188.120 ;
        RECT 126.275 188.060 126.565 188.105 ;
        RECT 129.570 188.060 129.710 188.260 ;
        RECT 131.335 188.215 131.625 188.260 ;
        RECT 132.660 188.215 132.950 188.260 ;
        RECT 130.400 188.105 130.720 188.120 ;
        RECT 126.275 187.920 129.710 188.060 ;
        RECT 126.275 187.875 126.565 187.920 ;
        RECT 130.335 187.875 130.720 188.105 ;
        RECT 131.410 188.060 131.550 188.215 ;
        RECT 146.500 188.200 146.820 188.460 ;
        RECT 135.000 188.060 135.320 188.120 ;
        RECT 136.840 188.060 137.160 188.120 ;
        RECT 131.410 187.920 137.160 188.060 ;
        RECT 130.400 187.860 130.720 187.875 ;
        RECT 135.000 187.860 135.320 187.920 ;
        RECT 136.840 187.860 137.160 187.920 ;
        RECT 137.300 188.060 137.620 188.120 ;
        RECT 138.235 188.060 138.525 188.105 ;
        RECT 137.300 187.920 138.525 188.060 ;
        RECT 137.300 187.860 137.620 187.920 ;
        RECT 138.235 187.875 138.525 187.920 ;
        RECT 151.100 188.060 151.420 188.120 ;
        RECT 152.955 188.060 153.245 188.105 ;
        RECT 151.100 187.920 153.245 188.060 ;
        RECT 151.100 187.860 151.420 187.920 ;
        RECT 152.955 187.875 153.245 187.920 ;
        RECT 22.690 187.240 157.810 187.720 ;
        RECT 31.040 187.040 31.360 187.100 ;
        RECT 24.690 186.900 33.570 187.040 ;
        RECT 24.690 186.405 24.830 186.900 ;
        RECT 31.040 186.840 31.360 186.900 ;
        RECT 32.895 186.515 33.185 186.745 ;
        RECT 33.430 186.700 33.570 186.900 ;
        RECT 48.980 186.840 49.300 187.100 ;
        RECT 52.675 187.040 52.965 187.085 ;
        RECT 54.960 187.040 55.280 187.100 ;
        RECT 52.675 186.900 55.280 187.040 ;
        RECT 52.675 186.855 52.965 186.900 ;
        RECT 54.960 186.840 55.280 186.900 ;
        RECT 57.260 186.840 57.580 187.100 ;
        RECT 67.840 187.040 68.160 187.100 ;
        RECT 68.300 187.040 68.620 187.100 ;
        RECT 64.250 186.900 68.620 187.040 ;
        RECT 33.430 186.560 34.030 186.700 ;
        RECT 25.980 186.405 26.300 186.420 ;
        RECT 24.615 186.175 24.905 186.405 ;
        RECT 25.950 186.175 26.300 186.405 ;
        RECT 32.970 186.360 33.110 186.515 ;
        RECT 33.340 186.360 33.660 186.420 ;
        RECT 32.970 186.220 33.660 186.360 ;
        RECT 25.980 186.160 26.300 186.175 ;
        RECT 33.340 186.160 33.660 186.220 ;
        RECT 25.495 186.020 25.785 186.065 ;
        RECT 26.685 186.020 26.975 186.065 ;
        RECT 29.205 186.020 29.495 186.065 ;
        RECT 25.495 185.880 29.495 186.020 ;
        RECT 25.495 185.835 25.785 185.880 ;
        RECT 26.685 185.835 26.975 185.880 ;
        RECT 29.205 185.835 29.495 185.880 ;
        RECT 25.100 185.680 25.390 185.725 ;
        RECT 27.200 185.680 27.490 185.725 ;
        RECT 28.770 185.680 29.060 185.725 ;
        RECT 25.100 185.540 29.060 185.680 ;
        RECT 25.100 185.495 25.390 185.540 ;
        RECT 27.200 185.495 27.490 185.540 ;
        RECT 28.770 185.495 29.060 185.540 ;
        RECT 31.500 185.480 31.820 185.740 ;
        RECT 31.960 185.140 32.280 185.400 ;
        RECT 32.880 185.140 33.200 185.400 ;
        RECT 33.890 185.340 34.030 186.560 ;
        RECT 35.195 186.360 35.485 186.405 ;
        RECT 34.810 186.220 35.485 186.360 ;
        RECT 34.810 185.740 34.950 186.220 ;
        RECT 35.195 186.175 35.485 186.220 ;
        RECT 36.115 186.360 36.405 186.405 ;
        RECT 36.560 186.360 36.880 186.420 ;
        RECT 36.115 186.220 36.880 186.360 ;
        RECT 36.115 186.175 36.405 186.220 ;
        RECT 36.560 186.160 36.880 186.220 ;
        RECT 37.480 186.360 37.800 186.420 ;
        RECT 38.875 186.360 39.165 186.405 ;
        RECT 37.480 186.220 39.165 186.360 ;
        RECT 37.480 186.160 37.800 186.220 ;
        RECT 38.875 186.175 39.165 186.220 ;
        RECT 44.840 186.160 45.160 186.420 ;
        RECT 45.315 186.175 45.605 186.405 ;
        RECT 46.235 186.360 46.525 186.405 ;
        RECT 47.615 186.360 47.905 186.405 ;
        RECT 49.070 186.360 49.210 186.840 ;
        RECT 46.235 186.220 49.210 186.360 ;
        RECT 51.295 186.360 51.585 186.405 ;
        RECT 55.420 186.360 55.740 186.420 ;
        RECT 57.350 186.405 57.490 186.840 ;
        RECT 64.250 186.700 64.390 186.900 ;
        RECT 67.840 186.840 68.160 186.900 ;
        RECT 68.300 186.840 68.620 186.900 ;
        RECT 80.260 186.840 80.580 187.100 ;
        RECT 83.035 187.040 83.325 187.085 ;
        RECT 84.400 187.040 84.720 187.100 ;
        RECT 83.035 186.900 84.720 187.040 ;
        RECT 83.035 186.855 83.325 186.900 ;
        RECT 84.400 186.840 84.720 186.900 ;
        RECT 87.620 186.840 87.940 187.100 ;
        RECT 98.660 186.840 98.980 187.100 ;
        RECT 99.120 186.840 99.440 187.100 ;
        RECT 103.735 186.855 104.025 187.085 ;
        RECT 61.030 186.560 64.390 186.700 ;
        RECT 51.295 186.220 55.740 186.360 ;
        RECT 46.235 186.175 46.525 186.220 ;
        RECT 47.615 186.175 47.905 186.220 ;
        RECT 51.295 186.175 51.585 186.220 ;
        RECT 45.390 185.740 45.530 186.175 ;
        RECT 55.420 186.160 55.740 186.220 ;
        RECT 55.895 186.360 56.185 186.405 ;
        RECT 56.355 186.360 56.645 186.405 ;
        RECT 55.895 186.220 56.645 186.360 ;
        RECT 55.895 186.175 56.185 186.220 ;
        RECT 56.355 186.175 56.645 186.220 ;
        RECT 57.275 186.175 57.565 186.405 ;
        RECT 57.720 186.160 58.040 186.420 ;
        RECT 61.030 186.405 61.170 186.560 ;
        RECT 60.955 186.175 61.245 186.405 ;
        RECT 61.415 186.175 61.705 186.405 ;
        RECT 50.375 186.020 50.665 186.065 ;
        RECT 50.820 186.020 51.140 186.080 ;
        RECT 54.515 186.020 54.805 186.065 ;
        RECT 50.375 185.880 51.140 186.020 ;
        RECT 50.375 185.835 50.665 185.880 ;
        RECT 50.820 185.820 51.140 185.880 ;
        RECT 51.830 185.880 54.805 186.020 ;
        RECT 34.720 185.480 35.040 185.740 ;
        RECT 45.300 185.480 45.620 185.740 ;
        RECT 35.640 185.340 35.960 185.400 ;
        RECT 33.890 185.200 35.960 185.340 ;
        RECT 35.640 185.140 35.960 185.200 ;
        RECT 37.020 185.140 37.340 185.400 ;
        RECT 37.940 185.140 38.260 185.400 ;
        RECT 47.140 185.140 47.460 185.400 ;
        RECT 48.060 185.340 48.380 185.400 ;
        RECT 51.830 185.340 51.970 185.880 ;
        RECT 54.515 185.835 54.805 185.880 ;
        RECT 54.960 185.820 55.280 186.080 ;
        RECT 61.490 186.020 61.630 186.175 ;
        RECT 61.860 186.160 62.180 186.420 ;
        RECT 64.250 186.405 64.390 186.560 ;
        RECT 64.635 186.700 64.925 186.745 ;
        RECT 75.660 186.700 75.980 186.760 ;
        RECT 64.635 186.560 75.980 186.700 ;
        RECT 64.635 186.515 64.925 186.560 ;
        RECT 75.660 186.500 75.980 186.560 ;
        RECT 76.580 186.700 76.900 186.760 ;
        RECT 77.975 186.700 78.265 186.745 ;
        RECT 80.350 186.700 80.490 186.840 ;
        RECT 81.180 186.700 81.500 186.760 ;
        RECT 84.875 186.700 85.165 186.745 ;
        RECT 85.320 186.700 85.640 186.760 ;
        RECT 87.710 186.700 87.850 186.840 ;
        RECT 98.200 186.700 98.520 186.760 ;
        RECT 76.580 186.560 85.640 186.700 ;
        RECT 76.580 186.500 76.900 186.560 ;
        RECT 77.975 186.515 78.265 186.560 ;
        RECT 81.180 186.500 81.500 186.560 ;
        RECT 84.875 186.515 85.165 186.560 ;
        RECT 85.320 186.500 85.640 186.560 ;
        RECT 85.870 186.560 87.850 186.700 ;
        RECT 97.370 186.560 98.520 186.700 ;
        RECT 62.795 186.175 63.085 186.405 ;
        RECT 64.175 186.175 64.465 186.405 ;
        RECT 62.320 186.020 62.640 186.080 ;
        RECT 61.490 185.880 62.640 186.020 ;
        RECT 62.870 186.020 63.010 186.175 ;
        RECT 65.080 186.160 65.400 186.420 ;
        RECT 66.015 186.360 66.305 186.405 ;
        RECT 70.155 186.360 70.445 186.405 ;
        RECT 66.015 186.220 70.445 186.360 ;
        RECT 66.015 186.175 66.305 186.220 ;
        RECT 70.155 186.175 70.445 186.220 ;
        RECT 70.600 186.360 70.920 186.420 ;
        RECT 72.915 186.360 73.205 186.405 ;
        RECT 70.600 186.220 73.205 186.360 ;
        RECT 70.600 186.160 70.920 186.220 ;
        RECT 72.915 186.175 73.205 186.220 ;
        RECT 77.040 186.160 77.360 186.420 ;
        RECT 77.515 186.360 77.805 186.405 ;
        RECT 78.420 186.360 78.740 186.420 ;
        RECT 77.515 186.220 78.740 186.360 ;
        RECT 77.515 186.175 77.805 186.220 ;
        RECT 78.420 186.160 78.740 186.220 ;
        RECT 78.895 186.360 79.185 186.405 ;
        RECT 79.355 186.360 79.645 186.405 ;
        RECT 78.895 186.220 79.645 186.360 ;
        RECT 78.895 186.175 79.185 186.220 ;
        RECT 79.355 186.175 79.645 186.220 ;
        RECT 80.260 186.360 80.580 186.420 ;
        RECT 83.020 186.360 83.340 186.420 ;
        RECT 83.955 186.360 84.245 186.405 ;
        RECT 80.260 186.220 84.245 186.360 ;
        RECT 80.260 186.160 80.580 186.220 ;
        RECT 83.020 186.160 83.340 186.220 ;
        RECT 83.955 186.175 84.245 186.220 ;
        RECT 84.400 186.160 84.720 186.420 ;
        RECT 85.870 186.405 86.010 186.560 ;
        RECT 85.795 186.175 86.085 186.405 ;
        RECT 86.715 186.360 87.005 186.405 ;
        RECT 87.160 186.360 87.480 186.420 ;
        RECT 86.715 186.220 87.480 186.360 ;
        RECT 86.715 186.175 87.005 186.220 ;
        RECT 87.160 186.160 87.480 186.220 ;
        RECT 91.300 186.360 91.620 186.420 ;
        RECT 97.370 186.405 97.510 186.560 ;
        RECT 98.200 186.500 98.520 186.560 ;
        RECT 91.775 186.360 92.065 186.405 ;
        RECT 91.300 186.220 92.065 186.360 ;
        RECT 91.300 186.160 91.620 186.220 ;
        RECT 91.775 186.175 92.065 186.220 ;
        RECT 97.295 186.175 97.585 186.405 ;
        RECT 97.740 186.160 98.060 186.420 ;
        RECT 98.750 186.405 98.890 186.840 ;
        RECT 99.210 186.405 99.350 186.840 ;
        RECT 103.810 186.420 103.950 186.855 ;
        RECT 107.400 186.840 107.720 187.100 ;
        RECT 109.845 187.040 110.135 187.085 ;
        RECT 113.380 187.040 113.700 187.100 ;
        RECT 109.845 186.900 113.700 187.040 ;
        RECT 109.845 186.855 110.135 186.900 ;
        RECT 113.380 186.840 113.700 186.900 ;
        RECT 117.520 186.840 117.840 187.100 ;
        RECT 126.260 187.040 126.580 187.100 ;
        RECT 128.560 187.040 128.880 187.100 ;
        RECT 129.035 187.040 129.325 187.085 ;
        RECT 126.260 186.900 129.325 187.040 ;
        RECT 126.260 186.840 126.580 186.900 ;
        RECT 98.675 186.175 98.965 186.405 ;
        RECT 99.135 186.175 99.425 186.405 ;
        RECT 103.720 186.360 104.040 186.420 ;
        RECT 104.655 186.360 104.945 186.405 ;
        RECT 103.720 186.220 104.945 186.360 ;
        RECT 107.490 186.360 107.630 186.840 ;
        RECT 108.795 186.515 109.085 186.745 ;
        RECT 117.610 186.700 117.750 186.840 ;
        RECT 117.610 186.560 119.130 186.700 ;
        RECT 107.875 186.360 108.165 186.405 ;
        RECT 107.490 186.220 108.165 186.360 ;
        RECT 103.720 186.160 104.040 186.220 ;
        RECT 104.655 186.175 104.945 186.220 ;
        RECT 107.875 186.175 108.165 186.220 ;
        RECT 66.475 186.020 66.765 186.065 ;
        RECT 62.870 185.880 66.765 186.020 ;
        RECT 62.320 185.820 62.640 185.880 ;
        RECT 66.475 185.835 66.765 185.880 ;
        RECT 69.220 185.820 69.540 186.080 ;
        RECT 77.130 186.020 77.270 186.160 ;
        RECT 80.350 186.020 80.490 186.160 ;
        RECT 77.130 185.880 80.490 186.020 ;
        RECT 82.560 186.020 82.880 186.080 ;
        RECT 91.390 186.020 91.530 186.160 ;
        RECT 82.560 185.880 91.530 186.020 ;
        RECT 99.580 186.020 99.900 186.080 ;
        RECT 101.435 186.020 101.725 186.065 ;
        RECT 106.940 186.020 107.260 186.080 ;
        RECT 108.870 186.020 109.010 186.515 ;
        RECT 118.990 186.420 119.130 186.560 ;
        RECT 117.520 186.405 117.840 186.420 ;
        RECT 117.520 186.175 117.870 186.405 ;
        RECT 117.520 186.160 117.840 186.175 ;
        RECT 118.900 186.160 119.220 186.420 ;
        RECT 124.435 186.360 124.725 186.405 ;
        RECT 124.435 186.220 126.490 186.360 ;
        RECT 124.435 186.175 124.725 186.220 ;
        RECT 99.580 185.880 101.725 186.020 ;
        RECT 82.560 185.820 82.880 185.880 ;
        RECT 99.580 185.820 99.900 185.880 ;
        RECT 101.435 185.835 101.725 185.880 ;
        RECT 105.650 185.880 109.010 186.020 ;
        RECT 114.325 186.020 114.615 186.065 ;
        RECT 116.845 186.020 117.135 186.065 ;
        RECT 118.035 186.020 118.325 186.065 ;
        RECT 114.325 185.880 118.325 186.020 ;
        RECT 52.215 185.680 52.505 185.725 ;
        RECT 52.215 185.540 56.570 185.680 ;
        RECT 52.215 185.495 52.505 185.540 ;
        RECT 54.590 185.400 54.730 185.540 ;
        RECT 48.060 185.200 51.970 185.340 ;
        RECT 48.060 185.140 48.380 185.200 ;
        RECT 54.500 185.140 54.820 185.400 ;
        RECT 56.430 185.385 56.570 185.540 ;
        RECT 58.640 185.480 58.960 185.740 ;
        RECT 61.860 185.680 62.180 185.740 ;
        RECT 65.080 185.680 65.400 185.740 ;
        RECT 61.860 185.540 65.400 185.680 ;
        RECT 61.860 185.480 62.180 185.540 ;
        RECT 65.080 185.480 65.400 185.540 ;
        RECT 89.475 185.680 89.765 185.725 ;
        RECT 90.840 185.680 91.160 185.740 ;
        RECT 89.475 185.540 91.160 185.680 ;
        RECT 89.475 185.495 89.765 185.540 ;
        RECT 90.840 185.480 91.160 185.540 ;
        RECT 96.360 185.480 96.680 185.740 ;
        RECT 102.800 185.480 103.120 185.740 ;
        RECT 103.260 185.680 103.580 185.740 ;
        RECT 105.650 185.725 105.790 185.880 ;
        RECT 106.940 185.820 107.260 185.880 ;
        RECT 114.325 185.835 114.615 185.880 ;
        RECT 116.845 185.835 117.135 185.880 ;
        RECT 118.035 185.835 118.325 185.880 ;
        RECT 105.575 185.680 105.865 185.725 ;
        RECT 103.260 185.540 105.865 185.680 ;
        RECT 103.260 185.480 103.580 185.540 ;
        RECT 104.270 185.400 104.410 185.540 ;
        RECT 105.575 185.495 105.865 185.540 ;
        RECT 107.415 185.680 107.705 185.725 ;
        RECT 107.860 185.680 108.180 185.740 ;
        RECT 126.350 185.725 126.490 186.220 ;
        RECT 107.415 185.540 108.180 185.680 ;
        RECT 107.415 185.495 107.705 185.540 ;
        RECT 107.860 185.480 108.180 185.540 ;
        RECT 114.760 185.680 115.050 185.725 ;
        RECT 116.330 185.680 116.620 185.725 ;
        RECT 118.430 185.680 118.720 185.725 ;
        RECT 114.760 185.540 118.720 185.680 ;
        RECT 114.760 185.495 115.050 185.540 ;
        RECT 116.330 185.495 116.620 185.540 ;
        RECT 118.430 185.495 118.720 185.540 ;
        RECT 126.275 185.495 126.565 185.725 ;
        RECT 56.355 185.155 56.645 185.385 ;
        RECT 60.020 185.140 60.340 185.400 ;
        RECT 63.255 185.340 63.545 185.385 ;
        RECT 63.700 185.340 64.020 185.400 ;
        RECT 63.255 185.200 64.020 185.340 ;
        RECT 63.255 185.155 63.545 185.200 ;
        RECT 63.700 185.140 64.020 185.200 ;
        RECT 76.120 185.140 76.440 185.400 ;
        RECT 88.095 185.340 88.385 185.385 ;
        RECT 88.540 185.340 88.860 185.400 ;
        RECT 88.095 185.200 88.860 185.340 ;
        RECT 88.095 185.155 88.385 185.200 ;
        RECT 88.540 185.140 88.860 185.200 ;
        RECT 89.000 185.140 89.320 185.400 ;
        RECT 91.315 185.340 91.605 185.385 ;
        RECT 92.680 185.340 93.000 185.400 ;
        RECT 91.315 185.200 93.000 185.340 ;
        RECT 91.315 185.155 91.605 185.200 ;
        RECT 92.680 185.140 93.000 185.200 ;
        RECT 104.180 185.140 104.500 185.400 ;
        RECT 109.700 185.140 110.020 185.400 ;
        RECT 110.620 185.140 110.940 185.400 ;
        RECT 112.000 185.140 112.320 185.400 ;
        RECT 123.500 185.140 123.820 185.400 ;
        RECT 126.810 185.340 126.950 186.900 ;
        RECT 128.560 186.840 128.880 186.900 ;
        RECT 129.035 186.855 129.325 186.900 ;
        RECT 132.240 186.840 132.560 187.100 ;
        RECT 134.095 187.040 134.385 187.085 ;
        RECT 136.395 187.040 136.685 187.085 ;
        RECT 134.095 186.900 136.685 187.040 ;
        RECT 134.095 186.855 134.385 186.900 ;
        RECT 136.395 186.855 136.685 186.900 ;
        RECT 141.440 186.840 141.760 187.100 ;
        RECT 147.435 187.040 147.725 187.085 ;
        RECT 147.435 186.900 151.330 187.040 ;
        RECT 147.435 186.855 147.725 186.900 ;
        RECT 127.115 186.700 127.405 186.745 ;
        RECT 127.640 186.700 127.960 186.760 ;
        RECT 127.115 186.560 127.960 186.700 ;
        RECT 127.115 186.515 127.405 186.560 ;
        RECT 127.640 186.500 127.960 186.560 ;
        RECT 128.115 186.700 128.405 186.745 ;
        RECT 128.115 186.560 129.250 186.700 ;
        RECT 128.115 186.515 128.405 186.560 ;
        RECT 128.575 186.360 128.865 186.405 ;
        RECT 127.270 186.220 128.865 186.360 ;
        RECT 129.110 186.360 129.250 186.560 ;
        RECT 129.480 186.500 129.800 186.760 ;
        RECT 129.110 186.220 129.710 186.360 ;
        RECT 127.270 186.080 127.410 186.220 ;
        RECT 128.575 186.175 128.865 186.220 ;
        RECT 127.180 185.820 127.500 186.080 ;
        RECT 129.570 186.020 129.710 186.220 ;
        RECT 129.940 186.160 130.260 186.420 ;
        RECT 131.795 186.360 132.085 186.405 ;
        RECT 132.330 186.360 132.470 186.840 ;
        RECT 139.615 186.700 139.905 186.745 ;
        RECT 141.900 186.700 142.220 186.760 ;
        RECT 139.615 186.560 142.220 186.700 ;
        RECT 139.615 186.515 139.905 186.560 ;
        RECT 141.900 186.500 142.220 186.560 ;
        RECT 144.660 186.700 144.980 186.760 ;
        RECT 146.515 186.700 146.805 186.745 ;
        RECT 148.655 186.700 148.945 186.745 ;
        RECT 144.660 186.560 146.805 186.700 ;
        RECT 144.660 186.500 144.980 186.560 ;
        RECT 146.515 186.515 146.805 186.560 ;
        RECT 147.050 186.560 148.945 186.700 ;
        RECT 131.795 186.220 132.470 186.360 ;
        RECT 134.080 186.360 134.400 186.420 ;
        RECT 136.855 186.360 137.145 186.405 ;
        RECT 134.080 186.220 137.145 186.360 ;
        RECT 131.795 186.175 132.085 186.220 ;
        RECT 134.080 186.160 134.400 186.220 ;
        RECT 136.855 186.175 137.145 186.220 ;
        RECT 137.300 186.160 137.620 186.420 ;
        RECT 138.695 186.360 138.985 186.405 ;
        RECT 137.850 186.220 138.985 186.360 ;
        RECT 133.160 186.020 133.480 186.080 ;
        RECT 137.850 186.020 137.990 186.220 ;
        RECT 138.695 186.175 138.985 186.220 ;
        RECT 140.075 186.175 140.365 186.405 ;
        RECT 140.535 186.360 140.825 186.405 ;
        RECT 141.440 186.360 141.760 186.420 ;
        RECT 140.535 186.220 141.760 186.360 ;
        RECT 140.535 186.175 140.825 186.220 ;
        RECT 140.150 186.020 140.290 186.175 ;
        RECT 141.440 186.160 141.760 186.220 ;
        RECT 145.580 186.160 145.900 186.420 ;
        RECT 146.040 186.360 146.360 186.420 ;
        RECT 147.050 186.360 147.190 186.560 ;
        RECT 148.655 186.515 148.945 186.560 ;
        RECT 149.720 186.500 150.040 186.760 ;
        RECT 151.190 186.405 151.330 186.900 ;
        RECT 146.040 186.220 147.190 186.360 ;
        RECT 146.040 186.160 146.360 186.220 ;
        RECT 151.115 186.175 151.405 186.405 ;
        RECT 129.570 185.880 133.480 186.020 ;
        RECT 129.570 185.400 129.710 185.880 ;
        RECT 133.160 185.820 133.480 185.880 ;
        RECT 135.550 185.880 137.990 186.020 ;
        RECT 138.310 185.880 140.290 186.020 ;
        RECT 144.200 186.020 144.520 186.080 ;
        RECT 144.675 186.020 144.965 186.065 ;
        RECT 145.670 186.020 145.810 186.160 ;
        RECT 150.640 186.020 150.960 186.080 ;
        RECT 144.200 185.880 150.960 186.020 ;
        RECT 135.550 185.740 135.690 185.880 ;
        RECT 135.460 185.480 135.780 185.740 ;
        RECT 137.760 185.680 138.080 185.740 ;
        RECT 138.310 185.725 138.450 185.880 ;
        RECT 144.200 185.820 144.520 185.880 ;
        RECT 144.675 185.835 144.965 185.880 ;
        RECT 150.640 185.820 150.960 185.880 ;
        RECT 138.235 185.680 138.525 185.725 ;
        RECT 137.760 185.540 138.525 185.680 ;
        RECT 137.760 185.480 138.080 185.540 ;
        RECT 138.235 185.495 138.525 185.540 ;
        RECT 146.130 185.540 148.570 185.680 ;
        RECT 127.195 185.340 127.485 185.385 ;
        RECT 126.810 185.200 127.485 185.340 ;
        RECT 127.195 185.155 127.485 185.200 ;
        RECT 129.480 185.140 129.800 185.400 ;
        RECT 131.320 185.340 131.640 185.400 ;
        RECT 132.255 185.340 132.545 185.385 ;
        RECT 131.320 185.200 132.545 185.340 ;
        RECT 131.320 185.140 131.640 185.200 ;
        RECT 132.255 185.155 132.545 185.200 ;
        RECT 142.820 185.340 143.140 185.400 ;
        RECT 146.130 185.340 146.270 185.540 ;
        RECT 142.820 185.200 146.270 185.340 ;
        RECT 146.515 185.340 146.805 185.385 ;
        RECT 146.960 185.340 147.280 185.400 ;
        RECT 146.515 185.200 147.280 185.340 ;
        RECT 142.820 185.140 143.140 185.200 ;
        RECT 146.515 185.155 146.805 185.200 ;
        RECT 146.960 185.140 147.280 185.200 ;
        RECT 147.420 185.340 147.740 185.400 ;
        RECT 147.895 185.340 148.185 185.385 ;
        RECT 147.420 185.200 148.185 185.340 ;
        RECT 148.430 185.340 148.570 185.540 ;
        RECT 148.815 185.340 149.105 185.385 ;
        RECT 148.430 185.200 149.105 185.340 ;
        RECT 147.420 185.140 147.740 185.200 ;
        RECT 147.895 185.155 148.185 185.200 ;
        RECT 148.815 185.155 149.105 185.200 ;
        RECT 150.180 185.140 150.500 185.400 ;
        RECT 22.690 184.520 157.010 185.000 ;
        RECT 25.980 184.320 26.300 184.380 ;
        RECT 26.915 184.320 27.205 184.365 ;
        RECT 25.980 184.180 27.205 184.320 ;
        RECT 25.980 184.120 26.300 184.180 ;
        RECT 26.915 184.135 27.205 184.180 ;
        RECT 31.960 184.120 32.280 184.380 ;
        RECT 34.275 184.320 34.565 184.365 ;
        RECT 42.540 184.320 42.860 184.380 ;
        RECT 32.510 184.180 42.860 184.320 ;
        RECT 32.050 183.640 32.190 184.120 ;
        RECT 27.910 183.500 32.190 183.640 ;
        RECT 27.910 183.345 28.050 183.500 ;
        RECT 27.835 183.115 28.125 183.345 ;
        RECT 31.500 183.100 31.820 183.360 ;
        RECT 31.960 183.100 32.280 183.360 ;
        RECT 31.590 182.960 31.730 183.100 ;
        RECT 32.510 182.960 32.650 184.180 ;
        RECT 34.275 184.135 34.565 184.180 ;
        RECT 42.540 184.120 42.860 184.180 ;
        RECT 55.420 184.320 55.740 184.380 ;
        RECT 56.355 184.320 56.645 184.365 ;
        RECT 59.575 184.320 59.865 184.365 ;
        RECT 69.220 184.320 69.540 184.380 ;
        RECT 55.420 184.180 59.865 184.320 ;
        RECT 55.420 184.120 55.740 184.180 ;
        RECT 56.355 184.135 56.645 184.180 ;
        RECT 59.575 184.135 59.865 184.180 ;
        RECT 62.870 184.180 69.540 184.320 ;
        RECT 32.895 183.980 33.185 184.025 ;
        RECT 34.720 183.980 35.040 184.040 ;
        RECT 32.895 183.840 35.040 183.980 ;
        RECT 32.895 183.795 33.185 183.840 ;
        RECT 34.720 183.780 35.040 183.840 ;
        RECT 36.600 183.980 36.890 184.025 ;
        RECT 38.700 183.980 38.990 184.025 ;
        RECT 40.270 183.980 40.560 184.025 ;
        RECT 36.600 183.840 40.560 183.980 ;
        RECT 36.600 183.795 36.890 183.840 ;
        RECT 38.700 183.795 38.990 183.840 ;
        RECT 40.270 183.795 40.560 183.840 ;
        RECT 45.340 183.980 45.630 184.025 ;
        RECT 47.440 183.980 47.730 184.025 ;
        RECT 49.010 183.980 49.300 184.025 ;
        RECT 45.340 183.840 49.300 183.980 ;
        RECT 45.340 183.795 45.630 183.840 ;
        RECT 47.440 183.795 47.730 183.840 ;
        RECT 49.010 183.795 49.300 183.840 ;
        RECT 54.960 183.980 55.280 184.040 ;
        RECT 62.335 183.980 62.625 184.025 ;
        RECT 54.960 183.840 62.625 183.980 ;
        RECT 54.960 183.780 55.280 183.840 ;
        RECT 36.995 183.640 37.285 183.685 ;
        RECT 38.185 183.640 38.475 183.685 ;
        RECT 40.705 183.640 40.995 183.685 ;
        RECT 36.995 183.500 40.995 183.640 ;
        RECT 36.995 183.455 37.285 183.500 ;
        RECT 38.185 183.455 38.475 183.500 ;
        RECT 40.705 183.455 40.995 183.500 ;
        RECT 45.735 183.640 46.025 183.685 ;
        RECT 46.925 183.640 47.215 183.685 ;
        RECT 49.445 183.640 49.735 183.685 ;
        RECT 45.735 183.500 49.735 183.640 ;
        RECT 45.735 183.455 46.025 183.500 ;
        RECT 46.925 183.455 47.215 183.500 ;
        RECT 49.445 183.455 49.735 183.500 ;
        RECT 51.370 183.500 57.490 183.640 ;
        RECT 35.640 183.300 35.960 183.360 ;
        RECT 36.115 183.300 36.405 183.345 ;
        RECT 44.855 183.300 45.145 183.345 ;
        RECT 51.370 183.300 51.510 183.500 ;
        RECT 57.350 183.345 57.490 183.500 ;
        RECT 57.810 183.345 57.950 183.840 ;
        RECT 62.335 183.795 62.625 183.840 ;
        RECT 58.180 183.640 58.500 183.700 ;
        RECT 58.655 183.640 58.945 183.685 ;
        RECT 58.180 183.500 58.945 183.640 ;
        RECT 58.180 183.440 58.500 183.500 ;
        RECT 58.655 183.455 58.945 183.500 ;
        RECT 62.870 183.345 63.010 184.180 ;
        RECT 69.220 184.120 69.540 184.180 ;
        RECT 77.515 184.320 77.805 184.365 ;
        RECT 82.560 184.320 82.880 184.380 ;
        RECT 77.515 184.180 82.880 184.320 ;
        RECT 77.515 184.135 77.805 184.180 ;
        RECT 82.560 184.120 82.880 184.180 ;
        RECT 94.535 184.320 94.825 184.365 ;
        RECT 97.740 184.320 98.060 184.380 ;
        RECT 94.535 184.180 98.060 184.320 ;
        RECT 94.535 184.135 94.825 184.180 ;
        RECT 97.740 184.120 98.060 184.180 ;
        RECT 109.700 184.320 110.020 184.380 ;
        RECT 111.095 184.320 111.385 184.365 ;
        RECT 109.700 184.180 111.385 184.320 ;
        RECT 109.700 184.120 110.020 184.180 ;
        RECT 111.095 184.135 111.385 184.180 ;
        RECT 112.015 184.320 112.305 184.365 ;
        RECT 112.460 184.320 112.780 184.380 ;
        RECT 112.015 184.180 112.780 184.320 ;
        RECT 112.015 184.135 112.305 184.180 ;
        RECT 63.740 183.980 64.030 184.025 ;
        RECT 65.840 183.980 66.130 184.025 ;
        RECT 67.410 183.980 67.700 184.025 ;
        RECT 63.740 183.840 67.700 183.980 ;
        RECT 63.740 183.795 64.030 183.840 ;
        RECT 65.840 183.795 66.130 183.840 ;
        RECT 67.410 183.795 67.700 183.840 ;
        RECT 71.100 183.980 71.390 184.025 ;
        RECT 73.200 183.980 73.490 184.025 ;
        RECT 74.770 183.980 75.060 184.025 ;
        RECT 71.100 183.840 75.060 183.980 ;
        RECT 71.100 183.795 71.390 183.840 ;
        RECT 73.200 183.795 73.490 183.840 ;
        RECT 74.770 183.795 75.060 183.840 ;
        RECT 78.460 183.980 78.750 184.025 ;
        RECT 80.560 183.980 80.850 184.025 ;
        RECT 82.130 183.980 82.420 184.025 ;
        RECT 78.460 183.840 82.420 183.980 ;
        RECT 78.460 183.795 78.750 183.840 ;
        RECT 80.560 183.795 80.850 183.840 ;
        RECT 82.130 183.795 82.420 183.840 ;
        RECT 84.875 183.980 85.165 184.025 ;
        RECT 85.780 183.980 86.100 184.040 ;
        RECT 88.540 183.980 88.860 184.040 ;
        RECT 84.875 183.840 88.860 183.980 ;
        RECT 84.875 183.795 85.165 183.840 ;
        RECT 85.780 183.780 86.100 183.840 ;
        RECT 88.540 183.780 88.860 183.840 ;
        RECT 98.660 183.980 98.950 184.025 ;
        RECT 100.230 183.980 100.520 184.025 ;
        RECT 102.330 183.980 102.620 184.025 ;
        RECT 112.090 183.980 112.230 184.135 ;
        RECT 112.460 184.120 112.780 184.180 ;
        RECT 114.315 184.320 114.605 184.365 ;
        RECT 117.520 184.320 117.840 184.380 ;
        RECT 114.315 184.180 117.840 184.320 ;
        RECT 114.315 184.135 114.605 184.180 ;
        RECT 117.520 184.120 117.840 184.180 ;
        RECT 127.640 184.320 127.960 184.380 ;
        RECT 128.575 184.320 128.865 184.365 ;
        RECT 127.640 184.180 128.865 184.320 ;
        RECT 127.640 184.120 127.960 184.180 ;
        RECT 128.575 184.135 128.865 184.180 ;
        RECT 131.320 184.120 131.640 184.380 ;
        RECT 132.240 184.120 132.560 184.380 ;
        RECT 134.080 184.120 134.400 184.380 ;
        RECT 134.540 184.320 134.860 184.380 ;
        RECT 135.475 184.320 135.765 184.365 ;
        RECT 134.540 184.180 135.765 184.320 ;
        RECT 134.540 184.120 134.860 184.180 ;
        RECT 135.475 184.135 135.765 184.180 ;
        RECT 137.315 184.320 137.605 184.365 ;
        RECT 137.760 184.320 138.080 184.380 ;
        RECT 137.315 184.180 138.080 184.320 ;
        RECT 137.315 184.135 137.605 184.180 ;
        RECT 137.760 184.120 138.080 184.180 ;
        RECT 139.615 184.320 139.905 184.365 ;
        RECT 141.440 184.320 141.760 184.380 ;
        RECT 139.615 184.180 141.760 184.320 ;
        RECT 139.615 184.135 139.905 184.180 ;
        RECT 141.440 184.120 141.760 184.180 ;
        RECT 142.835 184.320 143.125 184.365 ;
        RECT 144.660 184.320 144.980 184.380 ;
        RECT 146.960 184.320 147.280 184.380 ;
        RECT 142.835 184.180 144.980 184.320 ;
        RECT 142.835 184.135 143.125 184.180 ;
        RECT 144.660 184.120 144.980 184.180 ;
        RECT 145.210 184.180 147.280 184.320 ;
        RECT 98.660 183.840 102.620 183.980 ;
        RECT 98.660 183.795 98.950 183.840 ;
        RECT 100.230 183.795 100.520 183.840 ;
        RECT 102.330 183.795 102.620 183.840 ;
        RECT 110.250 183.840 112.230 183.980 ;
        RECT 121.700 183.980 121.990 184.025 ;
        RECT 123.800 183.980 124.090 184.025 ;
        RECT 125.370 183.980 125.660 184.025 ;
        RECT 121.700 183.840 125.660 183.980 ;
        RECT 64.135 183.640 64.425 183.685 ;
        RECT 65.325 183.640 65.615 183.685 ;
        RECT 67.845 183.640 68.135 183.685 ;
        RECT 64.135 183.500 68.135 183.640 ;
        RECT 64.135 183.455 64.425 183.500 ;
        RECT 65.325 183.455 65.615 183.500 ;
        RECT 67.845 183.455 68.135 183.500 ;
        RECT 71.495 183.640 71.785 183.685 ;
        RECT 72.685 183.640 72.975 183.685 ;
        RECT 75.205 183.640 75.495 183.685 ;
        RECT 71.495 183.500 75.495 183.640 ;
        RECT 71.495 183.455 71.785 183.500 ;
        RECT 72.685 183.455 72.975 183.500 ;
        RECT 75.205 183.455 75.495 183.500 ;
        RECT 78.855 183.640 79.145 183.685 ;
        RECT 80.045 183.640 80.335 183.685 ;
        RECT 82.565 183.640 82.855 183.685 ;
        RECT 78.855 183.500 82.855 183.640 ;
        RECT 78.855 183.455 79.145 183.500 ;
        RECT 80.045 183.455 80.335 183.500 ;
        RECT 82.565 183.455 82.855 183.500 ;
        RECT 86.255 183.640 86.545 183.685 ;
        RECT 98.225 183.640 98.515 183.685 ;
        RECT 100.745 183.640 101.035 183.685 ;
        RECT 101.935 183.640 102.225 183.685 ;
        RECT 86.255 183.500 93.830 183.640 ;
        RECT 86.255 183.455 86.545 183.500 ;
        RECT 54.975 183.300 55.265 183.345 ;
        RECT 55.895 183.300 56.185 183.345 ;
        RECT 35.640 183.160 45.145 183.300 ;
        RECT 35.640 183.100 35.960 183.160 ;
        RECT 36.115 183.115 36.405 183.160 ;
        RECT 44.855 183.115 45.145 183.160 ;
        RECT 48.150 183.160 51.510 183.300 ;
        RECT 51.830 183.160 56.185 183.300 ;
        RECT 31.590 182.820 32.650 182.960 ;
        RECT 33.355 182.960 33.645 183.005 ;
        RECT 36.560 182.960 36.880 183.020 ;
        RECT 33.355 182.820 36.880 182.960 ;
        RECT 33.355 182.775 33.645 182.820 ;
        RECT 36.560 182.760 36.880 182.820 ;
        RECT 37.450 182.960 37.740 183.005 ;
        RECT 37.940 182.960 38.260 183.020 ;
        RECT 46.220 183.005 46.540 183.020 ;
        RECT 37.450 182.820 38.260 182.960 ;
        RECT 37.450 182.775 37.740 182.820 ;
        RECT 37.940 182.760 38.260 182.820 ;
        RECT 46.190 182.775 46.540 183.005 ;
        RECT 46.220 182.760 46.540 182.775 ;
        RECT 32.420 182.620 32.740 182.680 ;
        RECT 34.260 182.665 34.580 182.680 ;
        RECT 34.260 182.620 34.645 182.665 ;
        RECT 32.420 182.480 35.015 182.620 ;
        RECT 32.420 182.420 32.740 182.480 ;
        RECT 34.260 182.435 34.645 182.480 ;
        RECT 34.260 182.420 34.580 182.435 ;
        RECT 35.180 182.420 35.500 182.680 ;
        RECT 36.650 182.620 36.790 182.760 ;
        RECT 48.150 182.680 48.290 183.160 ;
        RECT 43.015 182.620 43.305 182.665 ;
        RECT 48.060 182.620 48.380 182.680 ;
        RECT 36.650 182.480 48.380 182.620 ;
        RECT 43.015 182.435 43.305 182.480 ;
        RECT 48.060 182.420 48.380 182.480 ;
        RECT 48.520 182.620 48.840 182.680 ;
        RECT 50.820 182.620 51.140 182.680 ;
        RECT 51.830 182.665 51.970 183.160 ;
        RECT 54.975 183.115 55.265 183.160 ;
        RECT 55.895 183.115 56.185 183.160 ;
        RECT 57.275 183.115 57.565 183.345 ;
        RECT 57.735 183.115 58.025 183.345 ;
        RECT 60.035 183.115 60.325 183.345 ;
        RECT 62.795 183.115 63.085 183.345 ;
        RECT 63.255 183.300 63.545 183.345 ;
        RECT 70.615 183.300 70.905 183.345 ;
        RECT 74.740 183.300 75.060 183.360 ;
        RECT 77.975 183.300 78.265 183.345 ;
        RECT 63.255 183.160 78.265 183.300 ;
        RECT 63.255 183.115 63.545 183.160 ;
        RECT 70.615 183.115 70.905 183.160 ;
        RECT 60.110 182.960 60.250 183.115 ;
        RECT 74.740 183.100 75.060 183.160 ;
        RECT 77.975 183.115 78.265 183.160 ;
        RECT 85.795 183.115 86.085 183.345 ;
        RECT 86.715 183.300 87.005 183.345 ;
        RECT 88.080 183.300 88.400 183.360 ;
        RECT 86.715 183.160 88.400 183.300 ;
        RECT 86.715 183.115 87.005 183.160 ;
        RECT 63.700 182.960 64.020 183.020 ;
        RECT 64.480 182.960 64.770 183.005 ;
        RECT 60.110 182.820 63.470 182.960 ;
        RECT 51.755 182.620 52.045 182.665 ;
        RECT 48.520 182.480 52.045 182.620 ;
        RECT 48.520 182.420 48.840 182.480 ;
        RECT 50.820 182.420 51.140 182.480 ;
        RECT 51.755 182.435 52.045 182.480 ;
        RECT 52.200 182.420 52.520 182.680 ;
        RECT 63.330 182.620 63.470 182.820 ;
        RECT 63.700 182.820 64.770 182.960 ;
        RECT 63.700 182.760 64.020 182.820 ;
        RECT 64.480 182.775 64.770 182.820 ;
        RECT 71.950 182.960 72.240 183.005 ;
        RECT 76.120 182.960 76.440 183.020 ;
        RECT 79.340 183.005 79.660 183.020 ;
        RECT 71.950 182.820 76.440 182.960 ;
        RECT 71.950 182.775 72.240 182.820 ;
        RECT 76.120 182.760 76.440 182.820 ;
        RECT 79.310 182.775 79.660 183.005 ;
        RECT 85.870 182.960 86.010 183.115 ;
        RECT 88.080 183.100 88.400 183.160 ;
        RECT 88.540 183.300 88.860 183.360 ;
        RECT 90.395 183.300 90.685 183.345 ;
        RECT 88.540 183.160 90.685 183.300 ;
        RECT 88.540 183.100 88.860 183.160 ;
        RECT 90.395 183.115 90.685 183.160 ;
        RECT 90.840 183.100 91.160 183.360 ;
        RECT 91.760 183.100 92.080 183.360 ;
        RECT 93.690 183.345 93.830 183.500 ;
        RECT 98.225 183.500 102.225 183.640 ;
        RECT 98.225 183.455 98.515 183.500 ;
        RECT 100.745 183.455 101.035 183.500 ;
        RECT 101.935 183.455 102.225 183.500 ;
        RECT 102.815 183.640 103.105 183.685 ;
        RECT 105.100 183.640 105.420 183.700 ;
        RECT 102.815 183.500 105.420 183.640 ;
        RECT 102.815 183.455 103.105 183.500 ;
        RECT 105.100 183.440 105.420 183.500 ;
        RECT 93.155 183.300 93.445 183.345 ;
        RECT 92.310 183.160 93.445 183.300 ;
        RECT 90.930 182.960 91.070 183.100 ;
        RECT 85.870 182.820 91.070 182.960 ;
        RECT 79.340 182.760 79.660 182.775 ;
        RECT 70.155 182.620 70.445 182.665 ;
        RECT 70.600 182.620 70.920 182.680 ;
        RECT 63.330 182.480 70.920 182.620 ;
        RECT 70.155 182.435 70.445 182.480 ;
        RECT 70.600 182.420 70.920 182.480 ;
        RECT 87.620 182.420 87.940 182.680 ;
        RECT 89.000 182.620 89.320 182.680 ;
        RECT 92.310 182.620 92.450 183.160 ;
        RECT 93.155 183.115 93.445 183.160 ;
        RECT 93.615 183.115 93.905 183.345 ;
        RECT 109.240 183.100 109.560 183.360 ;
        RECT 110.250 183.345 110.390 183.840 ;
        RECT 121.700 183.795 121.990 183.840 ;
        RECT 123.800 183.795 124.090 183.840 ;
        RECT 125.370 183.795 125.660 183.840 ;
        RECT 112.000 183.640 112.320 183.700 ;
        RECT 118.900 183.640 119.220 183.700 ;
        RECT 121.215 183.640 121.505 183.685 ;
        RECT 112.000 183.500 112.690 183.640 ;
        RECT 112.000 183.440 112.320 183.500 ;
        RECT 110.175 183.115 110.465 183.345 ;
        RECT 110.620 183.100 110.940 183.360 ;
        RECT 112.550 183.345 112.690 183.500 ;
        RECT 118.900 183.500 121.505 183.640 ;
        RECT 118.900 183.440 119.220 183.500 ;
        RECT 121.215 183.455 121.505 183.500 ;
        RECT 122.095 183.640 122.385 183.685 ;
        RECT 123.285 183.640 123.575 183.685 ;
        RECT 125.805 183.640 126.095 183.685 ;
        RECT 131.410 183.640 131.550 184.120 ;
        RECT 134.170 183.640 134.310 184.120 ;
        RECT 142.360 183.980 142.680 184.040 ;
        RECT 143.740 183.980 144.060 184.040 ;
        RECT 145.210 183.980 145.350 184.180 ;
        RECT 146.960 184.120 147.280 184.180 ;
        RECT 148.355 184.320 148.645 184.365 ;
        RECT 149.720 184.320 150.040 184.380 ;
        RECT 148.355 184.180 150.040 184.320 ;
        RECT 148.355 184.135 148.645 184.180 ;
        RECT 149.720 184.120 150.040 184.180 ;
        RECT 142.360 183.840 144.060 183.980 ;
        RECT 142.360 183.780 142.680 183.840 ;
        RECT 143.740 183.780 144.060 183.840 ;
        RECT 144.750 183.840 145.350 183.980 ;
        RECT 151.100 183.980 151.390 184.025 ;
        RECT 152.670 183.980 152.960 184.025 ;
        RECT 154.770 183.980 155.060 184.025 ;
        RECT 151.100 183.840 155.060 183.980 ;
        RECT 137.300 183.640 137.620 183.700 ;
        RECT 144.750 183.640 144.890 183.840 ;
        RECT 151.100 183.795 151.390 183.840 ;
        RECT 152.670 183.795 152.960 183.840 ;
        RECT 154.770 183.795 155.060 183.840 ;
        RECT 122.095 183.500 126.095 183.640 ;
        RECT 122.095 183.455 122.385 183.500 ;
        RECT 123.285 183.455 123.575 183.500 ;
        RECT 125.805 183.455 126.095 183.500 ;
        RECT 129.110 183.500 130.630 183.640 ;
        RECT 131.410 183.500 132.010 183.640 ;
        RECT 134.170 183.500 137.070 183.640 ;
        RECT 129.110 183.360 129.250 183.500 ;
        RECT 112.475 183.115 112.765 183.345 ;
        RECT 113.395 183.115 113.685 183.345 ;
        RECT 92.695 182.960 92.985 183.005 ;
        RECT 99.120 182.960 99.440 183.020 ;
        RECT 92.695 182.820 99.440 182.960 ;
        RECT 92.695 182.775 92.985 182.820 ;
        RECT 99.120 182.760 99.440 182.820 ;
        RECT 101.420 183.005 101.740 183.020 ;
        RECT 101.420 182.775 101.770 183.005 ;
        RECT 110.710 182.960 110.850 183.100 ;
        RECT 113.470 182.960 113.610 183.115 ;
        RECT 129.020 183.100 129.340 183.360 ;
        RECT 129.495 183.300 129.785 183.345 ;
        RECT 129.940 183.300 130.260 183.360 ;
        RECT 130.490 183.345 130.630 183.500 ;
        RECT 129.495 183.160 130.260 183.300 ;
        RECT 129.495 183.115 129.785 183.160 ;
        RECT 110.710 182.820 113.610 182.960 ;
        RECT 122.550 182.960 122.840 183.005 ;
        RECT 123.500 182.960 123.820 183.020 ;
        RECT 129.570 182.960 129.710 183.115 ;
        RECT 129.940 183.100 130.260 183.160 ;
        RECT 130.415 183.115 130.705 183.345 ;
        RECT 130.875 183.300 131.165 183.345 ;
        RECT 131.320 183.300 131.640 183.360 ;
        RECT 131.870 183.345 132.010 183.500 ;
        RECT 130.875 183.160 131.640 183.300 ;
        RECT 130.875 183.115 131.165 183.160 ;
        RECT 131.320 183.100 131.640 183.160 ;
        RECT 131.795 183.115 132.085 183.345 ;
        RECT 135.000 183.100 135.320 183.360 ;
        RECT 136.930 183.300 137.070 183.500 ;
        RECT 137.300 183.500 140.290 183.640 ;
        RECT 137.300 183.440 137.620 183.500 ;
        RECT 140.150 183.345 140.290 183.500 ;
        RECT 142.450 183.500 144.890 183.640 ;
        RECT 145.135 183.640 145.425 183.685 ;
        RECT 150.665 183.640 150.955 183.685 ;
        RECT 153.185 183.640 153.475 183.685 ;
        RECT 154.375 183.640 154.665 183.685 ;
        RECT 145.135 183.500 147.190 183.640 ;
        RECT 142.450 183.345 142.590 183.500 ;
        RECT 145.135 183.455 145.425 183.500 ;
        RECT 147.050 183.360 147.190 183.500 ;
        RECT 150.665 183.500 154.665 183.640 ;
        RECT 150.665 183.455 150.955 183.500 ;
        RECT 153.185 183.455 153.475 183.500 ;
        RECT 154.375 183.455 154.665 183.500 ;
        RECT 139.155 183.300 139.445 183.345 ;
        RECT 136.930 183.160 139.445 183.300 ;
        RECT 139.155 183.115 139.445 183.160 ;
        RECT 140.075 183.115 140.365 183.345 ;
        RECT 142.375 183.115 142.665 183.345 ;
        RECT 142.820 183.300 143.140 183.360 ;
        RECT 143.755 183.300 144.045 183.345 ;
        RECT 142.820 183.160 144.045 183.300 ;
        RECT 122.550 182.820 123.820 182.960 ;
        RECT 122.550 182.775 122.840 182.820 ;
        RECT 101.420 182.760 101.740 182.775 ;
        RECT 123.500 182.760 123.820 182.820 ;
        RECT 128.190 182.820 129.710 182.960 ;
        RECT 128.190 182.680 128.330 182.820 ;
        RECT 142.450 182.680 142.590 183.115 ;
        RECT 142.820 183.100 143.140 183.160 ;
        RECT 143.755 183.115 144.045 183.160 ;
        RECT 144.675 183.300 144.965 183.345 ;
        RECT 146.040 183.300 146.360 183.360 ;
        RECT 144.675 183.160 146.360 183.300 ;
        RECT 144.675 183.115 144.965 183.160 ;
        RECT 146.040 183.100 146.360 183.160 ;
        RECT 146.960 183.100 147.280 183.360 ;
        RECT 151.100 183.300 151.420 183.360 ;
        RECT 155.255 183.300 155.545 183.345 ;
        RECT 151.100 183.160 155.545 183.300 ;
        RECT 151.100 183.100 151.420 183.160 ;
        RECT 155.255 183.115 155.545 183.160 ;
        RECT 153.860 183.005 154.180 183.020 ;
        RECT 153.860 182.775 154.210 183.005 ;
        RECT 153.860 182.760 154.180 182.775 ;
        RECT 89.000 182.480 92.450 182.620 ;
        RECT 89.000 182.420 89.320 182.480 ;
        RECT 95.900 182.420 96.220 182.680 ;
        RECT 128.100 182.420 128.420 182.680 ;
        RECT 141.440 182.420 141.760 182.680 ;
        RECT 142.360 182.420 142.680 182.680 ;
        RECT 146.975 182.620 147.265 182.665 ;
        RECT 147.420 182.620 147.740 182.680 ;
        RECT 146.975 182.480 147.740 182.620 ;
        RECT 146.975 182.435 147.265 182.480 ;
        RECT 147.420 182.420 147.740 182.480 ;
        RECT 147.880 182.420 148.200 182.680 ;
        RECT 22.690 181.800 157.810 182.280 ;
        RECT 35.180 181.400 35.500 181.660 ;
        RECT 37.020 181.400 37.340 181.660 ;
        RECT 37.480 181.600 37.800 181.660 ;
        RECT 38.875 181.600 39.165 181.645 ;
        RECT 37.480 181.460 39.165 181.600 ;
        RECT 37.480 181.400 37.800 181.460 ;
        RECT 38.875 181.415 39.165 181.460 ;
        RECT 45.775 181.600 46.065 181.645 ;
        RECT 46.220 181.600 46.540 181.660 ;
        RECT 45.775 181.460 46.540 181.600 ;
        RECT 45.775 181.415 46.065 181.460 ;
        RECT 46.220 181.400 46.540 181.460 ;
        RECT 47.140 181.400 47.460 181.660 ;
        RECT 52.200 181.400 52.520 181.660 ;
        RECT 66.475 181.600 66.765 181.645 ;
        RECT 69.220 181.600 69.540 181.660 ;
        RECT 66.475 181.460 69.540 181.600 ;
        RECT 66.475 181.415 66.765 181.460 ;
        RECT 69.220 181.400 69.540 181.460 ;
        RECT 78.895 181.600 79.185 181.645 ;
        RECT 79.340 181.600 79.660 181.660 ;
        RECT 87.620 181.600 87.940 181.660 ;
        RECT 78.895 181.460 79.660 181.600 ;
        RECT 78.895 181.415 79.185 181.460 ;
        RECT 79.340 181.400 79.660 181.460 ;
        RECT 81.730 181.460 87.940 181.600 ;
        RECT 25.980 180.720 26.300 180.980 ;
        RECT 31.040 180.720 31.360 180.980 ;
        RECT 31.960 180.720 32.280 180.980 ;
        RECT 35.270 180.920 35.410 181.400 ;
        RECT 37.110 181.260 37.250 181.400 ;
        RECT 37.955 181.260 38.245 181.305 ;
        RECT 47.230 181.260 47.370 181.400 ;
        RECT 37.110 181.120 38.245 181.260 ;
        RECT 37.955 181.075 38.245 181.120 ;
        RECT 43.550 181.120 47.370 181.260 ;
        RECT 36.115 180.920 36.405 180.965 ;
        RECT 35.270 180.780 36.405 180.920 ;
        RECT 36.115 180.735 36.405 180.780 ;
        RECT 42.080 180.920 42.400 180.980 ;
        RECT 43.550 180.965 43.690 181.120 ;
        RECT 42.555 180.920 42.845 180.965 ;
        RECT 42.080 180.780 42.845 180.920 ;
        RECT 36.190 180.580 36.330 180.735 ;
        RECT 42.080 180.720 42.400 180.780 ;
        RECT 42.555 180.735 42.845 180.780 ;
        RECT 43.475 180.735 43.765 180.965 ;
        RECT 43.935 180.735 44.225 180.965 ;
        RECT 44.395 180.920 44.685 180.965 ;
        RECT 52.290 180.920 52.430 181.400 ;
        RECT 60.020 181.260 60.340 181.320 ;
        RECT 60.800 181.260 61.090 181.305 ;
        RECT 60.020 181.120 61.090 181.260 ;
        RECT 60.020 181.060 60.340 181.120 ;
        RECT 60.800 181.075 61.090 181.120 ;
        RECT 69.680 181.260 70.000 181.320 ;
        RECT 80.275 181.260 80.565 181.305 ;
        RECT 69.680 181.120 80.565 181.260 ;
        RECT 69.680 181.060 70.000 181.120 ;
        RECT 80.275 181.075 80.565 181.120 ;
        RECT 44.395 180.780 52.430 180.920 ;
        RECT 54.975 180.920 55.265 180.965 ;
        RECT 54.975 180.780 65.310 180.920 ;
        RECT 44.395 180.735 44.685 180.780 ;
        RECT 54.975 180.735 55.265 180.780 ;
        RECT 44.010 180.580 44.150 180.735 ;
        RECT 65.170 180.640 65.310 180.780 ;
        RECT 79.815 180.735 80.105 180.965 ;
        RECT 80.735 180.920 81.025 180.965 ;
        RECT 81.180 180.920 81.500 180.980 ;
        RECT 81.730 180.965 81.870 181.460 ;
        RECT 87.620 181.400 87.940 181.460 ;
        RECT 88.080 181.600 88.400 181.660 ;
        RECT 89.475 181.600 89.765 181.645 ;
        RECT 88.080 181.460 89.765 181.600 ;
        RECT 88.080 181.400 88.400 181.460 ;
        RECT 89.475 181.415 89.765 181.460 ;
        RECT 89.935 181.600 90.225 181.645 ;
        RECT 90.840 181.600 91.160 181.660 ;
        RECT 89.935 181.460 91.160 181.600 ;
        RECT 89.935 181.415 90.225 181.460 ;
        RECT 90.840 181.400 91.160 181.460 ;
        RECT 94.060 181.600 94.380 181.660 ;
        RECT 104.180 181.600 104.500 181.660 ;
        RECT 94.060 181.460 104.500 181.600 ;
        RECT 94.060 181.400 94.380 181.460 ;
        RECT 104.180 181.400 104.500 181.460 ;
        RECT 109.700 181.400 110.020 181.660 ;
        RECT 118.440 181.400 118.760 181.660 ;
        RECT 120.280 181.600 120.600 181.660 ;
        RECT 122.580 181.600 122.900 181.660 ;
        RECT 141.455 181.600 141.745 181.645 ;
        RECT 142.360 181.600 142.680 181.660 ;
        RECT 120.280 181.460 124.190 181.600 ;
        RECT 120.280 181.400 120.600 181.460 ;
        RECT 122.580 181.400 122.900 181.460 ;
        RECT 88.540 181.060 88.860 181.320 ;
        RECT 94.520 181.060 94.840 181.320 ;
        RECT 96.835 181.075 97.125 181.305 ;
        RECT 97.280 181.260 97.600 181.320 ;
        RECT 97.835 181.260 98.125 181.305 ;
        RECT 97.280 181.120 98.125 181.260 ;
        RECT 104.270 181.260 104.410 181.400 ;
        RECT 104.270 181.120 109.470 181.260 ;
        RECT 80.735 180.780 81.500 180.920 ;
        RECT 80.735 180.735 81.025 180.780 ;
        RECT 36.190 180.440 44.150 180.580 ;
        RECT 54.040 180.580 54.360 180.640 ;
        RECT 59.575 180.580 59.865 180.625 ;
        RECT 54.040 180.440 59.865 180.580 ;
        RECT 54.040 180.380 54.360 180.440 ;
        RECT 59.575 180.395 59.865 180.440 ;
        RECT 60.455 180.580 60.745 180.625 ;
        RECT 61.645 180.580 61.935 180.625 ;
        RECT 64.165 180.580 64.455 180.625 ;
        RECT 60.455 180.440 64.455 180.580 ;
        RECT 60.455 180.395 60.745 180.440 ;
        RECT 61.645 180.395 61.935 180.440 ;
        RECT 64.165 180.395 64.455 180.440 ;
        RECT 65.080 180.580 65.400 180.640 ;
        RECT 69.695 180.580 69.985 180.625 ;
        RECT 65.080 180.440 69.985 180.580 ;
        RECT 79.890 180.580 80.030 180.735 ;
        RECT 81.180 180.720 81.500 180.780 ;
        RECT 81.655 180.735 81.945 180.965 ;
        RECT 85.780 180.720 86.100 180.980 ;
        RECT 90.380 180.720 90.700 180.980 ;
        RECT 96.910 180.920 97.050 181.075 ;
        RECT 97.280 181.060 97.600 181.120 ;
        RECT 97.835 181.075 98.125 181.120 ;
        RECT 101.880 180.920 102.200 180.980 ;
        RECT 96.910 180.780 102.200 180.920 ;
        RECT 101.880 180.720 102.200 180.780 ;
        RECT 103.275 180.735 103.565 180.965 ;
        RECT 104.195 180.920 104.485 180.965 ;
        RECT 105.100 180.920 105.420 180.980 ;
        RECT 108.780 180.920 109.100 180.980 ;
        RECT 104.195 180.780 109.100 180.920 ;
        RECT 104.195 180.735 104.485 180.780 ;
        RECT 91.315 180.580 91.605 180.625 ;
        RECT 91.760 180.580 92.080 180.640 ;
        RECT 103.350 180.580 103.490 180.735 ;
        RECT 105.100 180.720 105.420 180.780 ;
        RECT 108.780 180.720 109.100 180.780 ;
        RECT 104.640 180.580 104.960 180.640 ;
        RECT 79.890 180.440 80.490 180.580 ;
        RECT 65.080 180.380 65.400 180.440 ;
        RECT 69.695 180.395 69.985 180.440 ;
        RECT 60.060 180.240 60.350 180.285 ;
        RECT 62.160 180.240 62.450 180.285 ;
        RECT 63.730 180.240 64.020 180.285 ;
        RECT 60.060 180.100 64.020 180.240 ;
        RECT 60.060 180.055 60.350 180.100 ;
        RECT 62.160 180.055 62.450 180.100 ;
        RECT 63.730 180.055 64.020 180.100 ;
        RECT 80.350 179.960 80.490 180.440 ;
        RECT 91.315 180.440 97.050 180.580 ;
        RECT 103.350 180.440 104.960 180.580 ;
        RECT 109.330 180.580 109.470 181.120 ;
        RECT 109.790 180.920 109.930 181.400 ;
        RECT 111.540 181.260 111.860 181.320 ;
        RECT 115.695 181.260 115.985 181.305 ;
        RECT 111.540 181.120 115.985 181.260 ;
        RECT 118.530 181.260 118.670 181.400 ;
        RECT 121.660 181.260 121.980 181.320 ;
        RECT 124.050 181.305 124.190 181.460 ;
        RECT 141.455 181.460 142.680 181.600 ;
        RECT 141.455 181.415 141.745 181.460 ;
        RECT 142.360 181.400 142.680 181.460 ;
        RECT 142.820 181.600 143.140 181.660 ;
        RECT 144.215 181.600 144.505 181.645 ;
        RECT 142.820 181.460 144.505 181.600 ;
        RECT 142.820 181.400 143.140 181.460 ;
        RECT 144.215 181.415 144.505 181.460 ;
        RECT 147.880 181.600 148.200 181.660 ;
        RECT 153.860 181.600 154.180 181.660 ;
        RECT 154.335 181.600 154.625 181.645 ;
        RECT 147.880 181.460 153.630 181.600 ;
        RECT 147.880 181.400 148.200 181.460 ;
        RECT 118.530 181.120 123.270 181.260 ;
        RECT 111.540 181.060 111.860 181.120 ;
        RECT 115.695 181.075 115.985 181.120 ;
        RECT 121.660 181.060 121.980 181.120 ;
        RECT 112.015 180.920 112.305 180.965 ;
        RECT 109.790 180.780 112.305 180.920 ;
        RECT 112.015 180.735 112.305 180.780 ;
        RECT 116.155 180.920 116.445 180.965 ;
        RECT 118.455 180.920 118.745 180.965 ;
        RECT 116.155 180.780 118.745 180.920 ;
        RECT 116.155 180.735 116.445 180.780 ;
        RECT 118.455 180.735 118.745 180.780 ;
        RECT 120.280 180.920 120.600 180.980 ;
        RECT 123.130 180.965 123.270 181.120 ;
        RECT 123.975 181.075 124.265 181.305 ;
        RECT 150.180 181.260 150.500 181.320 ;
        RECT 149.810 181.120 150.500 181.260 ;
        RECT 121.215 180.920 121.505 180.965 ;
        RECT 120.280 180.780 121.505 180.920 ;
        RECT 120.280 180.720 120.600 180.780 ;
        RECT 121.215 180.735 121.505 180.780 ;
        RECT 123.055 180.735 123.345 180.965 ;
        RECT 123.515 180.920 123.805 180.965 ;
        RECT 124.420 180.920 124.740 180.980 ;
        RECT 149.810 180.965 149.950 181.120 ;
        RECT 150.180 181.060 150.500 181.120 ;
        RECT 150.640 181.260 150.960 181.320 ;
        RECT 152.035 181.260 152.325 181.305 ;
        RECT 150.640 181.120 152.325 181.260 ;
        RECT 150.640 181.060 150.960 181.120 ;
        RECT 152.035 181.075 152.325 181.120 ;
        RECT 123.515 180.780 124.740 180.920 ;
        RECT 123.515 180.735 123.805 180.780 ;
        RECT 124.420 180.720 124.740 180.780 ;
        RECT 124.895 180.920 125.185 180.965 ;
        RECT 126.275 180.920 126.565 180.965 ;
        RECT 124.895 180.780 126.565 180.920 ;
        RECT 124.895 180.735 125.185 180.780 ;
        RECT 126.275 180.735 126.565 180.780 ;
        RECT 149.780 180.735 150.070 180.965 ;
        RECT 151.100 180.720 151.420 180.980 ;
        RECT 151.560 180.920 151.880 180.980 ;
        RECT 152.955 180.920 153.245 180.965 ;
        RECT 151.560 180.780 153.245 180.920 ;
        RECT 153.490 180.920 153.630 181.460 ;
        RECT 153.860 181.460 154.625 181.600 ;
        RECT 153.860 181.400 154.180 181.460 ;
        RECT 154.335 181.415 154.625 181.460 ;
        RECT 155.255 180.920 155.545 180.965 ;
        RECT 153.490 180.780 155.545 180.920 ;
        RECT 151.560 180.720 151.880 180.780 ;
        RECT 152.955 180.735 153.245 180.780 ;
        RECT 155.255 180.735 155.545 180.780 ;
        RECT 109.715 180.580 110.005 180.625 ;
        RECT 109.330 180.440 110.005 180.580 ;
        RECT 91.315 180.395 91.605 180.440 ;
        RECT 91.760 180.380 92.080 180.440 ;
        RECT 89.000 180.240 89.320 180.300 ;
        RECT 92.695 180.240 92.985 180.285 ;
        RECT 93.140 180.240 93.460 180.300 ;
        RECT 94.980 180.240 95.300 180.300 ;
        RECT 89.000 180.100 92.450 180.240 ;
        RECT 89.000 180.040 89.320 180.100 ;
        RECT 25.075 179.900 25.365 179.945 ;
        RECT 25.520 179.900 25.840 179.960 ;
        RECT 25.075 179.760 25.840 179.900 ;
        RECT 25.075 179.715 25.365 179.760 ;
        RECT 25.520 179.700 25.840 179.760 ;
        RECT 32.880 179.700 33.200 179.960 ;
        RECT 37.955 179.900 38.245 179.945 ;
        RECT 42.080 179.900 42.400 179.960 ;
        RECT 37.955 179.760 42.400 179.900 ;
        RECT 37.955 179.715 38.245 179.760 ;
        RECT 42.080 179.700 42.400 179.760 ;
        RECT 54.500 179.700 54.820 179.960 ;
        RECT 66.920 179.700 67.240 179.960 ;
        RECT 70.600 179.900 70.920 179.960 ;
        RECT 75.200 179.900 75.520 179.960 ;
        RECT 70.600 179.760 75.520 179.900 ;
        RECT 70.600 179.700 70.920 179.760 ;
        RECT 75.200 179.700 75.520 179.760 ;
        RECT 80.260 179.700 80.580 179.960 ;
        RECT 87.160 179.900 87.480 179.960 ;
        RECT 88.540 179.900 88.860 179.960 ;
        RECT 89.920 179.900 90.240 179.960 ;
        RECT 87.160 179.760 90.240 179.900 ;
        RECT 92.310 179.900 92.450 180.100 ;
        RECT 92.695 180.100 95.300 180.240 ;
        RECT 92.695 180.055 92.985 180.100 ;
        RECT 93.140 180.040 93.460 180.100 ;
        RECT 94.980 180.040 95.300 180.100 ;
        RECT 96.910 179.960 97.050 180.440 ;
        RECT 104.640 180.380 104.960 180.440 ;
        RECT 109.715 180.395 110.005 180.440 ;
        RECT 129.495 180.580 129.785 180.625 ;
        RECT 129.940 180.580 130.260 180.640 ;
        RECT 129.495 180.440 130.260 180.580 ;
        RECT 129.495 180.395 129.785 180.440 ;
        RECT 129.940 180.380 130.260 180.440 ;
        RECT 132.700 180.380 133.020 180.640 ;
        RECT 138.680 180.580 139.000 180.640 ;
        RECT 139.155 180.580 139.445 180.625 ;
        RECT 138.680 180.440 139.445 180.580 ;
        RECT 138.680 180.380 139.000 180.440 ;
        RECT 139.155 180.395 139.445 180.440 ;
        RECT 146.525 180.580 146.815 180.625 ;
        RECT 149.045 180.580 149.335 180.625 ;
        RECT 150.235 180.580 150.525 180.625 ;
        RECT 146.525 180.440 150.525 180.580 ;
        RECT 146.525 180.395 146.815 180.440 ;
        RECT 149.045 180.395 149.335 180.440 ;
        RECT 150.235 180.395 150.525 180.440 ;
        RECT 134.540 180.040 134.860 180.300 ;
        RECT 140.995 180.240 141.285 180.285 ;
        RECT 143.280 180.240 143.600 180.300 ;
        RECT 140.995 180.100 143.600 180.240 ;
        RECT 140.995 180.055 141.285 180.100 ;
        RECT 143.280 180.040 143.600 180.100 ;
        RECT 146.960 180.240 147.250 180.285 ;
        RECT 148.530 180.240 148.820 180.285 ;
        RECT 150.630 180.240 150.920 180.285 ;
        RECT 146.960 180.100 150.920 180.240 ;
        RECT 146.960 180.055 147.250 180.100 ;
        RECT 148.530 180.055 148.820 180.100 ;
        RECT 150.630 180.055 150.920 180.100 ;
        RECT 94.060 179.900 94.380 179.960 ;
        RECT 94.535 179.900 94.825 179.945 ;
        RECT 92.310 179.760 94.825 179.900 ;
        RECT 87.160 179.700 87.480 179.760 ;
        RECT 88.540 179.700 88.860 179.760 ;
        RECT 89.920 179.700 90.240 179.760 ;
        RECT 94.060 179.700 94.380 179.760 ;
        RECT 94.535 179.715 94.825 179.760 ;
        RECT 95.455 179.900 95.745 179.945 ;
        RECT 95.900 179.900 96.220 179.960 ;
        RECT 95.455 179.760 96.220 179.900 ;
        RECT 95.455 179.715 95.745 179.760 ;
        RECT 95.900 179.700 96.220 179.760 ;
        RECT 96.820 179.700 97.140 179.960 ;
        RECT 97.755 179.900 98.045 179.945 ;
        RECT 98.200 179.900 98.520 179.960 ;
        RECT 97.755 179.760 98.520 179.900 ;
        RECT 97.755 179.715 98.045 179.760 ;
        RECT 98.200 179.700 98.520 179.760 ;
        RECT 98.660 179.700 98.980 179.960 ;
        RECT 103.260 179.700 103.580 179.960 ;
        RECT 110.620 179.700 110.940 179.960 ;
        RECT 122.120 179.700 122.440 179.960 ;
        RECT 135.000 179.700 135.320 179.960 ;
        RECT 147.420 179.900 147.740 179.960 ;
        RECT 153.875 179.900 154.165 179.945 ;
        RECT 147.420 179.760 154.165 179.900 ;
        RECT 147.420 179.700 147.740 179.760 ;
        RECT 153.875 179.715 154.165 179.760 ;
        RECT 22.690 179.080 157.010 179.560 ;
        RECT 31.055 178.880 31.345 178.925 ;
        RECT 31.960 178.880 32.280 178.940 ;
        RECT 31.055 178.740 32.280 178.880 ;
        RECT 31.055 178.695 31.345 178.740 ;
        RECT 31.960 178.680 32.280 178.740 ;
        RECT 32.435 178.880 32.725 178.925 ;
        RECT 32.880 178.880 33.200 178.940 ;
        RECT 32.435 178.740 33.200 178.880 ;
        RECT 32.435 178.695 32.725 178.740 ;
        RECT 32.880 178.680 33.200 178.740 ;
        RECT 35.180 178.880 35.500 178.940 ;
        RECT 37.035 178.880 37.325 178.925 ;
        RECT 43.920 178.880 44.240 178.940 ;
        RECT 35.180 178.740 44.240 178.880 ;
        RECT 35.180 178.680 35.500 178.740 ;
        RECT 37.035 178.695 37.325 178.740 ;
        RECT 43.920 178.680 44.240 178.740 ;
        RECT 51.755 178.880 52.045 178.925 ;
        RECT 54.500 178.880 54.820 178.940 ;
        RECT 51.755 178.740 54.820 178.880 ;
        RECT 51.755 178.695 52.045 178.740 ;
        RECT 54.500 178.680 54.820 178.740 ;
        RECT 56.355 178.880 56.645 178.925 ;
        RECT 61.875 178.880 62.165 178.925 ;
        RECT 65.080 178.880 65.400 178.940 ;
        RECT 56.355 178.740 65.400 178.880 ;
        RECT 56.355 178.695 56.645 178.740 ;
        RECT 61.875 178.695 62.165 178.740 ;
        RECT 65.080 178.680 65.400 178.740 ;
        RECT 74.740 178.680 75.060 178.940 ;
        RECT 89.935 178.695 90.225 178.925 ;
        RECT 90.380 178.880 90.700 178.940 ;
        RECT 91.775 178.880 92.065 178.925 ;
        RECT 90.380 178.740 92.065 178.880 ;
        RECT 24.640 178.540 24.930 178.585 ;
        RECT 26.740 178.540 27.030 178.585 ;
        RECT 28.310 178.540 28.600 178.585 ;
        RECT 24.640 178.400 28.600 178.540 ;
        RECT 24.640 178.355 24.930 178.400 ;
        RECT 26.740 178.355 27.030 178.400 ;
        RECT 28.310 178.355 28.600 178.400 ;
        RECT 31.515 178.355 31.805 178.585 ;
        RECT 25.035 178.200 25.325 178.245 ;
        RECT 26.225 178.200 26.515 178.245 ;
        RECT 28.745 178.200 29.035 178.245 ;
        RECT 31.590 178.200 31.730 178.355 ;
        RECT 25.035 178.060 29.035 178.200 ;
        RECT 25.035 178.015 25.325 178.060 ;
        RECT 26.225 178.015 26.515 178.060 ;
        RECT 28.745 178.015 29.035 178.060 ;
        RECT 29.290 178.060 31.730 178.200 ;
        RECT 32.050 178.200 32.190 178.680 ;
        RECT 34.260 178.540 34.580 178.600 ;
        RECT 36.115 178.540 36.405 178.585 ;
        RECT 34.260 178.400 36.405 178.540 ;
        RECT 34.260 178.340 34.580 178.400 ;
        RECT 36.115 178.355 36.405 178.400 ;
        RECT 42.540 178.540 42.860 178.600 ;
        RECT 42.540 178.400 46.450 178.540 ;
        RECT 42.540 178.340 42.860 178.400 ;
        RECT 45.300 178.200 45.620 178.260 ;
        RECT 45.775 178.200 46.065 178.245 ;
        RECT 32.050 178.060 38.170 178.200 ;
        RECT 24.155 177.675 24.445 177.905 ;
        RECT 29.290 177.860 29.430 178.060 ;
        RECT 37.020 177.860 37.340 177.920 ;
        RECT 26.070 177.720 29.430 177.860 ;
        RECT 31.590 177.720 37.340 177.860 ;
        RECT 24.230 177.180 24.370 177.675 ;
        RECT 26.070 177.580 26.210 177.720 ;
        RECT 25.520 177.565 25.840 177.580 ;
        RECT 25.490 177.520 25.840 177.565 ;
        RECT 25.325 177.380 25.840 177.520 ;
        RECT 25.490 177.335 25.840 177.380 ;
        RECT 25.520 177.320 25.840 177.335 ;
        RECT 25.980 177.320 26.300 177.580 ;
        RECT 29.200 177.520 29.520 177.580 ;
        RECT 31.590 177.520 31.730 177.720 ;
        RECT 36.805 177.660 37.340 177.720 ;
        RECT 38.030 177.860 38.170 178.060 ;
        RECT 45.300 178.060 46.065 178.200 ;
        RECT 46.310 178.200 46.450 178.400 ;
        RECT 48.520 178.340 48.840 178.600 ;
        RECT 52.200 178.540 52.520 178.600 ;
        RECT 64.620 178.540 64.910 178.585 ;
        RECT 66.190 178.540 66.480 178.585 ;
        RECT 68.290 178.540 68.580 178.585 ;
        RECT 52.200 178.400 55.650 178.540 ;
        RECT 52.200 178.340 52.520 178.400 ;
        RECT 51.295 178.200 51.585 178.245 ;
        RECT 46.310 178.060 55.190 178.200 ;
        RECT 45.300 178.000 45.620 178.060 ;
        RECT 45.775 178.015 46.065 178.060 ;
        RECT 51.295 178.015 51.585 178.060 ;
        RECT 43.475 177.860 43.765 177.905 ;
        RECT 48.995 177.860 49.285 177.905 ;
        RECT 38.030 177.720 49.285 177.860 ;
        RECT 35.640 177.520 35.960 177.580 ;
        RECT 29.200 177.380 31.730 177.520 ;
        RECT 32.050 177.380 35.960 177.520 ;
        RECT 36.805 177.550 37.120 177.660 ;
        RECT 38.030 177.565 38.170 177.720 ;
        RECT 43.475 177.675 43.765 177.720 ;
        RECT 48.995 177.675 49.285 177.720 ;
        RECT 53.890 177.860 54.180 177.905 ;
        RECT 54.500 177.860 54.820 177.920 ;
        RECT 55.050 177.905 55.190 178.060 ;
        RECT 53.890 177.720 54.820 177.860 ;
        RECT 53.890 177.675 54.180 177.720 ;
        RECT 54.500 177.660 54.820 177.720 ;
        RECT 54.975 177.675 55.265 177.905 ;
        RECT 55.510 177.860 55.650 178.400 ;
        RECT 64.620 178.400 68.580 178.540 ;
        RECT 74.830 178.540 74.970 178.680 ;
        RECT 78.920 178.540 79.210 178.585 ;
        RECT 81.020 178.540 81.310 178.585 ;
        RECT 82.590 178.540 82.880 178.585 ;
        RECT 74.830 178.400 78.650 178.540 ;
        RECT 64.620 178.355 64.910 178.400 ;
        RECT 66.190 178.355 66.480 178.400 ;
        RECT 68.290 178.355 68.580 178.400 ;
        RECT 78.510 178.245 78.650 178.400 ;
        RECT 78.920 178.400 82.880 178.540 ;
        RECT 90.010 178.540 90.150 178.695 ;
        RECT 90.380 178.680 90.700 178.740 ;
        RECT 91.775 178.695 92.065 178.740 ;
        RECT 94.520 178.680 94.840 178.940 ;
        RECT 94.980 178.680 95.300 178.940 ;
        RECT 95.915 178.880 96.205 178.925 ;
        RECT 97.740 178.880 98.060 178.940 ;
        RECT 95.915 178.740 98.060 178.880 ;
        RECT 95.915 178.695 96.205 178.740 ;
        RECT 97.740 178.680 98.060 178.740 ;
        RECT 98.660 178.880 98.980 178.940 ;
        RECT 100.975 178.880 101.265 178.925 ;
        RECT 98.660 178.740 101.265 178.880 ;
        RECT 98.660 178.680 98.980 178.740 ;
        RECT 100.975 178.695 101.265 178.740 ;
        RECT 101.420 178.680 101.740 178.940 ;
        RECT 101.880 178.680 102.200 178.940 ;
        RECT 127.180 178.880 127.500 178.940 ;
        RECT 140.520 178.880 140.840 178.940 ;
        RECT 102.430 178.740 140.840 178.880 ;
        RECT 91.300 178.540 91.620 178.600 ;
        RECT 90.010 178.400 91.620 178.540 ;
        RECT 78.920 178.355 79.210 178.400 ;
        RECT 81.020 178.355 81.310 178.400 ;
        RECT 82.590 178.355 82.880 178.400 ;
        RECT 91.300 178.340 91.620 178.400 ;
        RECT 92.220 178.540 92.540 178.600 ;
        RECT 94.060 178.540 94.380 178.600 ;
        RECT 92.220 178.400 94.380 178.540 ;
        RECT 92.220 178.340 92.540 178.400 ;
        RECT 94.060 178.340 94.380 178.400 ;
        RECT 64.185 178.200 64.475 178.245 ;
        RECT 66.705 178.200 66.995 178.245 ;
        RECT 67.895 178.200 68.185 178.245 ;
        RECT 64.185 178.060 68.185 178.200 ;
        RECT 64.185 178.015 64.475 178.060 ;
        RECT 66.705 178.015 66.995 178.060 ;
        RECT 67.895 178.015 68.185 178.060 ;
        RECT 68.775 178.200 69.065 178.245 ;
        RECT 68.775 178.060 75.430 178.200 ;
        RECT 68.775 178.015 69.065 178.060 ;
        RECT 75.290 177.920 75.430 178.060 ;
        RECT 78.435 178.015 78.725 178.245 ;
        RECT 79.315 178.200 79.605 178.245 ;
        RECT 80.505 178.200 80.795 178.245 ;
        RECT 83.025 178.200 83.315 178.245 ;
        RECT 79.315 178.060 83.315 178.200 ;
        RECT 79.315 178.015 79.605 178.060 ;
        RECT 80.505 178.015 80.795 178.060 ;
        RECT 83.025 178.015 83.315 178.060 ;
        RECT 87.160 178.200 87.480 178.260 ;
        RECT 89.000 178.200 89.320 178.260 ;
        RECT 90.840 178.200 91.160 178.260 ;
        RECT 92.680 178.200 93.000 178.260 ;
        RECT 95.440 178.200 95.760 178.260 ;
        RECT 87.160 178.060 89.320 178.200 ;
        RECT 87.160 178.000 87.480 178.060 ;
        RECT 89.000 178.000 89.320 178.060 ;
        RECT 89.550 178.060 93.000 178.200 ;
        RECT 57.720 177.860 58.040 177.920 ;
        RECT 55.510 177.720 58.040 177.860 ;
        RECT 36.805 177.505 37.095 177.550 ;
        RECT 29.200 177.320 29.520 177.380 ;
        RECT 32.050 177.180 32.190 177.380 ;
        RECT 35.640 177.320 35.960 177.380 ;
        RECT 37.955 177.335 38.245 177.565 ;
        RECT 45.315 177.520 45.605 177.565 ;
        RECT 46.695 177.520 46.985 177.565 ;
        RECT 45.315 177.380 46.985 177.520 ;
        RECT 45.315 177.335 45.605 177.380 ;
        RECT 46.695 177.335 46.985 177.380 ;
        RECT 47.615 177.520 47.905 177.565 ;
        RECT 48.060 177.520 48.380 177.580 ;
        RECT 47.615 177.380 48.380 177.520 ;
        RECT 47.615 177.335 47.905 177.380 ;
        RECT 48.060 177.320 48.380 177.380 ;
        RECT 24.230 177.040 32.190 177.180 ;
        RECT 32.435 177.180 32.725 177.225 ;
        RECT 33.340 177.180 33.660 177.240 ;
        RECT 32.435 177.040 33.660 177.180 ;
        RECT 32.435 176.995 32.725 177.040 ;
        RECT 33.340 176.980 33.660 177.040 ;
        RECT 43.920 176.980 44.240 177.240 ;
        RECT 44.380 176.980 44.700 177.240 ;
        RECT 47.140 176.980 47.460 177.240 ;
        RECT 49.455 177.180 49.745 177.225 ;
        RECT 53.595 177.180 53.885 177.225 ;
        RECT 54.040 177.180 54.360 177.240 ;
        RECT 49.455 177.040 54.360 177.180 ;
        RECT 49.455 176.995 49.745 177.040 ;
        RECT 53.595 176.995 53.885 177.040 ;
        RECT 54.040 176.980 54.360 177.040 ;
        RECT 54.515 177.180 54.805 177.225 ;
        RECT 55.510 177.180 55.650 177.720 ;
        RECT 57.720 177.660 58.040 177.720 ;
        RECT 58.655 177.860 58.945 177.905 ;
        RECT 59.100 177.860 59.420 177.920 ;
        RECT 70.140 177.860 70.460 177.920 ;
        RECT 58.655 177.720 59.420 177.860 ;
        RECT 58.655 177.675 58.945 177.720 ;
        RECT 59.100 177.660 59.420 177.720 ;
        RECT 68.850 177.720 70.460 177.860 ;
        RECT 58.180 177.320 58.500 177.580 ;
        RECT 63.240 177.520 63.560 177.580 ;
        RECT 67.440 177.520 67.730 177.565 ;
        RECT 63.240 177.380 67.730 177.520 ;
        RECT 63.240 177.320 63.560 177.380 ;
        RECT 67.440 177.335 67.730 177.380 ;
        RECT 54.515 177.040 55.650 177.180 ;
        RECT 54.515 176.995 54.805 177.040 ;
        RECT 57.260 176.980 57.580 177.240 ;
        RECT 64.160 177.180 64.480 177.240 ;
        RECT 68.850 177.180 68.990 177.720 ;
        RECT 70.140 177.660 70.460 177.720 ;
        RECT 70.600 177.660 70.920 177.920 ;
        RECT 71.980 177.660 72.300 177.920 ;
        RECT 72.455 177.675 72.745 177.905 ;
        RECT 71.060 177.320 71.380 177.580 ;
        RECT 71.520 177.520 71.840 177.580 ;
        RECT 72.530 177.520 72.670 177.675 ;
        RECT 75.200 177.660 75.520 177.920 ;
        RECT 89.550 177.905 89.690 178.060 ;
        RECT 90.840 178.000 91.160 178.060 ;
        RECT 92.680 178.000 93.000 178.060 ;
        RECT 93.690 178.060 95.760 178.200 ;
        RECT 89.475 177.675 89.765 177.905 ;
        RECT 89.920 177.860 90.240 177.920 ;
        RECT 93.690 177.905 93.830 178.060 ;
        RECT 95.440 178.000 95.760 178.060 ;
        RECT 95.900 178.000 96.220 178.260 ;
        RECT 93.615 177.860 93.905 177.905 ;
        RECT 89.920 177.720 93.905 177.860 ;
        RECT 95.990 177.860 96.130 178.000 ;
        RECT 97.295 177.860 97.585 177.905 ;
        RECT 95.990 177.720 97.585 177.860 ;
        RECT 97.830 177.860 97.970 178.680 ;
        RECT 98.215 178.540 98.505 178.585 ;
        RECT 101.510 178.540 101.650 178.680 ;
        RECT 98.215 178.400 101.650 178.540 ;
        RECT 98.215 178.355 98.505 178.400 ;
        RECT 102.430 178.200 102.570 178.740 ;
        RECT 127.180 178.680 127.500 178.740 ;
        RECT 140.520 178.680 140.840 178.740 ;
        RECT 142.835 178.880 143.125 178.925 ;
        RECT 143.740 178.880 144.060 178.940 ;
        RECT 149.260 178.880 149.580 178.940 ;
        RECT 142.835 178.740 144.060 178.880 ;
        RECT 142.835 178.695 143.125 178.740 ;
        RECT 143.740 178.680 144.060 178.740 ;
        RECT 144.290 178.740 149.580 178.880 ;
        RECT 113.880 178.540 114.170 178.585 ;
        RECT 115.980 178.540 116.270 178.585 ;
        RECT 117.550 178.540 117.840 178.585 ;
        RECT 102.890 178.400 103.950 178.540 ;
        RECT 102.890 178.260 103.030 178.400 ;
        RECT 100.130 178.060 102.570 178.200 ;
        RECT 100.130 177.905 100.270 178.060 ;
        RECT 102.800 178.000 103.120 178.260 ;
        RECT 103.260 178.000 103.580 178.260 ;
        RECT 103.810 178.200 103.950 178.400 ;
        RECT 113.880 178.400 117.840 178.540 ;
        RECT 113.880 178.355 114.170 178.400 ;
        RECT 115.980 178.355 116.270 178.400 ;
        RECT 117.550 178.355 117.840 178.400 ;
        RECT 121.240 178.540 121.530 178.585 ;
        RECT 123.340 178.540 123.630 178.585 ;
        RECT 124.910 178.540 125.200 178.585 ;
        RECT 121.240 178.400 125.200 178.540 ;
        RECT 121.240 178.355 121.530 178.400 ;
        RECT 123.340 178.355 123.630 178.400 ;
        RECT 124.910 178.355 125.200 178.400 ;
        RECT 127.655 178.540 127.945 178.585 ;
        RECT 129.940 178.540 130.260 178.600 ;
        RECT 127.655 178.400 130.260 178.540 ;
        RECT 127.655 178.355 127.945 178.400 ;
        RECT 129.940 178.340 130.260 178.400 ;
        RECT 133.635 178.540 133.925 178.585 ;
        RECT 137.775 178.540 138.065 178.585 ;
        RECT 133.635 178.400 138.065 178.540 ;
        RECT 133.635 178.355 133.925 178.400 ;
        RECT 137.775 178.355 138.065 178.400 ;
        RECT 141.440 178.540 141.760 178.600 ;
        RECT 144.290 178.540 144.430 178.740 ;
        RECT 149.260 178.680 149.580 178.740 ;
        RECT 146.960 178.540 147.280 178.600 ;
        RECT 141.440 178.400 144.430 178.540 ;
        RECT 141.440 178.340 141.760 178.400 ;
        RECT 105.115 178.200 105.405 178.245 ;
        RECT 103.810 178.060 105.405 178.200 ;
        RECT 105.115 178.015 105.405 178.060 ;
        RECT 114.275 178.200 114.565 178.245 ;
        RECT 115.465 178.200 115.755 178.245 ;
        RECT 117.985 178.200 118.275 178.245 ;
        RECT 114.275 178.060 118.275 178.200 ;
        RECT 114.275 178.015 114.565 178.060 ;
        RECT 115.465 178.015 115.755 178.060 ;
        RECT 117.985 178.015 118.275 178.060 ;
        RECT 118.900 178.200 119.220 178.260 ;
        RECT 120.755 178.200 121.045 178.245 ;
        RECT 118.900 178.060 121.045 178.200 ;
        RECT 118.900 178.000 119.220 178.060 ;
        RECT 120.755 178.015 121.045 178.060 ;
        RECT 121.635 178.200 121.925 178.245 ;
        RECT 122.825 178.200 123.115 178.245 ;
        RECT 125.345 178.200 125.635 178.245 ;
        RECT 121.635 178.060 125.635 178.200 ;
        RECT 121.635 178.015 121.925 178.060 ;
        RECT 122.825 178.015 123.115 178.060 ;
        RECT 125.345 178.015 125.635 178.060 ;
        RECT 129.020 178.000 129.340 178.260 ;
        RECT 130.415 178.200 130.705 178.245 ;
        RECT 132.700 178.200 133.020 178.260 ;
        RECT 136.380 178.200 136.700 178.260 ;
        RECT 130.415 178.060 136.700 178.200 ;
        RECT 130.415 178.015 130.705 178.060 ;
        RECT 132.700 178.000 133.020 178.060 ;
        RECT 136.380 178.000 136.700 178.060 ;
        RECT 136.855 178.200 137.145 178.245 ;
        RECT 136.855 178.060 142.130 178.200 ;
        RECT 136.855 178.015 137.145 178.060 ;
        RECT 100.055 177.860 100.345 177.905 ;
        RECT 97.830 177.720 100.345 177.860 ;
        RECT 71.520 177.380 72.670 177.520 ;
        RECT 79.770 177.520 80.060 177.565 ;
        RECT 84.400 177.520 84.720 177.580 ;
        RECT 79.770 177.380 84.720 177.520 ;
        RECT 71.520 177.320 71.840 177.380 ;
        RECT 79.770 177.335 80.060 177.380 ;
        RECT 84.400 177.320 84.720 177.380 ;
        RECT 64.160 177.040 68.990 177.180 ;
        RECT 64.160 176.980 64.480 177.040 ;
        RECT 69.220 176.980 69.540 177.240 ;
        RECT 75.675 177.180 75.965 177.225 ;
        RECT 78.880 177.180 79.200 177.240 ;
        RECT 75.675 177.040 79.200 177.180 ;
        RECT 75.675 176.995 75.965 177.040 ;
        RECT 78.880 176.980 79.200 177.040 ;
        RECT 85.320 177.180 85.640 177.240 ;
        RECT 89.550 177.180 89.690 177.675 ;
        RECT 89.920 177.660 90.240 177.720 ;
        RECT 93.615 177.675 93.905 177.720 ;
        RECT 97.295 177.675 97.585 177.720 ;
        RECT 100.055 177.675 100.345 177.720 ;
        RECT 101.420 177.660 101.740 177.920 ;
        RECT 103.735 177.675 104.025 177.905 ;
        RECT 106.495 177.675 106.785 177.905 ;
        RECT 92.220 177.520 92.540 177.580 ;
        RECT 92.695 177.520 92.985 177.565 ;
        RECT 96.835 177.520 97.125 177.565 ;
        RECT 92.220 177.380 92.985 177.520 ;
        RECT 92.220 177.320 92.540 177.380 ;
        RECT 92.695 177.335 92.985 177.380 ;
        RECT 93.690 177.380 97.125 177.520 ;
        RECT 103.810 177.520 103.950 177.675 ;
        RECT 104.655 177.520 104.945 177.565 ;
        RECT 103.810 177.380 104.945 177.520 ;
        RECT 106.570 177.520 106.710 177.675 ;
        RECT 106.940 177.660 107.260 177.920 ;
        RECT 110.620 177.660 110.940 177.920 ;
        RECT 113.395 177.860 113.685 177.905 ;
        RECT 118.990 177.860 119.130 178.000 ;
        RECT 122.120 177.905 122.440 177.920 ;
        RECT 122.090 177.860 122.440 177.905 ;
        RECT 113.395 177.720 119.130 177.860 ;
        RECT 121.925 177.720 122.440 177.860 ;
        RECT 129.110 177.860 129.250 178.000 ;
        RECT 133.160 177.860 133.480 177.920 ;
        RECT 129.110 177.720 133.480 177.860 ;
        RECT 113.395 177.675 113.685 177.720 ;
        RECT 122.090 177.675 122.440 177.720 ;
        RECT 122.120 177.660 122.440 177.675 ;
        RECT 133.160 177.660 133.480 177.720 ;
        RECT 135.000 177.660 135.320 177.920 ;
        RECT 135.460 177.660 135.780 177.920 ;
        RECT 137.300 177.660 137.620 177.920 ;
        RECT 140.075 177.860 140.365 177.905 ;
        RECT 140.520 177.860 140.840 177.920 ;
        RECT 140.075 177.720 140.840 177.860 ;
        RECT 140.075 177.675 140.365 177.720 ;
        RECT 140.520 177.660 140.840 177.720 ;
        RECT 140.995 177.675 141.285 177.905 ;
        RECT 110.710 177.520 110.850 177.660 ;
        RECT 114.620 177.520 114.910 177.565 ;
        RECT 106.570 177.380 110.390 177.520 ;
        RECT 110.710 177.380 114.910 177.520 ;
        RECT 93.690 177.240 93.830 177.380 ;
        RECT 96.835 177.335 97.125 177.380 ;
        RECT 104.655 177.335 104.945 177.380 ;
        RECT 85.320 177.040 89.690 177.180 ;
        RECT 85.320 176.980 85.640 177.040 ;
        RECT 93.600 176.980 93.920 177.240 ;
        RECT 95.900 177.225 96.220 177.240 ;
        RECT 95.835 176.995 96.220 177.225 ;
        RECT 95.900 176.980 96.220 176.995 ;
        RECT 98.200 177.180 98.520 177.240 ;
        RECT 99.135 177.180 99.425 177.225 ;
        RECT 99.580 177.180 99.900 177.240 ;
        RECT 98.200 177.040 99.900 177.180 ;
        RECT 104.730 177.180 104.870 177.335 ;
        RECT 106.020 177.180 106.340 177.240 ;
        RECT 104.730 177.040 106.340 177.180 ;
        RECT 98.200 176.980 98.520 177.040 ;
        RECT 99.135 176.995 99.425 177.040 ;
        RECT 99.580 176.980 99.900 177.040 ;
        RECT 106.020 176.980 106.340 177.040 ;
        RECT 106.480 177.180 106.800 177.240 ;
        RECT 107.875 177.180 108.165 177.225 ;
        RECT 106.480 177.040 108.165 177.180 ;
        RECT 110.250 177.180 110.390 177.380 ;
        RECT 114.620 177.335 114.910 177.380 ;
        RECT 128.100 177.320 128.420 177.580 ;
        RECT 112.460 177.180 112.780 177.240 ;
        RECT 110.250 177.040 112.780 177.180 ;
        RECT 106.480 176.980 106.800 177.040 ;
        RECT 107.875 176.995 108.165 177.040 ;
        RECT 112.460 176.980 112.780 177.040 ;
        RECT 118.440 177.180 118.760 177.240 ;
        RECT 120.280 177.180 120.600 177.240 ;
        RECT 118.440 177.040 120.600 177.180 ;
        RECT 118.440 176.980 118.760 177.040 ;
        RECT 120.280 176.980 120.600 177.040 ;
        RECT 134.080 177.180 134.400 177.240 ;
        RECT 134.555 177.180 134.845 177.225 ;
        RECT 134.080 177.040 134.845 177.180 ;
        RECT 134.080 176.980 134.400 177.040 ;
        RECT 134.555 176.995 134.845 177.040 ;
        RECT 138.680 177.180 139.000 177.240 ;
        RECT 139.155 177.180 139.445 177.225 ;
        RECT 138.680 177.040 139.445 177.180 ;
        RECT 141.070 177.180 141.210 177.675 ;
        RECT 141.440 177.660 141.760 177.920 ;
        RECT 141.990 177.520 142.130 178.060 ;
        RECT 144.290 177.905 144.430 178.400 ;
        RECT 145.670 178.400 147.280 178.540 ;
        RECT 145.670 177.905 145.810 178.400 ;
        RECT 146.960 178.340 147.280 178.400 ;
        RECT 148.380 178.540 148.670 178.585 ;
        RECT 150.480 178.540 150.770 178.585 ;
        RECT 152.050 178.540 152.340 178.585 ;
        RECT 148.380 178.400 152.340 178.540 ;
        RECT 148.380 178.355 148.670 178.400 ;
        RECT 150.480 178.355 150.770 178.400 ;
        RECT 152.050 178.355 152.340 178.400 ;
        RECT 148.775 178.200 149.065 178.245 ;
        RECT 149.965 178.200 150.255 178.245 ;
        RECT 152.485 178.200 152.775 178.245 ;
        RECT 146.130 178.060 148.570 178.200 ;
        RECT 146.130 177.905 146.270 178.060 ;
        RECT 144.215 177.675 144.505 177.905 ;
        RECT 145.135 177.675 145.425 177.905 ;
        RECT 145.595 177.675 145.885 177.905 ;
        RECT 146.055 177.675 146.345 177.905 ;
        RECT 147.420 177.860 147.740 177.920 ;
        RECT 147.895 177.860 148.185 177.905 ;
        RECT 147.420 177.720 148.185 177.860 ;
        RECT 148.430 177.860 148.570 178.060 ;
        RECT 148.775 178.060 152.775 178.200 ;
        RECT 148.775 178.015 149.065 178.060 ;
        RECT 149.965 178.015 150.255 178.060 ;
        RECT 152.485 178.015 152.775 178.060 ;
        RECT 148.430 177.720 152.250 177.860 ;
        RECT 142.675 177.520 142.965 177.565 ;
        RECT 141.990 177.380 142.965 177.520 ;
        RECT 142.675 177.335 142.965 177.380 ;
        RECT 143.740 177.320 144.060 177.580 ;
        RECT 145.210 177.520 145.350 177.675 ;
        RECT 147.420 177.660 147.740 177.720 ;
        RECT 147.895 177.675 148.185 177.720 ;
        RECT 146.960 177.520 147.280 177.580 ;
        RECT 149.120 177.520 149.410 177.565 ;
        RECT 145.210 177.380 147.280 177.520 ;
        RECT 146.960 177.320 147.280 177.380 ;
        RECT 147.510 177.380 149.410 177.520 ;
        RECT 147.510 177.225 147.650 177.380 ;
        RECT 149.120 177.335 149.410 177.380 ;
        RECT 152.110 177.240 152.250 177.720 ;
        RECT 141.915 177.180 142.205 177.225 ;
        RECT 141.070 177.040 142.205 177.180 ;
        RECT 138.680 176.980 139.000 177.040 ;
        RECT 139.155 176.995 139.445 177.040 ;
        RECT 141.915 176.995 142.205 177.040 ;
        RECT 147.435 176.995 147.725 177.225 ;
        RECT 152.020 176.980 152.340 177.240 ;
        RECT 154.780 176.980 155.100 177.240 ;
        RECT 22.690 176.360 157.810 176.840 ;
        RECT 35.180 176.160 35.500 176.220 ;
        RECT 34.810 176.020 35.500 176.160 ;
        RECT 30.135 175.820 30.425 175.865 ;
        RECT 31.040 175.820 31.360 175.880 ;
        RECT 30.135 175.680 31.360 175.820 ;
        RECT 30.135 175.635 30.425 175.680 ;
        RECT 25.995 175.295 26.285 175.525 ;
        RECT 26.070 174.800 26.210 175.295 ;
        RECT 29.200 175.280 29.520 175.540 ;
        RECT 30.210 175.480 30.350 175.635 ;
        RECT 31.040 175.620 31.360 175.680 ;
        RECT 32.435 175.820 32.725 175.865 ;
        RECT 33.800 175.820 34.120 175.880 ;
        RECT 34.810 175.865 34.950 176.020 ;
        RECT 35.180 175.960 35.500 176.020 ;
        RECT 35.640 175.960 35.960 176.220 ;
        RECT 44.855 176.160 45.145 176.205 ;
        RECT 54.960 176.160 55.280 176.220 ;
        RECT 44.855 176.020 54.730 176.160 ;
        RECT 44.855 175.975 45.145 176.020 ;
        RECT 32.435 175.680 34.120 175.820 ;
        RECT 32.435 175.635 32.725 175.680 ;
        RECT 33.800 175.620 34.120 175.680 ;
        RECT 34.735 175.635 35.025 175.865 ;
        RECT 35.730 175.820 35.870 175.960 ;
        RECT 43.920 175.820 44.240 175.880 ;
        RECT 48.075 175.820 48.365 175.865 ;
        RECT 50.360 175.820 50.680 175.880 ;
        RECT 35.730 175.680 36.330 175.820 ;
        RECT 30.595 175.480 30.885 175.525 ;
        RECT 30.210 175.340 30.885 175.480 ;
        RECT 30.595 175.295 30.885 175.340 ;
        RECT 28.295 175.140 28.585 175.185 ;
        RECT 34.810 175.140 34.950 175.635 ;
        RECT 36.190 175.525 36.330 175.680 ;
        RECT 43.920 175.680 44.610 175.820 ;
        RECT 43.920 175.620 44.240 175.680 ;
        RECT 37.480 175.525 37.800 175.540 ;
        RECT 44.470 175.525 44.610 175.680 ;
        RECT 48.075 175.680 50.680 175.820 ;
        RECT 54.590 175.820 54.730 176.020 ;
        RECT 54.960 176.020 57.950 176.160 ;
        RECT 54.960 175.960 55.280 176.020 ;
        RECT 57.810 175.820 57.950 176.020 ;
        RECT 58.180 175.960 58.500 176.220 ;
        RECT 58.730 176.020 62.090 176.160 ;
        RECT 58.730 175.820 58.870 176.020 ;
        RECT 54.590 175.680 57.490 175.820 ;
        RECT 57.810 175.680 58.870 175.820 ;
        RECT 61.950 175.820 62.090 176.020 ;
        RECT 63.240 175.960 63.560 176.220 ;
        RECT 66.935 176.160 67.225 176.205 ;
        RECT 71.520 176.160 71.840 176.220 ;
        RECT 66.935 176.020 71.840 176.160 ;
        RECT 66.935 175.975 67.225 176.020 ;
        RECT 67.010 175.820 67.150 175.975 ;
        RECT 71.520 175.960 71.840 176.020 ;
        RECT 71.980 176.160 72.300 176.220 ;
        RECT 74.755 176.160 75.045 176.205 ;
        RECT 71.980 176.020 75.045 176.160 ;
        RECT 71.980 175.960 72.300 176.020 ;
        RECT 74.755 175.975 75.045 176.020 ;
        RECT 78.435 175.975 78.725 176.205 ;
        RECT 78.880 176.160 79.200 176.220 ;
        RECT 85.320 176.160 85.640 176.220 ;
        RECT 78.880 176.020 81.410 176.160 ;
        RECT 71.060 175.820 71.380 175.880 ;
        RECT 61.950 175.680 67.150 175.820 ;
        RECT 68.160 175.680 71.380 175.820 ;
        RECT 48.075 175.635 48.365 175.680 ;
        RECT 50.360 175.620 50.680 175.680 ;
        RECT 35.560 175.480 35.850 175.525 ;
        RECT 28.295 175.000 34.950 175.140 ;
        RECT 35.270 175.340 35.850 175.480 ;
        RECT 28.295 174.955 28.585 175.000 ;
        RECT 33.355 174.800 33.645 174.845 ;
        RECT 26.070 174.660 33.645 174.800 ;
        RECT 33.355 174.615 33.645 174.660 ;
        RECT 25.075 174.460 25.365 174.505 ;
        RECT 25.520 174.460 25.840 174.520 ;
        RECT 25.075 174.320 25.840 174.460 ;
        RECT 25.075 174.275 25.365 174.320 ;
        RECT 25.520 174.260 25.840 174.320 ;
        RECT 32.435 174.460 32.725 174.505 ;
        RECT 33.815 174.460 34.105 174.505 ;
        RECT 32.435 174.320 34.105 174.460 ;
        RECT 35.270 174.460 35.410 175.340 ;
        RECT 35.560 175.295 35.850 175.340 ;
        RECT 36.115 175.295 36.405 175.525 ;
        RECT 37.450 175.295 37.800 175.525 ;
        RECT 44.395 175.295 44.685 175.525 ;
        RECT 37.480 175.280 37.800 175.295 ;
        RECT 46.220 175.280 46.540 175.540 ;
        RECT 50.820 175.280 51.140 175.540 ;
        RECT 51.295 175.295 51.585 175.525 ;
        RECT 52.200 175.480 52.520 175.540 ;
        RECT 52.675 175.480 52.965 175.525 ;
        RECT 52.200 175.340 52.965 175.480 ;
        RECT 36.995 175.140 37.285 175.185 ;
        RECT 38.185 175.140 38.475 175.185 ;
        RECT 40.705 175.140 40.995 175.185 ;
        RECT 36.995 175.000 40.995 175.140 ;
        RECT 51.370 175.140 51.510 175.295 ;
        RECT 52.200 175.280 52.520 175.340 ;
        RECT 52.675 175.295 52.965 175.340 ;
        RECT 54.040 175.280 54.360 175.540 ;
        RECT 54.960 175.280 55.280 175.540 ;
        RECT 55.510 175.525 55.650 175.680 ;
        RECT 57.350 175.530 57.490 175.680 ;
        RECT 57.350 175.525 57.950 175.530 ;
        RECT 55.435 175.295 55.725 175.525 ;
        RECT 55.895 175.480 56.185 175.525 ;
        RECT 55.895 175.340 56.570 175.480 ;
        RECT 55.895 175.295 56.185 175.340 ;
        RECT 51.370 175.000 56.090 175.140 ;
        RECT 36.995 174.955 37.285 175.000 ;
        RECT 38.185 174.955 38.475 175.000 ;
        RECT 40.705 174.955 40.995 175.000 ;
        RECT 36.600 174.800 36.890 174.845 ;
        RECT 38.700 174.800 38.990 174.845 ;
        RECT 40.270 174.800 40.560 174.845 ;
        RECT 36.600 174.660 40.560 174.800 ;
        RECT 36.600 174.615 36.890 174.660 ;
        RECT 38.700 174.615 38.990 174.660 ;
        RECT 40.270 174.615 40.560 174.660 ;
        RECT 43.015 174.800 43.305 174.845 ;
        RECT 44.380 174.800 44.700 174.860 ;
        RECT 49.915 174.800 50.205 174.845 ;
        RECT 52.660 174.800 52.980 174.860 ;
        RECT 43.015 174.660 47.370 174.800 ;
        RECT 43.015 174.615 43.305 174.660 ;
        RECT 37.020 174.460 37.340 174.520 ;
        RECT 35.270 174.320 37.340 174.460 ;
        RECT 32.435 174.275 32.725 174.320 ;
        RECT 33.815 174.275 34.105 174.320 ;
        RECT 37.020 174.260 37.340 174.320 ;
        RECT 37.940 174.460 38.260 174.520 ;
        RECT 43.090 174.460 43.230 174.615 ;
        RECT 44.380 174.600 44.700 174.660 ;
        RECT 37.940 174.320 43.230 174.460 ;
        RECT 47.230 174.460 47.370 174.660 ;
        RECT 49.915 174.660 52.980 174.800 ;
        RECT 49.915 174.615 50.205 174.660 ;
        RECT 52.660 174.600 52.980 174.660 ;
        RECT 53.210 174.660 54.730 174.800 ;
        RECT 51.740 174.460 52.060 174.520 ;
        RECT 47.230 174.320 52.060 174.460 ;
        RECT 37.940 174.260 38.260 174.320 ;
        RECT 51.740 174.260 52.060 174.320 ;
        RECT 52.200 174.260 52.520 174.520 ;
        RECT 53.210 174.505 53.350 174.660 ;
        RECT 54.590 174.520 54.730 174.660 ;
        RECT 53.135 174.275 53.425 174.505 ;
        RECT 54.500 174.260 54.820 174.520 ;
        RECT 55.950 174.460 56.090 175.000 ;
        RECT 56.430 174.800 56.570 175.340 ;
        RECT 56.815 175.295 57.105 175.525 ;
        RECT 57.350 175.390 58.190 175.525 ;
        RECT 57.810 175.340 58.190 175.390 ;
        RECT 57.900 175.295 58.190 175.340 ;
        RECT 59.560 175.480 59.880 175.540 ;
        RECT 60.035 175.480 60.325 175.525 ;
        RECT 60.955 175.480 61.245 175.525 ;
        RECT 59.560 175.340 61.245 175.480 ;
        RECT 56.890 175.140 57.030 175.295 ;
        RECT 59.560 175.280 59.880 175.340 ;
        RECT 60.035 175.295 60.325 175.340 ;
        RECT 60.955 175.295 61.245 175.340 ;
        RECT 61.875 175.295 62.165 175.525 ;
        RECT 57.260 175.140 57.580 175.200 ;
        RECT 56.890 175.000 57.580 175.140 ;
        RECT 57.260 174.940 57.580 175.000 ;
        RECT 60.480 175.140 60.800 175.200 ;
        RECT 61.950 175.140 62.090 175.295 ;
        RECT 64.160 175.280 64.480 175.540 ;
        RECT 64.620 175.280 64.940 175.540 ;
        RECT 65.095 175.295 65.385 175.525 ;
        RECT 66.015 175.480 66.305 175.525 ;
        RECT 66.920 175.480 67.240 175.540 ;
        RECT 68.160 175.480 68.300 175.680 ;
        RECT 71.060 175.620 71.380 175.680 ;
        RECT 72.610 175.820 72.900 175.865 ;
        RECT 78.510 175.820 78.650 175.975 ;
        RECT 78.880 175.960 79.200 176.020 ;
        RECT 72.610 175.680 78.650 175.820 ;
        RECT 72.610 175.635 72.900 175.680 ;
        RECT 66.015 175.340 67.240 175.480 ;
        RECT 66.015 175.295 66.305 175.340 ;
        RECT 60.480 175.000 62.090 175.140 ;
        RECT 62.780 175.140 63.100 175.200 ;
        RECT 65.170 175.140 65.310 175.295 ;
        RECT 66.920 175.280 67.240 175.340 ;
        RECT 67.470 175.340 68.300 175.480 ;
        RECT 70.140 175.480 70.460 175.540 ;
        RECT 73.835 175.480 74.125 175.525 ;
        RECT 74.740 175.480 75.060 175.540 ;
        RECT 79.355 175.480 79.645 175.525 ;
        RECT 70.140 175.340 73.590 175.480 ;
        RECT 67.470 175.140 67.610 175.340 ;
        RECT 70.140 175.280 70.460 175.340 ;
        RECT 62.780 175.000 67.610 175.140 ;
        RECT 69.245 175.140 69.535 175.185 ;
        RECT 71.765 175.140 72.055 175.185 ;
        RECT 72.955 175.140 73.245 175.185 ;
        RECT 69.245 175.000 73.245 175.140 ;
        RECT 73.450 175.140 73.590 175.340 ;
        RECT 73.835 175.340 75.060 175.480 ;
        RECT 73.835 175.295 74.125 175.340 ;
        RECT 74.740 175.280 75.060 175.340 ;
        RECT 75.290 175.340 79.645 175.480 ;
        RECT 75.290 175.140 75.430 175.340 ;
        RECT 79.355 175.295 79.645 175.340 ;
        RECT 79.815 175.295 80.105 175.525 ;
        RECT 80.275 175.480 80.565 175.525 ;
        RECT 80.720 175.480 81.040 175.540 ;
        RECT 81.270 175.525 81.410 176.020 ;
        RECT 83.570 176.020 85.640 176.160 ;
        RECT 83.570 175.525 83.710 176.020 ;
        RECT 85.320 175.960 85.640 176.020 ;
        RECT 90.395 175.975 90.685 176.205 ;
        RECT 93.155 176.160 93.445 176.205 ;
        RECT 95.455 176.160 95.745 176.205 ;
        RECT 93.155 176.020 95.745 176.160 ;
        RECT 93.155 175.975 93.445 176.020 ;
        RECT 95.455 175.975 95.745 176.020 ;
        RECT 84.415 175.820 84.705 175.865 ;
        RECT 86.255 175.820 86.545 175.865 ;
        RECT 84.415 175.680 86.545 175.820 ;
        RECT 84.415 175.635 84.705 175.680 ;
        RECT 86.255 175.635 86.545 175.680 ;
        RECT 88.540 175.620 88.860 175.880 ;
        RECT 89.580 175.820 89.870 175.865 ;
        RECT 90.470 175.820 90.610 175.975 ;
        RECT 95.900 175.960 96.220 176.220 ;
        RECT 96.360 175.960 96.680 176.220 ;
        RECT 97.280 175.960 97.600 176.220 ;
        RECT 101.420 176.205 101.740 176.220 ;
        RECT 101.400 176.160 101.740 176.205 ;
        RECT 101.225 176.020 101.740 176.160 ;
        RECT 101.400 175.975 101.740 176.020 ;
        RECT 101.420 175.960 101.740 175.975 ;
        RECT 102.800 175.960 103.120 176.220 ;
        RECT 106.020 175.960 106.340 176.220 ;
        RECT 106.480 175.960 106.800 176.220 ;
        RECT 106.940 175.960 107.260 176.220 ;
        RECT 110.175 176.160 110.465 176.205 ;
        RECT 108.410 176.020 110.465 176.160 ;
        RECT 95.990 175.820 96.130 175.960 ;
        RECT 89.580 175.680 90.150 175.820 ;
        RECT 90.470 175.680 96.130 175.820 ;
        RECT 96.450 175.820 96.590 175.960 ;
        RECT 101.895 175.820 102.185 175.865 ;
        RECT 106.570 175.820 106.710 175.960 ;
        RECT 96.450 175.680 100.730 175.820 ;
        RECT 89.580 175.635 89.870 175.680 ;
        RECT 80.275 175.340 81.040 175.480 ;
        RECT 80.275 175.295 80.565 175.340 ;
        RECT 77.515 175.140 77.805 175.185 ;
        RECT 73.450 175.000 75.430 175.140 ;
        RECT 76.670 175.000 77.805 175.140 ;
        RECT 60.480 174.940 60.800 175.000 ;
        RECT 62.780 174.940 63.100 175.000 ;
        RECT 69.245 174.955 69.535 175.000 ;
        RECT 71.765 174.955 72.055 175.000 ;
        RECT 72.955 174.955 73.245 175.000 ;
        RECT 59.560 174.800 59.880 174.860 ;
        RECT 61.415 174.800 61.705 174.845 ;
        RECT 56.430 174.660 58.410 174.800 ;
        RECT 58.270 174.520 58.410 174.660 ;
        RECT 59.560 174.660 61.705 174.800 ;
        RECT 59.560 174.600 59.880 174.660 ;
        RECT 61.415 174.615 61.705 174.660 ;
        RECT 69.680 174.800 69.970 174.845 ;
        RECT 71.250 174.800 71.540 174.845 ;
        RECT 73.350 174.800 73.640 174.845 ;
        RECT 69.680 174.660 73.640 174.800 ;
        RECT 69.680 174.615 69.970 174.660 ;
        RECT 71.250 174.615 71.540 174.660 ;
        RECT 73.350 174.615 73.640 174.660 ;
        RECT 76.670 174.520 76.810 175.000 ;
        RECT 77.515 174.955 77.805 175.000 ;
        RECT 79.890 174.800 80.030 175.295 ;
        RECT 80.720 175.280 81.040 175.340 ;
        RECT 81.195 175.295 81.485 175.525 ;
        RECT 83.495 175.295 83.785 175.525 ;
        RECT 83.955 175.295 84.245 175.525 ;
        RECT 84.875 175.480 85.165 175.525 ;
        RECT 89.000 175.480 89.320 175.540 ;
        RECT 84.875 175.340 89.320 175.480 ;
        RECT 84.875 175.295 85.165 175.340 ;
        RECT 83.035 175.140 83.325 175.185 ;
        RECT 84.030 175.140 84.170 175.295 ;
        RECT 89.000 175.280 89.320 175.340 ;
        RECT 90.010 175.140 90.150 175.680 ;
        RECT 90.855 175.480 91.145 175.525 ;
        RECT 90.855 175.340 94.750 175.480 ;
        RECT 90.855 175.295 91.145 175.340 ;
        RECT 91.300 175.140 91.620 175.200 ;
        RECT 83.035 175.000 86.010 175.140 ;
        RECT 90.010 175.000 91.620 175.140 ;
        RECT 83.035 174.955 83.325 175.000 ;
        RECT 83.940 174.800 84.260 174.860 ;
        RECT 79.890 174.660 84.260 174.800 ;
        RECT 83.940 174.600 84.260 174.660 ;
        RECT 85.870 174.520 86.010 175.000 ;
        RECT 91.300 174.940 91.620 175.000 ;
        RECT 93.600 174.940 93.920 175.200 ;
        RECT 94.610 175.140 94.750 175.340 ;
        RECT 94.980 175.280 95.300 175.540 ;
        RECT 95.915 175.480 96.205 175.525 ;
        RECT 96.820 175.480 97.140 175.540 ;
        RECT 95.915 175.340 97.140 175.480 ;
        RECT 95.915 175.295 96.205 175.340 ;
        RECT 96.820 175.280 97.140 175.340 ;
        RECT 97.740 175.280 98.060 175.540 ;
        RECT 100.590 175.525 100.730 175.680 ;
        RECT 101.895 175.680 106.710 175.820 ;
        RECT 107.030 175.820 107.170 175.960 ;
        RECT 108.410 175.820 108.550 176.020 ;
        RECT 110.175 175.975 110.465 176.020 ;
        RECT 111.095 175.975 111.385 176.205 ;
        RECT 112.460 176.160 112.780 176.220 ;
        RECT 114.315 176.160 114.605 176.205 ;
        RECT 112.460 176.020 114.605 176.160 ;
        RECT 107.030 175.680 108.550 175.820 ;
        RECT 111.170 175.820 111.310 175.975 ;
        RECT 112.460 175.960 112.780 176.020 ;
        RECT 114.315 175.975 114.605 176.020 ;
        RECT 133.160 175.960 133.480 176.220 ;
        RECT 134.540 176.160 134.860 176.220 ;
        RECT 135.015 176.160 135.305 176.205 ;
        RECT 134.540 176.020 135.305 176.160 ;
        RECT 134.540 175.960 134.860 176.020 ;
        RECT 135.015 175.975 135.305 176.020 ;
        RECT 116.600 175.820 116.920 175.880 ;
        RECT 111.170 175.680 116.920 175.820 ;
        RECT 101.895 175.635 102.185 175.680 ;
        RECT 100.515 175.295 100.805 175.525 ;
        RECT 100.975 175.480 101.265 175.525 ;
        RECT 100.975 175.340 102.110 175.480 ;
        RECT 100.975 175.295 101.265 175.340 ;
        RECT 101.970 175.200 102.110 175.340 ;
        RECT 103.720 175.280 104.040 175.540 ;
        RECT 104.195 175.295 104.485 175.525 ;
        RECT 97.280 175.140 97.600 175.200 ;
        RECT 94.610 175.000 97.600 175.140 ;
        RECT 97.280 174.940 97.600 175.000 ;
        RECT 101.880 174.940 102.200 175.200 ;
        RECT 88.095 174.800 88.385 174.845 ;
        RECT 92.220 174.800 92.540 174.860 ;
        RECT 88.095 174.660 92.540 174.800 ;
        RECT 88.095 174.615 88.385 174.660 ;
        RECT 92.220 174.600 92.540 174.660 ;
        RECT 92.695 174.615 92.985 174.845 ;
        RECT 94.075 174.800 94.365 174.845 ;
        RECT 98.215 174.800 98.505 174.845 ;
        RECT 94.075 174.660 98.505 174.800 ;
        RECT 103.810 174.800 103.950 175.280 ;
        RECT 104.270 175.140 104.410 175.295 ;
        RECT 104.640 175.280 104.960 175.540 ;
        RECT 105.100 175.480 105.420 175.540 ;
        RECT 105.575 175.480 105.865 175.525 ;
        RECT 105.100 175.340 105.865 175.480 ;
        RECT 105.100 175.280 105.420 175.340 ;
        RECT 105.575 175.295 105.865 175.340 ;
        RECT 107.400 175.280 107.720 175.540 ;
        RECT 108.410 175.525 108.550 175.680 ;
        RECT 116.600 175.620 116.920 175.680 ;
        RECT 107.875 175.295 108.165 175.525 ;
        RECT 108.335 175.295 108.625 175.525 ;
        RECT 109.255 175.295 109.545 175.525 ;
        RECT 111.080 175.480 111.370 175.525 ;
        RECT 111.540 175.480 111.860 175.540 ;
        RECT 111.080 175.340 111.860 175.480 ;
        RECT 111.080 175.295 111.370 175.340 ;
        RECT 107.490 175.140 107.630 175.280 ;
        RECT 104.270 175.000 107.630 175.140 ;
        RECT 107.950 174.800 108.090 175.295 ;
        RECT 109.330 175.140 109.470 175.295 ;
        RECT 111.540 175.280 111.860 175.340 ;
        RECT 112.000 175.480 112.320 175.540 ;
        RECT 112.935 175.480 113.225 175.525 ;
        RECT 113.840 175.480 114.160 175.540 ;
        RECT 112.000 175.340 114.160 175.480 ;
        RECT 112.000 175.280 112.320 175.340 ;
        RECT 112.935 175.295 113.225 175.340 ;
        RECT 113.840 175.280 114.160 175.340 ;
        RECT 118.455 175.480 118.745 175.525 ;
        RECT 118.900 175.480 119.220 175.540 ;
        RECT 119.820 175.525 120.140 175.540 ;
        RECT 118.455 175.340 119.220 175.480 ;
        RECT 118.455 175.295 118.745 175.340 ;
        RECT 118.900 175.280 119.220 175.340 ;
        RECT 119.790 175.295 120.140 175.525 ;
        RECT 119.820 175.280 120.140 175.295 ;
        RECT 128.100 175.480 128.420 175.540 ;
        RECT 129.955 175.480 130.245 175.525 ;
        RECT 128.100 175.340 130.245 175.480 ;
        RECT 128.100 175.280 128.420 175.340 ;
        RECT 129.955 175.295 130.245 175.340 ;
        RECT 132.715 175.480 133.005 175.525 ;
        RECT 133.250 175.480 133.390 175.960 ;
        RECT 132.715 175.340 133.390 175.480 ;
        RECT 135.090 175.480 135.230 175.975 ;
        RECT 137.300 175.960 137.620 176.220 ;
        RECT 138.220 175.960 138.540 176.220 ;
        RECT 139.580 176.160 139.870 176.205 ;
        RECT 141.440 176.160 141.760 176.220 ;
        RECT 139.580 176.020 141.760 176.160 ;
        RECT 139.580 175.975 139.870 176.020 ;
        RECT 141.440 175.960 141.760 176.020 ;
        RECT 144.200 176.160 144.520 176.220 ;
        RECT 146.960 176.160 147.280 176.220 ;
        RECT 147.435 176.160 147.725 176.205 ;
        RECT 144.200 176.020 145.350 176.160 ;
        RECT 144.200 175.960 144.520 176.020 ;
        RECT 135.475 175.480 135.765 175.525 ;
        RECT 135.090 175.340 135.765 175.480 ;
        RECT 132.715 175.295 133.005 175.340 ;
        RECT 135.475 175.295 135.765 175.340 ;
        RECT 135.935 175.295 136.225 175.525 ;
        RECT 136.380 175.480 136.700 175.540 ;
        RECT 136.855 175.480 137.145 175.525 ;
        RECT 136.380 175.340 137.145 175.480 ;
        RECT 109.330 175.000 112.230 175.140 ;
        RECT 103.810 174.660 108.090 174.800 ;
        RECT 94.075 174.615 94.365 174.660 ;
        RECT 98.215 174.615 98.505 174.660 ;
        RECT 56.800 174.460 57.120 174.520 ;
        RECT 57.275 174.460 57.565 174.505 ;
        RECT 55.950 174.320 57.565 174.460 ;
        RECT 56.800 174.260 57.120 174.320 ;
        RECT 57.275 174.275 57.565 174.320 ;
        RECT 58.180 174.460 58.500 174.520 ;
        RECT 76.580 174.460 76.900 174.520 ;
        RECT 58.180 174.320 76.900 174.460 ;
        RECT 58.180 174.260 58.500 174.320 ;
        RECT 76.580 174.260 76.900 174.320 ;
        RECT 85.320 174.260 85.640 174.520 ;
        RECT 85.780 174.260 86.100 174.520 ;
        RECT 86.255 174.460 86.545 174.505 ;
        RECT 87.160 174.460 87.480 174.520 ;
        RECT 86.255 174.320 87.480 174.460 ;
        RECT 86.255 174.275 86.545 174.320 ;
        RECT 87.160 174.260 87.480 174.320 ;
        RECT 89.475 174.460 89.765 174.505 ;
        RECT 90.840 174.460 91.160 174.520 ;
        RECT 89.475 174.320 91.160 174.460 ;
        RECT 92.770 174.460 92.910 174.615 ;
        RECT 112.090 174.520 112.230 175.000 ;
        RECT 113.380 174.940 113.700 175.200 ;
        RECT 119.335 175.140 119.625 175.185 ;
        RECT 120.525 175.140 120.815 175.185 ;
        RECT 123.045 175.140 123.335 175.185 ;
        RECT 119.335 175.000 123.335 175.140 ;
        RECT 119.335 174.955 119.625 175.000 ;
        RECT 120.525 174.955 120.815 175.000 ;
        RECT 123.045 174.955 123.335 175.000 ;
        RECT 129.035 175.140 129.325 175.185 ;
        RECT 132.255 175.140 132.545 175.185 ;
        RECT 134.080 175.140 134.400 175.200 ;
        RECT 136.010 175.140 136.150 175.295 ;
        RECT 136.380 175.280 136.700 175.340 ;
        RECT 136.855 175.295 137.145 175.340 ;
        RECT 129.035 175.000 129.435 175.140 ;
        RECT 132.255 175.000 136.150 175.140 ;
        RECT 129.035 174.955 129.325 175.000 ;
        RECT 132.255 174.955 132.545 175.000 ;
        RECT 115.235 174.800 115.525 174.845 ;
        RECT 118.440 174.800 118.760 174.860 ;
        RECT 115.235 174.660 118.760 174.800 ;
        RECT 115.235 174.615 115.525 174.660 ;
        RECT 118.440 174.600 118.760 174.660 ;
        RECT 118.940 174.800 119.230 174.845 ;
        RECT 121.040 174.800 121.330 174.845 ;
        RECT 122.610 174.800 122.900 174.845 ;
        RECT 118.940 174.660 122.900 174.800 ;
        RECT 118.940 174.615 119.230 174.660 ;
        RECT 121.040 174.615 121.330 174.660 ;
        RECT 122.610 174.615 122.900 174.660 ;
        RECT 125.355 174.800 125.645 174.845 ;
        RECT 129.110 174.800 129.250 174.955 ;
        RECT 134.080 174.940 134.400 175.000 ;
        RECT 125.355 174.660 134.310 174.800 ;
        RECT 125.355 174.615 125.645 174.660 ;
        RECT 95.900 174.460 96.220 174.520 ;
        RECT 92.770 174.320 96.220 174.460 ;
        RECT 89.475 174.275 89.765 174.320 ;
        RECT 90.840 174.260 91.160 174.320 ;
        RECT 95.900 174.260 96.220 174.320 ;
        RECT 112.000 174.260 112.320 174.520 ;
        RECT 126.260 174.260 126.580 174.520 ;
        RECT 129.940 174.460 130.260 174.520 ;
        RECT 134.170 174.505 134.310 174.660 ;
        RECT 130.415 174.460 130.705 174.505 ;
        RECT 129.940 174.320 130.705 174.460 ;
        RECT 129.940 174.260 130.260 174.320 ;
        RECT 130.415 174.275 130.705 174.320 ;
        RECT 134.095 174.460 134.385 174.505 ;
        RECT 137.390 174.460 137.530 175.960 ;
        RECT 138.310 175.480 138.450 175.960 ;
        RECT 139.155 175.820 139.445 175.865 ;
        RECT 143.740 175.820 144.060 175.880 ;
        RECT 139.155 175.680 144.060 175.820 ;
        RECT 139.155 175.635 139.445 175.680 ;
        RECT 143.740 175.620 144.060 175.680 ;
        RECT 144.675 175.635 144.965 175.865 ;
        RECT 145.210 175.820 145.350 176.020 ;
        RECT 146.960 176.020 147.725 176.160 ;
        RECT 146.960 175.960 147.280 176.020 ;
        RECT 147.435 175.975 147.725 176.020 ;
        RECT 152.020 175.960 152.340 176.220 ;
        RECT 154.780 175.960 155.100 176.220 ;
        RECT 145.675 175.820 145.965 175.865 ;
        RECT 154.870 175.820 155.010 175.960 ;
        RECT 145.210 175.680 145.965 175.820 ;
        RECT 145.675 175.635 145.965 175.680 ;
        RECT 146.130 175.680 155.010 175.820 ;
        RECT 138.695 175.480 138.985 175.525 ;
        RECT 138.310 175.340 138.985 175.480 ;
        RECT 138.695 175.295 138.985 175.340 ;
        RECT 140.075 175.480 140.365 175.525 ;
        RECT 143.295 175.480 143.585 175.525 ;
        RECT 144.750 175.480 144.890 175.635 ;
        RECT 146.130 175.480 146.270 175.680 ;
        RECT 140.075 175.340 143.050 175.480 ;
        RECT 140.075 175.295 140.365 175.340 ;
        RECT 137.775 175.140 138.065 175.185 ;
        RECT 141.900 175.140 142.220 175.200 ;
        RECT 137.775 175.000 142.220 175.140 ;
        RECT 142.910 175.140 143.050 175.340 ;
        RECT 143.295 175.340 146.270 175.480 ;
        RECT 147.895 175.480 148.185 175.525 ;
        RECT 149.735 175.480 150.025 175.525 ;
        RECT 147.895 175.340 150.025 175.480 ;
        RECT 143.295 175.295 143.585 175.340 ;
        RECT 147.895 175.295 148.185 175.340 ;
        RECT 149.735 175.295 150.025 175.340 ;
        RECT 150.655 175.480 150.945 175.525 ;
        RECT 151.100 175.480 151.420 175.540 ;
        RECT 154.870 175.525 155.010 175.680 ;
        RECT 150.655 175.340 151.420 175.480 ;
        RECT 150.655 175.295 150.945 175.340 ;
        RECT 145.120 175.140 145.440 175.200 ;
        RECT 142.910 175.000 145.440 175.140 ;
        RECT 137.775 174.955 138.065 175.000 ;
        RECT 141.900 174.940 142.220 175.000 ;
        RECT 145.120 174.940 145.440 175.000 ;
        RECT 146.515 174.800 146.805 174.845 ;
        RECT 147.970 174.800 148.110 175.295 ;
        RECT 149.810 175.140 149.950 175.295 ;
        RECT 151.100 175.280 151.420 175.340 ;
        RECT 154.795 175.295 155.085 175.525 ;
        RECT 149.810 175.000 152.250 175.140 ;
        RECT 146.515 174.660 148.110 174.800 ;
        RECT 146.515 174.615 146.805 174.660 ;
        RECT 152.110 174.520 152.250 175.000 ;
        RECT 134.095 174.320 137.530 174.460 ;
        RECT 134.095 174.275 134.385 174.320 ;
        RECT 142.820 174.260 143.140 174.520 ;
        RECT 145.595 174.460 145.885 174.505 ;
        RECT 149.720 174.460 150.040 174.520 ;
        RECT 145.595 174.320 150.040 174.460 ;
        RECT 145.595 174.275 145.885 174.320 ;
        RECT 149.720 174.260 150.040 174.320 ;
        RECT 150.180 174.260 150.500 174.520 ;
        RECT 152.020 174.260 152.340 174.520 ;
        RECT 22.690 173.640 157.010 174.120 ;
        RECT 31.055 173.440 31.345 173.485 ;
        RECT 35.180 173.440 35.500 173.500 ;
        RECT 31.055 173.300 35.500 173.440 ;
        RECT 31.055 173.255 31.345 173.300 ;
        RECT 35.180 173.240 35.500 173.300 ;
        RECT 37.480 173.240 37.800 173.500 ;
        RECT 45.775 173.440 46.065 173.485 ;
        RECT 46.220 173.440 46.540 173.500 ;
        RECT 45.775 173.300 46.540 173.440 ;
        RECT 45.775 173.255 46.065 173.300 ;
        RECT 24.640 173.100 24.930 173.145 ;
        RECT 26.740 173.100 27.030 173.145 ;
        RECT 28.310 173.100 28.600 173.145 ;
        RECT 24.640 172.960 28.600 173.100 ;
        RECT 24.640 172.915 24.930 172.960 ;
        RECT 26.740 172.915 27.030 172.960 ;
        RECT 28.310 172.915 28.600 172.960 ;
        RECT 43.460 173.100 43.780 173.160 ;
        RECT 45.315 173.100 45.605 173.145 ;
        RECT 43.460 172.960 45.605 173.100 ;
        RECT 43.460 172.900 43.780 172.960 ;
        RECT 45.315 172.915 45.605 172.960 ;
        RECT 25.035 172.760 25.325 172.805 ;
        RECT 26.225 172.760 26.515 172.805 ;
        RECT 28.745 172.760 29.035 172.805 ;
        RECT 25.035 172.620 29.035 172.760 ;
        RECT 25.035 172.575 25.325 172.620 ;
        RECT 26.225 172.575 26.515 172.620 ;
        RECT 28.745 172.575 29.035 172.620 ;
        RECT 24.140 172.220 24.460 172.480 ;
        RECT 25.520 172.465 25.840 172.480 ;
        RECT 25.490 172.420 25.840 172.465 ;
        RECT 25.325 172.280 25.840 172.420 ;
        RECT 25.490 172.235 25.840 172.280 ;
        RECT 25.520 172.220 25.840 172.235 ;
        RECT 36.560 172.220 36.880 172.480 ;
        RECT 37.940 172.220 38.260 172.480 ;
        RECT 43.475 172.420 43.765 172.465 ;
        RECT 45.850 172.420 45.990 173.255 ;
        RECT 46.220 173.240 46.540 173.300 ;
        RECT 52.200 173.240 52.520 173.500 ;
        RECT 52.660 173.440 52.980 173.500 ;
        RECT 54.500 173.440 54.820 173.500 ;
        RECT 52.660 173.300 54.820 173.440 ;
        RECT 52.660 173.240 52.980 173.300 ;
        RECT 54.500 173.240 54.820 173.300 ;
        RECT 60.480 173.240 60.800 173.500 ;
        RECT 69.220 173.240 69.540 173.500 ;
        RECT 71.060 173.440 71.380 173.500 ;
        RECT 71.060 173.300 76.350 173.440 ;
        RECT 71.060 173.240 71.380 173.300 ;
        RECT 43.475 172.280 45.990 172.420 ;
        RECT 47.600 172.465 47.920 172.480 ;
        RECT 47.600 172.420 47.930 172.465 ;
        RECT 47.600 172.280 48.115 172.420 ;
        RECT 43.475 172.235 43.765 172.280 ;
        RECT 47.600 172.235 47.930 172.280 ;
        RECT 47.600 172.220 47.920 172.235 ;
        RECT 33.340 171.880 33.660 172.140 ;
        RECT 34.275 172.080 34.565 172.125 ;
        RECT 38.030 172.080 38.170 172.220 ;
        RECT 34.275 171.940 38.170 172.080 ;
        RECT 43.935 172.080 44.225 172.125 ;
        RECT 43.935 171.940 45.070 172.080 ;
        RECT 34.275 171.895 34.565 171.940 ;
        RECT 43.935 171.895 44.225 171.940 ;
        RECT 44.930 171.800 45.070 171.940 ;
        RECT 45.760 171.880 46.080 172.140 ;
        RECT 46.680 171.880 47.000 172.140 ;
        RECT 47.155 171.895 47.445 172.125 ;
        RECT 52.290 172.080 52.430 173.240 ;
        RECT 57.720 173.100 58.040 173.160 ;
        RECT 58.195 173.100 58.485 173.145 ;
        RECT 57.720 172.960 58.485 173.100 ;
        RECT 57.720 172.900 58.040 172.960 ;
        RECT 58.195 172.915 58.485 172.960 ;
        RECT 61.030 172.960 68.530 173.100 ;
        RECT 56.430 172.620 59.790 172.760 ;
        RECT 56.430 172.465 56.570 172.620 ;
        RECT 59.650 172.480 59.790 172.620 ;
        RECT 61.030 172.480 61.170 172.960 ;
        RECT 68.390 172.805 68.530 172.960 ;
        RECT 65.555 172.760 65.845 172.805 ;
        RECT 62.410 172.620 65.845 172.760 ;
        RECT 56.355 172.235 56.645 172.465 ;
        RECT 56.800 172.220 57.120 172.480 ;
        RECT 57.720 172.420 58.040 172.480 ;
        RECT 58.655 172.420 58.945 172.465 ;
        RECT 57.720 172.280 58.945 172.420 ;
        RECT 57.720 172.220 58.040 172.280 ;
        RECT 58.655 172.235 58.945 172.280 ;
        RECT 59.100 172.220 59.420 172.480 ;
        RECT 59.560 172.220 59.880 172.480 ;
        RECT 60.940 172.220 61.260 172.480 ;
        RECT 62.410 172.465 62.550 172.620 ;
        RECT 65.555 172.575 65.845 172.620 ;
        RECT 68.315 172.575 68.605 172.805 ;
        RECT 62.335 172.235 62.625 172.465 ;
        RECT 62.780 172.420 63.100 172.480 ;
        RECT 63.255 172.420 63.545 172.465 ;
        RECT 62.780 172.280 63.545 172.420 ;
        RECT 62.780 172.220 63.100 172.280 ;
        RECT 63.255 172.235 63.545 172.280 ;
        RECT 64.160 172.220 64.480 172.480 ;
        RECT 57.275 172.080 57.565 172.125 ;
        RECT 59.190 172.080 59.330 172.220 ;
        RECT 52.290 171.940 56.110 172.080 ;
        RECT 35.180 171.540 35.500 171.800 ;
        RECT 37.480 171.740 37.800 171.800 ;
        RECT 42.555 171.740 42.845 171.785 ;
        RECT 37.480 171.600 42.845 171.740 ;
        RECT 37.480 171.540 37.800 171.600 ;
        RECT 42.555 171.555 42.845 171.600 ;
        RECT 44.380 171.540 44.700 171.800 ;
        RECT 44.840 171.540 45.160 171.800 ;
        RECT 46.220 171.740 46.540 171.800 ;
        RECT 47.230 171.740 47.370 171.895 ;
        RECT 46.220 171.600 47.370 171.740 ;
        RECT 54.960 171.740 55.280 171.800 ;
        RECT 55.435 171.740 55.725 171.785 ;
        RECT 54.960 171.600 55.725 171.740 ;
        RECT 55.970 171.740 56.110 171.940 ;
        RECT 57.275 171.940 59.330 172.080 ;
        RECT 63.715 172.080 64.005 172.125 ;
        RECT 66.460 172.080 66.780 172.140 ;
        RECT 63.715 171.940 66.780 172.080 ;
        RECT 69.310 172.080 69.450 173.240 ;
        RECT 70.180 173.100 70.470 173.145 ;
        RECT 72.280 173.100 72.570 173.145 ;
        RECT 73.850 173.100 74.140 173.145 ;
        RECT 70.180 172.960 74.140 173.100 ;
        RECT 76.210 173.100 76.350 173.300 ;
        RECT 76.580 173.240 76.900 173.500 ;
        RECT 80.720 173.440 81.040 173.500 ;
        RECT 77.130 173.300 81.040 173.440 ;
        RECT 77.130 173.100 77.270 173.300 ;
        RECT 80.720 173.240 81.040 173.300 ;
        RECT 84.400 173.240 84.720 173.500 ;
        RECT 85.320 173.240 85.640 173.500 ;
        RECT 92.220 173.240 92.540 173.500 ;
        RECT 94.075 173.440 94.365 173.485 ;
        RECT 97.740 173.440 98.060 173.500 ;
        RECT 94.075 173.300 98.060 173.440 ;
        RECT 94.075 173.255 94.365 173.300 ;
        RECT 76.210 172.960 77.270 173.100 ;
        RECT 77.540 173.100 77.830 173.145 ;
        RECT 79.640 173.100 79.930 173.145 ;
        RECT 81.210 173.100 81.500 173.145 ;
        RECT 77.540 172.960 81.500 173.100 ;
        RECT 70.180 172.915 70.470 172.960 ;
        RECT 72.280 172.915 72.570 172.960 ;
        RECT 73.850 172.915 74.140 172.960 ;
        RECT 77.540 172.915 77.830 172.960 ;
        RECT 79.640 172.915 79.930 172.960 ;
        RECT 81.210 172.915 81.500 172.960 ;
        RECT 70.575 172.760 70.865 172.805 ;
        RECT 71.765 172.760 72.055 172.805 ;
        RECT 74.285 172.760 74.575 172.805 ;
        RECT 70.575 172.620 74.575 172.760 ;
        RECT 70.575 172.575 70.865 172.620 ;
        RECT 71.765 172.575 72.055 172.620 ;
        RECT 74.285 172.575 74.575 172.620 ;
        RECT 77.935 172.760 78.225 172.805 ;
        RECT 79.125 172.760 79.415 172.805 ;
        RECT 81.645 172.760 81.935 172.805 ;
        RECT 77.935 172.620 81.935 172.760 ;
        RECT 77.935 172.575 78.225 172.620 ;
        RECT 79.125 172.575 79.415 172.620 ;
        RECT 81.645 172.575 81.935 172.620 ;
        RECT 69.695 172.420 69.985 172.465 ;
        RECT 75.200 172.420 75.520 172.480 ;
        RECT 85.410 172.465 85.550 173.240 ;
        RECT 89.000 173.100 89.320 173.160 ;
        RECT 89.000 172.960 92.450 173.100 ;
        RECT 89.000 172.900 89.320 172.960 ;
        RECT 85.780 172.760 86.100 172.820 ;
        RECT 85.780 172.620 91.530 172.760 ;
        RECT 85.780 172.560 86.100 172.620 ;
        RECT 91.390 172.465 91.530 172.620 ;
        RECT 92.310 172.465 92.450 172.960 ;
        RECT 93.600 172.900 93.920 173.160 ;
        RECT 93.690 172.465 93.830 172.900 ;
        RECT 77.055 172.420 77.345 172.465 ;
        RECT 69.695 172.280 77.345 172.420 ;
        RECT 69.695 172.235 69.985 172.280 ;
        RECT 75.200 172.220 75.520 172.280 ;
        RECT 77.055 172.235 77.345 172.280 ;
        RECT 85.335 172.235 85.625 172.465 ;
        RECT 90.395 172.235 90.685 172.465 ;
        RECT 91.315 172.235 91.605 172.465 ;
        RECT 92.235 172.235 92.525 172.465 ;
        RECT 93.615 172.235 93.905 172.465 ;
        RECT 70.920 172.080 71.210 172.125 ;
        RECT 69.310 171.940 71.210 172.080 ;
        RECT 57.275 171.895 57.565 171.940 ;
        RECT 63.715 171.895 64.005 171.940 ;
        RECT 66.460 171.880 66.780 171.940 ;
        RECT 70.920 171.895 71.210 171.940 ;
        RECT 78.390 172.080 78.680 172.125 ;
        RECT 79.340 172.080 79.660 172.140 ;
        RECT 90.470 172.080 90.610 172.235 ;
        RECT 94.150 172.080 94.290 173.255 ;
        RECT 97.740 173.240 98.060 173.300 ;
        RECT 98.675 173.440 98.965 173.485 ;
        RECT 99.120 173.440 99.440 173.500 ;
        RECT 98.675 173.300 99.440 173.440 ;
        RECT 98.675 173.255 98.965 173.300 ;
        RECT 99.120 173.240 99.440 173.300 ;
        RECT 112.000 173.440 112.320 173.500 ;
        RECT 114.775 173.440 115.065 173.485 ;
        RECT 112.000 173.300 115.065 173.440 ;
        RECT 112.000 173.240 112.320 173.300 ;
        RECT 114.775 173.255 115.065 173.300 ;
        RECT 119.820 173.240 120.140 173.500 ;
        RECT 121.660 173.240 121.980 173.500 ;
        RECT 126.260 173.240 126.580 173.500 ;
        RECT 142.835 173.440 143.125 173.485 ;
        RECT 143.740 173.440 144.060 173.500 ;
        RECT 142.835 173.300 144.060 173.440 ;
        RECT 142.835 173.255 143.125 173.300 ;
        RECT 143.740 173.240 144.060 173.300 ;
        RECT 95.900 172.900 96.220 173.160 ;
        RECT 112.460 172.900 112.780 173.160 ;
        RECT 95.990 172.420 96.130 172.900 ;
        RECT 112.550 172.760 112.690 172.900 ;
        RECT 112.550 172.620 114.990 172.760 ;
        RECT 96.375 172.420 96.665 172.465 ;
        RECT 95.990 172.280 96.665 172.420 ;
        RECT 96.375 172.235 96.665 172.280 ;
        RECT 97.280 172.420 97.600 172.480 ;
        RECT 97.755 172.420 98.045 172.465 ;
        RECT 97.280 172.280 98.045 172.420 ;
        RECT 97.280 172.220 97.600 172.280 ;
        RECT 97.755 172.235 98.045 172.280 ;
        RECT 113.395 172.235 113.685 172.465 ;
        RECT 78.390 171.940 79.660 172.080 ;
        RECT 78.390 171.895 78.680 171.940 ;
        RECT 79.340 171.880 79.660 171.940 ;
        RECT 84.030 171.940 94.290 172.080 ;
        RECT 59.115 171.740 59.405 171.785 ;
        RECT 55.970 171.600 59.405 171.740 ;
        RECT 46.220 171.540 46.540 171.600 ;
        RECT 54.960 171.540 55.280 171.600 ;
        RECT 55.435 171.555 55.725 171.600 ;
        RECT 59.115 171.555 59.405 171.600 ;
        RECT 65.080 171.540 65.400 171.800 ;
        RECT 84.030 171.785 84.170 171.940 ;
        RECT 113.470 171.800 113.610 172.235 ;
        RECT 113.840 172.220 114.160 172.480 ;
        RECT 114.850 172.465 114.990 172.620 ;
        RECT 114.775 172.235 115.065 172.465 ;
        RECT 117.980 172.420 118.300 172.480 ;
        RECT 120.755 172.420 121.045 172.465 ;
        RECT 121.750 172.420 121.890 173.240 ;
        RECT 117.980 172.280 121.890 172.420 ;
        RECT 117.980 172.220 118.300 172.280 ;
        RECT 120.755 172.235 121.045 172.280 ;
        RECT 122.120 172.220 122.440 172.480 ;
        RECT 122.595 172.420 122.885 172.465 ;
        RECT 126.350 172.420 126.490 173.240 ;
        RECT 148.840 173.100 149.130 173.145 ;
        RECT 150.940 173.100 151.230 173.145 ;
        RECT 152.510 173.100 152.800 173.145 ;
        RECT 148.840 172.960 152.800 173.100 ;
        RECT 148.840 172.915 149.130 172.960 ;
        RECT 150.940 172.915 151.230 172.960 ;
        RECT 152.510 172.915 152.800 172.960 ;
        RECT 133.160 172.760 133.480 172.820 ;
        RECT 135.015 172.760 135.305 172.805 ;
        RECT 149.235 172.760 149.525 172.805 ;
        RECT 150.425 172.760 150.715 172.805 ;
        RECT 152.945 172.760 153.235 172.805 ;
        RECT 133.160 172.620 135.305 172.760 ;
        RECT 133.160 172.560 133.480 172.620 ;
        RECT 135.015 172.575 135.305 172.620 ;
        RECT 141.070 172.620 149.030 172.760 ;
        RECT 122.595 172.280 126.490 172.420 ;
        RECT 122.595 172.235 122.885 172.280 ;
        RECT 129.020 172.220 129.340 172.480 ;
        RECT 129.480 172.420 129.800 172.480 ;
        RECT 129.955 172.420 130.245 172.465 ;
        RECT 141.070 172.420 141.210 172.620 ;
        RECT 148.890 172.480 149.030 172.620 ;
        RECT 149.235 172.620 153.235 172.760 ;
        RECT 149.235 172.575 149.525 172.620 ;
        RECT 150.425 172.575 150.715 172.620 ;
        RECT 152.945 172.575 153.235 172.620 ;
        RECT 129.480 172.280 141.210 172.420 ;
        RECT 142.360 172.420 142.680 172.480 ;
        RECT 143.755 172.420 144.045 172.465 ;
        RECT 142.360 172.280 144.045 172.420 ;
        RECT 129.480 172.220 129.800 172.280 ;
        RECT 129.955 172.235 130.245 172.280 ;
        RECT 142.360 172.220 142.680 172.280 ;
        RECT 143.755 172.235 144.045 172.280 ;
        RECT 144.215 172.235 144.505 172.465 ;
        RECT 117.060 172.080 117.380 172.140 ;
        RECT 121.215 172.080 121.505 172.125 ;
        RECT 117.060 171.940 121.505 172.080 ;
        RECT 117.060 171.880 117.380 171.940 ;
        RECT 121.215 171.895 121.505 171.940 ;
        RECT 121.675 172.080 121.965 172.125 ;
        RECT 122.210 172.080 122.350 172.220 ;
        RECT 121.675 171.940 122.350 172.080 ;
        RECT 130.400 172.080 130.720 172.140 ;
        RECT 132.255 172.080 132.545 172.125 ;
        RECT 130.400 171.940 132.545 172.080 ;
        RECT 121.675 171.895 121.965 171.940 ;
        RECT 130.400 171.880 130.720 171.940 ;
        RECT 132.255 171.895 132.545 171.940 ;
        RECT 141.900 172.080 142.220 172.140 ;
        RECT 144.290 172.080 144.430 172.235 ;
        RECT 144.660 172.220 144.980 172.480 ;
        RECT 147.420 172.420 147.740 172.480 ;
        RECT 148.355 172.420 148.645 172.465 ;
        RECT 146.130 172.280 148.645 172.420 ;
        RECT 141.900 171.940 144.430 172.080 ;
        RECT 141.900 171.880 142.220 171.940 ;
        RECT 83.955 171.555 84.245 171.785 ;
        RECT 87.620 171.540 87.940 171.800 ;
        RECT 93.600 171.740 93.920 171.800 ;
        RECT 94.980 171.740 95.300 171.800 ;
        RECT 96.835 171.740 97.125 171.785 ;
        RECT 93.600 171.600 97.125 171.740 ;
        RECT 93.600 171.540 93.920 171.600 ;
        RECT 94.980 171.540 95.300 171.600 ;
        RECT 96.835 171.555 97.125 171.600 ;
        RECT 113.380 171.540 113.700 171.800 ;
        RECT 117.520 171.740 117.840 171.800 ;
        RECT 118.900 171.740 119.220 171.800 ;
        RECT 117.520 171.600 119.220 171.740 ;
        RECT 117.520 171.540 117.840 171.600 ;
        RECT 118.900 171.540 119.220 171.600 ;
        RECT 129.495 171.740 129.785 171.785 ;
        RECT 130.860 171.740 131.180 171.800 ;
        RECT 129.495 171.600 131.180 171.740 ;
        RECT 129.495 171.555 129.785 171.600 ;
        RECT 130.860 171.540 131.180 171.600 ;
        RECT 137.300 171.740 137.620 171.800 ;
        RECT 146.130 171.740 146.270 172.280 ;
        RECT 147.420 172.220 147.740 172.280 ;
        RECT 148.355 172.235 148.645 172.280 ;
        RECT 148.800 172.220 149.120 172.480 ;
        RECT 147.880 172.080 148.200 172.140 ;
        RECT 149.580 172.080 149.870 172.125 ;
        RECT 147.880 171.940 149.870 172.080 ;
        RECT 147.880 171.880 148.200 171.940 ;
        RECT 149.580 171.895 149.870 171.940 ;
        RECT 137.300 171.600 146.270 171.740 ;
        RECT 151.100 171.740 151.420 171.800 ;
        RECT 155.255 171.740 155.545 171.785 ;
        RECT 151.100 171.600 155.545 171.740 ;
        RECT 137.300 171.540 137.620 171.600 ;
        RECT 151.100 171.540 151.420 171.600 ;
        RECT 155.255 171.555 155.545 171.600 ;
        RECT 22.690 170.920 157.810 171.400 ;
        RECT 32.895 170.720 33.185 170.765 ;
        RECT 33.340 170.720 33.660 170.780 ;
        RECT 32.895 170.580 33.660 170.720 ;
        RECT 32.895 170.535 33.185 170.580 ;
        RECT 33.340 170.520 33.660 170.580 ;
        RECT 33.800 170.720 34.120 170.780 ;
        RECT 35.195 170.720 35.485 170.765 ;
        RECT 33.800 170.580 35.485 170.720 ;
        RECT 33.800 170.520 34.120 170.580 ;
        RECT 35.195 170.535 35.485 170.580 ;
        RECT 36.115 170.720 36.405 170.765 ;
        RECT 36.560 170.720 36.880 170.780 ;
        RECT 37.480 170.765 37.800 170.780 ;
        RECT 37.415 170.720 37.800 170.765 ;
        RECT 36.115 170.580 36.880 170.720 ;
        RECT 36.115 170.535 36.405 170.580 ;
        RECT 36.560 170.520 36.880 170.580 ;
        RECT 37.110 170.580 37.800 170.720 ;
        RECT 31.975 170.040 32.265 170.085 ;
        RECT 34.260 170.040 34.580 170.100 ;
        RECT 37.110 170.040 37.250 170.580 ;
        RECT 37.415 170.535 37.800 170.580 ;
        RECT 37.480 170.520 37.800 170.535 ;
        RECT 44.380 170.520 44.700 170.780 ;
        RECT 45.315 170.720 45.605 170.765 ;
        RECT 47.140 170.720 47.460 170.780 ;
        RECT 45.315 170.580 47.460 170.720 ;
        RECT 45.315 170.535 45.605 170.580 ;
        RECT 47.140 170.520 47.460 170.580 ;
        RECT 54.500 170.720 54.820 170.780 ;
        RECT 60.495 170.720 60.785 170.765 ;
        RECT 60.940 170.720 61.260 170.780 ;
        RECT 54.500 170.580 57.030 170.720 ;
        RECT 54.500 170.520 54.820 170.580 ;
        RECT 37.940 170.380 38.260 170.440 ;
        RECT 38.415 170.380 38.705 170.425 ;
        RECT 37.940 170.240 38.705 170.380 ;
        RECT 37.940 170.180 38.260 170.240 ;
        RECT 38.415 170.195 38.705 170.240 ;
        RECT 43.935 170.380 44.225 170.425 ;
        RECT 44.470 170.380 44.610 170.520 ;
        RECT 55.435 170.380 55.725 170.425 ;
        RECT 56.355 170.380 56.645 170.425 ;
        RECT 43.935 170.240 45.990 170.380 ;
        RECT 43.935 170.195 44.225 170.240 ;
        RECT 45.850 170.100 45.990 170.240 ;
        RECT 55.435 170.240 56.645 170.380 ;
        RECT 55.435 170.195 55.725 170.240 ;
        RECT 56.355 170.195 56.645 170.240 ;
        RECT 31.975 169.900 37.250 170.040 ;
        RECT 39.795 170.040 40.085 170.085 ;
        RECT 40.240 170.040 40.560 170.100 ;
        RECT 39.795 169.900 40.560 170.040 ;
        RECT 31.975 169.855 32.265 169.900 ;
        RECT 34.260 169.840 34.580 169.900 ;
        RECT 39.795 169.855 40.085 169.900 ;
        RECT 40.240 169.840 40.560 169.900 ;
        RECT 43.460 169.840 43.780 170.100 ;
        RECT 44.395 170.040 44.685 170.085 ;
        RECT 44.840 170.040 45.160 170.100 ;
        RECT 44.395 169.900 45.160 170.040 ;
        RECT 44.395 169.855 44.685 169.900 ;
        RECT 44.840 169.840 45.160 169.900 ;
        RECT 45.760 169.840 46.080 170.100 ;
        RECT 48.995 170.040 49.285 170.085 ;
        RECT 50.360 170.040 50.680 170.100 ;
        RECT 48.995 169.900 50.680 170.040 ;
        RECT 48.995 169.855 49.285 169.900 ;
        RECT 50.360 169.840 50.680 169.900 ;
        RECT 54.040 169.840 54.360 170.100 ;
        RECT 54.960 170.040 55.280 170.100 ;
        RECT 55.895 170.040 56.185 170.085 ;
        RECT 56.890 170.040 57.030 170.580 ;
        RECT 60.495 170.580 61.260 170.720 ;
        RECT 60.495 170.535 60.785 170.580 ;
        RECT 60.940 170.520 61.260 170.580 ;
        RECT 69.680 170.720 70.000 170.780 ;
        RECT 71.980 170.720 72.300 170.780 ;
        RECT 69.680 170.580 72.300 170.720 ;
        RECT 69.680 170.520 70.000 170.580 ;
        RECT 71.980 170.520 72.300 170.580 ;
        RECT 79.430 170.580 81.410 170.720 ;
        RECT 57.275 170.380 57.565 170.425 ;
        RECT 58.640 170.380 58.960 170.440 ;
        RECT 57.275 170.240 58.960 170.380 ;
        RECT 57.275 170.195 57.565 170.240 ;
        RECT 58.640 170.180 58.960 170.240 ;
        RECT 65.080 170.380 65.400 170.440 ;
        RECT 66.060 170.380 66.350 170.425 ;
        RECT 65.080 170.240 66.350 170.380 ;
        RECT 65.080 170.180 65.400 170.240 ;
        RECT 66.060 170.195 66.350 170.240 ;
        RECT 68.300 170.180 68.620 170.440 ;
        RECT 75.660 170.380 75.980 170.440 ;
        RECT 77.500 170.380 77.820 170.440 ;
        RECT 70.230 170.240 72.670 170.380 ;
        RECT 70.230 170.100 70.370 170.240 ;
        RECT 54.960 169.900 55.650 170.040 ;
        RECT 54.960 169.840 55.280 169.900 ;
        RECT 31.040 169.500 31.360 169.760 ;
        RECT 37.020 169.500 37.340 169.760 ;
        RECT 55.510 169.745 55.650 169.900 ;
        RECT 55.895 169.900 57.030 170.040 ;
        RECT 55.895 169.855 56.185 169.900 ;
        RECT 69.220 169.840 69.540 170.100 ;
        RECT 69.680 169.840 70.000 170.100 ;
        RECT 70.140 169.840 70.460 170.100 ;
        RECT 70.600 169.840 70.920 170.100 ;
        RECT 71.060 170.040 71.380 170.100 ;
        RECT 71.535 170.040 71.825 170.085 ;
        RECT 71.060 169.900 71.825 170.040 ;
        RECT 71.060 169.840 71.380 169.900 ;
        RECT 71.535 169.855 71.825 169.900 ;
        RECT 71.980 169.840 72.300 170.100 ;
        RECT 72.530 170.085 72.670 170.240 ;
        RECT 75.660 170.240 77.820 170.380 ;
        RECT 75.660 170.180 75.980 170.240 ;
        RECT 77.500 170.180 77.820 170.240 ;
        RECT 77.975 170.380 78.265 170.425 ;
        RECT 79.430 170.380 79.570 170.580 ;
        RECT 80.735 170.380 81.025 170.425 ;
        RECT 77.975 170.240 79.570 170.380 ;
        RECT 79.890 170.240 81.025 170.380 ;
        RECT 77.975 170.195 78.265 170.240 ;
        RECT 79.890 170.100 80.030 170.240 ;
        RECT 80.735 170.195 81.025 170.240 ;
        RECT 81.270 170.100 81.410 170.580 ;
        RECT 93.600 170.520 93.920 170.780 ;
        RECT 96.375 170.720 96.665 170.765 ;
        RECT 97.280 170.720 97.600 170.780 ;
        RECT 96.375 170.580 97.600 170.720 ;
        RECT 96.375 170.535 96.665 170.580 ;
        RECT 97.280 170.520 97.600 170.580 ;
        RECT 100.515 170.720 100.805 170.765 ;
        RECT 102.800 170.720 103.120 170.780 ;
        RECT 104.640 170.720 104.960 170.780 ;
        RECT 100.515 170.580 104.960 170.720 ;
        RECT 100.515 170.535 100.805 170.580 ;
        RECT 102.800 170.520 103.120 170.580 ;
        RECT 104.640 170.520 104.960 170.580 ;
        RECT 116.600 170.520 116.920 170.780 ;
        RECT 129.020 170.520 129.340 170.780 ;
        RECT 131.320 170.720 131.640 170.780 ;
        RECT 129.570 170.580 131.640 170.720 ;
        RECT 105.100 170.380 105.420 170.440 ;
        RECT 106.080 170.380 106.370 170.425 ;
        RECT 105.100 170.240 106.370 170.380 ;
        RECT 105.100 170.180 105.420 170.240 ;
        RECT 106.080 170.195 106.370 170.240 ;
        RECT 72.455 169.855 72.745 170.085 ;
        RECT 75.200 169.840 75.520 170.100 ;
        RECT 77.055 169.855 77.345 170.085 ;
        RECT 78.895 169.855 79.185 170.085 ;
        RECT 55.435 169.515 55.725 169.745 ;
        RECT 62.805 169.700 63.095 169.745 ;
        RECT 65.325 169.700 65.615 169.745 ;
        RECT 66.515 169.700 66.805 169.745 ;
        RECT 62.805 169.560 66.805 169.700 ;
        RECT 62.805 169.515 63.095 169.560 ;
        RECT 65.325 169.515 65.615 169.560 ;
        RECT 66.515 169.515 66.805 169.560 ;
        RECT 67.395 169.700 67.685 169.745 ;
        RECT 75.290 169.700 75.430 169.840 ;
        RECT 67.395 169.560 75.430 169.700 ;
        RECT 77.130 169.700 77.270 169.855 ;
        RECT 78.970 169.700 79.110 169.855 ;
        RECT 79.800 169.840 80.120 170.100 ;
        RECT 80.260 169.840 80.580 170.100 ;
        RECT 81.180 169.840 81.500 170.100 ;
        RECT 82.115 170.040 82.405 170.085 ;
        RECT 87.620 170.040 87.940 170.100 ;
        RECT 91.300 170.040 91.620 170.100 ;
        RECT 94.075 170.040 94.365 170.085 ;
        RECT 82.115 169.900 87.940 170.040 ;
        RECT 82.115 169.855 82.405 169.900 ;
        RECT 87.620 169.840 87.940 169.900 ;
        RECT 89.090 169.900 94.365 170.040 ;
        RECT 82.575 169.700 82.865 169.745 ;
        RECT 77.130 169.560 77.730 169.700 ;
        RECT 78.970 169.560 82.865 169.700 ;
        RECT 67.395 169.515 67.685 169.560 ;
        RECT 33.355 169.360 33.645 169.405 ;
        RECT 36.575 169.360 36.865 169.405 ;
        RECT 37.110 169.360 37.250 169.500 ;
        RECT 42.540 169.360 42.860 169.420 ;
        RECT 33.355 169.220 37.250 169.360 ;
        RECT 37.570 169.220 42.860 169.360 ;
        RECT 33.355 169.175 33.645 169.220 ;
        RECT 36.575 169.175 36.865 169.220 ;
        RECT 35.180 168.820 35.500 169.080 ;
        RECT 37.570 169.065 37.710 169.220 ;
        RECT 42.540 169.160 42.860 169.220 ;
        RECT 54.515 169.360 54.805 169.405 ;
        RECT 58.180 169.360 58.500 169.420 ;
        RECT 54.515 169.220 58.500 169.360 ;
        RECT 54.515 169.175 54.805 169.220 ;
        RECT 58.180 169.160 58.500 169.220 ;
        RECT 63.240 169.360 63.530 169.405 ;
        RECT 64.810 169.360 65.100 169.405 ;
        RECT 66.910 169.360 67.200 169.405 ;
        RECT 63.240 169.220 67.200 169.360 ;
        RECT 77.590 169.360 77.730 169.560 ;
        RECT 82.575 169.515 82.865 169.560 ;
        RECT 83.940 169.700 84.260 169.760 ;
        RECT 85.335 169.700 85.625 169.745 ;
        RECT 83.940 169.560 85.625 169.700 ;
        RECT 83.940 169.500 84.260 169.560 ;
        RECT 85.335 169.515 85.625 169.560 ;
        RECT 80.260 169.360 80.580 169.420 ;
        RECT 77.590 169.220 80.580 169.360 ;
        RECT 63.240 169.175 63.530 169.220 ;
        RECT 64.810 169.175 65.100 169.220 ;
        RECT 66.910 169.175 67.200 169.220 ;
        RECT 80.260 169.160 80.580 169.220 ;
        RECT 37.495 168.835 37.785 169.065 ;
        RECT 37.940 169.020 38.260 169.080 ;
        RECT 38.875 169.020 39.165 169.065 ;
        RECT 37.940 168.880 39.165 169.020 ;
        RECT 37.940 168.820 38.260 168.880 ;
        RECT 38.875 168.835 39.165 168.880 ;
        RECT 47.600 169.020 47.920 169.080 ;
        RECT 49.455 169.020 49.745 169.065 ;
        RECT 47.600 168.880 49.745 169.020 ;
        RECT 47.600 168.820 47.920 168.880 ;
        RECT 49.455 168.835 49.745 168.880 ;
        RECT 51.280 168.820 51.600 169.080 ;
        RECT 57.260 168.820 57.580 169.080 ;
        RECT 73.375 169.020 73.665 169.065 ;
        RECT 75.660 169.020 75.980 169.080 ;
        RECT 73.375 168.880 75.980 169.020 ;
        RECT 73.375 168.835 73.665 168.880 ;
        RECT 75.660 168.820 75.980 168.880 ;
        RECT 76.120 168.820 76.440 169.080 ;
        RECT 79.340 168.820 79.660 169.080 ;
        RECT 85.410 169.020 85.550 169.515 ;
        RECT 89.090 169.420 89.230 169.900 ;
        RECT 91.300 169.840 91.620 169.900 ;
        RECT 94.075 169.855 94.365 169.900 ;
        RECT 109.240 170.040 109.560 170.100 ;
        RECT 110.995 170.040 111.285 170.085 ;
        RECT 109.240 169.900 111.285 170.040 ;
        RECT 116.690 170.040 116.830 170.520 ;
        RECT 129.570 170.380 129.710 170.580 ;
        RECT 131.320 170.520 131.640 170.580 ;
        RECT 133.160 170.720 133.480 170.780 ;
        RECT 136.395 170.720 136.685 170.765 ;
        RECT 133.160 170.580 136.685 170.720 ;
        RECT 133.160 170.520 133.480 170.580 ;
        RECT 136.395 170.535 136.685 170.580 ;
        RECT 138.695 170.720 138.985 170.765 ;
        RECT 141.900 170.720 142.220 170.780 ;
        RECT 138.695 170.580 142.220 170.720 ;
        RECT 138.695 170.535 138.985 170.580 ;
        RECT 141.900 170.520 142.220 170.580 ;
        RECT 142.360 170.720 142.680 170.780 ;
        RECT 148.735 170.720 149.025 170.765 ;
        RECT 150.180 170.720 150.500 170.780 ;
        RECT 142.360 170.580 148.110 170.720 ;
        RECT 142.360 170.520 142.680 170.580 ;
        RECT 130.860 170.425 131.180 170.440 ;
        RECT 123.130 170.240 129.710 170.380 ;
        RECT 123.130 170.085 123.270 170.240 ;
        RECT 130.720 170.195 131.180 170.425 ;
        RECT 142.820 170.380 143.140 170.440 ;
        RECT 130.860 170.180 131.180 170.195 ;
        RECT 139.690 170.240 143.140 170.380 ;
        RECT 119.835 170.040 120.125 170.085 ;
        RECT 123.055 170.040 123.345 170.085 ;
        RECT 116.690 169.900 120.125 170.040 ;
        RECT 109.240 169.840 109.560 169.900 ;
        RECT 110.995 169.855 111.285 169.900 ;
        RECT 119.835 169.855 120.125 169.900 ;
        RECT 120.370 169.900 123.345 170.040 ;
        RECT 102.825 169.700 103.115 169.745 ;
        RECT 105.345 169.700 105.635 169.745 ;
        RECT 106.535 169.700 106.825 169.745 ;
        RECT 102.825 169.560 106.825 169.700 ;
        RECT 102.825 169.515 103.115 169.560 ;
        RECT 105.345 169.515 105.635 169.560 ;
        RECT 106.535 169.515 106.825 169.560 ;
        RECT 107.415 169.700 107.705 169.745 ;
        RECT 109.700 169.700 110.020 169.760 ;
        RECT 107.415 169.560 110.020 169.700 ;
        RECT 107.415 169.515 107.705 169.560 ;
        RECT 109.700 169.500 110.020 169.560 ;
        RECT 110.595 169.700 110.885 169.745 ;
        RECT 111.785 169.700 112.075 169.745 ;
        RECT 114.305 169.700 114.595 169.745 ;
        RECT 110.595 169.560 114.595 169.700 ;
        RECT 110.595 169.515 110.885 169.560 ;
        RECT 111.785 169.515 112.075 169.560 ;
        RECT 114.305 169.515 114.595 169.560 ;
        RECT 89.000 169.160 89.320 169.420 ;
        RECT 95.455 169.360 95.745 169.405 ;
        RECT 91.850 169.220 95.745 169.360 ;
        RECT 91.850 169.065 91.990 169.220 ;
        RECT 95.455 169.175 95.745 169.220 ;
        RECT 103.260 169.360 103.550 169.405 ;
        RECT 104.830 169.360 105.120 169.405 ;
        RECT 106.930 169.360 107.220 169.405 ;
        RECT 103.260 169.220 107.220 169.360 ;
        RECT 103.260 169.175 103.550 169.220 ;
        RECT 104.830 169.175 105.120 169.220 ;
        RECT 106.930 169.175 107.220 169.220 ;
        RECT 110.200 169.360 110.490 169.405 ;
        RECT 112.300 169.360 112.590 169.405 ;
        RECT 113.870 169.360 114.160 169.405 ;
        RECT 120.370 169.360 120.510 169.900 ;
        RECT 123.055 169.855 123.345 169.900 ;
        RECT 127.195 170.040 127.485 170.085 ;
        RECT 129.940 170.040 130.260 170.100 ;
        RECT 139.690 170.085 139.830 170.240 ;
        RECT 142.820 170.180 143.140 170.240 ;
        RECT 144.660 170.380 144.980 170.440 ;
        RECT 147.435 170.380 147.725 170.425 ;
        RECT 144.660 170.240 147.725 170.380 ;
        RECT 144.660 170.180 144.980 170.240 ;
        RECT 147.435 170.195 147.725 170.240 ;
        RECT 138.235 170.040 138.525 170.085 ;
        RECT 127.195 169.900 130.260 170.040 ;
        RECT 127.195 169.855 127.485 169.900 ;
        RECT 129.940 169.840 130.260 169.900 ;
        RECT 137.850 169.900 138.525 170.040 ;
        RECT 121.660 169.700 121.980 169.760 ;
        RECT 126.735 169.700 127.025 169.745 ;
        RECT 121.660 169.560 127.025 169.700 ;
        RECT 121.660 169.500 121.980 169.560 ;
        RECT 126.735 169.515 127.025 169.560 ;
        RECT 129.480 169.500 129.800 169.760 ;
        RECT 130.375 169.700 130.665 169.745 ;
        RECT 131.565 169.700 131.855 169.745 ;
        RECT 134.085 169.700 134.375 169.745 ;
        RECT 130.375 169.560 134.375 169.700 ;
        RECT 130.375 169.515 130.665 169.560 ;
        RECT 131.565 169.515 131.855 169.560 ;
        RECT 134.085 169.515 134.375 169.560 ;
        RECT 137.850 169.700 137.990 169.900 ;
        RECT 138.235 169.855 138.525 169.900 ;
        RECT 139.155 170.040 139.445 170.085 ;
        RECT 139.615 170.040 139.905 170.085 ;
        RECT 139.155 169.900 139.905 170.040 ;
        RECT 139.155 169.855 139.445 169.900 ;
        RECT 139.615 169.855 139.905 169.900 ;
        RECT 140.535 169.855 140.825 170.085 ;
        RECT 140.995 169.855 141.285 170.085 ;
        RECT 141.455 170.040 141.745 170.085 ;
        RECT 141.900 170.040 142.220 170.100 ;
        RECT 141.455 169.900 142.220 170.040 ;
        RECT 141.455 169.855 141.745 169.900 ;
        RECT 140.610 169.700 140.750 169.855 ;
        RECT 137.850 169.560 140.750 169.700 ;
        RECT 141.070 169.700 141.210 169.855 ;
        RECT 141.900 169.840 142.220 169.900 ;
        RECT 145.580 169.840 145.900 170.100 ;
        RECT 146.975 170.040 147.265 170.085 ;
        RECT 147.970 170.040 148.110 170.580 ;
        RECT 148.735 170.580 150.500 170.720 ;
        RECT 148.735 170.535 149.025 170.580 ;
        RECT 150.180 170.520 150.500 170.580 ;
        RECT 151.100 170.520 151.420 170.780 ;
        RECT 149.260 170.380 149.580 170.440 ;
        RECT 149.735 170.380 150.025 170.425 ;
        RECT 149.260 170.240 150.025 170.380 ;
        RECT 149.260 170.180 149.580 170.240 ;
        RECT 149.735 170.195 150.025 170.240 ;
        RECT 151.190 170.380 151.330 170.520 ;
        RECT 152.955 170.380 153.245 170.425 ;
        RECT 151.190 170.240 153.245 170.380 ;
        RECT 151.190 170.085 151.330 170.240 ;
        RECT 152.955 170.195 153.245 170.240 ;
        RECT 146.975 169.900 148.110 170.040 ;
        RECT 146.975 169.855 147.265 169.900 ;
        RECT 151.115 169.855 151.405 170.085 ;
        RECT 152.020 169.840 152.340 170.100 ;
        RECT 154.335 169.855 154.625 170.085 ;
        RECT 142.360 169.700 142.680 169.760 ;
        RECT 141.070 169.560 142.680 169.700 ;
        RECT 110.200 169.220 114.160 169.360 ;
        RECT 110.200 169.175 110.490 169.220 ;
        RECT 112.300 169.175 112.590 169.220 ;
        RECT 113.870 169.175 114.160 169.220 ;
        RECT 114.390 169.220 120.510 169.360 ;
        RECT 91.775 169.020 92.065 169.065 ;
        RECT 85.410 168.880 92.065 169.020 ;
        RECT 91.775 168.835 92.065 168.880 ;
        RECT 94.980 169.020 95.300 169.080 ;
        RECT 114.390 169.020 114.530 169.220 ;
        RECT 94.980 168.880 114.530 169.020 ;
        RECT 114.760 169.020 115.080 169.080 ;
        RECT 117.075 169.020 117.365 169.065 ;
        RECT 114.760 168.880 117.365 169.020 ;
        RECT 129.570 169.020 129.710 169.500 ;
        RECT 129.980 169.360 130.270 169.405 ;
        RECT 132.080 169.360 132.370 169.405 ;
        RECT 133.650 169.360 133.940 169.405 ;
        RECT 129.980 169.220 133.940 169.360 ;
        RECT 129.980 169.175 130.270 169.220 ;
        RECT 132.080 169.175 132.370 169.220 ;
        RECT 133.650 169.175 133.940 169.220 ;
        RECT 137.850 169.080 137.990 169.560 ;
        RECT 142.360 169.500 142.680 169.560 ;
        RECT 143.280 169.700 143.600 169.760 ;
        RECT 145.135 169.700 145.425 169.745 ;
        RECT 143.280 169.560 145.425 169.700 ;
        RECT 143.280 169.500 143.600 169.560 ;
        RECT 145.135 169.515 145.425 169.560 ;
        RECT 148.340 169.700 148.660 169.760 ;
        RECT 154.410 169.700 154.550 169.855 ;
        RECT 148.340 169.560 154.550 169.700 ;
        RECT 148.340 169.500 148.660 169.560 ;
        RECT 153.875 169.360 154.165 169.405 ;
        RECT 148.890 169.220 154.165 169.360 ;
        RECT 137.300 169.020 137.620 169.080 ;
        RECT 129.570 168.880 137.620 169.020 ;
        RECT 94.980 168.820 95.300 168.880 ;
        RECT 114.760 168.820 115.080 168.880 ;
        RECT 117.075 168.835 117.365 168.880 ;
        RECT 137.300 168.820 137.620 168.880 ;
        RECT 137.760 168.820 138.080 169.080 ;
        RECT 144.215 169.020 144.505 169.065 ;
        RECT 145.120 169.020 145.440 169.080 ;
        RECT 144.215 168.880 145.440 169.020 ;
        RECT 144.215 168.835 144.505 168.880 ;
        RECT 145.120 168.820 145.440 168.880 ;
        RECT 146.960 169.020 147.280 169.080 ;
        RECT 148.890 169.065 149.030 169.220 ;
        RECT 153.875 169.175 154.165 169.220 ;
        RECT 147.895 169.020 148.185 169.065 ;
        RECT 146.960 168.880 148.185 169.020 ;
        RECT 146.960 168.820 147.280 168.880 ;
        RECT 147.895 168.835 148.185 168.880 ;
        RECT 148.815 168.835 149.105 169.065 ;
        RECT 150.640 168.820 150.960 169.080 ;
        RECT 154.780 168.820 155.100 169.080 ;
        RECT 22.690 168.200 157.010 168.680 ;
        RECT 31.040 167.800 31.360 168.060 ;
        RECT 32.420 167.800 32.740 168.060 ;
        RECT 34.720 168.000 35.040 168.060 ;
        RECT 42.540 168.000 42.860 168.060 ;
        RECT 47.140 168.000 47.460 168.060 ;
        RECT 53.595 168.000 53.885 168.045 ;
        RECT 32.970 167.860 53.885 168.000 ;
        RECT 24.640 167.660 24.930 167.705 ;
        RECT 26.740 167.660 27.030 167.705 ;
        RECT 28.310 167.660 28.600 167.705 ;
        RECT 24.640 167.520 28.600 167.660 ;
        RECT 31.130 167.660 31.270 167.800 ;
        RECT 32.970 167.660 33.110 167.860 ;
        RECT 34.720 167.800 35.040 167.860 ;
        RECT 42.540 167.800 42.860 167.860 ;
        RECT 47.140 167.800 47.460 167.860 ;
        RECT 53.595 167.815 53.885 167.860 ;
        RECT 61.860 168.000 62.180 168.060 ;
        RECT 65.555 168.000 65.845 168.045 ;
        RECT 61.860 167.860 65.845 168.000 ;
        RECT 61.860 167.800 62.180 167.860 ;
        RECT 65.555 167.815 65.845 167.860 ;
        RECT 79.800 168.000 80.120 168.060 ;
        RECT 88.540 168.000 88.860 168.060 ;
        RECT 89.935 168.000 90.225 168.045 ;
        RECT 79.800 167.860 88.310 168.000 ;
        RECT 79.800 167.800 80.120 167.860 ;
        RECT 31.130 167.520 33.110 167.660 ;
        RECT 33.340 167.660 33.660 167.720 ;
        RECT 34.275 167.660 34.565 167.705 ;
        RECT 33.340 167.520 34.565 167.660 ;
        RECT 24.640 167.475 24.930 167.520 ;
        RECT 26.740 167.475 27.030 167.520 ;
        RECT 28.310 167.475 28.600 167.520 ;
        RECT 33.340 167.460 33.660 167.520 ;
        RECT 34.275 167.475 34.565 167.520 ;
        RECT 37.520 167.660 37.810 167.705 ;
        RECT 39.620 167.660 39.910 167.705 ;
        RECT 41.190 167.660 41.480 167.705 ;
        RECT 37.520 167.520 41.480 167.660 ;
        RECT 37.520 167.475 37.810 167.520 ;
        RECT 39.620 167.475 39.910 167.520 ;
        RECT 41.190 167.475 41.480 167.520 ;
        RECT 43.460 167.660 43.780 167.720 ;
        RECT 43.935 167.660 44.225 167.705 ;
        RECT 43.460 167.520 46.910 167.660 ;
        RECT 43.460 167.460 43.780 167.520 ;
        RECT 43.935 167.475 44.225 167.520 ;
        RECT 24.140 167.120 24.460 167.380 ;
        RECT 25.035 167.320 25.325 167.365 ;
        RECT 26.225 167.320 26.515 167.365 ;
        RECT 28.745 167.320 29.035 167.365 ;
        RECT 25.035 167.180 29.035 167.320 ;
        RECT 25.035 167.135 25.325 167.180 ;
        RECT 26.225 167.135 26.515 167.180 ;
        RECT 28.745 167.135 29.035 167.180 ;
        RECT 37.915 167.320 38.205 167.365 ;
        RECT 39.105 167.320 39.395 167.365 ;
        RECT 41.625 167.320 41.915 167.365 ;
        RECT 45.775 167.320 46.065 167.365 ;
        RECT 37.915 167.180 41.915 167.320 ;
        RECT 37.915 167.135 38.205 167.180 ;
        RECT 39.105 167.135 39.395 167.180 ;
        RECT 41.625 167.135 41.915 167.180 ;
        RECT 44.930 167.180 46.065 167.320 ;
        RECT 44.930 167.040 45.070 167.180 ;
        RECT 45.775 167.135 46.065 167.180 ;
        RECT 37.020 166.780 37.340 167.040 ;
        RECT 44.840 166.780 45.160 167.040 ;
        RECT 45.300 166.780 45.620 167.040 ;
        RECT 46.770 167.025 46.910 167.520 ;
        RECT 52.215 167.475 52.505 167.705 ;
        RECT 53.120 167.660 53.440 167.720 ;
        RECT 80.260 167.660 80.580 167.720 ;
        RECT 53.120 167.520 66.690 167.660 ;
        RECT 50.835 167.320 51.125 167.365 ;
        RECT 51.280 167.320 51.600 167.380 ;
        RECT 50.835 167.180 51.600 167.320 ;
        RECT 52.290 167.320 52.430 167.475 ;
        RECT 53.120 167.460 53.440 167.520 ;
        RECT 59.560 167.320 59.880 167.380 ;
        RECT 52.290 167.180 54.730 167.320 ;
        RECT 50.835 167.135 51.125 167.180 ;
        RECT 51.280 167.120 51.600 167.180 ;
        RECT 46.235 166.980 46.525 167.025 ;
        RECT 45.850 166.840 46.525 166.980 ;
        RECT 25.490 166.640 25.780 166.685 ;
        RECT 25.980 166.640 26.300 166.700 ;
        RECT 25.490 166.500 26.300 166.640 ;
        RECT 25.490 166.455 25.780 166.500 ;
        RECT 25.980 166.440 26.300 166.500 ;
        RECT 38.370 166.455 38.660 166.685 ;
        RECT 31.500 166.100 31.820 166.360 ;
        RECT 32.435 166.300 32.725 166.345 ;
        RECT 33.800 166.300 34.120 166.360 ;
        RECT 35.640 166.300 35.960 166.360 ;
        RECT 32.435 166.160 35.960 166.300 ;
        RECT 32.435 166.115 32.725 166.160 ;
        RECT 33.800 166.100 34.120 166.160 ;
        RECT 35.640 166.100 35.960 166.160 ;
        RECT 37.940 166.300 38.260 166.360 ;
        RECT 38.490 166.300 38.630 166.455 ;
        RECT 37.940 166.160 38.630 166.300 ;
        RECT 37.940 166.100 38.260 166.160 ;
        RECT 44.380 166.100 44.700 166.360 ;
        RECT 45.390 166.300 45.530 166.780 ;
        RECT 45.850 166.700 45.990 166.840 ;
        RECT 46.235 166.795 46.525 166.840 ;
        RECT 46.695 166.980 46.985 167.025 ;
        RECT 47.600 166.980 47.920 167.040 ;
        RECT 46.695 166.840 47.920 166.980 ;
        RECT 46.695 166.795 46.985 166.840 ;
        RECT 47.600 166.780 47.920 166.840 ;
        RECT 48.980 166.780 49.300 167.040 ;
        RECT 50.375 166.980 50.665 167.025 ;
        RECT 50.375 166.840 52.890 166.980 ;
        RECT 50.375 166.795 50.665 166.840 ;
        RECT 45.760 166.440 46.080 166.700 ;
        RECT 51.280 166.685 51.600 166.700 ;
        RECT 51.280 166.455 51.710 166.685 ;
        RECT 51.280 166.440 51.600 166.455 ;
        RECT 52.750 166.360 52.890 166.840 ;
        RECT 54.590 166.640 54.730 167.180 ;
        RECT 56.890 167.180 59.880 167.320 ;
        RECT 54.960 166.780 55.280 167.040 ;
        RECT 55.420 166.980 55.740 167.040 ;
        RECT 56.355 166.980 56.645 167.025 ;
        RECT 55.420 166.840 56.645 166.980 ;
        RECT 55.420 166.780 55.740 166.840 ;
        RECT 56.355 166.795 56.645 166.840 ;
        RECT 56.890 166.685 57.030 167.180 ;
        RECT 59.560 167.120 59.880 167.180 ;
        RECT 57.275 166.795 57.565 167.025 ;
        RECT 57.735 166.980 58.025 167.025 ;
        RECT 58.640 166.980 58.960 167.040 ;
        RECT 66.550 167.025 66.690 167.520 ;
        RECT 80.260 167.520 83.250 167.660 ;
        RECT 80.260 167.460 80.580 167.520 ;
        RECT 67.395 167.320 67.685 167.365 ;
        RECT 69.220 167.320 69.540 167.380 ;
        RECT 82.100 167.320 82.420 167.380 ;
        RECT 83.110 167.365 83.250 167.520 ;
        RECT 67.395 167.180 82.420 167.320 ;
        RECT 67.395 167.135 67.685 167.180 ;
        RECT 69.220 167.120 69.540 167.180 ;
        RECT 82.100 167.120 82.420 167.180 ;
        RECT 83.035 167.135 83.325 167.365 ;
        RECT 88.170 167.320 88.310 167.860 ;
        RECT 88.540 167.860 90.225 168.000 ;
        RECT 88.540 167.800 88.860 167.860 ;
        RECT 89.935 167.815 90.225 167.860 ;
        RECT 105.100 168.000 105.420 168.060 ;
        RECT 106.035 168.000 106.325 168.045 ;
        RECT 105.100 167.860 106.325 168.000 ;
        RECT 105.100 167.800 105.420 167.860 ;
        RECT 106.035 167.815 106.325 167.860 ;
        RECT 109.240 167.800 109.560 168.060 ;
        RECT 113.380 168.000 113.700 168.060 ;
        RECT 113.855 168.000 114.145 168.045 ;
        RECT 113.380 167.860 114.145 168.000 ;
        RECT 113.380 167.800 113.700 167.860 ;
        RECT 113.855 167.815 114.145 167.860 ;
        RECT 117.535 168.000 117.825 168.045 ;
        RECT 122.120 168.000 122.440 168.060 ;
        RECT 139.155 168.000 139.445 168.045 ;
        RECT 117.535 167.860 122.440 168.000 ;
        RECT 117.535 167.815 117.825 167.860 ;
        RECT 122.120 167.800 122.440 167.860 ;
        RECT 126.350 167.860 139.445 168.000 ;
        RECT 89.475 167.660 89.765 167.705 ;
        RECT 91.300 167.660 91.620 167.720 ;
        RECT 116.600 167.660 116.920 167.720 ;
        RECT 119.400 167.660 119.690 167.705 ;
        RECT 121.500 167.660 121.790 167.705 ;
        RECT 123.070 167.660 123.360 167.705 ;
        RECT 89.475 167.520 91.620 167.660 ;
        RECT 89.475 167.475 89.765 167.520 ;
        RECT 91.300 167.460 91.620 167.520 ;
        RECT 105.190 167.520 119.130 167.660 ;
        RECT 102.355 167.320 102.645 167.365 ;
        RECT 102.800 167.320 103.120 167.380 ;
        RECT 88.170 167.180 102.110 167.320 ;
        RECT 57.735 166.840 58.960 166.980 ;
        RECT 57.735 166.795 58.025 166.840 ;
        RECT 56.815 166.640 57.105 166.685 ;
        RECT 54.590 166.500 57.105 166.640 ;
        RECT 57.350 166.640 57.490 166.795 ;
        RECT 58.640 166.780 58.960 166.840 ;
        RECT 66.475 166.795 66.765 167.025 ;
        RECT 67.855 166.795 68.145 167.025 ;
        RECT 70.140 166.980 70.460 167.040 ;
        RECT 71.075 166.980 71.365 167.025 ;
        RECT 70.140 166.840 71.365 166.980 ;
        RECT 59.100 166.640 59.420 166.700 ;
        RECT 57.350 166.500 59.420 166.640 ;
        RECT 67.930 166.640 68.070 166.795 ;
        RECT 70.140 166.780 70.460 166.840 ;
        RECT 71.075 166.795 71.365 166.840 ;
        RECT 74.280 166.780 74.600 167.040 ;
        RECT 77.960 166.980 78.280 167.040 ;
        RECT 82.575 166.980 82.865 167.025 ;
        RECT 77.960 166.840 82.865 166.980 ;
        RECT 77.960 166.780 78.280 166.840 ;
        RECT 82.575 166.795 82.865 166.840 ;
        RECT 83.495 166.795 83.785 167.025 ;
        RECT 69.680 166.640 70.000 166.700 ;
        RECT 74.370 166.640 74.510 166.780 ;
        RECT 82.100 166.640 82.420 166.700 ;
        RECT 83.570 166.640 83.710 166.795 ;
        RECT 84.400 166.780 84.720 167.040 ;
        RECT 89.000 166.980 89.320 167.040 ;
        RECT 89.935 166.980 90.225 167.025 ;
        RECT 89.000 166.840 90.225 166.980 ;
        RECT 89.000 166.780 89.320 166.840 ;
        RECT 89.935 166.795 90.225 166.840 ;
        RECT 90.395 166.980 90.685 167.025 ;
        RECT 93.140 166.980 93.460 167.040 ;
        RECT 90.395 166.840 93.460 166.980 ;
        RECT 90.395 166.795 90.685 166.840 ;
        RECT 93.140 166.780 93.460 166.840 ;
        RECT 94.980 166.780 95.300 167.040 ;
        RECT 67.930 166.500 74.510 166.640 ;
        RECT 74.830 166.500 76.350 166.640 ;
        RECT 56.815 166.455 57.105 166.500 ;
        RECT 59.100 166.440 59.420 166.500 ;
        RECT 69.680 166.440 70.000 166.500 ;
        RECT 48.060 166.300 48.380 166.360 ;
        RECT 45.390 166.160 48.380 166.300 ;
        RECT 48.060 166.100 48.380 166.160 ;
        RECT 52.660 166.100 52.980 166.360 ;
        RECT 55.435 166.300 55.725 166.345 ;
        RECT 57.260 166.300 57.580 166.360 ;
        RECT 55.435 166.160 57.580 166.300 ;
        RECT 55.435 166.115 55.725 166.160 ;
        RECT 57.260 166.100 57.580 166.160 ;
        RECT 68.300 166.100 68.620 166.360 ;
        RECT 71.520 166.300 71.840 166.360 ;
        RECT 74.830 166.300 74.970 166.500 ;
        RECT 71.520 166.160 74.970 166.300 ;
        RECT 71.520 166.100 71.840 166.160 ;
        RECT 75.200 166.100 75.520 166.360 ;
        RECT 76.210 166.300 76.350 166.500 ;
        RECT 82.100 166.500 83.710 166.640 ;
        RECT 87.160 166.640 87.480 166.700 ;
        RECT 87.635 166.640 87.925 166.685 ;
        RECT 87.160 166.500 87.925 166.640 ;
        RECT 82.100 166.440 82.420 166.500 ;
        RECT 87.160 166.440 87.480 166.500 ;
        RECT 87.635 166.455 87.925 166.500 ;
        RECT 91.315 166.640 91.605 166.685 ;
        RECT 92.680 166.640 93.000 166.700 ;
        RECT 95.070 166.640 95.210 166.780 ;
        RECT 91.315 166.500 95.210 166.640 ;
        RECT 101.970 166.640 102.110 167.180 ;
        RECT 102.355 167.180 103.120 167.320 ;
        RECT 102.355 167.135 102.645 167.180 ;
        RECT 102.800 167.120 103.120 167.180 ;
        RECT 105.190 166.640 105.330 167.520 ;
        RECT 116.600 167.460 116.920 167.520 ;
        RECT 105.575 167.320 105.865 167.365 ;
        RECT 111.080 167.320 111.400 167.380 ;
        RECT 114.760 167.320 115.080 167.380 ;
        RECT 105.575 167.180 109.010 167.320 ;
        RECT 105.575 167.135 105.865 167.180 ;
        RECT 106.940 166.980 107.260 167.040 ;
        RECT 108.870 167.025 109.010 167.180 ;
        RECT 110.710 167.180 111.400 167.320 ;
        RECT 106.940 166.840 108.550 166.980 ;
        RECT 106.940 166.780 107.260 166.840 ;
        RECT 107.415 166.640 107.705 166.685 ;
        RECT 101.970 166.500 107.705 166.640 ;
        RECT 91.315 166.455 91.605 166.500 ;
        RECT 92.680 166.440 93.000 166.500 ;
        RECT 107.415 166.455 107.705 166.500 ;
        RECT 107.875 166.455 108.165 166.685 ;
        RECT 108.410 166.640 108.550 166.840 ;
        RECT 108.795 166.795 109.085 167.025 ;
        RECT 109.240 166.980 109.560 167.040 ;
        RECT 110.710 167.025 110.850 167.180 ;
        RECT 111.080 167.120 111.400 167.180 ;
        RECT 112.090 167.180 115.080 167.320 ;
        RECT 118.990 167.320 119.130 167.520 ;
        RECT 119.400 167.520 123.360 167.660 ;
        RECT 119.400 167.475 119.690 167.520 ;
        RECT 121.500 167.475 121.790 167.520 ;
        RECT 123.070 167.475 123.360 167.520 ;
        RECT 119.795 167.320 120.085 167.365 ;
        RECT 120.985 167.320 121.275 167.365 ;
        RECT 123.505 167.320 123.795 167.365 ;
        RECT 118.990 167.180 119.590 167.320 ;
        RECT 112.090 167.025 112.230 167.180 ;
        RECT 114.760 167.120 115.080 167.180 ;
        RECT 110.175 166.980 110.465 167.025 ;
        RECT 109.240 166.840 110.465 166.980 ;
        RECT 109.240 166.780 109.560 166.840 ;
        RECT 110.175 166.795 110.465 166.840 ;
        RECT 110.635 166.795 110.925 167.025 ;
        RECT 112.015 166.795 112.305 167.025 ;
        RECT 114.315 166.795 114.605 167.025 ;
        RECT 109.330 166.640 109.470 166.780 ;
        RECT 108.410 166.500 109.470 166.640 ;
        RECT 111.095 166.455 111.385 166.685 ;
        RECT 114.390 166.640 114.530 166.795 ;
        RECT 115.220 166.780 115.540 167.040 ;
        RECT 115.680 166.780 116.000 167.040 ;
        RECT 116.600 166.780 116.920 167.040 ;
        RECT 117.060 166.980 117.380 167.040 ;
        RECT 118.915 166.980 119.205 167.025 ;
        RECT 117.060 166.840 119.205 166.980 ;
        RECT 119.450 166.980 119.590 167.180 ;
        RECT 119.795 167.180 123.795 167.320 ;
        RECT 119.795 167.135 120.085 167.180 ;
        RECT 120.985 167.135 121.275 167.180 ;
        RECT 123.505 167.135 123.795 167.180 ;
        RECT 126.350 167.025 126.490 167.860 ;
        RECT 139.155 167.815 139.445 167.860 ;
        RECT 144.660 168.000 144.980 168.060 ;
        RECT 146.055 168.000 146.345 168.045 ;
        RECT 144.660 167.860 146.345 168.000 ;
        RECT 144.660 167.800 144.980 167.860 ;
        RECT 146.055 167.815 146.345 167.860 ;
        RECT 147.880 167.800 148.200 168.060 ;
        RECT 148.340 167.800 148.660 168.060 ;
        RECT 129.980 167.660 130.270 167.705 ;
        RECT 132.080 167.660 132.370 167.705 ;
        RECT 133.650 167.660 133.940 167.705 ;
        RECT 129.980 167.520 133.940 167.660 ;
        RECT 129.980 167.475 130.270 167.520 ;
        RECT 132.080 167.475 132.370 167.520 ;
        RECT 133.650 167.475 133.940 167.520 ;
        RECT 136.395 167.660 136.685 167.705 ;
        RECT 137.760 167.660 138.080 167.720 ;
        RECT 136.395 167.520 138.080 167.660 ;
        RECT 136.395 167.475 136.685 167.520 ;
        RECT 137.760 167.460 138.080 167.520 ;
        RECT 141.900 167.660 142.220 167.720 ;
        RECT 144.200 167.660 144.520 167.720 ;
        RECT 141.900 167.520 144.520 167.660 ;
        RECT 141.900 167.460 142.220 167.520 ;
        RECT 144.200 167.460 144.520 167.520 ;
        RECT 151.100 167.660 151.390 167.705 ;
        RECT 152.670 167.660 152.960 167.705 ;
        RECT 154.770 167.660 155.060 167.705 ;
        RECT 151.100 167.520 155.060 167.660 ;
        RECT 151.100 167.475 151.390 167.520 ;
        RECT 152.670 167.475 152.960 167.520 ;
        RECT 154.770 167.475 155.060 167.520 ;
        RECT 129.480 167.120 129.800 167.380 ;
        RECT 130.375 167.320 130.665 167.365 ;
        RECT 131.565 167.320 131.855 167.365 ;
        RECT 134.085 167.320 134.375 167.365 ;
        RECT 130.375 167.180 134.375 167.320 ;
        RECT 130.375 167.135 130.665 167.180 ;
        RECT 131.565 167.135 131.855 167.180 ;
        RECT 134.085 167.135 134.375 167.180 ;
        RECT 147.420 167.120 147.740 167.380 ;
        RECT 150.665 167.320 150.955 167.365 ;
        RECT 153.185 167.320 153.475 167.365 ;
        RECT 154.375 167.320 154.665 167.365 ;
        RECT 150.665 167.180 154.665 167.320 ;
        RECT 150.665 167.135 150.955 167.180 ;
        RECT 153.185 167.135 153.475 167.180 ;
        RECT 154.375 167.135 154.665 167.180 ;
        RECT 119.450 166.840 120.970 166.980 ;
        RECT 117.060 166.780 117.380 166.840 ;
        RECT 118.915 166.795 119.205 166.840 ;
        RECT 116.140 166.640 116.460 166.700 ;
        RECT 114.390 166.500 116.460 166.640 ;
        RECT 85.780 166.300 86.100 166.360 ;
        RECT 76.210 166.160 86.100 166.300 ;
        RECT 85.780 166.100 86.100 166.160 ;
        RECT 88.080 166.300 88.400 166.360 ;
        RECT 88.635 166.300 88.925 166.345 ;
        RECT 88.080 166.160 88.925 166.300 ;
        RECT 88.080 166.100 88.400 166.160 ;
        RECT 88.635 166.115 88.925 166.160 ;
        RECT 103.260 166.300 103.580 166.360 ;
        RECT 105.100 166.300 105.420 166.360 ;
        RECT 103.260 166.160 105.420 166.300 ;
        RECT 107.950 166.300 108.090 166.455 ;
        RECT 108.320 166.300 108.640 166.360 ;
        RECT 111.170 166.300 111.310 166.455 ;
        RECT 116.140 166.440 116.460 166.500 ;
        RECT 119.360 166.640 119.680 166.700 ;
        RECT 120.140 166.640 120.430 166.685 ;
        RECT 119.360 166.500 120.430 166.640 ;
        RECT 120.830 166.640 120.970 166.840 ;
        RECT 126.275 166.795 126.565 167.025 ;
        RECT 127.655 166.980 127.945 167.025 ;
        RECT 126.810 166.840 127.945 166.980 ;
        RECT 126.810 166.700 126.950 166.840 ;
        RECT 127.655 166.795 127.945 166.840 ;
        RECT 128.100 166.780 128.420 167.040 ;
        RECT 141.915 166.795 142.205 167.025 ;
        RECT 126.720 166.640 127.040 166.700 ;
        RECT 120.830 166.500 127.040 166.640 ;
        RECT 119.360 166.440 119.680 166.500 ;
        RECT 120.140 166.455 120.430 166.500 ;
        RECT 126.720 166.440 127.040 166.500 ;
        RECT 127.180 166.440 127.500 166.700 ;
        RECT 130.720 166.640 131.010 166.685 ;
        RECT 130.260 166.500 131.010 166.640 ;
        RECT 107.950 166.160 111.310 166.300 ;
        RECT 125.815 166.300 126.105 166.345 ;
        RECT 128.560 166.300 128.880 166.360 ;
        RECT 125.815 166.160 128.880 166.300 ;
        RECT 103.260 166.100 103.580 166.160 ;
        RECT 105.100 166.100 105.420 166.160 ;
        RECT 108.320 166.100 108.640 166.160 ;
        RECT 125.815 166.115 126.105 166.160 ;
        RECT 128.560 166.100 128.880 166.160 ;
        RECT 129.035 166.300 129.325 166.345 ;
        RECT 130.260 166.300 130.400 166.500 ;
        RECT 130.720 166.455 131.010 166.500 ;
        RECT 137.760 166.640 138.080 166.700 ;
        RECT 141.990 166.640 142.130 166.795 ;
        RECT 142.820 166.780 143.140 167.040 ;
        RECT 143.755 166.980 144.045 167.025 ;
        RECT 143.370 166.840 144.045 166.980 ;
        RECT 143.370 166.700 143.510 166.840 ;
        RECT 143.755 166.795 144.045 166.840 ;
        RECT 144.200 166.780 144.520 167.040 ;
        RECT 144.675 166.795 144.965 167.025 ;
        RECT 137.760 166.500 142.130 166.640 ;
        RECT 137.760 166.440 138.080 166.500 ;
        RECT 143.280 166.440 143.600 166.700 ;
        RECT 144.750 166.640 144.890 166.795 ;
        RECT 146.960 166.780 147.280 167.040 ;
        RECT 147.510 166.980 147.650 167.120 ;
        RECT 152.480 166.980 152.800 167.040 ;
        RECT 155.255 166.980 155.545 167.025 ;
        RECT 147.510 166.840 155.545 166.980 ;
        RECT 152.480 166.780 152.800 166.840 ;
        RECT 155.255 166.795 155.545 166.840 ;
        RECT 150.640 166.640 150.960 166.700 ;
        RECT 144.750 166.500 150.960 166.640 ;
        RECT 129.035 166.160 130.400 166.300 ;
        RECT 142.360 166.300 142.680 166.360 ;
        RECT 144.750 166.300 144.890 166.500 ;
        RECT 150.640 166.440 150.960 166.500 ;
        RECT 153.860 166.685 154.180 166.700 ;
        RECT 153.860 166.455 154.210 166.685 ;
        RECT 153.860 166.440 154.180 166.455 ;
        RECT 142.360 166.160 144.890 166.300 ;
        RECT 129.035 166.115 129.325 166.160 ;
        RECT 142.360 166.100 142.680 166.160 ;
        RECT 22.690 165.480 157.810 165.960 ;
        RECT 25.980 165.080 26.300 165.340 ;
        RECT 31.500 165.280 31.820 165.340 ;
        RECT 28.830 165.140 31.820 165.280 ;
        RECT 26.915 164.600 27.205 164.645 ;
        RECT 28.830 164.600 28.970 165.140 ;
        RECT 31.500 165.080 31.820 165.140 ;
        RECT 31.975 165.280 32.265 165.325 ;
        RECT 32.420 165.280 32.740 165.340 ;
        RECT 34.720 165.280 35.040 165.340 ;
        RECT 31.975 165.140 32.740 165.280 ;
        RECT 31.975 165.095 32.265 165.140 ;
        RECT 32.420 165.080 32.740 165.140 ;
        RECT 32.970 165.140 35.040 165.280 ;
        RECT 32.970 164.985 33.110 165.140 ;
        RECT 34.720 165.080 35.040 165.140 ;
        RECT 35.640 165.280 35.960 165.340 ;
        RECT 39.335 165.280 39.625 165.325 ;
        RECT 35.640 165.140 39.625 165.280 ;
        RECT 35.640 165.080 35.960 165.140 ;
        RECT 39.335 165.095 39.625 165.140 ;
        RECT 40.240 165.080 40.560 165.340 ;
        RECT 48.075 165.280 48.365 165.325 ;
        RECT 48.980 165.280 49.300 165.340 ;
        RECT 48.075 165.140 50.590 165.280 ;
        RECT 48.075 165.095 48.365 165.140 ;
        RECT 48.980 165.080 49.300 165.140 ;
        RECT 32.895 164.755 33.185 164.985 ;
        RECT 33.815 164.940 34.105 164.985 ;
        RECT 34.260 164.940 34.580 165.000 ;
        RECT 33.815 164.800 37.710 164.940 ;
        RECT 33.815 164.755 34.105 164.800 ;
        RECT 34.260 164.740 34.580 164.800 ;
        RECT 37.570 164.645 37.710 164.800 ;
        RECT 26.915 164.460 28.970 164.600 ;
        RECT 37.495 164.600 37.785 164.645 ;
        RECT 37.495 164.460 37.895 164.600 ;
        RECT 26.915 164.415 27.205 164.460 ;
        RECT 37.495 164.415 37.785 164.460 ;
        RECT 45.775 164.415 46.065 164.645 ;
        RECT 47.600 164.600 47.920 164.660 ;
        RECT 48.995 164.600 49.285 164.645 ;
        RECT 47.600 164.460 49.285 164.600 ;
        RECT 45.850 164.260 45.990 164.415 ;
        RECT 47.600 164.400 47.920 164.460 ;
        RECT 48.995 164.415 49.285 164.460 ;
        RECT 49.900 164.260 50.220 164.320 ;
        RECT 45.850 164.120 50.220 164.260 ;
        RECT 50.450 164.260 50.590 165.140 ;
        RECT 51.280 165.080 51.600 165.340 ;
        RECT 51.740 165.080 52.060 165.340 ;
        RECT 52.215 165.280 52.505 165.325 ;
        RECT 52.660 165.280 52.980 165.340 ;
        RECT 52.215 165.140 52.980 165.280 ;
        RECT 52.215 165.095 52.505 165.140 ;
        RECT 52.660 165.080 52.980 165.140 ;
        RECT 57.260 165.080 57.580 165.340 ;
        RECT 57.735 165.280 58.025 165.325 ;
        RECT 58.180 165.280 58.500 165.340 ;
        RECT 57.735 165.140 58.500 165.280 ;
        RECT 57.735 165.095 58.025 165.140 ;
        RECT 58.180 165.080 58.500 165.140 ;
        RECT 70.600 165.080 70.920 165.340 ;
        RECT 83.940 165.080 84.260 165.340 ;
        RECT 92.695 165.280 92.985 165.325 ;
        RECT 93.140 165.280 93.460 165.340 ;
        RECT 92.695 165.140 93.460 165.280 ;
        RECT 92.695 165.095 92.985 165.140 ;
        RECT 93.140 165.080 93.460 165.140 ;
        RECT 102.800 165.280 103.120 165.340 ;
        RECT 108.320 165.280 108.640 165.340 ;
        RECT 115.680 165.280 116.000 165.340 ;
        RECT 102.800 165.140 110.390 165.280 ;
        RECT 102.800 165.080 103.120 165.140 ;
        RECT 108.320 165.080 108.640 165.140 ;
        RECT 51.830 164.645 51.970 165.080 ;
        RECT 51.755 164.415 52.045 164.645 ;
        RECT 53.135 164.415 53.425 164.645 ;
        RECT 53.580 164.600 53.900 164.660 ;
        RECT 57.350 164.645 57.490 165.080 ;
        RECT 76.120 164.940 76.440 165.000 ;
        RECT 110.250 164.985 110.390 165.140 ;
        RECT 115.680 165.140 117.290 165.280 ;
        RECT 115.680 165.080 116.000 165.140 ;
        RECT 78.280 164.940 78.570 164.985 ;
        RECT 76.120 164.800 78.570 164.940 ;
        RECT 76.120 164.740 76.440 164.800 ;
        RECT 78.280 164.755 78.570 164.800 ;
        RECT 97.830 164.800 99.810 164.940 ;
        RECT 55.435 164.600 55.725 164.645 ;
        RECT 53.580 164.460 55.725 164.600 ;
        RECT 53.210 164.260 53.350 164.415 ;
        RECT 53.580 164.400 53.900 164.460 ;
        RECT 55.435 164.415 55.725 164.460 ;
        RECT 57.275 164.415 57.565 164.645 ;
        RECT 57.720 164.400 58.040 164.660 ;
        RECT 58.640 164.400 58.960 164.660 ;
        RECT 59.560 164.400 59.880 164.660 ;
        RECT 63.700 164.600 64.020 164.660 ;
        RECT 64.535 164.600 64.825 164.645 ;
        RECT 63.700 164.460 64.825 164.600 ;
        RECT 63.700 164.400 64.020 164.460 ;
        RECT 64.535 164.415 64.825 164.460 ;
        RECT 75.200 164.600 75.520 164.660 ;
        RECT 77.040 164.600 77.360 164.660 ;
        RECT 75.200 164.460 77.360 164.600 ;
        RECT 75.200 164.400 75.520 164.460 ;
        RECT 77.040 164.400 77.360 164.460 ;
        RECT 90.840 164.645 91.160 164.660 ;
        RECT 90.840 164.415 91.190 164.645 ;
        RECT 97.830 164.600 97.970 164.800 ;
        RECT 99.670 164.645 99.810 164.800 ;
        RECT 100.590 164.800 105.790 164.940 ;
        RECT 94.610 164.460 97.970 164.600 ;
        RECT 98.315 164.600 98.605 164.645 ;
        RECT 99.595 164.600 99.885 164.645 ;
        RECT 98.315 164.460 99.350 164.600 ;
        RECT 90.840 164.400 91.160 164.415 ;
        RECT 50.450 164.120 53.350 164.260 ;
        RECT 54.960 164.260 55.280 164.320 ;
        RECT 56.355 164.260 56.645 164.305 ;
        RECT 57.810 164.260 57.950 164.400 ;
        RECT 54.960 164.120 56.110 164.260 ;
        RECT 49.900 164.060 50.220 164.120 ;
        RECT 54.960 164.060 55.280 164.120 ;
        RECT 47.140 163.720 47.460 163.980 ;
        RECT 53.120 163.720 53.440 163.980 ;
        RECT 54.500 163.920 54.820 163.980 ;
        RECT 55.435 163.920 55.725 163.965 ;
        RECT 54.500 163.780 55.725 163.920 ;
        RECT 55.970 163.920 56.110 164.120 ;
        RECT 56.355 164.120 57.950 164.260 ;
        RECT 60.020 164.260 60.340 164.320 ;
        RECT 63.255 164.260 63.545 164.305 ;
        RECT 60.020 164.120 63.545 164.260 ;
        RECT 56.355 164.075 56.645 164.120 ;
        RECT 60.020 164.060 60.340 164.120 ;
        RECT 63.255 164.075 63.545 164.120 ;
        RECT 64.135 164.260 64.425 164.305 ;
        RECT 65.325 164.260 65.615 164.305 ;
        RECT 67.845 164.260 68.135 164.305 ;
        RECT 73.375 164.260 73.665 164.305 ;
        RECT 64.135 164.120 68.135 164.260 ;
        RECT 64.135 164.075 64.425 164.120 ;
        RECT 65.325 164.075 65.615 164.120 ;
        RECT 67.845 164.075 68.135 164.120 ;
        RECT 70.690 164.120 73.665 164.260 ;
        RECT 60.940 163.920 61.260 163.980 ;
        RECT 55.970 163.780 61.260 163.920 ;
        RECT 54.500 163.720 54.820 163.780 ;
        RECT 55.435 163.735 55.725 163.780 ;
        RECT 60.940 163.720 61.260 163.780 ;
        RECT 63.740 163.920 64.030 163.965 ;
        RECT 65.840 163.920 66.130 163.965 ;
        RECT 67.410 163.920 67.700 163.965 ;
        RECT 63.740 163.780 67.700 163.920 ;
        RECT 63.740 163.735 64.030 163.780 ;
        RECT 65.840 163.735 66.130 163.780 ;
        RECT 67.410 163.735 67.700 163.780 ;
        RECT 70.140 163.720 70.460 163.980 ;
        RECT 39.335 163.580 39.625 163.625 ;
        RECT 44.380 163.580 44.700 163.640 ;
        RECT 39.335 163.440 44.700 163.580 ;
        RECT 39.335 163.395 39.625 163.440 ;
        RECT 44.380 163.380 44.700 163.440 ;
        RECT 50.360 163.580 50.680 163.640 ;
        RECT 70.230 163.580 70.370 163.720 ;
        RECT 70.690 163.640 70.830 164.120 ;
        RECT 73.375 164.075 73.665 164.120 ;
        RECT 77.935 164.260 78.225 164.305 ;
        RECT 79.125 164.260 79.415 164.305 ;
        RECT 81.645 164.260 81.935 164.305 ;
        RECT 77.935 164.120 81.935 164.260 ;
        RECT 77.935 164.075 78.225 164.120 ;
        RECT 79.125 164.075 79.415 164.120 ;
        RECT 81.645 164.075 81.935 164.120 ;
        RECT 87.645 164.260 87.935 164.305 ;
        RECT 90.165 164.260 90.455 164.305 ;
        RECT 91.355 164.260 91.645 164.305 ;
        RECT 87.645 164.120 91.645 164.260 ;
        RECT 87.645 164.075 87.935 164.120 ;
        RECT 90.165 164.075 90.455 164.120 ;
        RECT 91.355 164.075 91.645 164.120 ;
        RECT 92.235 164.075 92.525 164.305 ;
        RECT 77.540 163.920 77.830 163.965 ;
        RECT 79.640 163.920 79.930 163.965 ;
        RECT 81.210 163.920 81.500 163.965 ;
        RECT 77.540 163.780 81.500 163.920 ;
        RECT 77.540 163.735 77.830 163.780 ;
        RECT 79.640 163.735 79.930 163.780 ;
        RECT 81.210 163.735 81.500 163.780 ;
        RECT 88.080 163.920 88.370 163.965 ;
        RECT 89.650 163.920 89.940 163.965 ;
        RECT 91.750 163.920 92.040 163.965 ;
        RECT 88.080 163.780 92.040 163.920 ;
        RECT 88.080 163.735 88.370 163.780 ;
        RECT 89.650 163.735 89.940 163.780 ;
        RECT 91.750 163.735 92.040 163.780 ;
        RECT 50.360 163.440 70.370 163.580 ;
        RECT 50.360 163.380 50.680 163.440 ;
        RECT 70.600 163.380 70.920 163.640 ;
        RECT 85.335 163.580 85.625 163.625 ;
        RECT 89.000 163.580 89.320 163.640 ;
        RECT 85.335 163.440 89.320 163.580 ;
        RECT 92.310 163.580 92.450 164.075 ;
        RECT 94.610 163.580 94.750 164.460 ;
        RECT 98.315 164.415 98.605 164.460 ;
        RECT 95.005 164.260 95.295 164.305 ;
        RECT 97.525 164.260 97.815 164.305 ;
        RECT 98.715 164.260 99.005 164.305 ;
        RECT 95.005 164.120 99.005 164.260 ;
        RECT 99.210 164.260 99.350 164.460 ;
        RECT 99.595 164.460 99.995 164.600 ;
        RECT 99.595 164.415 99.885 164.460 ;
        RECT 100.590 164.320 100.730 164.800 ;
        RECT 101.895 164.415 102.185 164.645 ;
        RECT 99.210 164.120 100.270 164.260 ;
        RECT 95.005 164.075 95.295 164.120 ;
        RECT 97.525 164.075 97.815 164.120 ;
        RECT 98.715 164.075 99.005 164.120 ;
        RECT 95.440 163.920 95.730 163.965 ;
        RECT 97.010 163.920 97.300 163.965 ;
        RECT 99.110 163.920 99.400 163.965 ;
        RECT 95.440 163.780 99.400 163.920 ;
        RECT 100.130 163.920 100.270 164.120 ;
        RECT 100.500 164.060 100.820 164.320 ;
        RECT 101.420 164.260 101.740 164.320 ;
        RECT 101.970 164.260 102.110 164.415 ;
        RECT 102.800 164.400 103.120 164.660 ;
        RECT 103.260 164.400 103.580 164.660 ;
        RECT 104.180 164.400 104.500 164.660 ;
        RECT 105.650 164.645 105.790 164.800 ;
        RECT 110.175 164.755 110.465 164.985 ;
        RECT 115.770 164.940 115.910 165.080 ;
        RECT 113.470 164.800 115.910 164.940 ;
        RECT 104.655 164.415 104.945 164.645 ;
        RECT 105.575 164.600 105.865 164.645 ;
        RECT 108.780 164.600 109.100 164.660 ;
        RECT 109.255 164.600 109.545 164.645 ;
        RECT 105.575 164.460 108.090 164.600 ;
        RECT 105.575 164.415 105.865 164.460 ;
        RECT 101.420 164.120 102.110 164.260 ;
        RECT 101.420 164.060 101.740 164.120 ;
        RECT 103.735 163.920 104.025 163.965 ;
        RECT 100.130 163.780 104.025 163.920 ;
        RECT 95.440 163.735 95.730 163.780 ;
        RECT 97.010 163.735 97.300 163.780 ;
        RECT 99.110 163.735 99.400 163.780 ;
        RECT 103.735 163.735 104.025 163.780 ;
        RECT 98.660 163.580 98.980 163.640 ;
        RECT 92.310 163.440 98.980 163.580 ;
        RECT 85.335 163.395 85.625 163.440 ;
        RECT 89.000 163.380 89.320 163.440 ;
        RECT 98.660 163.380 98.980 163.440 ;
        RECT 100.960 163.580 101.280 163.640 ;
        RECT 104.730 163.580 104.870 164.415 ;
        RECT 105.115 164.075 105.405 164.305 ;
        RECT 105.190 163.920 105.330 164.075 ;
        RECT 106.940 163.920 107.260 163.980 ;
        RECT 105.190 163.780 107.260 163.920 ;
        RECT 107.950 163.920 108.090 164.460 ;
        RECT 108.780 164.460 109.545 164.600 ;
        RECT 108.780 164.400 109.100 164.460 ;
        RECT 109.255 164.415 109.545 164.460 ;
        RECT 109.715 164.415 110.005 164.645 ;
        RECT 111.095 164.600 111.385 164.645 ;
        RECT 112.935 164.600 113.225 164.645 ;
        RECT 111.095 164.460 113.225 164.600 ;
        RECT 111.095 164.415 111.385 164.460 ;
        RECT 112.935 164.415 113.225 164.460 ;
        RECT 109.790 164.260 109.930 164.415 ;
        RECT 113.470 164.320 113.610 164.800 ;
        RECT 115.220 164.600 115.540 164.660 ;
        RECT 117.150 164.645 117.290 165.140 ;
        RECT 117.980 165.080 118.300 165.340 ;
        RECT 119.360 165.080 119.680 165.340 ;
        RECT 121.660 165.280 121.980 165.340 ;
        RECT 142.360 165.280 142.680 165.340 ;
        RECT 121.660 165.140 142.680 165.280 ;
        RECT 121.660 165.080 121.980 165.140 ;
        RECT 142.360 165.080 142.680 165.140 ;
        RECT 153.860 165.280 154.180 165.340 ;
        RECT 154.335 165.280 154.625 165.325 ;
        RECT 153.860 165.140 154.625 165.280 ;
        RECT 153.860 165.080 154.180 165.140 ;
        RECT 154.335 165.095 154.625 165.140 ;
        RECT 149.260 164.940 149.580 165.000 ;
        RECT 152.035 164.940 152.325 164.985 ;
        RECT 120.215 164.800 128.330 164.940 ;
        RECT 117.075 164.600 117.365 164.645 ;
        RECT 115.220 164.460 116.830 164.600 ;
        RECT 115.220 164.400 115.540 164.460 ;
        RECT 110.160 164.260 110.480 164.320 ;
        RECT 112.460 164.260 112.780 164.320 ;
        RECT 109.790 164.120 112.780 164.260 ;
        RECT 110.160 164.060 110.480 164.120 ;
        RECT 112.460 164.060 112.780 164.120 ;
        RECT 113.380 164.060 113.700 164.320 ;
        RECT 116.140 164.060 116.460 164.320 ;
        RECT 116.690 164.260 116.830 164.460 ;
        RECT 117.075 164.460 117.475 164.600 ;
        RECT 117.075 164.415 117.365 164.460 ;
        RECT 117.995 164.415 118.285 164.645 ;
        RECT 119.360 164.600 119.680 164.660 ;
        RECT 120.215 164.645 120.355 164.800 ;
        RECT 128.190 164.660 128.330 164.800 ;
        RECT 148.430 164.800 152.325 164.940 ;
        RECT 120.175 164.600 120.465 164.645 ;
        RECT 119.360 164.460 120.465 164.600 ;
        RECT 118.070 164.260 118.210 164.415 ;
        RECT 119.360 164.400 119.680 164.460 ;
        RECT 120.175 164.415 120.465 164.460 ;
        RECT 120.755 164.415 121.045 164.645 ;
        RECT 121.215 164.415 121.505 164.645 ;
        RECT 122.135 164.600 122.425 164.645 ;
        RECT 126.275 164.600 126.565 164.645 ;
        RECT 122.135 164.460 126.565 164.600 ;
        RECT 122.135 164.415 122.425 164.460 ;
        RECT 126.275 164.415 126.565 164.460 ;
        RECT 116.690 164.120 118.210 164.260 ;
        RECT 115.680 163.920 116.000 163.980 ;
        RECT 107.950 163.780 116.000 163.920 ;
        RECT 106.940 163.720 107.260 163.780 ;
        RECT 115.680 163.720 116.000 163.780 ;
        RECT 119.820 163.920 120.140 163.980 ;
        RECT 120.850 163.920 120.990 164.415 ;
        RECT 121.290 164.260 121.430 164.415 ;
        RECT 126.720 164.400 127.040 164.660 ;
        RECT 127.180 164.400 127.500 164.660 ;
        RECT 128.100 164.400 128.420 164.660 ;
        RECT 128.560 164.600 128.880 164.660 ;
        RECT 129.035 164.600 129.325 164.645 ;
        RECT 141.900 164.600 142.220 164.660 ;
        RECT 148.430 164.645 148.570 164.800 ;
        RECT 149.260 164.740 149.580 164.800 ;
        RECT 152.035 164.755 152.325 164.800 ;
        RECT 153.115 164.940 153.405 164.985 ;
        RECT 154.780 164.940 155.100 165.000 ;
        RECT 153.115 164.800 155.100 164.940 ;
        RECT 153.115 164.755 153.405 164.800 ;
        RECT 154.780 164.740 155.100 164.800 ;
        RECT 128.560 164.460 142.220 164.600 ;
        RECT 128.560 164.400 128.880 164.460 ;
        RECT 129.035 164.415 129.325 164.460 ;
        RECT 141.900 164.400 142.220 164.460 ;
        RECT 144.215 164.600 144.505 164.645 ;
        RECT 144.675 164.600 144.965 164.645 ;
        RECT 144.215 164.460 144.965 164.600 ;
        RECT 144.215 164.415 144.505 164.460 ;
        RECT 144.675 164.415 144.965 164.460 ;
        RECT 148.355 164.415 148.645 164.645 ;
        RECT 150.195 164.415 150.485 164.645 ;
        RECT 150.655 164.600 150.945 164.645 ;
        RECT 150.655 164.460 152.250 164.600 ;
        RECT 150.655 164.415 150.945 164.460 ;
        RECT 126.810 164.260 126.950 164.400 ;
        RECT 121.290 164.120 126.950 164.260 ;
        RECT 124.420 163.920 124.740 163.980 ;
        RECT 119.820 163.780 124.740 163.920 ;
        RECT 119.820 163.720 120.140 163.780 ;
        RECT 124.420 163.720 124.740 163.780 ;
        RECT 100.960 163.440 104.870 163.580 ;
        RECT 108.335 163.580 108.625 163.625 ;
        RECT 109.240 163.580 109.560 163.640 ;
        RECT 108.335 163.440 109.560 163.580 ;
        RECT 100.960 163.380 101.280 163.440 ;
        RECT 108.335 163.395 108.625 163.440 ;
        RECT 109.240 163.380 109.560 163.440 ;
        RECT 125.340 163.580 125.660 163.640 ;
        RECT 127.270 163.580 127.410 164.400 ;
        RECT 134.540 164.060 134.860 164.320 ;
        RECT 137.760 164.060 138.080 164.320 ;
        RECT 147.420 164.060 147.740 164.320 ;
        RECT 129.020 163.920 129.340 163.980 ;
        RECT 135.015 163.920 135.305 163.965 ;
        RECT 129.020 163.780 135.305 163.920 ;
        RECT 129.020 163.720 129.340 163.780 ;
        RECT 135.015 163.735 135.305 163.780 ;
        RECT 141.900 163.920 142.220 163.980 ;
        RECT 143.755 163.920 144.045 163.965 ;
        RECT 150.270 163.920 150.410 164.415 ;
        RECT 141.900 163.780 150.410 163.920 ;
        RECT 141.900 163.720 142.220 163.780 ;
        RECT 143.755 163.735 144.045 163.780 ;
        RECT 152.110 163.640 152.250 164.460 ;
        RECT 155.255 164.415 155.545 164.645 ;
        RECT 153.875 163.920 154.165 163.965 ;
        RECT 155.330 163.920 155.470 164.415 ;
        RECT 153.875 163.780 155.470 163.920 ;
        RECT 153.875 163.735 154.165 163.780 ;
        RECT 125.340 163.440 127.410 163.580 ;
        RECT 127.640 163.580 127.960 163.640 ;
        RECT 131.335 163.580 131.625 163.625 ;
        RECT 127.640 163.440 131.625 163.580 ;
        RECT 125.340 163.380 125.660 163.440 ;
        RECT 127.640 163.380 127.960 163.440 ;
        RECT 131.335 163.395 131.625 163.440 ;
        RECT 149.260 163.380 149.580 163.640 ;
        RECT 152.020 163.580 152.340 163.640 ;
        RECT 152.955 163.580 153.245 163.625 ;
        RECT 152.020 163.440 153.245 163.580 ;
        RECT 152.020 163.380 152.340 163.440 ;
        RECT 152.955 163.395 153.245 163.440 ;
        RECT 22.690 162.760 157.010 163.240 ;
        RECT 38.860 162.560 39.180 162.620 ;
        RECT 39.335 162.560 39.625 162.605 ;
        RECT 37.570 162.420 39.625 162.560 ;
        RECT 37.570 162.280 37.710 162.420 ;
        RECT 38.860 162.360 39.180 162.420 ;
        RECT 39.335 162.375 39.625 162.420 ;
        RECT 41.175 162.560 41.465 162.605 ;
        RECT 46.220 162.560 46.540 162.620 ;
        RECT 41.175 162.420 46.540 162.560 ;
        RECT 41.175 162.375 41.465 162.420 ;
        RECT 46.220 162.360 46.540 162.420 ;
        RECT 49.900 162.560 50.220 162.620 ;
        RECT 54.960 162.560 55.280 162.620 ;
        RECT 49.900 162.420 55.280 162.560 ;
        RECT 49.900 162.360 50.220 162.420 ;
        RECT 54.960 162.360 55.280 162.420 ;
        RECT 58.640 162.360 58.960 162.620 ;
        RECT 59.115 162.375 59.405 162.605 ;
        RECT 26.455 162.220 26.745 162.265 ;
        RECT 26.455 162.080 28.050 162.220 ;
        RECT 26.455 162.035 26.745 162.080 ;
        RECT 27.375 161.880 27.665 161.925 ;
        RECT 25.150 161.740 27.665 161.880 ;
        RECT 25.150 161.585 25.290 161.740 ;
        RECT 27.375 161.695 27.665 161.740 ;
        RECT 27.910 161.600 28.050 162.080 ;
        RECT 37.480 162.020 37.800 162.280 ;
        RECT 54.515 162.220 54.805 162.265 ;
        RECT 58.730 162.220 58.870 162.360 ;
        RECT 54.515 162.080 58.870 162.220 ;
        RECT 54.515 162.035 54.805 162.080 ;
        RECT 28.295 161.880 28.585 161.925 ;
        RECT 45.760 161.880 46.080 161.940 ;
        RECT 47.600 161.880 47.920 161.940 ;
        RECT 28.295 161.740 32.190 161.880 ;
        RECT 28.295 161.695 28.585 161.740 ;
        RECT 32.050 161.600 32.190 161.740 ;
        RECT 37.570 161.740 39.550 161.880 ;
        RECT 25.075 161.355 25.365 161.585 ;
        RECT 26.915 161.540 27.205 161.585 ;
        RECT 26.070 161.400 27.205 161.540 ;
        RECT 25.150 160.920 25.290 161.355 ;
        RECT 25.060 160.660 25.380 160.920 ;
        RECT 25.535 160.860 25.825 160.905 ;
        RECT 26.070 160.860 26.210 161.400 ;
        RECT 26.915 161.355 27.205 161.400 ;
        RECT 27.820 161.340 28.140 161.600 ;
        RECT 31.040 161.540 31.360 161.600 ;
        RECT 31.515 161.540 31.805 161.585 ;
        RECT 31.040 161.400 31.805 161.540 ;
        RECT 31.040 161.340 31.360 161.400 ;
        RECT 31.515 161.355 31.805 161.400 ;
        RECT 26.455 161.200 26.745 161.245 ;
        RECT 28.295 161.200 28.585 161.245 ;
        RECT 26.455 161.060 28.585 161.200 ;
        RECT 31.590 161.200 31.730 161.355 ;
        RECT 31.960 161.340 32.280 161.600 ;
        RECT 32.435 161.540 32.725 161.585 ;
        RECT 33.800 161.540 34.120 161.600 ;
        RECT 32.435 161.400 34.120 161.540 ;
        RECT 32.435 161.355 32.725 161.400 ;
        RECT 33.800 161.340 34.120 161.400 ;
        RECT 37.020 161.540 37.340 161.600 ;
        RECT 37.570 161.585 37.710 161.740 ;
        RECT 37.495 161.540 37.785 161.585 ;
        RECT 37.020 161.400 37.785 161.540 ;
        RECT 37.020 161.340 37.340 161.400 ;
        RECT 37.495 161.355 37.785 161.400 ;
        RECT 38.860 161.340 39.180 161.600 ;
        RECT 39.410 161.585 39.550 161.740 ;
        RECT 44.470 161.740 47.920 161.880 ;
        RECT 44.470 161.585 44.610 161.740 ;
        RECT 45.760 161.680 46.080 161.740 ;
        RECT 47.600 161.680 47.920 161.740 ;
        RECT 58.640 161.880 58.960 161.940 ;
        RECT 59.190 161.880 59.330 162.375 ;
        RECT 60.940 162.360 61.260 162.620 ;
        RECT 63.700 162.360 64.020 162.620 ;
        RECT 80.275 162.560 80.565 162.605 ;
        RECT 81.180 162.560 81.500 162.620 ;
        RECT 80.275 162.420 81.500 162.560 ;
        RECT 80.275 162.375 80.565 162.420 ;
        RECT 81.180 162.360 81.500 162.420 ;
        RECT 88.080 162.360 88.400 162.620 ;
        RECT 90.840 162.360 91.160 162.620 ;
        RECT 100.055 162.560 100.345 162.605 ;
        RECT 103.260 162.560 103.580 162.620 ;
        RECT 116.600 162.560 116.920 162.620 ;
        RECT 100.055 162.420 103.580 162.560 ;
        RECT 100.055 162.375 100.345 162.420 ;
        RECT 103.260 162.360 103.580 162.420 ;
        RECT 105.650 162.420 116.920 162.560 ;
        RECT 61.030 162.220 61.170 162.360 ;
        RECT 70.155 162.220 70.445 162.265 ;
        RECT 70.600 162.220 70.920 162.280 ;
        RECT 61.030 162.080 70.920 162.220 ;
        RECT 70.155 162.035 70.445 162.080 ;
        RECT 70.600 162.020 70.920 162.080 ;
        RECT 72.900 162.220 73.190 162.265 ;
        RECT 74.470 162.220 74.760 162.265 ;
        RECT 76.570 162.220 76.860 162.265 ;
        RECT 100.960 162.220 101.280 162.280 ;
        RECT 72.900 162.080 76.860 162.220 ;
        RECT 72.900 162.035 73.190 162.080 ;
        RECT 74.470 162.035 74.760 162.080 ;
        RECT 76.570 162.035 76.860 162.080 ;
        RECT 84.490 162.080 101.280 162.220 ;
        RECT 84.490 161.940 84.630 162.080 ;
        RECT 100.960 162.020 101.280 162.080 ;
        RECT 101.420 162.220 101.740 162.280 ;
        RECT 105.650 162.220 105.790 162.420 ;
        RECT 116.600 162.360 116.920 162.420 ;
        RECT 119.360 162.360 119.680 162.620 ;
        RECT 127.640 162.360 127.960 162.620 ;
        RECT 137.760 162.360 138.080 162.620 ;
        RECT 142.375 162.560 142.665 162.605 ;
        RECT 143.280 162.560 143.600 162.620 ;
        RECT 142.375 162.420 143.600 162.560 ;
        RECT 142.375 162.375 142.665 162.420 ;
        RECT 143.280 162.360 143.600 162.420 ;
        RECT 145.135 162.560 145.425 162.605 ;
        RECT 145.580 162.560 145.900 162.620 ;
        RECT 145.135 162.420 145.900 162.560 ;
        RECT 145.135 162.375 145.425 162.420 ;
        RECT 145.580 162.360 145.900 162.420 ;
        RECT 147.420 162.360 147.740 162.620 ;
        RECT 148.340 162.360 148.660 162.620 ;
        RECT 152.480 162.560 152.800 162.620 ;
        RECT 152.955 162.560 153.245 162.605 ;
        RECT 152.480 162.420 153.245 162.560 ;
        RECT 152.480 162.360 152.800 162.420 ;
        RECT 152.955 162.375 153.245 162.420 ;
        RECT 101.420 162.080 105.790 162.220 ;
        RECT 106.020 162.220 106.310 162.265 ;
        RECT 107.590 162.220 107.880 162.265 ;
        RECT 109.690 162.220 109.980 162.265 ;
        RECT 106.020 162.080 109.980 162.220 ;
        RECT 101.420 162.020 101.740 162.080 ;
        RECT 106.020 162.035 106.310 162.080 ;
        RECT 107.590 162.035 107.880 162.080 ;
        RECT 109.690 162.035 109.980 162.080 ;
        RECT 111.540 162.220 111.860 162.280 ;
        RECT 115.220 162.220 115.540 162.280 ;
        RECT 116.155 162.220 116.445 162.265 ;
        RECT 111.540 162.080 119.590 162.220 ;
        RECT 111.540 162.020 111.860 162.080 ;
        RECT 115.220 162.020 115.540 162.080 ;
        RECT 116.155 162.035 116.445 162.080 ;
        RECT 67.840 161.880 68.160 161.940 ;
        RECT 71.060 161.880 71.380 161.940 ;
        RECT 71.980 161.880 72.300 161.940 ;
        RECT 58.640 161.740 59.330 161.880 ;
        RECT 65.630 161.740 72.300 161.880 ;
        RECT 58.640 161.680 58.960 161.740 ;
        RECT 39.335 161.355 39.625 161.585 ;
        RECT 39.795 161.355 40.085 161.585 ;
        RECT 44.395 161.355 44.685 161.585 ;
        RECT 38.415 161.200 38.705 161.245 ;
        RECT 39.870 161.200 40.010 161.355 ;
        RECT 44.840 161.340 45.160 161.600 ;
        RECT 54.960 161.540 55.280 161.600 ;
        RECT 55.435 161.540 55.725 161.585 ;
        RECT 54.960 161.400 55.725 161.540 ;
        RECT 54.960 161.340 55.280 161.400 ;
        RECT 55.435 161.355 55.725 161.400 ;
        RECT 56.815 161.540 57.105 161.585 ;
        RECT 56.815 161.400 58.410 161.540 ;
        RECT 56.815 161.355 57.105 161.400 ;
        RECT 31.590 161.060 40.010 161.200 ;
        RECT 45.775 161.200 46.065 161.245 ;
        RECT 47.140 161.200 47.460 161.260 ;
        RECT 45.775 161.060 47.460 161.200 ;
        RECT 26.455 161.015 26.745 161.060 ;
        RECT 28.295 161.015 28.585 161.060 ;
        RECT 38.415 161.015 38.705 161.060 ;
        RECT 45.775 161.015 46.065 161.060 ;
        RECT 47.140 161.000 47.460 161.060 ;
        RECT 56.355 161.200 56.645 161.245 ;
        RECT 57.720 161.200 58.040 161.260 ;
        RECT 56.355 161.060 58.040 161.200 ;
        RECT 56.355 161.015 56.645 161.060 ;
        RECT 57.720 161.000 58.040 161.060 ;
        RECT 58.270 160.920 58.410 161.400 ;
        RECT 59.575 161.355 59.865 161.585 ;
        RECT 64.160 161.540 64.480 161.600 ;
        RECT 65.630 161.585 65.770 161.740 ;
        RECT 67.840 161.680 68.160 161.740 ;
        RECT 71.060 161.680 71.380 161.740 ;
        RECT 71.980 161.680 72.300 161.740 ;
        RECT 72.465 161.880 72.755 161.925 ;
        RECT 74.985 161.880 75.275 161.925 ;
        RECT 76.175 161.880 76.465 161.925 ;
        RECT 72.465 161.740 76.465 161.880 ;
        RECT 72.465 161.695 72.755 161.740 ;
        RECT 74.985 161.695 75.275 161.740 ;
        RECT 76.175 161.695 76.465 161.740 ;
        RECT 84.400 161.680 84.720 161.940 ;
        RECT 93.140 161.880 93.460 161.940 ;
        RECT 94.075 161.880 94.365 161.925 ;
        RECT 90.010 161.740 94.365 161.880 ;
        RECT 64.635 161.540 64.925 161.585 ;
        RECT 64.160 161.400 64.925 161.540 ;
        RECT 59.650 160.920 59.790 161.355 ;
        RECT 64.160 161.340 64.480 161.400 ;
        RECT 64.635 161.355 64.925 161.400 ;
        RECT 65.555 161.355 65.845 161.585 ;
        RECT 66.475 161.540 66.765 161.585 ;
        RECT 68.300 161.540 68.620 161.600 ;
        RECT 66.475 161.400 68.620 161.540 ;
        RECT 66.475 161.355 66.765 161.400 ;
        RECT 68.300 161.340 68.620 161.400 ;
        RECT 75.660 161.585 75.980 161.600 ;
        RECT 75.660 161.355 76.010 161.585 ;
        RECT 77.040 161.540 77.360 161.600 ;
        RECT 78.880 161.540 79.200 161.600 ;
        RECT 77.040 161.400 79.200 161.540 ;
        RECT 75.660 161.340 75.980 161.355 ;
        RECT 77.040 161.340 77.360 161.400 ;
        RECT 78.880 161.340 79.200 161.400 ;
        RECT 81.195 161.355 81.485 161.585 ;
        RECT 65.095 161.200 65.385 161.245 ;
        RECT 66.000 161.200 66.320 161.260 ;
        RECT 69.220 161.200 69.540 161.260 ;
        RECT 74.740 161.200 75.060 161.260 ;
        RECT 65.095 161.060 75.060 161.200 ;
        RECT 81.270 161.200 81.410 161.355 ;
        RECT 82.100 161.340 82.420 161.600 ;
        RECT 82.575 161.540 82.865 161.585 ;
        RECT 84.490 161.540 84.630 161.680 ;
        RECT 82.575 161.400 84.630 161.540 ;
        RECT 82.575 161.355 82.865 161.400 ;
        RECT 89.000 161.340 89.320 161.600 ;
        RECT 90.010 161.585 90.150 161.740 ;
        RECT 93.140 161.680 93.460 161.740 ;
        RECT 94.075 161.695 94.365 161.740 ;
        RECT 99.135 161.880 99.425 161.925 ;
        RECT 105.585 161.880 105.875 161.925 ;
        RECT 108.105 161.880 108.395 161.925 ;
        RECT 109.295 161.880 109.585 161.925 ;
        RECT 99.135 161.740 104.870 161.880 ;
        RECT 99.135 161.695 99.425 161.740 ;
        RECT 89.935 161.355 90.225 161.585 ;
        RECT 90.395 161.355 90.685 161.585 ;
        RECT 83.940 161.200 84.260 161.260 ;
        RECT 81.270 161.060 84.260 161.200 ;
        RECT 90.470 161.200 90.610 161.355 ;
        RECT 91.760 161.340 92.080 161.600 ;
        RECT 97.295 161.540 97.585 161.585 ;
        RECT 98.675 161.540 98.965 161.585 ;
        RECT 97.295 161.400 98.965 161.540 ;
        RECT 97.295 161.355 97.585 161.400 ;
        RECT 98.675 161.355 98.965 161.400 ;
        RECT 90.840 161.200 91.160 161.260 ;
        RECT 99.210 161.200 99.350 161.695 ;
        RECT 90.470 161.060 99.350 161.200 ;
        RECT 65.095 161.015 65.385 161.060 ;
        RECT 66.000 161.000 66.320 161.060 ;
        RECT 69.220 161.000 69.540 161.060 ;
        RECT 74.740 161.000 75.060 161.060 ;
        RECT 83.940 161.000 84.260 161.060 ;
        RECT 90.840 161.000 91.160 161.060 ;
        RECT 28.755 160.860 29.045 160.905 ;
        RECT 25.535 160.720 29.045 160.860 ;
        RECT 25.535 160.675 25.825 160.720 ;
        RECT 28.755 160.675 29.045 160.720 ;
        RECT 33.340 160.660 33.660 160.920 ;
        RECT 36.560 160.660 36.880 160.920 ;
        RECT 44.380 160.660 44.700 160.920 ;
        RECT 57.260 160.660 57.580 160.920 ;
        RECT 58.180 160.660 58.500 160.920 ;
        RECT 59.560 160.660 59.880 160.920 ;
        RECT 84.030 160.860 84.170 161.000 ;
        RECT 91.300 160.860 91.620 160.920 ;
        RECT 84.030 160.720 91.620 160.860 ;
        RECT 91.300 160.660 91.620 160.720 ;
        RECT 91.760 160.860 92.080 160.920 ;
        RECT 100.500 160.860 100.820 160.920 ;
        RECT 91.760 160.720 100.820 160.860 ;
        RECT 91.760 160.660 92.080 160.720 ;
        RECT 100.500 160.660 100.820 160.720 ;
        RECT 103.275 160.860 103.565 160.905 ;
        RECT 104.180 160.860 104.500 160.920 ;
        RECT 103.275 160.720 104.500 160.860 ;
        RECT 104.730 160.860 104.870 161.740 ;
        RECT 105.585 161.740 109.585 161.880 ;
        RECT 105.585 161.695 105.875 161.740 ;
        RECT 108.105 161.695 108.395 161.740 ;
        RECT 109.295 161.695 109.585 161.740 ;
        RECT 115.680 161.880 116.000 161.940 ;
        RECT 115.680 161.740 118.670 161.880 ;
        RECT 115.680 161.680 116.000 161.740 ;
        RECT 109.700 161.540 110.020 161.600 ;
        RECT 110.175 161.540 110.465 161.585 ;
        RECT 109.700 161.400 110.465 161.540 ;
        RECT 109.700 161.340 110.020 161.400 ;
        RECT 110.175 161.355 110.465 161.400 ;
        RECT 116.600 161.540 116.920 161.600 ;
        RECT 118.530 161.585 118.670 161.740 ;
        RECT 119.450 161.585 119.590 162.080 ;
        RECT 127.730 161.880 127.870 162.360 ;
        RECT 129.520 162.220 129.810 162.265 ;
        RECT 131.620 162.220 131.910 162.265 ;
        RECT 133.190 162.220 133.480 162.265 ;
        RECT 129.520 162.080 133.480 162.220 ;
        RECT 129.520 162.035 129.810 162.080 ;
        RECT 131.620 162.035 131.910 162.080 ;
        RECT 133.190 162.035 133.480 162.080 ;
        RECT 135.935 162.220 136.225 162.265 ;
        RECT 137.850 162.220 137.990 162.360 ;
        RECT 135.935 162.080 137.990 162.220 ;
        RECT 135.935 162.035 136.225 162.080 ;
        RECT 125.890 161.740 127.870 161.880 ;
        RECT 129.915 161.880 130.205 161.925 ;
        RECT 131.105 161.880 131.395 161.925 ;
        RECT 133.625 161.880 133.915 161.925 ;
        RECT 137.850 161.880 137.990 162.080 ;
        RECT 144.675 162.220 144.965 162.265 ;
        RECT 147.510 162.220 147.650 162.360 ;
        RECT 144.675 162.080 147.650 162.220 ;
        RECT 144.675 162.035 144.965 162.080 ;
        RECT 129.915 161.740 133.915 161.880 ;
        RECT 125.890 161.585 126.030 161.740 ;
        RECT 129.915 161.695 130.205 161.740 ;
        RECT 131.105 161.695 131.395 161.740 ;
        RECT 133.625 161.695 133.915 161.740 ;
        RECT 137.390 161.740 137.990 161.880 ;
        RECT 139.615 161.880 139.905 161.925 ;
        RECT 140.060 161.880 140.380 161.940 ;
        RECT 148.430 161.880 148.570 162.360 ;
        RECT 139.615 161.740 148.570 161.880 ;
        RECT 117.075 161.540 117.365 161.585 ;
        RECT 116.600 161.400 117.365 161.540 ;
        RECT 116.600 161.340 116.920 161.400 ;
        RECT 117.075 161.355 117.365 161.400 ;
        RECT 118.455 161.355 118.745 161.585 ;
        RECT 119.375 161.355 119.665 161.585 ;
        RECT 125.815 161.355 126.105 161.585 ;
        RECT 126.720 161.340 127.040 161.600 ;
        RECT 127.655 161.540 127.945 161.585 ;
        RECT 128.100 161.540 128.420 161.600 ;
        RECT 137.390 161.585 137.530 161.740 ;
        RECT 139.615 161.695 139.905 161.740 ;
        RECT 140.060 161.680 140.380 161.740 ;
        RECT 127.655 161.400 128.420 161.540 ;
        RECT 127.655 161.355 127.945 161.400 ;
        RECT 128.100 161.340 128.420 161.400 ;
        RECT 129.035 161.355 129.325 161.585 ;
        RECT 137.315 161.355 137.605 161.585 ;
        RECT 137.775 161.540 138.065 161.585 ;
        RECT 139.140 161.540 139.460 161.600 ;
        RECT 141.900 161.585 142.220 161.600 ;
        RECT 137.775 161.400 139.460 161.540 ;
        RECT 137.775 161.355 138.065 161.400 ;
        RECT 108.950 161.200 109.240 161.245 ;
        RECT 110.620 161.200 110.940 161.260 ;
        RECT 108.950 161.060 110.940 161.200 ;
        RECT 108.950 161.015 109.240 161.060 ;
        RECT 110.620 161.000 110.940 161.060 ;
        RECT 117.995 161.200 118.285 161.245 ;
        RECT 126.810 161.200 126.950 161.340 ;
        RECT 117.995 161.060 126.950 161.200 ;
        RECT 117.995 161.015 118.285 161.060 ;
        RECT 127.195 161.015 127.485 161.245 ;
        RECT 121.660 160.860 121.980 160.920 ;
        RECT 104.730 160.720 121.980 160.860 ;
        RECT 103.275 160.675 103.565 160.720 ;
        RECT 104.180 160.660 104.500 160.720 ;
        RECT 121.660 160.660 121.980 160.720 ;
        RECT 122.120 160.860 122.440 160.920 ;
        RECT 127.270 160.860 127.410 161.015 ;
        RECT 122.120 160.720 127.410 160.860 ;
        RECT 122.120 160.660 122.440 160.720 ;
        RECT 128.560 160.660 128.880 160.920 ;
        RECT 129.110 160.860 129.250 161.355 ;
        RECT 139.140 161.340 139.460 161.400 ;
        RECT 141.750 161.355 142.220 161.585 ;
        RECT 141.900 161.340 142.220 161.355 ;
        RECT 146.500 161.340 146.820 161.600 ;
        RECT 129.480 161.200 129.800 161.260 ;
        RECT 130.260 161.200 130.550 161.245 ;
        RECT 129.480 161.060 130.550 161.200 ;
        RECT 129.480 161.000 129.800 161.060 ;
        RECT 130.260 161.015 130.550 161.060 ;
        RECT 134.540 161.000 134.860 161.260 ;
        RECT 142.835 161.015 143.125 161.245 ;
        RECT 131.320 160.860 131.640 160.920 ;
        RECT 129.110 160.720 131.640 160.860 ;
        RECT 134.630 160.860 134.770 161.000 ;
        RECT 141.455 160.860 141.745 160.905 ;
        RECT 142.910 160.860 143.050 161.015 ;
        RECT 134.630 160.720 143.050 160.860 ;
        RECT 131.320 160.660 131.640 160.720 ;
        RECT 141.455 160.675 141.745 160.720 ;
        RECT 22.690 160.040 157.810 160.520 ;
        RECT 33.340 159.640 33.660 159.900 ;
        RECT 37.020 159.840 37.340 159.900 ;
        RECT 44.855 159.840 45.145 159.885 ;
        RECT 37.020 159.700 45.145 159.840 ;
        RECT 37.020 159.640 37.340 159.700 ;
        RECT 44.855 159.655 45.145 159.700 ;
        RECT 45.300 159.840 45.620 159.900 ;
        RECT 47.155 159.840 47.445 159.885 ;
        RECT 45.300 159.700 47.445 159.840 ;
        RECT 45.300 159.640 45.620 159.700 ;
        RECT 47.155 159.655 47.445 159.700 ;
        RECT 54.960 159.840 55.280 159.900 ;
        RECT 55.435 159.840 55.725 159.885 ;
        RECT 54.960 159.700 55.725 159.840 ;
        RECT 54.960 159.640 55.280 159.700 ;
        RECT 55.435 159.655 55.725 159.700 ;
        RECT 24.140 159.160 24.460 159.220 ;
        RECT 28.755 159.160 29.045 159.205 ;
        RECT 24.140 159.020 29.045 159.160 ;
        RECT 33.430 159.160 33.570 159.640 ;
        RECT 36.100 159.500 36.420 159.560 ;
        RECT 37.495 159.500 37.785 159.545 ;
        RECT 36.100 159.360 49.670 159.500 ;
        RECT 36.100 159.300 36.420 159.360 ;
        RECT 37.495 159.315 37.785 159.360 ;
        RECT 49.530 159.220 49.670 159.360 ;
        RECT 39.235 159.160 39.525 159.205 ;
        RECT 33.430 159.020 39.525 159.160 ;
        RECT 24.140 158.960 24.460 159.020 ;
        RECT 28.755 158.975 29.045 159.020 ;
        RECT 39.235 158.975 39.525 159.020 ;
        RECT 46.465 159.160 46.755 159.205 ;
        RECT 47.615 159.160 47.905 159.205 ;
        RECT 48.980 159.160 49.300 159.220 ;
        RECT 46.465 159.020 47.370 159.160 ;
        RECT 46.465 158.975 46.755 159.020 ;
        RECT 27.820 158.620 28.140 158.880 ;
        RECT 28.830 158.820 28.970 158.975 ;
        RECT 37.940 158.820 38.260 158.880 ;
        RECT 28.830 158.680 38.260 158.820 ;
        RECT 37.940 158.620 38.260 158.680 ;
        RECT 38.835 158.820 39.125 158.865 ;
        RECT 40.025 158.820 40.315 158.865 ;
        RECT 42.545 158.820 42.835 158.865 ;
        RECT 38.835 158.680 42.835 158.820 ;
        RECT 47.230 158.820 47.370 159.020 ;
        RECT 47.615 159.020 49.300 159.160 ;
        RECT 47.615 158.975 47.905 159.020 ;
        RECT 48.980 158.960 49.300 159.020 ;
        RECT 49.440 158.960 49.760 159.220 ;
        RECT 55.510 159.160 55.650 159.655 ;
        RECT 57.260 159.640 57.580 159.900 ;
        RECT 59.100 159.640 59.420 159.900 ;
        RECT 71.980 159.840 72.300 159.900 ;
        RECT 75.675 159.840 75.965 159.885 ;
        RECT 71.980 159.700 75.965 159.840 ;
        RECT 71.980 159.640 72.300 159.700 ;
        RECT 75.675 159.655 75.965 159.700 ;
        RECT 82.100 159.840 82.420 159.900 ;
        RECT 82.100 159.700 89.690 159.840 ;
        RECT 82.100 159.640 82.420 159.700 ;
        RECT 57.350 159.500 57.490 159.640 ;
        RECT 58.320 159.500 58.610 159.545 ;
        RECT 57.350 159.360 58.610 159.500 ;
        RECT 58.320 159.315 58.610 159.360 ;
        RECT 86.240 159.300 86.560 159.560 ;
        RECT 55.895 159.160 56.185 159.205 ;
        RECT 55.510 159.020 56.185 159.160 ;
        RECT 55.895 158.975 56.185 159.020 ;
        RECT 57.260 158.960 57.580 159.220 ;
        RECT 65.195 159.160 65.485 159.205 ;
        RECT 66.000 159.160 66.320 159.220 ;
        RECT 65.195 159.020 66.320 159.160 ;
        RECT 65.195 158.975 65.485 159.020 ;
        RECT 66.000 158.960 66.320 159.020 ;
        RECT 69.680 159.160 70.000 159.220 ;
        RECT 72.500 159.160 72.790 159.205 ;
        RECT 69.680 159.020 72.790 159.160 ;
        RECT 69.680 158.960 70.000 159.020 ;
        RECT 72.500 158.975 72.790 159.020 ;
        RECT 74.740 158.960 75.060 159.220 ;
        RECT 78.880 158.960 79.200 159.220 ;
        RECT 80.735 158.975 81.025 159.205 ;
        RECT 81.195 158.975 81.485 159.205 ;
        RECT 82.115 159.160 82.405 159.205 ;
        RECT 83.495 159.160 83.785 159.205 ;
        RECT 82.115 159.020 83.785 159.160 ;
        RECT 86.330 159.160 86.470 159.300 ;
        RECT 87.175 159.160 87.465 159.205 ;
        RECT 86.330 159.020 87.465 159.160 ;
        RECT 89.550 159.160 89.690 159.700 ;
        RECT 89.935 159.655 90.225 159.885 ;
        RECT 91.300 159.840 91.620 159.900 ;
        RECT 101.420 159.840 101.740 159.900 ;
        RECT 91.300 159.700 101.740 159.840 ;
        RECT 90.010 159.500 90.150 159.655 ;
        RECT 91.300 159.640 91.620 159.700 ;
        RECT 101.420 159.640 101.740 159.700 ;
        RECT 109.240 159.640 109.560 159.900 ;
        RECT 116.140 159.840 116.460 159.900 ;
        RECT 116.615 159.840 116.905 159.885 ;
        RECT 116.140 159.700 116.905 159.840 ;
        RECT 116.140 159.640 116.460 159.700 ;
        RECT 116.615 159.655 116.905 159.700 ;
        RECT 128.560 159.840 128.880 159.900 ;
        RECT 134.540 159.840 134.860 159.900 ;
        RECT 136.395 159.840 136.685 159.885 ;
        RECT 128.560 159.700 130.400 159.840 ;
        RECT 128.560 159.640 128.880 159.700 ;
        RECT 90.855 159.500 91.145 159.545 ;
        RECT 90.010 159.360 91.145 159.500 ;
        RECT 90.855 159.315 91.145 159.360 ;
        RECT 92.695 159.500 92.985 159.545 ;
        RECT 109.330 159.500 109.470 159.640 ;
        RECT 110.940 159.500 111.230 159.545 ;
        RECT 92.695 159.360 103.490 159.500 ;
        RECT 109.330 159.360 111.230 159.500 ;
        RECT 92.695 159.315 92.985 159.360 ;
        RECT 92.770 159.160 92.910 159.315 ;
        RECT 103.350 159.220 103.490 159.360 ;
        RECT 110.940 159.315 111.230 159.360 ;
        RECT 112.000 159.500 112.320 159.560 ;
        RECT 122.120 159.500 122.440 159.560 ;
        RECT 129.480 159.500 129.800 159.560 ;
        RECT 112.000 159.360 122.440 159.500 ;
        RECT 112.000 159.300 112.320 159.360 ;
        RECT 122.120 159.300 122.440 159.360 ;
        RECT 126.350 159.360 128.790 159.500 ;
        RECT 89.550 159.020 92.910 159.160 ;
        RECT 95.455 159.160 95.745 159.205 ;
        RECT 95.900 159.160 96.220 159.220 ;
        RECT 95.455 159.020 96.220 159.160 ;
        RECT 82.115 158.975 82.405 159.020 ;
        RECT 83.495 158.975 83.785 159.020 ;
        RECT 87.175 158.975 87.465 159.020 ;
        RECT 95.455 158.975 95.745 159.020 ;
        RECT 47.230 158.680 47.830 158.820 ;
        RECT 38.835 158.635 39.125 158.680 ;
        RECT 40.025 158.635 40.315 158.680 ;
        RECT 42.545 158.635 42.835 158.680 ;
        RECT 38.440 158.480 38.730 158.525 ;
        RECT 40.540 158.480 40.830 158.525 ;
        RECT 42.110 158.480 42.400 158.525 ;
        RECT 38.440 158.340 42.400 158.480 ;
        RECT 38.440 158.295 38.730 158.340 ;
        RECT 40.540 158.295 40.830 158.340 ;
        RECT 42.110 158.295 42.400 158.340 ;
        RECT 47.690 158.200 47.830 158.680 ;
        RECT 53.135 158.635 53.425 158.865 ;
        RECT 57.735 158.820 58.025 158.865 ;
        RECT 58.180 158.820 58.500 158.880 ;
        RECT 57.735 158.680 58.500 158.820 ;
        RECT 57.735 158.635 58.025 158.680 ;
        RECT 25.075 158.140 25.365 158.185 ;
        RECT 25.520 158.140 25.840 158.200 ;
        RECT 25.075 158.000 25.840 158.140 ;
        RECT 25.075 157.955 25.365 158.000 ;
        RECT 25.520 157.940 25.840 158.000 ;
        RECT 45.300 157.940 45.620 158.200 ;
        RECT 47.600 158.140 47.920 158.200 ;
        RECT 53.210 158.140 53.350 158.635 ;
        RECT 58.180 158.620 58.500 158.680 ;
        RECT 61.885 158.820 62.175 158.865 ;
        RECT 64.405 158.820 64.695 158.865 ;
        RECT 65.595 158.820 65.885 158.865 ;
        RECT 61.885 158.680 65.885 158.820 ;
        RECT 61.885 158.635 62.175 158.680 ;
        RECT 64.405 158.635 64.695 158.680 ;
        RECT 65.595 158.635 65.885 158.680 ;
        RECT 66.475 158.820 66.765 158.865 ;
        RECT 68.760 158.820 69.080 158.880 ;
        RECT 66.475 158.680 69.080 158.820 ;
        RECT 66.475 158.635 66.765 158.680 ;
        RECT 68.760 158.620 69.080 158.680 ;
        RECT 69.245 158.820 69.535 158.865 ;
        RECT 71.765 158.820 72.055 158.865 ;
        RECT 72.955 158.820 73.245 158.865 ;
        RECT 69.245 158.680 73.245 158.820 ;
        RECT 69.245 158.635 69.535 158.680 ;
        RECT 71.765 158.635 72.055 158.680 ;
        RECT 72.955 158.635 73.245 158.680 ;
        RECT 73.835 158.820 74.125 158.865 ;
        RECT 78.970 158.820 79.110 158.960 ;
        RECT 73.835 158.680 79.110 158.820 ;
        RECT 73.835 158.635 74.125 158.680 ;
        RECT 54.960 158.480 55.280 158.540 ;
        RECT 62.320 158.480 62.610 158.525 ;
        RECT 63.890 158.480 64.180 158.525 ;
        RECT 65.990 158.480 66.280 158.525 ;
        RECT 54.960 158.340 62.090 158.480 ;
        RECT 54.960 158.280 55.280 158.340 ;
        RECT 59.100 158.140 59.420 158.200 ;
        RECT 47.600 158.000 59.420 158.140 ;
        RECT 47.600 157.940 47.920 158.000 ;
        RECT 59.100 157.940 59.420 158.000 ;
        RECT 59.560 157.940 59.880 158.200 ;
        RECT 61.950 158.140 62.090 158.340 ;
        RECT 62.320 158.340 66.280 158.480 ;
        RECT 62.320 158.295 62.610 158.340 ;
        RECT 63.890 158.295 64.180 158.340 ;
        RECT 65.990 158.295 66.280 158.340 ;
        RECT 69.680 158.480 69.970 158.525 ;
        RECT 71.250 158.480 71.540 158.525 ;
        RECT 73.350 158.480 73.640 158.525 ;
        RECT 69.680 158.340 73.640 158.480 ;
        RECT 80.810 158.480 80.950 158.975 ;
        RECT 81.270 158.820 81.410 158.975 ;
        RECT 95.900 158.960 96.220 159.020 ;
        RECT 96.375 159.160 96.665 159.205 ;
        RECT 96.835 159.160 97.125 159.205 ;
        RECT 96.375 159.020 97.125 159.160 ;
        RECT 96.375 158.975 96.665 159.020 ;
        RECT 96.835 158.975 97.125 159.020 ;
        RECT 103.260 158.960 103.580 159.220 ;
        RECT 109.255 159.160 109.545 159.205 ;
        RECT 110.160 159.160 110.480 159.220 ;
        RECT 109.255 159.020 110.480 159.160 ;
        RECT 109.255 158.975 109.545 159.020 ;
        RECT 110.160 158.960 110.480 159.020 ;
        RECT 112.460 159.160 112.780 159.220 ;
        RECT 115.680 159.160 116.000 159.220 ;
        RECT 112.460 159.020 116.000 159.160 ;
        RECT 112.460 158.960 112.780 159.020 ;
        RECT 115.680 158.960 116.000 159.020 ;
        RECT 117.980 158.960 118.300 159.220 ;
        RECT 123.515 159.160 123.805 159.205 ;
        RECT 124.880 159.160 125.200 159.220 ;
        RECT 126.350 159.205 126.490 159.360 ;
        RECT 128.650 159.220 128.790 159.360 ;
        RECT 129.110 159.360 129.800 159.500 ;
        RECT 130.260 159.500 130.400 159.700 ;
        RECT 134.540 159.700 136.685 159.840 ;
        RECT 134.540 159.640 134.860 159.700 ;
        RECT 136.395 159.655 136.685 159.700 ;
        RECT 139.140 159.640 139.460 159.900 ;
        RECT 140.060 159.640 140.380 159.900 ;
        RECT 144.215 159.840 144.505 159.885 ;
        RECT 147.420 159.840 147.740 159.900 ;
        RECT 144.215 159.700 147.740 159.840 ;
        RECT 144.215 159.655 144.505 159.700 ;
        RECT 147.420 159.640 147.740 159.700 ;
        RECT 149.260 159.640 149.580 159.900 ;
        RECT 152.020 159.640 152.340 159.900 ;
        RECT 154.780 159.640 155.100 159.900 ;
        RECT 130.720 159.500 131.010 159.545 ;
        RECT 130.260 159.360 131.010 159.500 ;
        RECT 123.515 159.020 125.200 159.160 ;
        RECT 123.515 158.975 123.805 159.020 ;
        RECT 124.880 158.960 125.200 159.020 ;
        RECT 126.275 158.975 126.565 159.205 ;
        RECT 126.720 159.160 127.040 159.220 ;
        RECT 127.195 159.160 127.485 159.205 ;
        RECT 126.720 159.020 127.485 159.160 ;
        RECT 126.720 158.960 127.040 159.020 ;
        RECT 127.195 158.975 127.485 159.020 ;
        RECT 127.655 158.975 127.945 159.205 ;
        RECT 83.020 158.820 83.340 158.880 ;
        RECT 81.270 158.680 83.340 158.820 ;
        RECT 83.020 158.620 83.340 158.680 ;
        RECT 88.080 158.820 88.400 158.880 ;
        RECT 88.555 158.820 88.845 158.865 ;
        RECT 88.080 158.680 88.845 158.820 ;
        RECT 88.080 158.620 88.400 158.680 ;
        RECT 88.555 158.635 88.845 158.680 ;
        RECT 94.535 158.820 94.825 158.865 ;
        RECT 109.700 158.820 110.020 158.880 ;
        RECT 94.535 158.680 95.670 158.820 ;
        RECT 94.535 158.635 94.825 158.680 ;
        RECT 95.530 158.480 95.670 158.680 ;
        RECT 101.970 158.680 110.020 158.820 ;
        RECT 80.810 158.340 95.670 158.480 ;
        RECT 69.680 158.295 69.970 158.340 ;
        RECT 71.250 158.295 71.540 158.340 ;
        RECT 73.350 158.295 73.640 158.340 ;
        RECT 95.530 158.200 95.670 158.340 ;
        RECT 97.755 158.480 98.045 158.525 ;
        RECT 99.580 158.480 99.900 158.540 ;
        RECT 97.755 158.340 99.900 158.480 ;
        RECT 97.755 158.295 98.045 158.340 ;
        RECT 99.580 158.280 99.900 158.340 ;
        RECT 66.920 158.140 67.240 158.200 ;
        RECT 61.950 158.000 67.240 158.140 ;
        RECT 66.920 157.940 67.240 158.000 ;
        RECT 81.640 158.140 81.960 158.200 ;
        RECT 82.575 158.140 82.865 158.185 ;
        RECT 81.640 158.000 82.865 158.140 ;
        RECT 81.640 157.940 81.960 158.000 ;
        RECT 82.575 157.955 82.865 158.000 ;
        RECT 89.015 158.140 89.305 158.185 ;
        RECT 90.380 158.140 90.700 158.200 ;
        RECT 89.015 158.000 90.700 158.140 ;
        RECT 89.015 157.955 89.305 158.000 ;
        RECT 90.380 157.940 90.700 158.000 ;
        RECT 95.440 157.940 95.760 158.200 ;
        RECT 99.120 158.140 99.440 158.200 ;
        RECT 101.970 158.185 102.110 158.680 ;
        RECT 109.700 158.620 110.020 158.680 ;
        RECT 110.595 158.820 110.885 158.865 ;
        RECT 111.785 158.820 112.075 158.865 ;
        RECT 114.305 158.820 114.595 158.865 ;
        RECT 110.595 158.680 114.595 158.820 ;
        RECT 115.770 158.820 115.910 158.960 ;
        RECT 121.200 158.820 121.520 158.880 ;
        RECT 127.730 158.820 127.870 158.975 ;
        RECT 128.100 158.960 128.420 159.220 ;
        RECT 128.560 158.960 128.880 159.220 ;
        RECT 115.770 158.680 127.870 158.820 ;
        RECT 110.595 158.635 110.885 158.680 ;
        RECT 111.785 158.635 112.075 158.680 ;
        RECT 114.305 158.635 114.595 158.680 ;
        RECT 121.200 158.620 121.520 158.680 ;
        RECT 103.260 158.280 103.580 158.540 ;
        RECT 129.110 158.525 129.250 159.360 ;
        RECT 129.480 159.300 129.800 159.360 ;
        RECT 130.720 159.315 131.010 159.360 ;
        RECT 139.230 159.160 139.370 159.640 ;
        RECT 140.995 159.500 141.285 159.545 ;
        RECT 145.580 159.500 145.900 159.560 ;
        RECT 140.995 159.360 145.900 159.500 ;
        RECT 149.350 159.500 149.490 159.640 ;
        RECT 149.780 159.500 150.070 159.545 ;
        RECT 149.350 159.360 150.070 159.500 ;
        RECT 140.995 159.315 141.285 159.360 ;
        RECT 145.580 159.300 145.900 159.360 ;
        RECT 149.780 159.315 150.070 159.360 ;
        RECT 150.640 159.300 150.960 159.560 ;
        RECT 139.615 159.160 139.905 159.205 ;
        RECT 139.230 159.020 139.905 159.160 ;
        RECT 139.615 158.975 139.905 159.020 ;
        RECT 129.495 158.635 129.785 158.865 ;
        RECT 130.375 158.820 130.665 158.865 ;
        RECT 131.565 158.820 131.855 158.865 ;
        RECT 134.085 158.820 134.375 158.865 ;
        RECT 130.375 158.680 134.375 158.820 ;
        RECT 130.375 158.635 130.665 158.680 ;
        RECT 131.565 158.635 131.855 158.680 ;
        RECT 134.085 158.635 134.375 158.680 ;
        RECT 146.525 158.820 146.815 158.865 ;
        RECT 149.045 158.820 149.335 158.865 ;
        RECT 150.235 158.820 150.525 158.865 ;
        RECT 146.525 158.680 150.525 158.820 ;
        RECT 150.730 158.820 150.870 159.300 ;
        RECT 151.115 159.160 151.405 159.205 ;
        RECT 152.480 159.160 152.800 159.220 ;
        RECT 151.115 159.020 152.800 159.160 ;
        RECT 151.115 158.975 151.405 159.020 ;
        RECT 152.480 158.960 152.800 159.020 ;
        RECT 152.955 159.160 153.245 159.205 ;
        RECT 153.400 159.160 153.720 159.220 ;
        RECT 152.955 159.020 153.720 159.160 ;
        RECT 152.955 158.975 153.245 159.020 ;
        RECT 153.400 158.960 153.720 159.020 ;
        RECT 153.875 159.160 154.165 159.205 ;
        RECT 154.335 159.160 154.625 159.205 ;
        RECT 153.875 159.020 154.625 159.160 ;
        RECT 153.875 158.975 154.165 159.020 ;
        RECT 154.335 158.975 154.625 159.020 ;
        RECT 154.780 159.160 155.100 159.220 ;
        RECT 155.255 159.160 155.545 159.205 ;
        RECT 154.780 159.020 155.545 159.160 ;
        RECT 153.950 158.820 154.090 158.975 ;
        RECT 154.780 158.960 155.100 159.020 ;
        RECT 155.255 158.975 155.545 159.020 ;
        RECT 150.730 158.680 154.090 158.820 ;
        RECT 146.525 158.635 146.815 158.680 ;
        RECT 149.045 158.635 149.335 158.680 ;
        RECT 150.235 158.635 150.525 158.680 ;
        RECT 110.200 158.480 110.490 158.525 ;
        RECT 112.300 158.480 112.590 158.525 ;
        RECT 113.870 158.480 114.160 158.525 ;
        RECT 110.200 158.340 114.160 158.480 ;
        RECT 110.200 158.295 110.490 158.340 ;
        RECT 112.300 158.295 112.590 158.340 ;
        RECT 113.870 158.295 114.160 158.340 ;
        RECT 129.035 158.295 129.325 158.525 ;
        RECT 101.895 158.140 102.185 158.185 ;
        RECT 99.120 158.000 102.185 158.140 ;
        RECT 103.350 158.140 103.490 158.280 ;
        RECT 113.380 158.140 113.700 158.200 ;
        RECT 103.350 158.000 113.700 158.140 ;
        RECT 99.120 157.940 99.440 158.000 ;
        RECT 101.895 157.955 102.185 158.000 ;
        RECT 113.380 157.940 113.700 158.000 ;
        RECT 116.600 158.140 116.920 158.200 ;
        RECT 117.075 158.140 117.365 158.185 ;
        RECT 116.600 158.000 117.365 158.140 ;
        RECT 116.600 157.940 116.920 158.000 ;
        RECT 117.075 157.955 117.365 158.000 ;
        RECT 124.420 157.940 124.740 158.200 ;
        RECT 129.570 158.140 129.710 158.635 ;
        RECT 129.980 158.480 130.270 158.525 ;
        RECT 132.080 158.480 132.370 158.525 ;
        RECT 133.650 158.480 133.940 158.525 ;
        RECT 129.980 158.340 133.940 158.480 ;
        RECT 129.980 158.295 130.270 158.340 ;
        RECT 132.080 158.295 132.370 158.340 ;
        RECT 133.650 158.295 133.940 158.340 ;
        RECT 140.995 158.480 141.285 158.525 ;
        RECT 142.820 158.480 143.140 158.540 ;
        RECT 140.995 158.340 143.140 158.480 ;
        RECT 140.995 158.295 141.285 158.340 ;
        RECT 142.820 158.280 143.140 158.340 ;
        RECT 146.960 158.480 147.250 158.525 ;
        RECT 148.530 158.480 148.820 158.525 ;
        RECT 150.630 158.480 150.920 158.525 ;
        RECT 146.960 158.340 150.920 158.480 ;
        RECT 146.960 158.295 147.250 158.340 ;
        RECT 148.530 158.295 148.820 158.340 ;
        RECT 150.630 158.295 150.920 158.340 ;
        RECT 131.320 158.140 131.640 158.200 ;
        RECT 129.570 158.000 131.640 158.140 ;
        RECT 131.320 157.940 131.640 158.000 ;
        RECT 22.690 157.320 157.010 157.800 ;
        RECT 31.040 156.920 31.360 157.180 ;
        RECT 33.800 156.920 34.120 157.180 ;
        RECT 34.275 157.120 34.565 157.165 ;
        RECT 36.560 157.120 36.880 157.180 ;
        RECT 34.275 156.980 36.880 157.120 ;
        RECT 34.275 156.935 34.565 156.980 ;
        RECT 36.560 156.920 36.880 156.980 ;
        RECT 37.035 157.120 37.325 157.165 ;
        RECT 37.480 157.120 37.800 157.180 ;
        RECT 37.035 156.980 37.800 157.120 ;
        RECT 37.035 156.935 37.325 156.980 ;
        RECT 24.640 156.780 24.930 156.825 ;
        RECT 26.740 156.780 27.030 156.825 ;
        RECT 28.310 156.780 28.600 156.825 ;
        RECT 24.640 156.640 28.600 156.780 ;
        RECT 24.640 156.595 24.930 156.640 ;
        RECT 26.740 156.595 27.030 156.640 ;
        RECT 28.310 156.595 28.600 156.640 ;
        RECT 25.035 156.440 25.325 156.485 ;
        RECT 26.225 156.440 26.515 156.485 ;
        RECT 28.745 156.440 29.035 156.485 ;
        RECT 25.035 156.300 29.035 156.440 ;
        RECT 25.035 156.255 25.325 156.300 ;
        RECT 26.225 156.255 26.515 156.300 ;
        RECT 28.745 156.255 29.035 156.300 ;
        RECT 24.140 155.900 24.460 156.160 ;
        RECT 25.520 156.145 25.840 156.160 ;
        RECT 25.490 156.100 25.840 156.145 ;
        RECT 25.325 155.960 25.840 156.100 ;
        RECT 25.490 155.915 25.840 155.960 ;
        RECT 25.520 155.900 25.840 155.915 ;
        RECT 31.130 155.760 31.270 156.920 ;
        RECT 33.890 156.780 34.030 156.920 ;
        RECT 35.195 156.780 35.485 156.825 ;
        RECT 37.110 156.780 37.250 156.935 ;
        RECT 37.480 156.920 37.800 156.980 ;
        RECT 37.940 156.920 38.260 157.180 ;
        RECT 44.840 157.120 45.160 157.180 ;
        RECT 54.515 157.120 54.805 157.165 ;
        RECT 44.840 156.980 54.805 157.120 ;
        RECT 44.840 156.920 45.160 156.980 ;
        RECT 54.515 156.935 54.805 156.980 ;
        RECT 56.815 157.120 57.105 157.165 ;
        RECT 57.260 157.120 57.580 157.180 ;
        RECT 56.815 156.980 57.580 157.120 ;
        RECT 56.815 156.935 57.105 156.980 ;
        RECT 33.890 156.640 35.485 156.780 ;
        RECT 35.195 156.595 35.485 156.640 ;
        RECT 36.650 156.640 37.250 156.780 ;
        RECT 36.650 156.500 36.790 156.640 ;
        RECT 36.560 156.240 36.880 156.500 ;
        RECT 38.030 156.440 38.170 156.920 ;
        RECT 38.900 156.780 39.190 156.825 ;
        RECT 41.000 156.780 41.290 156.825 ;
        RECT 42.570 156.780 42.860 156.825 ;
        RECT 38.900 156.640 42.860 156.780 ;
        RECT 38.900 156.595 39.190 156.640 ;
        RECT 41.000 156.595 41.290 156.640 ;
        RECT 42.570 156.595 42.860 156.640 ;
        RECT 45.315 156.780 45.605 156.825 ;
        RECT 47.600 156.780 47.920 156.840 ;
        RECT 45.315 156.640 47.920 156.780 ;
        RECT 45.315 156.595 45.605 156.640 ;
        RECT 47.600 156.580 47.920 156.640 ;
        RECT 48.100 156.780 48.390 156.825 ;
        RECT 50.200 156.780 50.490 156.825 ;
        RECT 51.770 156.780 52.060 156.825 ;
        RECT 48.100 156.640 52.060 156.780 ;
        RECT 48.100 156.595 48.390 156.640 ;
        RECT 50.200 156.595 50.490 156.640 ;
        RECT 51.770 156.595 52.060 156.640 ;
        RECT 38.415 156.440 38.705 156.485 ;
        RECT 38.030 156.300 38.705 156.440 ;
        RECT 38.415 156.255 38.705 156.300 ;
        RECT 39.295 156.440 39.585 156.485 ;
        RECT 40.485 156.440 40.775 156.485 ;
        RECT 43.005 156.440 43.295 156.485 ;
        RECT 48.495 156.440 48.785 156.485 ;
        RECT 49.685 156.440 49.975 156.485 ;
        RECT 52.205 156.440 52.495 156.485 ;
        RECT 39.295 156.300 43.295 156.440 ;
        RECT 39.295 156.255 39.585 156.300 ;
        RECT 40.485 156.255 40.775 156.300 ;
        RECT 43.005 156.255 43.295 156.300 ;
        RECT 45.850 156.300 47.370 156.440 ;
        RECT 31.500 156.100 31.820 156.160 ;
        RECT 32.435 156.100 32.725 156.145 ;
        RECT 42.080 156.100 42.400 156.160 ;
        RECT 45.850 156.100 45.990 156.300 ;
        RECT 47.230 156.145 47.370 156.300 ;
        RECT 48.495 156.300 52.495 156.440 ;
        RECT 48.495 156.255 48.785 156.300 ;
        RECT 49.685 156.255 49.975 156.300 ;
        RECT 52.205 156.255 52.495 156.300 ;
        RECT 31.500 155.960 38.170 156.100 ;
        RECT 31.500 155.900 31.820 155.960 ;
        RECT 32.435 155.915 32.725 155.960 ;
        RECT 37.020 155.805 37.340 155.820 ;
        RECT 36.115 155.760 36.405 155.805 ;
        RECT 31.130 155.620 36.405 155.760 ;
        RECT 36.115 155.575 36.405 155.620 ;
        RECT 37.020 155.575 37.405 155.805 ;
        RECT 37.020 155.560 37.340 155.575 ;
        RECT 34.260 155.220 34.580 155.480 ;
        RECT 38.030 155.465 38.170 155.960 ;
        RECT 42.080 155.960 45.990 156.100 ;
        RECT 42.080 155.900 42.400 155.960 ;
        RECT 46.235 155.915 46.525 156.145 ;
        RECT 47.155 155.915 47.445 156.145 ;
        RECT 47.615 156.100 47.905 156.145 ;
        RECT 51.280 156.100 51.600 156.160 ;
        RECT 47.615 155.960 51.600 156.100 ;
        RECT 54.590 156.100 54.730 156.935 ;
        RECT 57.260 156.920 57.580 156.980 ;
        RECT 58.655 157.120 58.945 157.165 ;
        RECT 59.560 157.120 59.880 157.180 ;
        RECT 62.780 157.120 63.100 157.180 ;
        RECT 90.840 157.120 91.160 157.180 ;
        RECT 58.655 156.980 62.090 157.120 ;
        RECT 58.655 156.935 58.945 156.980 ;
        RECT 59.560 156.920 59.880 156.980 ;
        RECT 61.950 156.485 62.090 156.980 ;
        RECT 62.780 156.980 91.160 157.120 ;
        RECT 62.780 156.920 63.100 156.980 ;
        RECT 90.840 156.920 91.160 156.980 ;
        RECT 92.695 157.120 92.985 157.165 ;
        RECT 94.060 157.120 94.380 157.180 ;
        RECT 92.695 156.980 94.380 157.120 ;
        RECT 92.695 156.935 92.985 156.980 ;
        RECT 94.060 156.920 94.380 156.980 ;
        RECT 94.610 156.980 109.470 157.120 ;
        RECT 72.020 156.780 72.310 156.825 ;
        RECT 74.120 156.780 74.410 156.825 ;
        RECT 75.690 156.780 75.980 156.825 ;
        RECT 72.020 156.640 75.980 156.780 ;
        RECT 72.020 156.595 72.310 156.640 ;
        RECT 74.120 156.595 74.410 156.640 ;
        RECT 75.690 156.595 75.980 156.640 ;
        RECT 79.380 156.780 79.670 156.825 ;
        RECT 81.480 156.780 81.770 156.825 ;
        RECT 83.050 156.780 83.340 156.825 ;
        RECT 92.220 156.780 92.540 156.840 ;
        RECT 94.610 156.780 94.750 156.980 ;
        RECT 79.380 156.640 83.340 156.780 ;
        RECT 79.380 156.595 79.670 156.640 ;
        RECT 81.480 156.595 81.770 156.640 ;
        RECT 83.050 156.595 83.340 156.640 ;
        RECT 85.410 156.640 94.750 156.780 ;
        RECT 96.820 156.780 97.110 156.825 ;
        RECT 98.390 156.780 98.680 156.825 ;
        RECT 100.490 156.780 100.780 156.825 ;
        RECT 96.820 156.640 100.780 156.780 ;
        RECT 61.875 156.255 62.165 156.485 ;
        RECT 66.920 156.240 67.240 156.500 ;
        RECT 68.760 156.440 69.080 156.500 ;
        RECT 71.060 156.440 71.380 156.500 ;
        RECT 71.535 156.440 71.825 156.485 ;
        RECT 68.760 156.300 71.825 156.440 ;
        RECT 68.760 156.240 69.080 156.300 ;
        RECT 71.060 156.240 71.380 156.300 ;
        RECT 71.535 156.255 71.825 156.300 ;
        RECT 72.415 156.440 72.705 156.485 ;
        RECT 73.605 156.440 73.895 156.485 ;
        RECT 76.125 156.440 76.415 156.485 ;
        RECT 72.415 156.300 76.415 156.440 ;
        RECT 72.415 156.255 72.705 156.300 ;
        RECT 73.605 156.255 73.895 156.300 ;
        RECT 76.125 156.255 76.415 156.300 ;
        RECT 78.880 156.240 79.200 156.500 ;
        RECT 79.775 156.440 80.065 156.485 ;
        RECT 80.965 156.440 81.255 156.485 ;
        RECT 83.485 156.440 83.775 156.485 ;
        RECT 79.775 156.300 83.775 156.440 ;
        RECT 79.775 156.255 80.065 156.300 ;
        RECT 80.965 156.255 81.255 156.300 ;
        RECT 83.485 156.255 83.775 156.300 ;
        RECT 58.640 156.100 58.960 156.160 ;
        RECT 59.115 156.100 59.405 156.145 ;
        RECT 54.590 155.960 59.405 156.100 ;
        RECT 47.615 155.915 47.905 155.960 ;
        RECT 39.780 155.805 40.100 155.820 ;
        RECT 39.750 155.575 40.100 155.805 ;
        RECT 39.780 155.560 40.100 155.575 ;
        RECT 46.310 155.480 46.450 155.915 ;
        RECT 51.280 155.900 51.600 155.960 ;
        RECT 58.640 155.900 58.960 155.960 ;
        RECT 59.115 155.915 59.405 155.960 ;
        RECT 80.230 156.100 80.520 156.145 ;
        RECT 81.640 156.100 81.960 156.160 ;
        RECT 80.230 155.960 81.960 156.100 ;
        RECT 80.230 155.915 80.520 155.960 ;
        RECT 81.640 155.900 81.960 155.960 ;
        RECT 46.695 155.760 46.985 155.805 ;
        RECT 48.840 155.760 49.130 155.805 ;
        RECT 46.695 155.620 49.130 155.760 ;
        RECT 46.695 155.575 46.985 155.620 ;
        RECT 48.840 155.575 49.130 155.620 ;
        RECT 66.920 155.760 67.240 155.820 ;
        RECT 72.870 155.760 73.160 155.805 ;
        RECT 75.200 155.760 75.520 155.820 ;
        RECT 66.920 155.620 70.830 155.760 ;
        RECT 66.920 155.560 67.240 155.620 ;
        RECT 37.955 155.235 38.245 155.465 ;
        RECT 46.220 155.220 46.540 155.480 ;
        RECT 65.080 155.220 65.400 155.480 ;
        RECT 70.140 155.220 70.460 155.480 ;
        RECT 70.690 155.420 70.830 155.620 ;
        RECT 72.870 155.620 75.520 155.760 ;
        RECT 72.870 155.575 73.160 155.620 ;
        RECT 75.200 155.560 75.520 155.620 ;
        RECT 76.580 155.760 76.900 155.820 ;
        RECT 85.410 155.760 85.550 156.640 ;
        RECT 92.220 156.580 92.540 156.640 ;
        RECT 96.820 156.595 97.110 156.640 ;
        RECT 98.390 156.595 98.680 156.640 ;
        RECT 100.490 156.595 100.780 156.640 ;
        RECT 86.240 156.440 86.560 156.500 ;
        RECT 90.840 156.440 91.160 156.500 ;
        RECT 86.240 156.300 91.160 156.440 ;
        RECT 86.240 156.240 86.560 156.300 ;
        RECT 88.080 156.100 88.400 156.160 ;
        RECT 88.630 156.145 88.770 156.300 ;
        RECT 90.840 156.240 91.160 156.300 ;
        RECT 91.315 156.440 91.605 156.485 ;
        RECT 91.760 156.440 92.080 156.500 ;
        RECT 96.385 156.440 96.675 156.485 ;
        RECT 98.905 156.440 99.195 156.485 ;
        RECT 100.095 156.440 100.385 156.485 ;
        RECT 91.315 156.300 92.080 156.440 ;
        RECT 91.315 156.255 91.605 156.300 ;
        RECT 91.760 156.240 92.080 156.300 ;
        RECT 92.310 156.300 94.290 156.440 ;
        RECT 76.580 155.620 85.550 155.760 ;
        RECT 85.870 155.960 88.400 156.100 ;
        RECT 76.580 155.560 76.900 155.620 ;
        RECT 75.660 155.420 75.980 155.480 ;
        RECT 70.690 155.280 75.980 155.420 ;
        RECT 75.660 155.220 75.980 155.280 ;
        RECT 78.435 155.420 78.725 155.465 ;
        RECT 82.560 155.420 82.880 155.480 ;
        RECT 78.435 155.280 82.880 155.420 ;
        RECT 78.435 155.235 78.725 155.280 ;
        RECT 82.560 155.220 82.880 155.280 ;
        RECT 85.320 155.420 85.640 155.480 ;
        RECT 85.870 155.465 86.010 155.960 ;
        RECT 88.080 155.900 88.400 155.960 ;
        RECT 88.555 155.915 88.845 156.145 ;
        RECT 90.380 156.100 90.700 156.160 ;
        RECT 92.310 156.100 92.450 156.300 ;
        RECT 90.380 155.960 92.450 156.100 ;
        RECT 90.380 155.900 90.700 155.960 ;
        RECT 92.925 155.930 93.215 155.975 ;
        RECT 85.795 155.420 86.085 155.465 ;
        RECT 85.320 155.280 86.085 155.420 ;
        RECT 88.170 155.420 88.310 155.900 ;
        RECT 91.775 155.760 92.065 155.805 ;
        RECT 91.390 155.620 92.065 155.760 ;
        RECT 92.850 155.760 93.215 155.930 ;
        RECT 92.850 155.620 93.370 155.760 ;
        RECT 91.390 155.420 91.530 155.620 ;
        RECT 91.775 155.575 92.065 155.620 ;
        RECT 93.230 155.480 93.370 155.620 ;
        RECT 94.150 155.480 94.290 156.300 ;
        RECT 96.385 156.300 100.385 156.440 ;
        RECT 96.385 156.255 96.675 156.300 ;
        RECT 98.905 156.255 99.195 156.300 ;
        RECT 100.095 156.255 100.385 156.300 ;
        RECT 104.180 156.240 104.500 156.500 ;
        RECT 109.330 156.440 109.470 156.980 ;
        RECT 110.620 156.920 110.940 157.180 ;
        RECT 119.820 157.120 120.140 157.180 ;
        RECT 111.170 156.980 120.140 157.120 ;
        RECT 111.170 156.440 111.310 156.980 ;
        RECT 119.820 156.920 120.140 156.980 ;
        RECT 114.800 156.780 115.090 156.825 ;
        RECT 116.900 156.780 117.190 156.825 ;
        RECT 118.470 156.780 118.760 156.825 ;
        RECT 123.960 156.780 124.280 156.840 ;
        RECT 114.800 156.640 118.760 156.780 ;
        RECT 114.800 156.595 115.090 156.640 ;
        RECT 116.900 156.595 117.190 156.640 ;
        RECT 118.470 156.595 118.760 156.640 ;
        RECT 119.450 156.640 124.280 156.780 ;
        RECT 109.330 156.300 111.310 156.440 ;
        RECT 115.195 156.440 115.485 156.485 ;
        RECT 116.385 156.440 116.675 156.485 ;
        RECT 118.905 156.440 119.195 156.485 ;
        RECT 115.195 156.300 119.195 156.440 ;
        RECT 100.975 156.100 101.265 156.145 ;
        RECT 99.210 155.960 101.265 156.100 ;
        RECT 99.210 155.820 99.350 155.960 ;
        RECT 100.975 155.915 101.265 155.960 ;
        RECT 107.415 156.100 107.705 156.145 ;
        RECT 107.875 156.100 108.165 156.145 ;
        RECT 107.415 155.960 108.165 156.100 ;
        RECT 107.415 155.915 107.705 155.960 ;
        RECT 107.875 155.915 108.165 155.960 ;
        RECT 108.320 156.100 108.640 156.160 ;
        RECT 109.330 156.145 109.470 156.300 ;
        RECT 115.195 156.255 115.485 156.300 ;
        RECT 116.385 156.255 116.675 156.300 ;
        RECT 118.905 156.255 119.195 156.300 ;
        RECT 108.795 156.100 109.085 156.145 ;
        RECT 108.320 155.960 109.085 156.100 ;
        RECT 108.320 155.900 108.640 155.960 ;
        RECT 108.795 155.915 109.085 155.960 ;
        RECT 109.255 155.915 109.545 156.145 ;
        RECT 109.700 155.900 110.020 156.160 ;
        RECT 112.460 155.900 112.780 156.160 ;
        RECT 114.315 156.100 114.605 156.145 ;
        RECT 114.760 156.100 115.080 156.160 ;
        RECT 119.450 156.100 119.590 156.640 ;
        RECT 123.960 156.580 124.280 156.640 ;
        RECT 127.180 156.780 127.470 156.825 ;
        RECT 128.750 156.780 129.040 156.825 ;
        RECT 130.850 156.780 131.140 156.825 ;
        RECT 127.180 156.640 131.140 156.780 ;
        RECT 127.180 156.595 127.470 156.640 ;
        RECT 128.750 156.595 129.040 156.640 ;
        RECT 130.850 156.595 131.140 156.640 ;
        RECT 148.840 156.780 149.130 156.825 ;
        RECT 150.940 156.780 151.230 156.825 ;
        RECT 152.510 156.780 152.800 156.825 ;
        RECT 148.840 156.640 152.800 156.780 ;
        RECT 148.840 156.595 149.130 156.640 ;
        RECT 150.940 156.595 151.230 156.640 ;
        RECT 152.510 156.595 152.800 156.640 ;
        RECT 126.745 156.440 127.035 156.485 ;
        RECT 129.265 156.440 129.555 156.485 ;
        RECT 130.455 156.440 130.745 156.485 ;
        RECT 122.670 156.300 124.190 156.440 ;
        RECT 122.670 156.145 122.810 156.300 ;
        RECT 124.050 156.160 124.190 156.300 ;
        RECT 126.745 156.300 130.745 156.440 ;
        RECT 126.745 156.255 127.035 156.300 ;
        RECT 129.265 156.255 129.555 156.300 ;
        RECT 130.455 156.255 130.745 156.300 ;
        RECT 149.235 156.440 149.525 156.485 ;
        RECT 150.425 156.440 150.715 156.485 ;
        RECT 152.945 156.440 153.235 156.485 ;
        RECT 149.235 156.300 153.235 156.440 ;
        RECT 149.235 156.255 149.525 156.300 ;
        RECT 150.425 156.255 150.715 156.300 ;
        RECT 152.945 156.255 153.235 156.300 ;
        RECT 114.315 155.960 115.080 156.100 ;
        RECT 114.315 155.915 114.605 155.960 ;
        RECT 114.760 155.900 115.080 155.960 ;
        RECT 115.310 155.960 119.590 156.100 ;
        RECT 99.120 155.560 99.440 155.820 ;
        RECT 99.580 155.805 99.900 155.820 ;
        RECT 99.580 155.760 99.930 155.805 ;
        RECT 112.550 155.760 112.690 155.900 ;
        RECT 115.310 155.760 115.450 155.960 ;
        RECT 122.595 155.915 122.885 156.145 ;
        RECT 123.515 155.915 123.805 156.145 ;
        RECT 99.580 155.620 100.095 155.760 ;
        RECT 112.550 155.620 115.450 155.760 ;
        RECT 115.650 155.760 115.940 155.805 ;
        RECT 116.600 155.760 116.920 155.820 ;
        RECT 121.675 155.760 121.965 155.805 ;
        RECT 115.650 155.620 116.920 155.760 ;
        RECT 99.580 155.575 99.930 155.620 ;
        RECT 115.650 155.575 115.940 155.620 ;
        RECT 99.580 155.560 99.900 155.575 ;
        RECT 116.600 155.560 116.920 155.620 ;
        RECT 118.070 155.620 121.965 155.760 ;
        RECT 88.170 155.280 91.530 155.420 ;
        RECT 85.320 155.220 85.640 155.280 ;
        RECT 85.795 155.235 86.085 155.280 ;
        RECT 93.140 155.220 93.460 155.480 ;
        RECT 93.600 155.220 93.920 155.480 ;
        RECT 94.060 155.420 94.380 155.480 ;
        RECT 96.360 155.420 96.680 155.480 ;
        RECT 94.060 155.280 96.680 155.420 ;
        RECT 94.060 155.220 94.380 155.280 ;
        RECT 96.360 155.220 96.680 155.280 ;
        RECT 117.520 155.420 117.840 155.480 ;
        RECT 118.070 155.420 118.210 155.620 ;
        RECT 121.675 155.575 121.965 155.620 ;
        RECT 123.590 155.760 123.730 155.915 ;
        RECT 123.960 155.900 124.280 156.160 ;
        RECT 124.420 156.100 124.740 156.160 ;
        RECT 130.000 156.100 130.290 156.145 ;
        RECT 124.420 155.960 130.290 156.100 ;
        RECT 124.420 155.900 124.740 155.960 ;
        RECT 130.000 155.915 130.290 155.960 ;
        RECT 131.320 156.100 131.640 156.160 ;
        RECT 135.000 156.100 135.320 156.160 ;
        RECT 131.320 155.960 135.320 156.100 ;
        RECT 131.320 155.900 131.640 155.960 ;
        RECT 135.000 155.900 135.320 155.960 ;
        RECT 138.220 155.900 138.540 156.160 ;
        RECT 148.355 156.100 148.645 156.145 ;
        RECT 151.100 156.100 151.420 156.160 ;
        RECT 152.480 156.100 152.800 156.160 ;
        RECT 148.355 155.960 152.800 156.100 ;
        RECT 148.355 155.915 148.645 155.960 ;
        RECT 151.100 155.900 151.420 155.960 ;
        RECT 152.480 155.900 152.800 155.960 ;
        RECT 147.880 155.760 148.200 155.820 ;
        RECT 149.580 155.760 149.870 155.805 ;
        RECT 123.590 155.620 131.090 155.760 ;
        RECT 117.520 155.280 118.210 155.420 ;
        RECT 121.215 155.420 121.505 155.465 ;
        RECT 123.590 155.420 123.730 155.620 ;
        RECT 130.950 155.480 131.090 155.620 ;
        RECT 147.880 155.620 149.870 155.760 ;
        RECT 147.880 155.560 148.200 155.620 ;
        RECT 149.580 155.575 149.870 155.620 ;
        RECT 121.215 155.280 123.730 155.420 ;
        RECT 124.435 155.420 124.725 155.465 ;
        RECT 130.400 155.420 130.720 155.480 ;
        RECT 124.435 155.280 130.720 155.420 ;
        RECT 117.520 155.220 117.840 155.280 ;
        RECT 121.215 155.235 121.505 155.280 ;
        RECT 124.435 155.235 124.725 155.280 ;
        RECT 130.400 155.220 130.720 155.280 ;
        RECT 130.860 155.220 131.180 155.480 ;
        RECT 137.300 155.220 137.620 155.480 ;
        RECT 155.240 155.220 155.560 155.480 ;
        RECT 22.690 154.600 157.810 155.080 ;
        RECT 39.335 154.400 39.625 154.445 ;
        RECT 39.780 154.400 40.100 154.460 ;
        RECT 39.335 154.260 40.100 154.400 ;
        RECT 39.335 154.215 39.625 154.260 ;
        RECT 39.780 154.200 40.100 154.260 ;
        RECT 41.555 154.400 41.845 154.445 ;
        RECT 45.300 154.400 45.620 154.460 ;
        RECT 41.555 154.260 45.620 154.400 ;
        RECT 41.555 154.215 41.845 154.260 ;
        RECT 45.300 154.200 45.620 154.260 ;
        RECT 46.220 154.400 46.540 154.460 ;
        RECT 46.695 154.400 46.985 154.445 ;
        RECT 46.220 154.260 46.985 154.400 ;
        RECT 46.220 154.200 46.540 154.260 ;
        RECT 46.695 154.215 46.985 154.260 ;
        RECT 58.180 154.200 58.500 154.460 ;
        RECT 62.320 154.400 62.640 154.460 ;
        RECT 64.620 154.400 64.940 154.460 ;
        RECT 62.320 154.260 64.940 154.400 ;
        RECT 62.320 154.200 62.640 154.260 ;
        RECT 64.620 154.200 64.940 154.260 ;
        RECT 65.080 154.200 65.400 154.460 ;
        RECT 66.000 154.200 66.320 154.460 ;
        RECT 66.475 154.400 66.765 154.445 ;
        RECT 69.680 154.400 70.000 154.460 ;
        RECT 66.475 154.260 70.000 154.400 ;
        RECT 66.475 154.215 66.765 154.260 ;
        RECT 69.680 154.200 70.000 154.260 ;
        RECT 71.995 154.400 72.285 154.445 ;
        RECT 74.740 154.400 75.060 154.460 ;
        RECT 71.995 154.260 75.060 154.400 ;
        RECT 71.995 154.215 72.285 154.260 ;
        RECT 74.740 154.200 75.060 154.260 ;
        RECT 75.200 154.200 75.520 154.460 ;
        RECT 83.020 154.200 83.340 154.460 ;
        RECT 84.860 154.200 85.180 154.460 ;
        RECT 85.320 154.200 85.640 154.460 ;
        RECT 90.840 154.400 91.160 154.460 ;
        RECT 93.140 154.400 93.460 154.460 ;
        RECT 90.840 154.260 93.460 154.400 ;
        RECT 90.840 154.200 91.160 154.260 ;
        RECT 93.140 154.200 93.460 154.260 ;
        RECT 95.900 154.200 96.220 154.460 ;
        RECT 97.740 154.400 98.060 154.460 ;
        RECT 97.740 154.260 105.330 154.400 ;
        RECT 97.740 154.200 98.060 154.260 ;
        RECT 34.260 154.060 34.580 154.120 ;
        RECT 42.080 154.060 42.400 154.120 ;
        RECT 42.555 154.060 42.845 154.105 ;
        RECT 52.660 154.060 52.980 154.120 ;
        RECT 65.170 154.060 65.310 154.200 ;
        RECT 34.260 153.920 41.390 154.060 ;
        RECT 34.260 153.860 34.580 153.920 ;
        RECT 26.900 153.520 27.220 153.780 ;
        RECT 40.255 153.720 40.545 153.765 ;
        RECT 41.250 153.720 41.390 153.920 ;
        RECT 42.080 153.920 42.845 154.060 ;
        RECT 42.080 153.860 42.400 153.920 ;
        RECT 42.555 153.875 42.845 153.920 ;
        RECT 44.470 153.920 52.980 154.060 ;
        RECT 44.470 153.720 44.610 153.920 ;
        RECT 52.660 153.860 52.980 153.920 ;
        RECT 63.330 153.920 65.310 154.060 ;
        RECT 67.855 154.060 68.145 154.105 ;
        RECT 76.580 154.060 76.900 154.120 ;
        RECT 84.950 154.060 85.090 154.200 ;
        RECT 67.855 153.920 76.900 154.060 ;
        RECT 40.255 153.580 40.930 153.720 ;
        RECT 41.250 153.580 44.610 153.720 ;
        RECT 40.255 153.535 40.545 153.580 ;
        RECT 40.790 153.085 40.930 153.580 ;
        RECT 44.840 153.520 45.160 153.780 ;
        RECT 50.375 153.720 50.665 153.765 ;
        RECT 54.515 153.720 54.805 153.765 ;
        RECT 50.375 153.580 54.805 153.720 ;
        RECT 50.375 153.535 50.665 153.580 ;
        RECT 54.515 153.535 54.805 153.580 ;
        RECT 59.100 153.720 59.420 153.780 ;
        RECT 63.330 153.765 63.470 153.920 ;
        RECT 67.855 153.875 68.145 153.920 ;
        RECT 76.580 153.860 76.900 153.920 ;
        RECT 84.490 153.920 85.090 154.060 ;
        RECT 96.360 154.060 96.680 154.120 ;
        RECT 98.215 154.060 98.505 154.105 ;
        RECT 96.360 153.920 98.505 154.060 ;
        RECT 60.495 153.720 60.785 153.765 ;
        RECT 59.100 153.580 60.785 153.720 ;
        RECT 59.100 153.520 59.420 153.580 ;
        RECT 60.495 153.535 60.785 153.580 ;
        RECT 63.255 153.535 63.545 153.765 ;
        RECT 64.175 153.720 64.465 153.765 ;
        RECT 63.790 153.580 64.465 153.720 ;
        RECT 45.315 153.380 45.605 153.425 ;
        RECT 47.140 153.380 47.460 153.440 ;
        RECT 50.835 153.380 51.125 153.425 ;
        RECT 45.315 153.240 51.125 153.380 ;
        RECT 45.315 153.195 45.605 153.240 ;
        RECT 47.140 153.180 47.460 153.240 ;
        RECT 50.835 153.195 51.125 153.240 ;
        RECT 40.715 152.855 41.005 153.085 ;
        RECT 50.910 153.040 51.050 153.195 ;
        RECT 57.720 153.180 58.040 153.440 ;
        RECT 62.780 153.180 63.100 153.440 ;
        RECT 62.870 153.040 63.010 153.180 ;
        RECT 50.910 152.900 63.010 153.040 ;
        RECT 25.520 152.700 25.840 152.760 ;
        RECT 25.995 152.700 26.285 152.745 ;
        RECT 25.520 152.560 26.285 152.700 ;
        RECT 25.520 152.500 25.840 152.560 ;
        RECT 25.995 152.515 26.285 152.560 ;
        RECT 41.635 152.700 41.925 152.745 ;
        RECT 44.380 152.700 44.700 152.760 ;
        RECT 41.635 152.560 44.700 152.700 ;
        RECT 41.635 152.515 41.925 152.560 ;
        RECT 44.380 152.500 44.700 152.560 ;
        RECT 51.740 152.500 52.060 152.760 ;
        RECT 54.960 152.700 55.280 152.760 ;
        RECT 59.115 152.700 59.405 152.745 ;
        RECT 54.960 152.560 59.405 152.700 ;
        RECT 63.790 152.700 63.930 153.580 ;
        RECT 64.175 153.535 64.465 153.580 ;
        RECT 64.620 153.520 64.940 153.780 ;
        RECT 65.095 153.720 65.385 153.765 ;
        RECT 67.395 153.720 67.685 153.765 ;
        RECT 65.095 153.580 67.685 153.720 ;
        RECT 65.095 153.535 65.385 153.580 ;
        RECT 67.395 153.535 67.685 153.580 ;
        RECT 65.170 153.380 65.310 153.535 ;
        RECT 64.250 153.240 65.310 153.380 ;
        RECT 67.470 153.380 67.610 153.535 ;
        RECT 68.300 153.520 68.620 153.780 ;
        RECT 69.235 153.720 69.525 153.765 ;
        RECT 70.140 153.720 70.460 153.780 ;
        RECT 69.235 153.580 70.460 153.720 ;
        RECT 69.235 153.535 69.525 153.580 ;
        RECT 70.140 153.520 70.460 153.580 ;
        RECT 73.835 153.535 74.125 153.765 ;
        RECT 69.695 153.380 69.985 153.425 ;
        RECT 67.470 153.240 73.130 153.380 ;
        RECT 64.250 153.100 64.390 153.240 ;
        RECT 69.695 153.195 69.985 153.240 ;
        RECT 64.160 152.840 64.480 153.100 ;
        RECT 67.840 152.840 68.160 153.100 ;
        RECT 72.990 153.085 73.130 153.240 ;
        RECT 71.535 152.855 71.825 153.085 ;
        RECT 72.915 152.855 73.205 153.085 ;
        RECT 73.910 153.040 74.050 153.535 ;
        RECT 76.120 153.520 76.440 153.780 ;
        RECT 77.040 153.520 77.360 153.780 ;
        RECT 77.975 153.720 78.265 153.765 ;
        RECT 78.435 153.720 78.725 153.765 ;
        RECT 77.975 153.580 78.725 153.720 ;
        RECT 77.975 153.535 78.265 153.580 ;
        RECT 78.435 153.535 78.725 153.580 ;
        RECT 81.655 153.720 81.945 153.765 ;
        RECT 82.560 153.720 82.880 153.780 ;
        RECT 81.655 153.580 82.880 153.720 ;
        RECT 81.655 153.535 81.945 153.580 ;
        RECT 82.560 153.520 82.880 153.580 ;
        RECT 84.490 153.380 84.630 153.920 ;
        RECT 96.360 153.860 96.680 153.920 ;
        RECT 98.215 153.875 98.505 153.920 ;
        RECT 84.860 153.520 85.180 153.780 ;
        RECT 88.080 153.720 88.400 153.780 ;
        RECT 88.555 153.720 88.845 153.765 ;
        RECT 88.080 153.580 88.845 153.720 ;
        RECT 88.080 153.520 88.400 153.580 ;
        RECT 88.555 153.535 88.845 153.580 ;
        RECT 90.840 153.520 91.160 153.780 ;
        RECT 94.250 153.720 94.540 153.765 ;
        RECT 96.450 153.720 96.590 153.860 ;
        RECT 94.250 153.580 96.590 153.720 ;
        RECT 100.040 153.720 100.360 153.780 ;
        RECT 101.435 153.720 101.725 153.765 ;
        RECT 100.040 153.580 101.725 153.720 ;
        RECT 94.250 153.535 94.540 153.580 ;
        RECT 100.040 153.520 100.360 153.580 ;
        RECT 101.435 153.535 101.725 153.580 ;
        RECT 104.640 153.520 104.960 153.780 ;
        RECT 105.190 153.720 105.330 154.260 ;
        RECT 105.575 154.215 105.865 154.445 ;
        RECT 114.760 154.400 115.080 154.460 ;
        RECT 116.600 154.400 116.920 154.460 ;
        RECT 114.760 154.260 116.920 154.400 ;
        RECT 105.650 154.060 105.790 154.215 ;
        RECT 114.760 154.200 115.080 154.260 ;
        RECT 116.600 154.200 116.920 154.260 ;
        RECT 117.075 154.400 117.365 154.445 ;
        RECT 117.520 154.400 117.840 154.460 ;
        RECT 117.075 154.260 117.840 154.400 ;
        RECT 117.075 154.215 117.365 154.260 ;
        RECT 117.520 154.200 117.840 154.260 ;
        RECT 117.980 154.400 118.300 154.460 ;
        RECT 118.915 154.400 119.205 154.445 ;
        RECT 117.980 154.260 119.205 154.400 ;
        RECT 117.980 154.200 118.300 154.260 ;
        RECT 118.915 154.215 119.205 154.260 ;
        RECT 124.880 154.400 125.200 154.460 ;
        RECT 126.275 154.400 126.565 154.445 ;
        RECT 124.880 154.260 126.565 154.400 ;
        RECT 124.880 154.200 125.200 154.260 ;
        RECT 126.275 154.215 126.565 154.260 ;
        RECT 107.260 154.060 107.550 154.105 ;
        RECT 105.650 153.920 107.550 154.060 ;
        RECT 107.260 153.875 107.550 153.920 ;
        RECT 110.160 154.060 110.480 154.120 ;
        RECT 134.555 154.060 134.845 154.105 ;
        RECT 146.500 154.060 146.820 154.120 ;
        RECT 110.160 153.920 146.820 154.060 ;
        RECT 110.160 153.860 110.480 153.920 ;
        RECT 134.555 153.875 134.845 153.920 ;
        RECT 146.500 153.860 146.820 153.920 ;
        RECT 116.615 153.720 116.905 153.765 ;
        RECT 118.900 153.720 119.220 153.780 ;
        RECT 105.190 153.580 111.310 153.720 ;
        RECT 85.795 153.380 86.085 153.425 ;
        RECT 93.140 153.380 93.460 153.440 ;
        RECT 98.675 153.380 98.965 153.425 ;
        RECT 84.490 153.240 98.965 153.380 ;
        RECT 85.795 153.195 86.085 153.240 ;
        RECT 93.140 153.180 93.460 153.240 ;
        RECT 98.675 153.195 98.965 153.240 ;
        RECT 106.035 153.195 106.325 153.425 ;
        RECT 106.915 153.380 107.205 153.425 ;
        RECT 108.105 153.380 108.395 153.425 ;
        RECT 110.625 153.380 110.915 153.425 ;
        RECT 106.915 153.240 110.915 153.380 ;
        RECT 106.915 153.195 107.205 153.240 ;
        RECT 108.105 153.195 108.395 153.240 ;
        RECT 110.625 153.195 110.915 153.240 ;
        RECT 90.380 153.040 90.700 153.100 ;
        RECT 73.910 152.900 90.700 153.040 ;
        RECT 67.930 152.700 68.070 152.840 ;
        RECT 63.790 152.560 68.070 152.700 ;
        RECT 71.610 152.700 71.750 152.855 ;
        RECT 90.380 152.840 90.700 152.900 ;
        RECT 74.740 152.700 75.060 152.760 ;
        RECT 71.610 152.560 75.060 152.700 ;
        RECT 54.960 152.500 55.280 152.560 ;
        RECT 59.115 152.515 59.405 152.560 ;
        RECT 74.740 152.500 75.060 152.560 ;
        RECT 75.660 152.700 75.980 152.760 ;
        RECT 92.680 152.700 93.000 152.760 ;
        RECT 75.660 152.560 93.000 152.700 ;
        RECT 75.660 152.500 75.980 152.560 ;
        RECT 92.680 152.500 93.000 152.560 ;
        RECT 93.155 152.700 93.445 152.745 ;
        RECT 94.980 152.700 95.300 152.760 ;
        RECT 93.155 152.560 95.300 152.700 ;
        RECT 93.155 152.515 93.445 152.560 ;
        RECT 94.980 152.500 95.300 152.560 ;
        RECT 100.500 152.500 100.820 152.760 ;
        RECT 106.110 152.700 106.250 153.195 ;
        RECT 106.520 153.040 106.810 153.085 ;
        RECT 108.620 153.040 108.910 153.085 ;
        RECT 110.190 153.040 110.480 153.085 ;
        RECT 106.520 152.900 110.480 153.040 ;
        RECT 111.170 153.040 111.310 153.580 ;
        RECT 116.615 153.580 119.220 153.720 ;
        RECT 116.615 153.535 116.905 153.580 ;
        RECT 118.900 153.520 119.220 153.580 ;
        RECT 120.280 153.520 120.600 153.780 ;
        RECT 120.740 153.720 121.060 153.780 ;
        RECT 122.595 153.720 122.885 153.765 ;
        RECT 120.740 153.580 122.885 153.720 ;
        RECT 120.740 153.520 121.060 153.580 ;
        RECT 122.595 153.535 122.885 153.580 ;
        RECT 123.975 153.535 124.265 153.765 ;
        RECT 116.155 153.380 116.445 153.425 ;
        RECT 117.980 153.380 118.300 153.440 ;
        RECT 116.155 153.240 118.300 153.380 ;
        RECT 116.155 153.195 116.445 153.240 ;
        RECT 117.980 153.180 118.300 153.240 ;
        RECT 121.200 153.180 121.520 153.440 ;
        RECT 124.050 153.040 124.190 153.535 ;
        RECT 124.420 153.520 124.740 153.780 ;
        RECT 125.355 153.720 125.645 153.765 ;
        RECT 128.115 153.720 128.405 153.765 ;
        RECT 125.355 153.580 128.405 153.720 ;
        RECT 125.355 153.535 125.645 153.580 ;
        RECT 128.115 153.535 128.405 153.580 ;
        RECT 130.860 153.520 131.180 153.780 ;
        RECT 155.240 153.520 155.560 153.780 ;
        RECT 125.800 153.380 126.120 153.440 ;
        RECT 128.575 153.380 128.865 153.425 ;
        RECT 125.800 153.240 128.865 153.380 ;
        RECT 125.800 153.180 126.120 153.240 ;
        RECT 128.575 153.195 128.865 153.240 ;
        RECT 129.020 153.180 129.340 153.440 ;
        RECT 130.400 153.040 130.720 153.100 ;
        RECT 131.780 153.040 132.100 153.100 ;
        RECT 111.170 152.900 122.350 153.040 ;
        RECT 124.050 152.900 132.100 153.040 ;
        RECT 106.520 152.855 106.810 152.900 ;
        RECT 108.620 152.855 108.910 152.900 ;
        RECT 110.190 152.855 110.480 152.900 ;
        RECT 109.700 152.700 110.020 152.760 ;
        RECT 106.110 152.560 110.020 152.700 ;
        RECT 109.700 152.500 110.020 152.560 ;
        RECT 112.920 152.500 113.240 152.760 ;
        RECT 119.360 152.500 119.680 152.760 ;
        RECT 121.660 152.500 121.980 152.760 ;
        RECT 122.210 152.700 122.350 152.900 ;
        RECT 130.400 152.840 130.720 152.900 ;
        RECT 131.780 152.840 132.100 152.900 ;
        RECT 125.340 152.700 125.660 152.760 ;
        RECT 122.210 152.560 125.660 152.700 ;
        RECT 125.340 152.500 125.660 152.560 ;
        RECT 131.335 152.700 131.625 152.745 ;
        RECT 133.160 152.700 133.480 152.760 ;
        RECT 131.335 152.560 133.480 152.700 ;
        RECT 131.335 152.515 131.625 152.560 ;
        RECT 133.160 152.500 133.480 152.560 ;
        RECT 135.000 152.700 135.320 152.760 ;
        RECT 141.915 152.700 142.205 152.745 ;
        RECT 147.420 152.700 147.740 152.760 ;
        RECT 135.000 152.560 147.740 152.700 ;
        RECT 135.000 152.500 135.320 152.560 ;
        RECT 141.915 152.515 142.205 152.560 ;
        RECT 147.420 152.500 147.740 152.560 ;
        RECT 152.020 152.500 152.340 152.760 ;
        RECT 22.690 151.880 157.010 152.360 ;
        RECT 42.080 151.480 42.400 151.740 ;
        RECT 66.000 151.480 66.320 151.740 ;
        RECT 75.200 151.680 75.520 151.740 ;
        RECT 77.040 151.680 77.360 151.740 ;
        RECT 80.260 151.680 80.580 151.740 ;
        RECT 82.575 151.680 82.865 151.725 ;
        RECT 87.160 151.680 87.480 151.740 ;
        RECT 66.550 151.540 75.520 151.680 ;
        RECT 24.640 151.340 24.930 151.385 ;
        RECT 26.740 151.340 27.030 151.385 ;
        RECT 28.310 151.340 28.600 151.385 ;
        RECT 24.640 151.200 28.600 151.340 ;
        RECT 24.640 151.155 24.930 151.200 ;
        RECT 26.740 151.155 27.030 151.200 ;
        RECT 28.310 151.155 28.600 151.200 ;
        RECT 25.035 151.000 25.325 151.045 ;
        RECT 26.225 151.000 26.515 151.045 ;
        RECT 28.745 151.000 29.035 151.045 ;
        RECT 42.170 151.000 42.310 151.480 ;
        RECT 64.620 151.340 64.940 151.400 ;
        RECT 66.550 151.340 66.690 151.540 ;
        RECT 75.200 151.480 75.520 151.540 ;
        RECT 75.795 151.540 87.480 151.680 ;
        RECT 75.795 151.340 75.935 151.540 ;
        RECT 77.040 151.480 77.360 151.540 ;
        RECT 80.260 151.480 80.580 151.540 ;
        RECT 82.575 151.495 82.865 151.540 ;
        RECT 87.160 151.480 87.480 151.540 ;
        RECT 90.380 151.480 90.700 151.740 ;
        RECT 91.315 151.680 91.605 151.725 ;
        RECT 93.600 151.680 93.920 151.740 ;
        RECT 96.360 151.680 96.680 151.740 ;
        RECT 91.315 151.540 96.680 151.680 ;
        RECT 91.315 151.495 91.605 151.540 ;
        RECT 93.600 151.480 93.920 151.540 ;
        RECT 96.360 151.480 96.680 151.540 ;
        RECT 98.675 151.680 98.965 151.725 ;
        RECT 100.040 151.680 100.360 151.740 ;
        RECT 98.675 151.540 100.360 151.680 ;
        RECT 98.675 151.495 98.965 151.540 ;
        RECT 100.040 151.480 100.360 151.540 ;
        RECT 104.640 151.680 104.960 151.740 ;
        RECT 106.495 151.680 106.785 151.725 ;
        RECT 104.640 151.540 106.785 151.680 ;
        RECT 104.640 151.480 104.960 151.540 ;
        RECT 106.495 151.495 106.785 151.540 ;
        RECT 116.600 151.680 116.920 151.740 ;
        RECT 120.295 151.680 120.585 151.725 ;
        RECT 116.600 151.540 120.585 151.680 ;
        RECT 116.600 151.480 116.920 151.540 ;
        RECT 120.295 151.495 120.585 151.540 ;
        RECT 137.315 151.680 137.605 151.725 ;
        RECT 137.760 151.680 138.080 151.740 ;
        RECT 137.315 151.540 138.080 151.680 ;
        RECT 137.315 151.495 137.605 151.540 ;
        RECT 137.760 151.480 138.080 151.540 ;
        RECT 138.220 151.480 138.540 151.740 ;
        RECT 146.055 151.680 146.345 151.725 ;
        RECT 147.880 151.680 148.200 151.740 ;
        RECT 146.055 151.540 148.200 151.680 ;
        RECT 146.055 151.495 146.345 151.540 ;
        RECT 147.880 151.480 148.200 151.540 ;
        RECT 81.180 151.340 81.500 151.400 ;
        RECT 94.980 151.340 95.300 151.400 ;
        RECT 64.620 151.200 66.690 151.340 ;
        RECT 69.310 151.200 75.935 151.340 ;
        RECT 76.210 151.200 81.500 151.340 ;
        RECT 64.620 151.140 64.940 151.200 ;
        RECT 66.920 151.000 67.240 151.060 ;
        RECT 25.035 150.860 29.035 151.000 ;
        RECT 25.035 150.815 25.325 150.860 ;
        RECT 26.225 150.815 26.515 150.860 ;
        RECT 28.745 150.815 29.035 150.860 ;
        RECT 41.250 150.860 43.690 151.000 ;
        RECT 24.140 150.460 24.460 150.720 ;
        RECT 25.520 150.705 25.840 150.720 ;
        RECT 25.490 150.660 25.840 150.705 ;
        RECT 25.325 150.520 25.840 150.660 ;
        RECT 25.490 150.475 25.840 150.520 ;
        RECT 25.520 150.460 25.840 150.475 ;
        RECT 32.880 150.460 33.200 150.720 ;
        RECT 33.815 150.660 34.105 150.705 ;
        RECT 34.260 150.660 34.580 150.720 ;
        RECT 33.815 150.520 34.580 150.660 ;
        RECT 33.815 150.475 34.105 150.520 ;
        RECT 34.260 150.460 34.580 150.520 ;
        RECT 35.640 150.660 35.960 150.720 ;
        RECT 37.495 150.660 37.785 150.705 ;
        RECT 35.640 150.520 37.785 150.660 ;
        RECT 35.640 150.460 35.960 150.520 ;
        RECT 37.495 150.475 37.785 150.520 ;
        RECT 40.255 150.660 40.545 150.705 ;
        RECT 40.700 150.660 41.020 150.720 ;
        RECT 40.255 150.520 41.020 150.660 ;
        RECT 40.255 150.475 40.545 150.520 ;
        RECT 40.700 150.460 41.020 150.520 ;
        RECT 36.560 150.320 36.880 150.380 ;
        RECT 41.250 150.320 41.390 150.860 ;
        RECT 41.635 150.660 41.925 150.705 ;
        RECT 41.635 150.520 42.770 150.660 ;
        RECT 41.635 150.475 41.925 150.520 ;
        RECT 31.130 150.180 36.880 150.320 ;
        RECT 25.060 149.980 25.380 150.040 ;
        RECT 31.130 150.025 31.270 150.180 ;
        RECT 36.560 150.120 36.880 150.180 ;
        RECT 38.490 150.180 41.390 150.320 ;
        RECT 42.630 150.320 42.770 150.520 ;
        RECT 43.000 150.460 43.320 150.720 ;
        RECT 43.550 150.705 43.690 150.860 ;
        RECT 62.870 150.860 67.240 151.000 ;
        RECT 43.475 150.475 43.765 150.705 ;
        RECT 48.995 150.660 49.285 150.705 ;
        RECT 50.360 150.660 50.680 150.720 ;
        RECT 44.010 150.520 48.750 150.660 ;
        RECT 44.010 150.320 44.150 150.520 ;
        RECT 42.630 150.180 44.150 150.320 ;
        RECT 31.055 149.980 31.345 150.025 ;
        RECT 25.060 149.840 31.345 149.980 ;
        RECT 25.060 149.780 25.380 149.840 ;
        RECT 31.055 149.795 31.345 149.840 ;
        RECT 33.355 149.980 33.645 150.025 ;
        RECT 33.800 149.980 34.120 150.040 ;
        RECT 38.490 150.025 38.630 150.180 ;
        RECT 44.840 150.120 45.160 150.380 ;
        RECT 45.300 150.120 45.620 150.380 ;
        RECT 33.355 149.840 34.120 149.980 ;
        RECT 33.355 149.795 33.645 149.840 ;
        RECT 33.800 149.780 34.120 149.840 ;
        RECT 38.415 149.795 38.705 150.025 ;
        RECT 41.160 149.980 41.480 150.040 ;
        RECT 42.095 149.980 42.385 150.025 ;
        RECT 41.160 149.840 42.385 149.980 ;
        RECT 44.930 149.980 45.070 150.120 ;
        RECT 45.775 149.980 46.065 150.025 ;
        RECT 44.930 149.840 46.065 149.980 ;
        RECT 48.610 149.980 48.750 150.520 ;
        RECT 48.995 150.520 50.680 150.660 ;
        RECT 48.995 150.475 49.285 150.520 ;
        RECT 50.360 150.460 50.680 150.520 ;
        RECT 51.280 150.660 51.600 150.720 ;
        RECT 58.195 150.660 58.485 150.705 ;
        RECT 60.020 150.660 60.340 150.720 ;
        RECT 51.280 150.520 60.340 150.660 ;
        RECT 51.280 150.460 51.600 150.520 ;
        RECT 58.195 150.475 58.485 150.520 ;
        RECT 60.020 150.460 60.340 150.520 ;
        RECT 62.320 150.660 62.640 150.720 ;
        RECT 62.870 150.705 63.010 150.860 ;
        RECT 66.920 150.800 67.240 150.860 ;
        RECT 62.795 150.660 63.085 150.705 ;
        RECT 62.320 150.520 63.085 150.660 ;
        RECT 62.320 150.460 62.640 150.520 ;
        RECT 62.795 150.475 63.085 150.520 ;
        RECT 63.240 150.460 63.560 150.720 ;
        RECT 63.700 150.460 64.020 150.720 ;
        RECT 64.175 150.660 64.465 150.705 ;
        RECT 64.620 150.660 64.940 150.720 ;
        RECT 64.175 150.520 64.940 150.660 ;
        RECT 64.175 150.475 64.465 150.520 ;
        RECT 64.620 150.460 64.940 150.520 ;
        RECT 67.855 150.475 68.145 150.705 ;
        RECT 68.775 150.660 69.065 150.705 ;
        RECT 69.310 150.660 69.450 151.200 ;
        RECT 76.210 151.060 76.350 151.200 ;
        RECT 81.180 151.140 81.500 151.200 ;
        RECT 89.550 151.200 95.300 151.340 ;
        RECT 76.120 151.000 76.440 151.060 ;
        RECT 89.550 151.000 89.690 151.200 ;
        RECT 94.980 151.140 95.300 151.200 ;
        RECT 95.900 151.140 96.220 151.400 ;
        RECT 99.620 151.340 99.910 151.385 ;
        RECT 101.720 151.340 102.010 151.385 ;
        RECT 103.290 151.340 103.580 151.385 ;
        RECT 112.920 151.340 113.240 151.400 ;
        RECT 133.620 151.340 133.940 151.400 ;
        RECT 99.620 151.200 103.580 151.340 ;
        RECT 99.620 151.155 99.910 151.200 ;
        RECT 101.720 151.155 102.010 151.200 ;
        RECT 103.290 151.155 103.580 151.200 ;
        RECT 112.550 151.200 133.940 151.340 ;
        RECT 71.610 150.860 76.440 151.000 ;
        RECT 68.775 150.520 69.450 150.660 ;
        RECT 69.695 150.660 69.985 150.705 ;
        RECT 71.610 150.660 71.750 150.860 ;
        RECT 76.120 150.800 76.440 150.860 ;
        RECT 80.810 150.860 81.870 151.000 ;
        RECT 69.695 150.520 71.750 150.660 ;
        RECT 68.775 150.475 69.065 150.520 ;
        RECT 69.695 150.475 69.985 150.520 ;
        RECT 49.440 150.320 49.760 150.380 ;
        RECT 49.440 150.180 64.390 150.320 ;
        RECT 49.440 150.120 49.760 150.180 ;
        RECT 64.250 150.040 64.390 150.180 ;
        RECT 65.095 150.135 65.385 150.365 ;
        RECT 60.940 149.980 61.260 150.040 ;
        RECT 48.610 149.840 61.260 149.980 ;
        RECT 41.160 149.780 41.480 149.840 ;
        RECT 42.095 149.795 42.385 149.840 ;
        RECT 45.775 149.795 46.065 149.840 ;
        RECT 60.940 149.780 61.260 149.840 ;
        RECT 61.860 149.780 62.180 150.040 ;
        RECT 64.160 149.780 64.480 150.040 ;
        RECT 64.620 149.980 64.940 150.040 ;
        RECT 65.170 149.980 65.310 150.135 ;
        RECT 64.620 149.840 65.310 149.980 ;
        RECT 65.540 149.980 65.860 150.040 ;
        RECT 66.095 149.980 66.385 150.025 ;
        RECT 65.540 149.840 66.385 149.980 ;
        RECT 64.620 149.780 64.940 149.840 ;
        RECT 65.540 149.780 65.860 149.840 ;
        RECT 66.095 149.795 66.385 149.840 ;
        RECT 66.920 149.780 67.240 150.040 ;
        RECT 67.930 149.980 68.070 150.475 ;
        RECT 71.980 150.460 72.300 150.720 ;
        RECT 72.440 150.460 72.760 150.720 ;
        RECT 74.295 150.660 74.585 150.705 ;
        RECT 75.200 150.660 75.520 150.720 ;
        RECT 75.675 150.660 75.965 150.705 ;
        RECT 74.295 150.520 75.965 150.660 ;
        RECT 74.295 150.475 74.585 150.520 ;
        RECT 75.200 150.460 75.520 150.520 ;
        RECT 75.675 150.475 75.965 150.520 ;
        RECT 78.895 150.660 79.185 150.705 ;
        RECT 79.355 150.660 79.645 150.705 ;
        RECT 80.810 150.660 80.950 150.860 ;
        RECT 78.895 150.520 79.645 150.660 ;
        RECT 78.895 150.475 79.185 150.520 ;
        RECT 79.355 150.475 79.645 150.520 ;
        RECT 79.890 150.520 80.950 150.660 ;
        RECT 69.220 150.120 69.540 150.380 ;
        RECT 79.890 150.320 80.030 150.520 ;
        RECT 81.180 150.460 81.500 150.720 ;
        RECT 81.730 150.660 81.870 150.860 ;
        RECT 84.950 150.860 89.690 151.000 ;
        RECT 83.020 150.660 83.340 150.720 ;
        RECT 81.730 150.520 83.340 150.660 ;
        RECT 83.020 150.460 83.340 150.520 ;
        RECT 83.495 150.660 83.785 150.705 ;
        RECT 83.940 150.660 84.260 150.720 ;
        RECT 84.950 150.705 85.090 150.860 ;
        RECT 83.495 150.520 84.260 150.660 ;
        RECT 83.495 150.475 83.785 150.520 ;
        RECT 83.940 150.460 84.260 150.520 ;
        RECT 84.415 150.475 84.705 150.705 ;
        RECT 84.855 150.475 85.145 150.705 ;
        RECT 87.620 150.660 87.940 150.720 ;
        RECT 89.550 150.705 89.690 150.860 ;
        RECT 93.155 151.000 93.445 151.045 ;
        RECT 94.535 151.000 94.825 151.045 ;
        RECT 95.990 151.000 96.130 151.140 ;
        RECT 93.155 150.860 96.590 151.000 ;
        RECT 93.155 150.815 93.445 150.860 ;
        RECT 94.535 150.815 94.825 150.860 ;
        RECT 88.095 150.660 88.385 150.705 ;
        RECT 87.620 150.520 89.230 150.660 ;
        RECT 70.690 150.180 80.030 150.320 ;
        RECT 69.680 149.980 70.000 150.040 ;
        RECT 70.690 150.025 70.830 150.180 ;
        RECT 80.260 150.120 80.580 150.380 ;
        RECT 80.735 150.135 81.025 150.365 ;
        RECT 67.930 149.840 70.000 149.980 ;
        RECT 69.680 149.780 70.000 149.840 ;
        RECT 70.615 149.795 70.905 150.025 ;
        RECT 71.075 149.980 71.365 150.025 ;
        RECT 71.520 149.980 71.840 150.040 ;
        RECT 71.075 149.840 71.840 149.980 ;
        RECT 71.075 149.795 71.365 149.840 ;
        RECT 71.520 149.780 71.840 149.840 ;
        RECT 75.660 149.980 75.980 150.040 ;
        RECT 79.800 149.980 80.120 150.040 ;
        RECT 80.810 149.980 80.950 150.135 ;
        RECT 75.660 149.840 80.950 149.980 ;
        RECT 81.180 149.980 81.500 150.040 ;
        RECT 82.115 149.980 82.405 150.025 ;
        RECT 81.180 149.840 82.405 149.980 ;
        RECT 84.490 149.980 84.630 150.475 ;
        RECT 87.620 150.460 87.940 150.520 ;
        RECT 88.095 150.475 88.385 150.520 ;
        RECT 89.090 150.320 89.230 150.520 ;
        RECT 89.475 150.475 89.765 150.705 ;
        RECT 95.915 150.475 96.205 150.705 ;
        RECT 94.520 150.320 94.840 150.380 ;
        RECT 94.995 150.320 95.285 150.365 ;
        RECT 89.090 150.180 95.285 150.320 ;
        RECT 94.520 150.120 94.840 150.180 ;
        RECT 94.995 150.135 95.285 150.180 ;
        RECT 87.620 149.980 87.940 150.040 ;
        RECT 84.490 149.840 87.940 149.980 ;
        RECT 75.660 149.780 75.980 149.840 ;
        RECT 79.800 149.780 80.120 149.840 ;
        RECT 81.180 149.780 81.500 149.840 ;
        RECT 82.115 149.795 82.405 149.840 ;
        RECT 87.620 149.780 87.940 149.840 ;
        RECT 88.095 149.980 88.385 150.025 ;
        RECT 88.540 149.980 88.860 150.040 ;
        RECT 88.095 149.840 88.860 149.980 ;
        RECT 88.095 149.795 88.385 149.840 ;
        RECT 88.540 149.780 88.860 149.840 ;
        RECT 91.300 149.980 91.620 150.040 ;
        RECT 95.440 149.980 95.760 150.040 ;
        RECT 95.990 149.980 96.130 150.475 ;
        RECT 96.450 150.320 96.590 150.860 ;
        RECT 96.820 150.800 97.140 151.060 ;
        RECT 99.120 151.000 99.440 151.060 ;
        RECT 97.370 150.860 99.440 151.000 ;
        RECT 97.370 150.720 97.510 150.860 ;
        RECT 99.120 150.800 99.440 150.860 ;
        RECT 100.015 151.000 100.305 151.045 ;
        RECT 101.205 151.000 101.495 151.045 ;
        RECT 103.725 151.000 104.015 151.045 ;
        RECT 100.015 150.860 104.015 151.000 ;
        RECT 100.015 150.815 100.305 150.860 ;
        RECT 101.205 150.815 101.495 150.860 ;
        RECT 103.725 150.815 104.015 150.860 ;
        RECT 109.240 150.800 109.560 151.060 ;
        RECT 112.550 151.045 112.690 151.200 ;
        RECT 112.920 151.140 113.240 151.200 ;
        RECT 133.620 151.140 133.940 151.200 ;
        RECT 145.135 151.155 145.425 151.385 ;
        RECT 149.720 151.340 150.010 151.385 ;
        RECT 151.290 151.340 151.580 151.385 ;
        RECT 153.390 151.340 153.680 151.385 ;
        RECT 149.720 151.200 153.680 151.340 ;
        RECT 149.720 151.155 150.010 151.200 ;
        RECT 151.290 151.155 151.580 151.200 ;
        RECT 153.390 151.155 153.680 151.200 ;
        RECT 112.475 150.815 112.765 151.045 ;
        RECT 117.980 151.000 118.300 151.060 ;
        RECT 125.815 151.000 126.105 151.045 ;
        RECT 129.020 151.000 129.340 151.060 ;
        RECT 117.980 150.860 129.340 151.000 ;
        RECT 117.980 150.800 118.300 150.860 ;
        RECT 125.815 150.815 126.105 150.860 ;
        RECT 129.020 150.800 129.340 150.860 ;
        RECT 130.400 150.800 130.720 151.060 ;
        RECT 142.835 150.815 143.125 151.045 ;
        RECT 97.280 150.460 97.600 150.720 ;
        RECT 97.740 150.460 98.060 150.720 ;
        RECT 100.500 150.705 100.820 150.720 ;
        RECT 100.470 150.660 100.820 150.705 ;
        RECT 100.305 150.520 100.820 150.660 ;
        RECT 100.470 150.475 100.820 150.520 ;
        RECT 100.500 150.460 100.820 150.475 ;
        RECT 107.860 150.660 108.180 150.720 ;
        RECT 108.795 150.660 109.085 150.705 ;
        RECT 107.860 150.520 109.085 150.660 ;
        RECT 107.860 150.460 108.180 150.520 ;
        RECT 108.795 150.475 109.085 150.520 ;
        RECT 110.160 150.460 110.480 150.720 ;
        RECT 111.540 150.460 111.860 150.720 ;
        RECT 118.440 150.660 118.760 150.720 ;
        RECT 125.355 150.660 125.645 150.705 ;
        RECT 118.440 150.520 125.645 150.660 ;
        RECT 118.440 150.460 118.760 150.520 ;
        RECT 125.355 150.475 125.645 150.520 ;
        RECT 131.320 150.460 131.640 150.720 ;
        RECT 132.240 150.460 132.560 150.720 ;
        RECT 132.700 150.460 133.020 150.720 ;
        RECT 134.555 150.475 134.845 150.705 ;
        RECT 135.935 150.660 136.225 150.705 ;
        RECT 140.060 150.660 140.380 150.720 ;
        RECT 135.935 150.520 140.380 150.660 ;
        RECT 135.935 150.475 136.225 150.520 ;
        RECT 108.335 150.320 108.625 150.365 ;
        RECT 110.250 150.320 110.390 150.460 ;
        RECT 113.855 150.320 114.145 150.365 ;
        RECT 119.820 150.320 120.140 150.380 ;
        RECT 96.450 150.180 102.570 150.320 ;
        RECT 102.430 150.040 102.570 150.180 ;
        RECT 108.335 150.180 109.885 150.320 ;
        RECT 110.250 150.180 120.140 150.320 ;
        RECT 134.630 150.320 134.770 150.475 ;
        RECT 140.060 150.460 140.380 150.520 ;
        RECT 141.455 150.660 141.745 150.705 ;
        RECT 142.360 150.660 142.680 150.720 ;
        RECT 142.910 150.660 143.050 150.815 ;
        RECT 141.455 150.520 143.050 150.660 ;
        RECT 141.455 150.475 141.745 150.520 ;
        RECT 142.360 150.460 142.680 150.520 ;
        RECT 143.295 150.475 143.585 150.705 ;
        RECT 145.210 150.660 145.350 151.155 ;
        RECT 149.285 151.000 149.575 151.045 ;
        RECT 151.805 151.000 152.095 151.045 ;
        RECT 152.995 151.000 153.285 151.045 ;
        RECT 149.285 150.860 153.285 151.000 ;
        RECT 149.285 150.815 149.575 150.860 ;
        RECT 151.805 150.815 152.095 150.860 ;
        RECT 152.995 150.815 153.285 150.860 ;
        RECT 145.595 150.660 145.885 150.705 ;
        RECT 145.210 150.520 145.885 150.660 ;
        RECT 145.595 150.475 145.885 150.520 ;
        RECT 146.040 150.660 146.360 150.720 ;
        RECT 146.515 150.660 146.805 150.705 ;
        RECT 146.040 150.520 146.805 150.660 ;
        RECT 136.395 150.320 136.685 150.365 ;
        RECT 136.840 150.320 137.160 150.380 ;
        RECT 134.630 150.180 136.150 150.320 ;
        RECT 108.335 150.135 108.625 150.180 ;
        RECT 91.300 149.840 96.130 149.980 ;
        RECT 102.340 149.980 102.660 150.040 ;
        RECT 106.035 149.980 106.325 150.025 ;
        RECT 102.340 149.840 106.325 149.980 ;
        RECT 109.745 149.980 109.885 150.180 ;
        RECT 113.855 150.135 114.145 150.180 ;
        RECT 119.820 150.120 120.140 150.180 ;
        RECT 110.635 149.980 110.925 150.025 ;
        RECT 109.745 149.840 110.925 149.980 ;
        RECT 91.300 149.780 91.620 149.840 ;
        RECT 95.440 149.780 95.760 149.840 ;
        RECT 102.340 149.780 102.660 149.840 ;
        RECT 106.035 149.795 106.325 149.840 ;
        RECT 110.635 149.795 110.925 149.840 ;
        RECT 122.120 149.980 122.440 150.040 ;
        RECT 123.055 149.980 123.345 150.025 ;
        RECT 122.120 149.840 123.345 149.980 ;
        RECT 122.120 149.780 122.440 149.840 ;
        RECT 123.055 149.795 123.345 149.840 ;
        RECT 124.880 149.780 125.200 150.040 ;
        RECT 134.080 149.780 134.400 150.040 ;
        RECT 135.460 149.780 135.780 150.040 ;
        RECT 136.010 149.980 136.150 150.180 ;
        RECT 136.395 150.180 137.160 150.320 ;
        RECT 136.395 150.135 136.685 150.180 ;
        RECT 136.840 150.120 137.160 150.180 ;
        RECT 137.475 150.320 137.765 150.365 ;
        RECT 139.155 150.320 139.445 150.365 ;
        RECT 137.475 150.180 139.445 150.320 ;
        RECT 143.370 150.320 143.510 150.475 ;
        RECT 146.040 150.460 146.360 150.520 ;
        RECT 146.515 150.475 146.805 150.520 ;
        RECT 148.800 150.660 149.120 150.720 ;
        RECT 151.100 150.660 151.420 150.720 ;
        RECT 153.875 150.660 154.165 150.705 ;
        RECT 148.800 150.520 154.165 150.660 ;
        RECT 148.800 150.460 149.120 150.520 ;
        RECT 151.100 150.460 151.420 150.520 ;
        RECT 153.875 150.475 154.165 150.520 ;
        RECT 149.260 150.320 149.580 150.380 ;
        RECT 152.540 150.320 152.830 150.365 ;
        RECT 143.370 150.180 147.650 150.320 ;
        RECT 137.475 150.135 137.765 150.180 ;
        RECT 139.155 150.135 139.445 150.180 ;
        RECT 140.995 149.980 141.285 150.025 ;
        RECT 143.280 149.980 143.600 150.040 ;
        RECT 136.010 149.840 143.600 149.980 ;
        RECT 140.995 149.795 141.285 149.840 ;
        RECT 143.280 149.780 143.600 149.840 ;
        RECT 144.200 149.980 144.520 150.040 ;
        RECT 146.975 149.980 147.265 150.025 ;
        RECT 144.200 149.840 147.265 149.980 ;
        RECT 147.510 149.980 147.650 150.180 ;
        RECT 149.260 150.180 152.830 150.320 ;
        RECT 149.260 150.120 149.580 150.180 ;
        RECT 152.540 150.135 152.830 150.180 ;
        RECT 152.020 149.980 152.340 150.040 ;
        RECT 147.510 149.840 152.340 149.980 ;
        RECT 144.200 149.780 144.520 149.840 ;
        RECT 146.975 149.795 147.265 149.840 ;
        RECT 152.020 149.780 152.340 149.840 ;
        RECT 22.690 149.160 157.810 149.640 ;
        RECT 26.900 148.960 27.220 149.020 ;
        RECT 27.375 148.960 27.665 149.005 ;
        RECT 26.900 148.820 27.665 148.960 ;
        RECT 26.900 148.760 27.220 148.820 ;
        RECT 27.375 148.775 27.665 148.820 ;
        RECT 29.660 148.960 29.980 149.020 ;
        RECT 32.880 148.960 33.200 149.020 ;
        RECT 29.660 148.820 33.200 148.960 ;
        RECT 29.660 148.760 29.980 148.820 ;
        RECT 32.880 148.760 33.200 148.820 ;
        RECT 45.300 148.960 45.620 149.020 ;
        RECT 47.155 148.960 47.445 149.005 ;
        RECT 45.300 148.820 47.445 148.960 ;
        RECT 45.300 148.760 45.620 148.820 ;
        RECT 47.155 148.775 47.445 148.820 ;
        RECT 57.720 148.960 58.040 149.020 ;
        RECT 60.495 148.960 60.785 149.005 ;
        RECT 57.720 148.820 60.785 148.960 ;
        RECT 57.720 148.760 58.040 148.820 ;
        RECT 60.495 148.775 60.785 148.820 ;
        RECT 63.715 148.960 64.005 149.005 ;
        RECT 66.000 148.960 66.320 149.020 ;
        RECT 63.715 148.820 66.320 148.960 ;
        RECT 63.715 148.775 64.005 148.820 ;
        RECT 33.310 148.620 33.600 148.665 ;
        RECT 33.800 148.620 34.120 148.680 ;
        RECT 60.570 148.620 60.710 148.775 ;
        RECT 66.000 148.760 66.320 148.820 ;
        RECT 66.920 148.760 67.240 149.020 ;
        RECT 71.535 148.960 71.825 149.005 ;
        RECT 70.690 148.820 71.825 148.960 ;
        RECT 63.240 148.620 63.560 148.680 ;
        RECT 24.230 148.480 32.190 148.620 ;
        RECT 24.230 148.340 24.370 148.480 ;
        RECT 24.140 148.080 24.460 148.340 ;
        RECT 25.060 148.080 25.380 148.340 ;
        RECT 30.595 148.280 30.885 148.325 ;
        RECT 31.040 148.280 31.360 148.340 ;
        RECT 32.050 148.325 32.190 148.480 ;
        RECT 33.310 148.480 34.120 148.620 ;
        RECT 33.310 148.435 33.600 148.480 ;
        RECT 33.800 148.420 34.120 148.480 ;
        RECT 39.870 148.480 51.050 148.620 ;
        RECT 60.570 148.480 63.560 148.620 ;
        RECT 39.870 148.325 40.010 148.480 ;
        RECT 41.160 148.325 41.480 148.340 ;
        RECT 30.595 148.140 31.360 148.280 ;
        RECT 30.595 148.095 30.885 148.140 ;
        RECT 31.040 148.080 31.360 148.140 ;
        RECT 31.975 148.095 32.265 148.325 ;
        RECT 39.795 148.095 40.085 148.325 ;
        RECT 41.130 148.280 41.480 148.325 ;
        RECT 40.965 148.140 41.480 148.280 ;
        RECT 41.130 148.095 41.480 148.140 ;
        RECT 41.160 148.080 41.480 148.095 ;
        RECT 47.140 148.080 47.460 148.340 ;
        RECT 50.910 148.325 51.050 148.480 ;
        RECT 63.240 148.420 63.560 148.480 ;
        RECT 48.075 148.095 48.365 148.325 ;
        RECT 50.835 148.280 51.125 148.325 ;
        RECT 51.280 148.280 51.600 148.340 ;
        RECT 52.200 148.325 52.520 148.340 ;
        RECT 52.170 148.280 52.520 148.325 ;
        RECT 50.835 148.140 51.600 148.280 ;
        RECT 52.005 148.140 52.520 148.280 ;
        RECT 50.835 148.095 51.125 148.140 ;
        RECT 31.515 147.755 31.805 147.985 ;
        RECT 32.855 147.940 33.145 147.985 ;
        RECT 34.045 147.940 34.335 147.985 ;
        RECT 36.565 147.940 36.855 147.985 ;
        RECT 32.855 147.800 36.855 147.940 ;
        RECT 32.855 147.755 33.145 147.800 ;
        RECT 34.045 147.755 34.335 147.800 ;
        RECT 36.565 147.755 36.855 147.800 ;
        RECT 40.675 147.940 40.965 147.985 ;
        RECT 41.865 147.940 42.155 147.985 ;
        RECT 44.385 147.940 44.675 147.985 ;
        RECT 40.675 147.800 44.675 147.940 ;
        RECT 48.150 147.940 48.290 148.095 ;
        RECT 51.280 148.080 51.600 148.140 ;
        RECT 52.170 148.095 52.520 148.140 ;
        RECT 60.035 148.095 60.325 148.325 ;
        RECT 60.955 148.095 61.245 148.325 ;
        RECT 62.335 148.280 62.625 148.325 ;
        RECT 62.780 148.280 63.100 148.340 ;
        RECT 62.335 148.140 63.100 148.280 ;
        RECT 62.335 148.095 62.625 148.140 ;
        RECT 52.200 148.080 52.520 148.095 ;
        RECT 51.715 147.940 52.005 147.985 ;
        RECT 52.905 147.940 53.195 147.985 ;
        RECT 55.425 147.940 55.715 147.985 ;
        RECT 48.150 147.800 51.050 147.940 ;
        RECT 40.675 147.755 40.965 147.800 ;
        RECT 41.865 147.755 42.155 147.800 ;
        RECT 44.385 147.755 44.675 147.800 ;
        RECT 26.900 147.400 27.220 147.660 ;
        RECT 31.590 147.260 31.730 147.755 ;
        RECT 32.460 147.600 32.750 147.645 ;
        RECT 34.560 147.600 34.850 147.645 ;
        RECT 36.130 147.600 36.420 147.645 ;
        RECT 32.460 147.460 36.420 147.600 ;
        RECT 32.460 147.415 32.750 147.460 ;
        RECT 34.560 147.415 34.850 147.460 ;
        RECT 36.130 147.415 36.420 147.460 ;
        RECT 40.280 147.600 40.570 147.645 ;
        RECT 42.380 147.600 42.670 147.645 ;
        RECT 43.950 147.600 44.240 147.645 ;
        RECT 48.980 147.600 49.300 147.660 ;
        RECT 40.280 147.460 44.240 147.600 ;
        RECT 40.280 147.415 40.570 147.460 ;
        RECT 42.380 147.415 42.670 147.460 ;
        RECT 43.950 147.415 44.240 147.460 ;
        RECT 44.470 147.460 49.300 147.600 ;
        RECT 37.940 147.260 38.260 147.320 ;
        RECT 38.875 147.260 39.165 147.305 ;
        RECT 31.590 147.120 39.165 147.260 ;
        RECT 37.940 147.060 38.260 147.120 ;
        RECT 38.875 147.075 39.165 147.120 ;
        RECT 40.700 147.260 41.020 147.320 ;
        RECT 44.470 147.260 44.610 147.460 ;
        RECT 48.980 147.400 49.300 147.460 ;
        RECT 40.700 147.120 44.610 147.260 ;
        RECT 46.695 147.260 46.985 147.305 ;
        RECT 50.360 147.260 50.680 147.320 ;
        RECT 46.695 147.120 50.680 147.260 ;
        RECT 50.910 147.260 51.050 147.800 ;
        RECT 51.715 147.800 55.715 147.940 ;
        RECT 51.715 147.755 52.005 147.800 ;
        RECT 52.905 147.755 53.195 147.800 ;
        RECT 55.425 147.755 55.715 147.800 ;
        RECT 51.320 147.600 51.610 147.645 ;
        RECT 53.420 147.600 53.710 147.645 ;
        RECT 54.990 147.600 55.280 147.645 ;
        RECT 51.320 147.460 55.280 147.600 ;
        RECT 60.110 147.600 60.250 148.095 ;
        RECT 61.030 147.940 61.170 148.095 ;
        RECT 62.780 148.080 63.100 148.140 ;
        RECT 63.700 148.280 64.020 148.340 ;
        RECT 67.010 148.280 67.150 148.760 ;
        RECT 69.850 148.620 70.140 148.665 ;
        RECT 70.690 148.620 70.830 148.820 ;
        RECT 71.535 148.775 71.825 148.820 ;
        RECT 75.200 148.760 75.520 149.020 ;
        RECT 81.640 148.960 81.960 149.020 ;
        RECT 88.540 148.960 88.860 149.020 ;
        RECT 81.640 148.820 88.860 148.960 ;
        RECT 81.640 148.760 81.960 148.820 ;
        RECT 88.540 148.760 88.860 148.820 ;
        RECT 91.300 148.960 91.620 149.020 ;
        RECT 93.155 148.960 93.445 149.005 ;
        RECT 91.300 148.820 93.445 148.960 ;
        RECT 91.300 148.760 91.620 148.820 ;
        RECT 93.155 148.775 93.445 148.820 ;
        RECT 97.740 148.960 98.060 149.020 ;
        RECT 100.515 148.960 100.805 149.005 ;
        RECT 97.740 148.820 100.805 148.960 ;
        RECT 97.740 148.760 98.060 148.820 ;
        RECT 100.515 148.775 100.805 148.820 ;
        RECT 102.340 148.960 102.660 149.020 ;
        RECT 102.815 148.960 103.105 149.005 ;
        RECT 107.860 148.960 108.180 149.020 ;
        RECT 102.340 148.820 103.105 148.960 ;
        RECT 102.340 148.760 102.660 148.820 ;
        RECT 102.815 148.775 103.105 148.820 ;
        RECT 103.350 148.820 108.180 148.960 ;
        RECT 92.695 148.620 92.985 148.665 ;
        RECT 94.520 148.620 94.840 148.680 ;
        RECT 103.350 148.620 103.490 148.820 ;
        RECT 107.860 148.760 108.180 148.820 ;
        RECT 122.120 148.760 122.440 149.020 ;
        RECT 123.515 148.960 123.805 149.005 ;
        RECT 124.880 148.960 125.200 149.020 ;
        RECT 123.515 148.820 125.200 148.960 ;
        RECT 123.515 148.775 123.805 148.820 ;
        RECT 124.880 148.760 125.200 148.820 ;
        RECT 129.480 148.960 129.800 149.020 ;
        RECT 129.480 148.820 131.550 148.960 ;
        RECT 129.480 148.760 129.800 148.820 ;
        RECT 109.700 148.620 110.020 148.680 ;
        RECT 116.600 148.620 116.920 148.680 ;
        RECT 69.850 148.480 70.830 148.620 ;
        RECT 71.150 148.480 82.330 148.620 ;
        RECT 69.850 148.435 70.140 148.480 ;
        RECT 71.150 148.340 71.290 148.480 ;
        RECT 82.190 148.340 82.330 148.480 ;
        RECT 88.630 148.480 91.530 148.620 ;
        RECT 63.700 148.140 65.770 148.280 ;
        RECT 67.010 148.140 70.830 148.280 ;
        RECT 63.700 148.080 64.020 148.140 ;
        RECT 63.790 147.940 63.930 148.080 ;
        RECT 61.030 147.800 63.930 147.940 ;
        RECT 60.940 147.600 61.260 147.660 ;
        RECT 60.110 147.460 61.260 147.600 ;
        RECT 51.320 147.415 51.610 147.460 ;
        RECT 53.420 147.415 53.710 147.460 ;
        RECT 54.990 147.415 55.280 147.460 ;
        RECT 60.940 147.400 61.260 147.460 ;
        RECT 61.400 147.600 61.720 147.660 ;
        RECT 61.875 147.600 62.165 147.645 ;
        RECT 65.080 147.600 65.400 147.660 ;
        RECT 61.400 147.460 65.400 147.600 ;
        RECT 61.400 147.400 61.720 147.460 ;
        RECT 61.875 147.415 62.165 147.460 ;
        RECT 65.080 147.400 65.400 147.460 ;
        RECT 54.500 147.260 54.820 147.320 ;
        RECT 50.910 147.120 54.820 147.260 ;
        RECT 40.700 147.060 41.020 147.120 ;
        RECT 46.695 147.075 46.985 147.120 ;
        RECT 50.360 147.060 50.680 147.120 ;
        RECT 54.500 147.060 54.820 147.120 ;
        RECT 59.100 147.060 59.420 147.320 ;
        RECT 64.175 147.260 64.465 147.305 ;
        RECT 65.630 147.260 65.770 148.140 ;
        RECT 66.485 147.940 66.775 147.985 ;
        RECT 69.005 147.940 69.295 147.985 ;
        RECT 70.195 147.940 70.485 147.985 ;
        RECT 66.485 147.800 70.485 147.940 ;
        RECT 70.690 147.940 70.830 148.140 ;
        RECT 71.060 148.080 71.380 148.340 ;
        RECT 80.720 148.325 81.040 148.340 ;
        RECT 72.455 148.095 72.745 148.325 ;
        RECT 80.720 148.095 81.125 148.325 ;
        RECT 72.530 147.940 72.670 148.095 ;
        RECT 80.720 148.080 81.040 148.095 ;
        RECT 82.100 148.080 82.420 148.340 ;
        RECT 82.560 148.080 82.880 148.340 ;
        RECT 88.630 148.325 88.770 148.480 ;
        RECT 88.555 148.095 88.845 148.325 ;
        RECT 89.475 148.280 89.765 148.325 ;
        RECT 91.390 148.280 91.530 148.480 ;
        RECT 92.695 148.480 103.490 148.620 ;
        RECT 106.570 148.480 116.920 148.620 ;
        RECT 92.695 148.435 92.985 148.480 ;
        RECT 94.520 148.420 94.840 148.480 ;
        RECT 96.820 148.280 97.140 148.340 ;
        RECT 89.475 148.140 91.070 148.280 ;
        RECT 91.390 148.140 97.140 148.280 ;
        RECT 89.475 148.095 89.765 148.140 ;
        RECT 70.690 147.800 72.670 147.940 ;
        RECT 77.525 147.940 77.815 147.985 ;
        RECT 80.045 147.940 80.335 147.985 ;
        RECT 81.235 147.940 81.525 147.985 ;
        RECT 77.525 147.800 81.525 147.940 ;
        RECT 66.485 147.755 66.775 147.800 ;
        RECT 69.005 147.755 69.295 147.800 ;
        RECT 70.195 147.755 70.485 147.800 ;
        RECT 77.525 147.755 77.815 147.800 ;
        RECT 80.045 147.755 80.335 147.800 ;
        RECT 81.235 147.755 81.525 147.800 ;
        RECT 66.920 147.600 67.210 147.645 ;
        RECT 68.490 147.600 68.780 147.645 ;
        RECT 70.590 147.600 70.880 147.645 ;
        RECT 66.920 147.460 70.880 147.600 ;
        RECT 66.920 147.415 67.210 147.460 ;
        RECT 68.490 147.415 68.780 147.460 ;
        RECT 70.590 147.415 70.880 147.460 ;
        RECT 71.060 147.600 71.380 147.660 ;
        RECT 71.980 147.600 72.300 147.660 ;
        RECT 90.930 147.645 91.070 148.140 ;
        RECT 92.770 148.000 92.910 148.140 ;
        RECT 96.820 148.080 97.140 148.140 ;
        RECT 102.355 148.280 102.645 148.325 ;
        RECT 102.355 148.140 104.870 148.280 ;
        RECT 102.355 148.095 102.645 148.140 ;
        RECT 92.680 147.740 93.000 148.000 ;
        RECT 93.140 147.940 93.460 148.000 ;
        RECT 93.615 147.940 93.905 147.985 ;
        RECT 103.275 147.940 103.565 147.985 ;
        RECT 93.140 147.800 103.565 147.940 ;
        RECT 93.140 147.740 93.460 147.800 ;
        RECT 93.615 147.755 93.905 147.800 ;
        RECT 103.275 147.755 103.565 147.800 ;
        RECT 77.960 147.600 78.250 147.645 ;
        RECT 79.530 147.600 79.820 147.645 ;
        RECT 81.630 147.600 81.920 147.645 ;
        RECT 71.060 147.460 74.050 147.600 ;
        RECT 71.060 147.400 71.380 147.460 ;
        RECT 71.980 147.400 72.300 147.460 ;
        RECT 66.460 147.260 66.780 147.320 ;
        RECT 72.440 147.260 72.760 147.320 ;
        RECT 64.175 147.120 72.760 147.260 ;
        RECT 73.910 147.260 74.050 147.460 ;
        RECT 77.960 147.460 81.920 147.600 ;
        RECT 77.960 147.415 78.250 147.460 ;
        RECT 79.530 147.415 79.820 147.460 ;
        RECT 81.630 147.415 81.920 147.460 ;
        RECT 90.855 147.415 91.145 147.645 ;
        RECT 83.035 147.260 83.325 147.305 ;
        RECT 73.910 147.120 83.325 147.260 ;
        RECT 64.175 147.075 64.465 147.120 ;
        RECT 66.460 147.060 66.780 147.120 ;
        RECT 72.440 147.060 72.760 147.120 ;
        RECT 83.035 147.075 83.325 147.120 ;
        RECT 90.395 147.260 90.685 147.305 ;
        RECT 91.300 147.260 91.620 147.320 ;
        RECT 90.395 147.120 91.620 147.260 ;
        RECT 104.730 147.260 104.870 148.140 ;
        RECT 105.100 148.080 105.420 148.340 ;
        RECT 106.570 148.325 106.710 148.480 ;
        RECT 109.700 148.420 110.020 148.480 ;
        RECT 114.850 148.325 114.990 148.480 ;
        RECT 116.600 148.420 116.920 148.480 ;
        RECT 121.660 148.420 121.980 148.680 ;
        RECT 106.495 148.095 106.785 148.325 ;
        RECT 107.775 148.280 108.065 148.325 ;
        RECT 107.030 148.140 108.065 148.280 ;
        RECT 107.030 147.940 107.170 148.140 ;
        RECT 107.775 148.095 108.065 148.140 ;
        RECT 114.775 148.095 115.065 148.325 ;
        RECT 116.110 148.280 116.400 148.325 ;
        RECT 121.750 148.280 121.890 148.420 ;
        RECT 116.110 148.140 121.890 148.280 ;
        RECT 122.210 148.280 122.350 148.760 ;
        RECT 131.410 148.620 131.550 148.820 ;
        RECT 132.700 148.760 133.020 149.020 ;
        RECT 135.460 148.760 135.780 149.020 ;
        RECT 140.060 148.960 140.380 149.020 ;
        RECT 141.455 148.960 141.745 149.005 ;
        RECT 142.835 148.960 143.125 149.005 ;
        RECT 140.060 148.820 143.125 148.960 ;
        RECT 140.060 148.760 140.380 148.820 ;
        RECT 141.455 148.775 141.745 148.820 ;
        RECT 142.835 148.775 143.125 148.820 ;
        RECT 143.280 148.960 143.600 149.020 ;
        RECT 143.280 148.820 147.650 148.960 ;
        RECT 143.280 148.760 143.600 148.820 ;
        RECT 135.550 148.620 135.690 148.760 ;
        RECT 124.050 148.480 130.630 148.620 ;
        RECT 123.055 148.280 123.345 148.325 ;
        RECT 122.210 148.140 123.345 148.280 ;
        RECT 116.110 148.095 116.400 148.140 ;
        RECT 123.055 148.095 123.345 148.140 ;
        RECT 106.110 147.800 107.170 147.940 ;
        RECT 107.375 147.940 107.665 147.985 ;
        RECT 108.565 147.940 108.855 147.985 ;
        RECT 111.085 147.940 111.375 147.985 ;
        RECT 107.375 147.800 111.375 147.940 ;
        RECT 106.110 147.645 106.250 147.800 ;
        RECT 107.375 147.755 107.665 147.800 ;
        RECT 108.565 147.755 108.855 147.800 ;
        RECT 111.085 147.755 111.375 147.800 ;
        RECT 115.655 147.940 115.945 147.985 ;
        RECT 116.845 147.940 117.135 147.985 ;
        RECT 119.365 147.940 119.655 147.985 ;
        RECT 115.655 147.800 119.655 147.940 ;
        RECT 115.655 147.755 115.945 147.800 ;
        RECT 116.845 147.755 117.135 147.800 ;
        RECT 119.365 147.755 119.655 147.800 ;
        RECT 121.200 147.940 121.520 148.000 ;
        RECT 124.050 147.940 124.190 148.480 ;
        RECT 124.420 148.080 124.740 148.340 ;
        RECT 130.490 148.325 130.630 148.480 ;
        RECT 131.410 148.480 135.690 148.620 ;
        RECT 135.890 148.620 136.180 148.665 ;
        RECT 137.300 148.620 137.620 148.680 ;
        RECT 135.890 148.480 137.620 148.620 ;
        RECT 129.495 148.095 129.785 148.325 ;
        RECT 130.415 148.095 130.705 148.325 ;
        RECT 121.200 147.800 124.190 147.940 ;
        RECT 121.200 147.740 121.520 147.800 ;
        RECT 125.340 147.740 125.660 148.000 ;
        RECT 106.035 147.415 106.325 147.645 ;
        RECT 106.980 147.600 107.270 147.645 ;
        RECT 109.080 147.600 109.370 147.645 ;
        RECT 110.650 147.600 110.940 147.645 ;
        RECT 115.260 147.600 115.550 147.645 ;
        RECT 117.360 147.600 117.650 147.645 ;
        RECT 118.930 147.600 119.220 147.645 ;
        RECT 106.980 147.460 110.940 147.600 ;
        RECT 106.980 147.415 107.270 147.460 ;
        RECT 109.080 147.415 109.370 147.460 ;
        RECT 110.650 147.415 110.940 147.460 ;
        RECT 111.170 147.460 114.070 147.600 ;
        RECT 111.170 147.320 111.310 147.460 ;
        RECT 111.080 147.260 111.400 147.320 ;
        RECT 104.730 147.120 111.400 147.260 ;
        RECT 90.395 147.075 90.685 147.120 ;
        RECT 91.300 147.060 91.620 147.120 ;
        RECT 111.080 147.060 111.400 147.120 ;
        RECT 113.380 147.060 113.700 147.320 ;
        RECT 113.930 147.260 114.070 147.460 ;
        RECT 115.260 147.460 119.220 147.600 ;
        RECT 121.290 147.600 121.430 147.740 ;
        RECT 121.675 147.600 121.965 147.645 ;
        RECT 121.290 147.460 121.965 147.600 ;
        RECT 129.570 147.600 129.710 148.095 ;
        RECT 130.860 148.080 131.180 148.340 ;
        RECT 131.410 148.325 131.550 148.480 ;
        RECT 135.890 148.435 136.180 148.480 ;
        RECT 137.300 148.420 137.620 148.480 ;
        RECT 144.200 148.420 144.520 148.680 ;
        RECT 146.975 148.435 147.265 148.665 ;
        RECT 131.335 148.095 131.625 148.325 ;
        RECT 134.555 148.280 134.845 148.325 ;
        RECT 135.000 148.280 135.320 148.340 ;
        RECT 134.555 148.140 135.320 148.280 ;
        RECT 134.555 148.095 134.845 148.140 ;
        RECT 135.000 148.080 135.320 148.140 ;
        RECT 141.440 148.280 141.760 148.340 ;
        RECT 143.755 148.295 144.045 148.325 ;
        RECT 142.910 148.280 144.045 148.295 ;
        RECT 141.440 148.155 144.045 148.280 ;
        RECT 141.440 148.140 143.050 148.155 ;
        RECT 141.440 148.080 141.760 148.140 ;
        RECT 143.755 148.095 144.045 148.155 ;
        RECT 135.435 147.940 135.725 147.985 ;
        RECT 136.625 147.940 136.915 147.985 ;
        RECT 139.145 147.940 139.435 147.985 ;
        RECT 135.435 147.800 139.435 147.940 ;
        RECT 135.435 147.755 135.725 147.800 ;
        RECT 136.625 147.755 136.915 147.800 ;
        RECT 139.145 147.755 139.435 147.800 ;
        RECT 141.915 147.940 142.205 147.985 ;
        RECT 142.360 147.940 142.680 148.000 ;
        RECT 144.290 147.940 144.430 148.420 ;
        RECT 141.915 147.800 144.430 147.940 ;
        RECT 141.915 147.755 142.205 147.800 ;
        RECT 142.360 147.740 142.680 147.800 ;
        RECT 134.080 147.600 134.400 147.660 ;
        RECT 129.570 147.460 134.400 147.600 ;
        RECT 115.260 147.415 115.550 147.460 ;
        RECT 117.360 147.415 117.650 147.460 ;
        RECT 118.930 147.415 119.220 147.460 ;
        RECT 121.675 147.415 121.965 147.460 ;
        RECT 134.080 147.400 134.400 147.460 ;
        RECT 135.040 147.600 135.330 147.645 ;
        RECT 137.140 147.600 137.430 147.645 ;
        RECT 138.710 147.600 139.000 147.645 ;
        RECT 135.040 147.460 139.000 147.600 ;
        RECT 135.040 147.415 135.330 147.460 ;
        RECT 137.140 147.415 137.430 147.460 ;
        RECT 138.710 147.415 139.000 147.460 ;
        RECT 144.200 147.600 144.520 147.660 ;
        RECT 144.675 147.600 144.965 147.645 ;
        RECT 145.135 147.600 145.425 147.645 ;
        RECT 147.050 147.600 147.190 148.435 ;
        RECT 147.510 147.940 147.650 148.820 ;
        RECT 147.895 148.775 148.185 149.005 ;
        RECT 147.970 148.280 148.110 148.775 ;
        RECT 149.260 148.760 149.580 149.020 ;
        RECT 148.355 148.280 148.645 148.325 ;
        RECT 147.970 148.140 148.645 148.280 ;
        RECT 148.355 148.095 148.645 148.140 ;
        RECT 155.240 147.940 155.560 148.000 ;
        RECT 147.510 147.800 155.560 147.940 ;
        RECT 155.240 147.740 155.560 147.800 ;
        RECT 144.200 147.460 145.425 147.600 ;
        RECT 144.200 147.400 144.520 147.460 ;
        RECT 144.675 147.415 144.965 147.460 ;
        RECT 145.135 147.415 145.425 147.460 ;
        RECT 145.570 147.460 147.190 147.600 ;
        RECT 118.440 147.260 118.760 147.320 ;
        RECT 113.930 147.120 118.760 147.260 ;
        RECT 118.440 147.060 118.760 147.120 ;
        RECT 122.120 147.060 122.440 147.320 ;
        RECT 125.800 147.260 126.120 147.320 ;
        RECT 130.860 147.260 131.180 147.320 ;
        RECT 125.800 147.120 131.180 147.260 ;
        RECT 125.800 147.060 126.120 147.120 ;
        RECT 130.860 147.060 131.180 147.120 ;
        RECT 143.740 147.260 144.060 147.320 ;
        RECT 145.570 147.260 145.710 147.460 ;
        RECT 143.740 147.120 145.710 147.260 ;
        RECT 143.740 147.060 144.060 147.120 ;
        RECT 146.960 147.060 147.280 147.320 ;
        RECT 22.690 146.440 157.010 146.920 ;
        RECT 33.815 146.240 34.105 146.285 ;
        RECT 34.260 146.240 34.580 146.300 ;
        RECT 52.200 146.240 52.520 146.300 ;
        RECT 52.675 146.240 52.965 146.285 ;
        RECT 33.815 146.100 34.580 146.240 ;
        RECT 33.815 146.055 34.105 146.100 ;
        RECT 34.260 146.040 34.580 146.100 ;
        RECT 35.730 146.100 45.990 146.240 ;
        RECT 35.730 145.960 35.870 146.100 ;
        RECT 31.960 145.700 32.280 145.960 ;
        RECT 35.180 145.900 35.500 145.960 ;
        RECT 33.430 145.760 35.500 145.900 ;
        RECT 29.660 145.360 29.980 145.620 ;
        RECT 32.050 145.560 32.190 145.700 ;
        RECT 33.430 145.605 33.570 145.760 ;
        RECT 35.180 145.700 35.500 145.760 ;
        RECT 35.640 145.700 35.960 145.960 ;
        RECT 37.020 145.900 37.340 145.960 ;
        RECT 37.940 145.900 38.260 145.960 ;
        RECT 45.850 145.945 45.990 146.100 ;
        RECT 52.200 146.100 52.965 146.240 ;
        RECT 52.200 146.040 52.520 146.100 ;
        RECT 52.675 146.055 52.965 146.100 ;
        RECT 56.355 146.240 56.645 146.285 ;
        RECT 61.860 146.240 62.180 146.300 ;
        RECT 56.355 146.100 62.180 146.240 ;
        RECT 56.355 146.055 56.645 146.100 ;
        RECT 61.860 146.040 62.180 146.100 ;
        RECT 69.680 146.240 70.000 146.300 ;
        RECT 71.995 146.240 72.285 146.285 ;
        RECT 69.680 146.100 72.285 146.240 ;
        RECT 69.680 146.040 70.000 146.100 ;
        RECT 71.995 146.055 72.285 146.100 ;
        RECT 82.100 146.040 82.420 146.300 ;
        RECT 95.440 146.040 95.760 146.300 ;
        RECT 99.135 146.240 99.425 146.285 ;
        RECT 100.960 146.240 101.280 146.300 ;
        RECT 99.135 146.100 101.280 146.240 ;
        RECT 99.135 146.055 99.425 146.100 ;
        RECT 100.960 146.040 101.280 146.100 ;
        RECT 105.100 146.240 105.420 146.300 ;
        RECT 108.795 146.240 109.085 146.285 ;
        RECT 118.440 146.240 118.760 146.300 ;
        RECT 105.100 146.100 109.085 146.240 ;
        RECT 105.100 146.040 105.420 146.100 ;
        RECT 108.795 146.055 109.085 146.100 ;
        RECT 116.230 146.100 118.760 146.240 ;
        RECT 37.020 145.760 40.010 145.900 ;
        RECT 37.020 145.700 37.340 145.760 ;
        RECT 37.940 145.700 38.260 145.760 ;
        RECT 39.870 145.605 40.010 145.760 ;
        RECT 45.775 145.715 46.065 145.945 ;
        RECT 58.195 145.900 58.485 145.945 ;
        RECT 59.100 145.900 59.420 145.960 ;
        RECT 64.620 145.900 64.940 145.960 ;
        RECT 49.990 145.760 55.190 145.900 ;
        RECT 33.300 145.560 33.590 145.605 ;
        RECT 32.050 145.420 33.590 145.560 ;
        RECT 33.300 145.375 33.590 145.420 ;
        RECT 34.275 145.560 34.565 145.605 ;
        RECT 34.275 145.420 38.170 145.560 ;
        RECT 34.275 145.375 34.565 145.420 ;
        RECT 26.900 145.020 27.220 145.280 ;
        RECT 29.215 145.220 29.505 145.265 ;
        RECT 29.750 145.220 29.890 145.360 ;
        RECT 29.215 145.080 29.890 145.220 ;
        RECT 31.040 145.220 31.360 145.280 ;
        RECT 31.040 145.080 32.145 145.220 ;
        RECT 29.215 145.035 29.505 145.080 ;
        RECT 31.040 145.020 31.360 145.080 ;
        RECT 26.990 144.880 27.130 145.020 ;
        RECT 32.005 144.880 32.145 145.080 ;
        RECT 34.350 144.880 34.490 145.375 ;
        RECT 38.030 145.280 38.170 145.420 ;
        RECT 39.795 145.375 40.085 145.605 ;
        RECT 34.735 145.220 35.025 145.265 ;
        RECT 37.035 145.220 37.325 145.265 ;
        RECT 34.735 145.080 37.325 145.220 ;
        RECT 34.735 145.035 35.025 145.080 ;
        RECT 37.035 145.035 37.325 145.080 ;
        RECT 37.940 145.020 38.260 145.280 ;
        RECT 44.395 145.220 44.685 145.265 ;
        RECT 45.300 145.220 45.620 145.280 ;
        RECT 44.395 145.080 45.620 145.220 ;
        RECT 44.395 145.035 44.685 145.080 ;
        RECT 45.300 145.020 45.620 145.080 ;
        RECT 48.980 145.220 49.300 145.280 ;
        RECT 49.990 145.220 50.130 145.760 ;
        RECT 50.375 145.560 50.665 145.605 ;
        RECT 54.500 145.560 54.820 145.620 ;
        RECT 50.375 145.420 54.820 145.560 ;
        RECT 55.050 145.560 55.190 145.760 ;
        RECT 58.195 145.760 59.420 145.900 ;
        RECT 58.195 145.715 58.485 145.760 ;
        RECT 59.100 145.700 59.420 145.760 ;
        RECT 63.330 145.760 64.940 145.900 ;
        RECT 55.050 145.420 62.550 145.560 ;
        RECT 50.375 145.375 50.665 145.420 ;
        RECT 54.500 145.360 54.820 145.420 ;
        RECT 62.410 145.280 62.550 145.420 ;
        RECT 48.980 145.080 50.130 145.220 ;
        RECT 51.740 145.220 52.060 145.280 ;
        RECT 52.215 145.220 52.505 145.265 ;
        RECT 51.740 145.080 52.505 145.220 ;
        RECT 48.980 145.020 49.300 145.080 ;
        RECT 51.740 145.020 52.060 145.080 ;
        RECT 52.215 145.035 52.505 145.080 ;
        RECT 53.135 145.220 53.425 145.265 ;
        RECT 53.580 145.220 53.900 145.280 ;
        RECT 53.135 145.080 53.900 145.220 ;
        RECT 53.135 145.035 53.425 145.080 ;
        RECT 53.580 145.020 53.900 145.080 ;
        RECT 62.320 145.020 62.640 145.280 ;
        RECT 56.355 144.880 56.645 144.925 ;
        RECT 63.330 144.880 63.470 145.760 ;
        RECT 64.620 145.700 64.940 145.760 ;
        RECT 65.080 145.900 65.400 145.960 ;
        RECT 67.840 145.900 68.160 145.960 ;
        RECT 65.080 145.760 68.160 145.900 ;
        RECT 65.080 145.700 65.400 145.760 ;
        RECT 67.840 145.700 68.160 145.760 ;
        RECT 89.040 145.900 89.330 145.945 ;
        RECT 91.140 145.900 91.430 145.945 ;
        RECT 92.710 145.900 93.000 145.945 ;
        RECT 89.040 145.760 93.000 145.900 ;
        RECT 89.040 145.715 89.330 145.760 ;
        RECT 91.140 145.715 91.430 145.760 ;
        RECT 92.710 145.715 93.000 145.760 ;
        RECT 63.715 145.560 64.005 145.605 ;
        RECT 68.300 145.560 68.620 145.620 ;
        RECT 75.200 145.560 75.520 145.620 ;
        RECT 63.715 145.420 68.620 145.560 ;
        RECT 63.715 145.375 64.005 145.420 ;
        RECT 68.300 145.360 68.620 145.420 ;
        RECT 69.770 145.420 75.520 145.560 ;
        RECT 64.620 145.020 64.940 145.280 ;
        RECT 65.080 145.020 65.400 145.280 ;
        RECT 66.935 145.220 67.225 145.265 ;
        RECT 69.770 145.220 69.910 145.420 ;
        RECT 75.200 145.360 75.520 145.420 ;
        RECT 89.435 145.560 89.725 145.605 ;
        RECT 90.625 145.560 90.915 145.605 ;
        RECT 93.145 145.560 93.435 145.605 ;
        RECT 89.435 145.420 93.435 145.560 ;
        RECT 89.435 145.375 89.725 145.420 ;
        RECT 90.625 145.375 90.915 145.420 ;
        RECT 93.145 145.375 93.435 145.420 ;
        RECT 94.980 145.560 95.300 145.620 ;
        RECT 94.980 145.420 100.730 145.560 ;
        RECT 94.980 145.360 95.300 145.420 ;
        RECT 66.935 145.080 69.910 145.220 ;
        RECT 66.935 145.035 67.225 145.080 ;
        RECT 70.140 145.020 70.460 145.280 ;
        RECT 75.675 145.220 75.965 145.265 ;
        RECT 77.960 145.220 78.280 145.280 ;
        RECT 75.675 145.080 78.280 145.220 ;
        RECT 75.675 145.035 75.965 145.080 ;
        RECT 26.990 144.740 31.730 144.880 ;
        RECT 32.005 144.740 34.490 144.880 ;
        RECT 54.590 144.740 63.470 144.880 ;
        RECT 64.160 144.880 64.480 144.940 ;
        RECT 75.750 144.880 75.890 145.035 ;
        RECT 77.960 145.020 78.280 145.080 ;
        RECT 86.240 145.220 86.560 145.280 ;
        RECT 88.555 145.220 88.845 145.265 ;
        RECT 97.280 145.220 97.600 145.280 ;
        RECT 86.240 145.080 97.600 145.220 ;
        RECT 86.240 145.020 86.560 145.080 ;
        RECT 88.555 145.035 88.845 145.080 ;
        RECT 97.280 145.020 97.600 145.080 ;
        RECT 97.755 145.220 98.045 145.265 ;
        RECT 98.215 145.220 98.505 145.265 ;
        RECT 97.755 145.080 98.505 145.220 ;
        RECT 97.755 145.035 98.045 145.080 ;
        RECT 98.215 145.035 98.505 145.080 ;
        RECT 64.160 144.740 75.890 144.880 ;
        RECT 89.890 144.880 90.180 144.925 ;
        RECT 90.840 144.880 91.160 144.940 ;
        RECT 89.890 144.740 91.160 144.880 ;
        RECT 31.590 144.600 31.730 144.740 ;
        RECT 54.590 144.600 54.730 144.740 ;
        RECT 56.355 144.695 56.645 144.740 ;
        RECT 64.160 144.680 64.480 144.740 ;
        RECT 89.890 144.695 90.180 144.740 ;
        RECT 90.840 144.680 91.160 144.740 ;
        RECT 95.440 144.680 95.760 144.940 ;
        RECT 95.900 144.680 96.220 144.940 ;
        RECT 96.835 144.695 97.125 144.925 ;
        RECT 100.590 144.880 100.730 145.420 ;
        RECT 101.050 145.220 101.190 146.040 ;
        RECT 107.415 145.560 107.705 145.605 ;
        RECT 109.240 145.560 109.560 145.620 ;
        RECT 116.230 145.605 116.370 146.100 ;
        RECT 118.440 146.040 118.760 146.100 ;
        RECT 118.915 146.240 119.205 146.285 ;
        RECT 120.740 146.240 121.060 146.300 ;
        RECT 124.880 146.240 125.200 146.300 ;
        RECT 118.915 146.100 121.060 146.240 ;
        RECT 118.915 146.055 119.205 146.100 ;
        RECT 120.740 146.040 121.060 146.100 ;
        RECT 121.290 146.100 125.200 146.240 ;
        RECT 121.290 145.900 121.430 146.100 ;
        RECT 124.880 146.040 125.200 146.100 ;
        RECT 125.340 146.240 125.660 146.300 ;
        RECT 128.575 146.240 128.865 146.285 ;
        RECT 125.340 146.100 128.865 146.240 ;
        RECT 125.340 146.040 125.660 146.100 ;
        RECT 128.575 146.055 128.865 146.100 ;
        RECT 116.690 145.760 121.430 145.900 ;
        RECT 122.160 145.900 122.450 145.945 ;
        RECT 124.260 145.900 124.550 145.945 ;
        RECT 125.830 145.900 126.120 145.945 ;
        RECT 122.160 145.760 126.120 145.900 ;
        RECT 112.015 145.560 112.305 145.605 ;
        RECT 116.155 145.560 116.445 145.605 ;
        RECT 107.415 145.420 116.445 145.560 ;
        RECT 107.415 145.375 107.705 145.420 ;
        RECT 109.240 145.360 109.560 145.420 ;
        RECT 112.015 145.375 112.305 145.420 ;
        RECT 116.155 145.375 116.445 145.420 ;
        RECT 103.735 145.220 104.025 145.265 ;
        RECT 104.180 145.220 104.500 145.280 ;
        RECT 101.050 145.080 104.500 145.220 ;
        RECT 103.735 145.035 104.025 145.080 ;
        RECT 104.180 145.020 104.500 145.080 ;
        RECT 106.035 145.035 106.325 145.265 ;
        RECT 111.095 145.220 111.385 145.265 ;
        RECT 112.460 145.220 112.780 145.280 ;
        RECT 111.095 145.080 112.780 145.220 ;
        RECT 111.095 145.035 111.385 145.080 ;
        RECT 106.110 144.880 106.250 145.035 ;
        RECT 112.460 145.020 112.780 145.080 ;
        RECT 116.690 144.925 116.830 145.760 ;
        RECT 122.160 145.715 122.450 145.760 ;
        RECT 124.260 145.715 124.550 145.760 ;
        RECT 125.830 145.715 126.120 145.760 ;
        RECT 117.060 145.560 117.380 145.620 ;
        RECT 121.675 145.560 121.965 145.605 ;
        RECT 117.060 145.420 121.965 145.560 ;
        RECT 117.060 145.360 117.380 145.420 ;
        RECT 121.675 145.375 121.965 145.420 ;
        RECT 122.555 145.560 122.845 145.605 ;
        RECT 123.745 145.560 124.035 145.605 ;
        RECT 126.265 145.560 126.555 145.605 ;
        RECT 122.555 145.420 126.555 145.560 ;
        RECT 122.555 145.375 122.845 145.420 ;
        RECT 123.745 145.375 124.035 145.420 ;
        RECT 126.265 145.375 126.555 145.420 ;
        RECT 119.360 145.020 119.680 145.280 ;
        RECT 122.120 145.220 122.440 145.280 ;
        RECT 122.955 145.220 123.245 145.265 ;
        RECT 122.120 145.080 123.245 145.220 ;
        RECT 122.120 145.020 122.440 145.080 ;
        RECT 122.955 145.035 123.245 145.080 ;
        RECT 100.590 144.740 106.250 144.880 ;
        RECT 28.280 144.340 28.600 144.600 ;
        RECT 28.740 144.340 29.060 144.600 ;
        RECT 31.500 144.340 31.820 144.600 ;
        RECT 54.500 144.340 54.820 144.600 ;
        RECT 54.960 144.540 55.280 144.600 ;
        RECT 55.435 144.540 55.725 144.585 ;
        RECT 54.960 144.400 55.725 144.540 ;
        RECT 54.960 144.340 55.280 144.400 ;
        RECT 55.435 144.355 55.725 144.400 ;
        RECT 63.240 144.540 63.560 144.600 ;
        RECT 66.000 144.540 66.320 144.600 ;
        RECT 63.240 144.400 66.320 144.540 ;
        RECT 63.240 144.340 63.560 144.400 ;
        RECT 66.000 144.340 66.320 144.400 ;
        RECT 67.380 144.340 67.700 144.600 ;
        RECT 95.530 144.540 95.670 144.680 ;
        RECT 96.910 144.540 97.050 144.695 ;
        RECT 103.810 144.600 103.950 144.740 ;
        RECT 116.615 144.695 116.905 144.925 ;
        RECT 117.075 144.880 117.365 144.925 ;
        RECT 119.450 144.880 119.590 145.020 ;
        RECT 117.075 144.740 119.590 144.880 ;
        RECT 128.650 144.880 128.790 146.055 ;
        RECT 131.320 146.040 131.640 146.300 ;
        RECT 132.240 146.240 132.560 146.300 ;
        RECT 132.715 146.240 133.005 146.285 ;
        RECT 132.240 146.100 133.005 146.240 ;
        RECT 132.240 146.040 132.560 146.100 ;
        RECT 132.715 146.055 133.005 146.100 ;
        RECT 133.620 146.040 133.940 146.300 ;
        RECT 134.080 146.240 134.400 146.300 ;
        RECT 136.395 146.240 136.685 146.285 ;
        RECT 134.080 146.100 136.685 146.240 ;
        RECT 134.080 146.040 134.400 146.100 ;
        RECT 136.395 146.055 136.685 146.100 ;
        RECT 137.760 146.240 138.080 146.300 ;
        RECT 138.235 146.240 138.525 146.285 ;
        RECT 140.520 146.240 140.840 146.300 ;
        RECT 137.760 146.100 140.840 146.240 ;
        RECT 137.760 146.040 138.080 146.100 ;
        RECT 138.235 146.055 138.525 146.100 ;
        RECT 140.520 146.040 140.840 146.100 ;
        RECT 140.995 146.240 141.285 146.285 ;
        RECT 146.960 146.240 147.280 146.300 ;
        RECT 140.995 146.100 147.280 146.240 ;
        RECT 140.995 146.055 141.285 146.100 ;
        RECT 146.960 146.040 147.280 146.100 ;
        RECT 131.410 145.900 131.550 146.040 ;
        RECT 133.175 145.900 133.465 145.945 ;
        RECT 131.410 145.760 133.465 145.900 ;
        RECT 133.710 145.900 133.850 146.040 ;
        RECT 135.475 145.900 135.765 145.945 ;
        RECT 133.710 145.760 135.765 145.900 ;
        RECT 133.175 145.715 133.465 145.760 ;
        RECT 135.475 145.715 135.765 145.760 ;
        RECT 141.440 145.700 141.760 145.960 ;
        RECT 142.360 145.700 142.680 145.960 ;
        RECT 148.840 145.900 149.130 145.945 ;
        RECT 150.940 145.900 151.230 145.945 ;
        RECT 152.510 145.900 152.800 145.945 ;
        RECT 148.840 145.760 152.800 145.900 ;
        RECT 148.840 145.715 149.130 145.760 ;
        RECT 150.940 145.715 151.230 145.760 ;
        RECT 152.510 145.715 152.800 145.760 ;
        RECT 136.855 145.560 137.145 145.605 ;
        RECT 141.530 145.560 141.670 145.700 ;
        RECT 131.410 145.420 134.770 145.560 ;
        RECT 129.480 145.220 129.800 145.280 ;
        RECT 131.410 145.265 131.550 145.420 ;
        RECT 134.630 145.265 134.770 145.420 ;
        RECT 135.550 145.420 137.145 145.560 ;
        RECT 135.550 145.280 135.690 145.420 ;
        RECT 136.855 145.375 137.145 145.420 ;
        RECT 140.150 145.420 141.670 145.560 ;
        RECT 129.955 145.220 130.245 145.265 ;
        RECT 129.480 145.080 130.245 145.220 ;
        RECT 129.480 145.020 129.800 145.080 ;
        RECT 129.955 145.035 130.245 145.080 ;
        RECT 131.335 145.035 131.625 145.265 ;
        RECT 131.795 145.220 132.085 145.265 ;
        RECT 134.095 145.220 134.385 145.265 ;
        RECT 131.795 145.080 134.385 145.220 ;
        RECT 131.795 145.035 132.085 145.080 ;
        RECT 134.095 145.035 134.385 145.080 ;
        RECT 134.555 145.035 134.845 145.265 ;
        RECT 128.650 144.740 130.630 144.880 ;
        RECT 117.075 144.695 117.365 144.740 ;
        RECT 95.530 144.400 97.050 144.540 ;
        RECT 103.720 144.340 104.040 144.600 ;
        RECT 110.620 144.340 110.940 144.600 ;
        RECT 113.380 144.540 113.700 144.600 ;
        RECT 125.800 144.540 126.120 144.600 ;
        RECT 113.380 144.400 126.120 144.540 ;
        RECT 130.490 144.540 130.630 144.740 ;
        RECT 130.860 144.680 131.180 144.940 ;
        RECT 131.870 144.540 132.010 145.035 ;
        RECT 134.630 144.880 134.770 145.035 ;
        RECT 135.460 145.020 135.780 145.280 ;
        RECT 135.920 145.020 136.240 145.280 ;
        RECT 136.380 145.220 136.700 145.280 ;
        RECT 140.150 145.265 140.290 145.420 ;
        RECT 139.615 145.220 139.905 145.265 ;
        RECT 136.380 145.080 139.905 145.220 ;
        RECT 136.380 145.020 136.700 145.080 ;
        RECT 139.615 145.035 139.905 145.080 ;
        RECT 140.075 145.035 140.365 145.265 ;
        RECT 140.520 145.020 140.840 145.280 ;
        RECT 141.455 145.035 141.745 145.265 ;
        RECT 142.450 145.220 142.590 145.700 ;
        RECT 149.235 145.560 149.525 145.605 ;
        RECT 150.425 145.560 150.715 145.605 ;
        RECT 152.945 145.560 153.235 145.605 ;
        RECT 149.235 145.420 153.235 145.560 ;
        RECT 149.235 145.375 149.525 145.420 ;
        RECT 150.425 145.375 150.715 145.420 ;
        RECT 152.945 145.375 153.235 145.420 ;
        RECT 142.835 145.220 143.125 145.265 ;
        RECT 142.450 145.080 143.125 145.220 ;
        RECT 142.835 145.035 143.125 145.080 ;
        RECT 148.355 145.220 148.645 145.265 ;
        RECT 148.800 145.220 149.120 145.280 ;
        RECT 148.355 145.080 149.120 145.220 ;
        RECT 148.355 145.035 148.645 145.080 ;
        RECT 141.530 144.880 141.670 145.035 ;
        RECT 148.800 145.020 149.120 145.080 ;
        RECT 149.720 144.925 150.040 144.940 ;
        RECT 142.375 144.880 142.665 144.925 ;
        RECT 134.630 144.740 142.665 144.880 ;
        RECT 142.375 144.695 142.665 144.740 ;
        RECT 149.690 144.695 150.040 144.925 ;
        RECT 149.720 144.680 150.040 144.695 ;
        RECT 130.490 144.400 132.010 144.540 ;
        RECT 145.120 144.540 145.440 144.600 ;
        RECT 155.255 144.540 155.545 144.585 ;
        RECT 145.120 144.400 155.545 144.540 ;
        RECT 113.380 144.340 113.700 144.400 ;
        RECT 125.800 144.340 126.120 144.400 ;
        RECT 145.120 144.340 145.440 144.400 ;
        RECT 155.255 144.355 155.545 144.400 ;
        RECT 22.690 143.720 157.810 144.200 ;
        RECT 28.740 143.520 29.060 143.580 ;
        RECT 31.515 143.520 31.805 143.565 ;
        RECT 43.000 143.520 43.320 143.580 ;
        RECT 44.380 143.520 44.700 143.580 ;
        RECT 47.155 143.520 47.445 143.565 ;
        RECT 28.740 143.380 31.805 143.520 ;
        RECT 28.740 143.320 29.060 143.380 ;
        RECT 31.515 143.335 31.805 143.380 ;
        RECT 37.110 143.380 40.010 143.520 ;
        RECT 37.110 143.240 37.250 143.380 ;
        RECT 37.020 142.980 37.340 143.240 ;
        RECT 37.480 143.180 37.800 143.240 ;
        RECT 39.335 143.180 39.625 143.225 ;
        RECT 37.480 143.040 39.625 143.180 ;
        RECT 37.480 142.980 37.800 143.040 ;
        RECT 39.335 142.995 39.625 143.040 ;
        RECT 24.140 142.640 24.460 142.900 ;
        RECT 25.490 142.840 25.780 142.885 ;
        RECT 26.900 142.840 27.220 142.900 ;
        RECT 25.490 142.700 27.220 142.840 ;
        RECT 25.490 142.655 25.780 142.700 ;
        RECT 26.900 142.640 27.220 142.700 ;
        RECT 34.735 142.840 35.025 142.885 ;
        RECT 34.735 142.700 37.710 142.840 ;
        RECT 34.735 142.655 35.025 142.700 ;
        RECT 25.035 142.500 25.325 142.545 ;
        RECT 26.225 142.500 26.515 142.545 ;
        RECT 28.745 142.500 29.035 142.545 ;
        RECT 25.035 142.360 29.035 142.500 ;
        RECT 25.035 142.315 25.325 142.360 ;
        RECT 26.225 142.315 26.515 142.360 ;
        RECT 28.745 142.315 29.035 142.360 ;
        RECT 24.640 142.160 24.930 142.205 ;
        RECT 26.740 142.160 27.030 142.205 ;
        RECT 28.310 142.160 28.600 142.205 ;
        RECT 24.640 142.020 28.600 142.160 ;
        RECT 24.640 141.975 24.930 142.020 ;
        RECT 26.740 141.975 27.030 142.020 ;
        RECT 28.310 141.975 28.600 142.020 ;
        RECT 31.055 142.160 31.345 142.205 ;
        RECT 33.800 142.160 34.120 142.220 ;
        RECT 34.810 142.160 34.950 142.655 ;
        RECT 36.575 142.315 36.865 142.545 ;
        RECT 31.055 142.020 34.950 142.160 ;
        RECT 31.055 141.975 31.345 142.020 ;
        RECT 33.800 141.960 34.120 142.020 ;
        RECT 36.650 141.880 36.790 142.315 ;
        RECT 37.020 142.300 37.340 142.560 ;
        RECT 37.570 142.545 37.710 142.700 ;
        RECT 37.940 142.640 38.260 142.900 ;
        RECT 39.870 142.840 40.010 143.380 ;
        RECT 43.000 143.380 47.445 143.520 ;
        RECT 43.000 143.320 43.320 143.380 ;
        RECT 44.380 143.320 44.700 143.380 ;
        RECT 47.155 143.335 47.445 143.380 ;
        RECT 58.655 143.520 58.945 143.565 ;
        RECT 61.400 143.520 61.720 143.580 ;
        RECT 58.655 143.380 61.720 143.520 ;
        RECT 58.655 143.335 58.945 143.380 ;
        RECT 61.400 143.320 61.720 143.380 ;
        RECT 62.335 143.520 62.625 143.565 ;
        RECT 63.240 143.520 63.560 143.580 ;
        RECT 62.335 143.380 63.560 143.520 ;
        RECT 62.335 143.335 62.625 143.380 ;
        RECT 63.240 143.320 63.560 143.380 ;
        RECT 64.175 143.520 64.465 143.565 ;
        RECT 65.540 143.520 65.860 143.580 ;
        RECT 64.175 143.380 65.860 143.520 ;
        RECT 64.175 143.335 64.465 143.380 ;
        RECT 65.540 143.320 65.860 143.380 ;
        RECT 67.380 143.320 67.700 143.580 ;
        RECT 68.300 143.320 68.620 143.580 ;
        RECT 75.200 143.520 75.520 143.580 ;
        RECT 79.355 143.520 79.645 143.565 ;
        RECT 75.200 143.380 79.645 143.520 ;
        RECT 75.200 143.320 75.520 143.380 ;
        RECT 79.355 143.335 79.645 143.380 ;
        RECT 85.780 143.520 86.100 143.580 ;
        RECT 91.760 143.520 92.080 143.580 ;
        RECT 85.780 143.380 88.310 143.520 ;
        RECT 85.780 143.320 86.100 143.380 ;
        RECT 45.300 143.180 45.620 143.240 ;
        RECT 67.470 143.180 67.610 143.320 ;
        RECT 45.300 143.040 61.170 143.180 ;
        RECT 45.300 142.980 45.620 143.040 ;
        RECT 40.715 142.840 41.005 142.885 ;
        RECT 39.870 142.700 41.005 142.840 ;
        RECT 40.715 142.655 41.005 142.700 ;
        RECT 43.000 142.640 43.320 142.900 ;
        RECT 44.840 142.640 45.160 142.900 ;
        RECT 45.390 142.840 45.530 142.980 ;
        RECT 45.775 142.840 46.065 142.885 ;
        RECT 45.390 142.700 46.065 142.840 ;
        RECT 45.775 142.655 46.065 142.700 ;
        RECT 46.695 142.840 46.985 142.885 ;
        RECT 48.075 142.840 48.365 142.885 ;
        RECT 46.695 142.700 48.365 142.840 ;
        RECT 46.695 142.655 46.985 142.700 ;
        RECT 48.075 142.655 48.365 142.700 ;
        RECT 51.280 142.840 51.600 142.900 ;
        RECT 53.120 142.885 53.440 142.900 ;
        RECT 51.755 142.840 52.045 142.885 ;
        RECT 51.280 142.700 52.045 142.840 ;
        RECT 51.280 142.640 51.600 142.700 ;
        RECT 51.755 142.655 52.045 142.700 ;
        RECT 53.090 142.655 53.440 142.885 ;
        RECT 53.120 142.640 53.440 142.655 ;
        RECT 37.495 142.500 37.785 142.545 ;
        RECT 39.795 142.500 40.085 142.545 ;
        RECT 37.495 142.360 40.085 142.500 ;
        RECT 37.495 142.315 37.785 142.360 ;
        RECT 39.795 142.315 40.085 142.360 ;
        RECT 52.635 142.500 52.925 142.545 ;
        RECT 53.825 142.500 54.115 142.545 ;
        RECT 56.345 142.500 56.635 142.545 ;
        RECT 52.635 142.360 56.635 142.500 ;
        RECT 52.635 142.315 52.925 142.360 ;
        RECT 53.825 142.315 54.115 142.360 ;
        RECT 56.345 142.315 56.635 142.360 ;
        RECT 38.875 142.160 39.165 142.205 ;
        RECT 40.700 142.160 41.020 142.220 ;
        RECT 38.875 142.020 41.020 142.160 ;
        RECT 38.875 141.975 39.165 142.020 ;
        RECT 40.700 141.960 41.020 142.020 ;
        RECT 41.635 142.160 41.925 142.205 ;
        RECT 46.680 142.160 47.000 142.220 ;
        RECT 41.635 142.020 47.000 142.160 ;
        RECT 41.635 141.975 41.925 142.020 ;
        RECT 46.680 141.960 47.000 142.020 ;
        RECT 52.240 142.160 52.530 142.205 ;
        RECT 54.340 142.160 54.630 142.205 ;
        RECT 55.910 142.160 56.200 142.205 ;
        RECT 52.240 142.020 56.200 142.160 ;
        RECT 61.030 142.160 61.170 143.040 ;
        RECT 61.490 143.040 67.610 143.180 ;
        RECT 61.490 142.885 61.630 143.040 ;
        RECT 61.415 142.655 61.705 142.885 ;
        RECT 61.875 142.840 62.165 142.885 ;
        RECT 62.320 142.840 62.640 142.900 ;
        RECT 61.875 142.700 62.640 142.840 ;
        RECT 61.875 142.655 62.165 142.700 ;
        RECT 62.320 142.640 62.640 142.700 ;
        RECT 63.255 142.840 63.545 142.885 ;
        RECT 63.700 142.840 64.020 142.900 ;
        RECT 63.255 142.700 64.020 142.840 ;
        RECT 63.255 142.655 63.545 142.700 ;
        RECT 63.700 142.640 64.020 142.700 ;
        RECT 64.620 142.640 64.940 142.900 ;
        RECT 65.540 142.640 65.860 142.900 ;
        RECT 66.000 142.640 66.320 142.900 ;
        RECT 66.460 142.840 66.780 142.900 ;
        RECT 68.390 142.885 68.530 143.320 ;
        RECT 88.170 143.225 88.310 143.380 ;
        RECT 90.930 143.380 92.080 143.520 ;
        RECT 78.895 143.180 79.185 143.225 ;
        RECT 88.095 143.180 88.385 143.225 ;
        RECT 89.920 143.180 90.240 143.240 ;
        RECT 68.850 143.040 69.910 143.180 ;
        RECT 68.850 142.900 68.990 143.040 ;
        RECT 67.395 142.840 67.685 142.885 ;
        RECT 66.460 142.700 67.685 142.840 ;
        RECT 66.460 142.640 66.780 142.700 ;
        RECT 67.395 142.655 67.685 142.700 ;
        RECT 68.315 142.655 68.605 142.885 ;
        RECT 68.760 142.640 69.080 142.900 ;
        RECT 69.770 142.885 69.910 143.040 ;
        RECT 71.150 143.040 74.050 143.180 ;
        RECT 71.150 142.885 71.290 143.040 ;
        RECT 69.235 142.655 69.525 142.885 ;
        RECT 69.695 142.655 69.985 142.885 ;
        RECT 71.075 142.655 71.365 142.885 ;
        RECT 64.710 142.500 64.850 142.640 ;
        RECT 69.310 142.500 69.450 142.655 ;
        RECT 71.520 142.640 71.840 142.900 ;
        RECT 64.710 142.360 69.450 142.500 ;
        RECT 70.155 142.500 70.445 142.545 ;
        RECT 70.600 142.500 70.920 142.560 ;
        RECT 70.155 142.360 70.920 142.500 ;
        RECT 70.155 142.315 70.445 142.360 ;
        RECT 70.600 142.300 70.920 142.360 ;
        RECT 66.000 142.160 66.320 142.220 ;
        RECT 71.610 142.160 71.750 142.640 ;
        RECT 61.030 142.020 65.770 142.160 ;
        RECT 52.240 141.975 52.530 142.020 ;
        RECT 54.340 141.975 54.630 142.020 ;
        RECT 55.910 141.975 56.200 142.020 ;
        RECT 65.630 141.880 65.770 142.020 ;
        RECT 66.000 142.020 71.750 142.160 ;
        RECT 73.910 142.160 74.050 143.040 ;
        RECT 78.895 143.040 86.930 143.180 ;
        RECT 78.895 142.995 79.185 143.040 ;
        RECT 74.280 142.840 74.600 142.900 ;
        RECT 83.020 142.840 83.340 142.900 ;
        RECT 84.920 142.840 85.210 142.885 ;
        RECT 74.280 142.700 76.350 142.840 ;
        RECT 74.280 142.640 74.600 142.700 ;
        RECT 75.675 142.315 75.965 142.545 ;
        RECT 74.280 142.160 74.600 142.220 ;
        RECT 73.910 142.020 74.600 142.160 ;
        RECT 66.000 141.960 66.320 142.020 ;
        RECT 74.280 141.960 74.600 142.020 ;
        RECT 75.750 141.880 75.890 142.315 ;
        RECT 36.560 141.820 36.880 141.880 ;
        RECT 39.335 141.820 39.625 141.865 ;
        RECT 36.560 141.680 39.625 141.820 ;
        RECT 36.560 141.620 36.880 141.680 ;
        RECT 39.335 141.635 39.625 141.680 ;
        RECT 42.080 141.620 42.400 141.880 ;
        RECT 59.560 141.820 59.880 141.880 ;
        RECT 60.955 141.820 61.245 141.865 ;
        RECT 59.560 141.680 61.245 141.820 ;
        RECT 59.560 141.620 59.880 141.680 ;
        RECT 60.955 141.635 61.245 141.680 ;
        RECT 65.540 141.620 65.860 141.880 ;
        RECT 66.935 141.820 67.225 141.865 ;
        RECT 71.060 141.820 71.380 141.880 ;
        RECT 66.935 141.680 71.380 141.820 ;
        RECT 66.935 141.635 67.225 141.680 ;
        RECT 71.060 141.620 71.380 141.680 ;
        RECT 71.520 141.820 71.840 141.880 ;
        RECT 71.995 141.820 72.285 141.865 ;
        RECT 71.520 141.680 72.285 141.820 ;
        RECT 71.520 141.620 71.840 141.680 ;
        RECT 71.995 141.635 72.285 141.680 ;
        RECT 75.660 141.620 75.980 141.880 ;
        RECT 76.210 141.820 76.350 142.700 ;
        RECT 83.020 142.700 85.210 142.840 ;
        RECT 83.020 142.640 83.340 142.700 ;
        RECT 84.920 142.655 85.210 142.700 ;
        RECT 86.240 142.640 86.560 142.900 ;
        RECT 86.790 142.885 86.930 143.040 ;
        RECT 88.095 143.040 90.240 143.180 ;
        RECT 88.095 142.995 88.385 143.040 ;
        RECT 89.920 142.980 90.240 143.040 ;
        RECT 86.715 142.655 87.005 142.885 ;
        RECT 87.160 142.840 87.480 142.900 ;
        RECT 87.635 142.840 87.925 142.885 ;
        RECT 87.160 142.700 87.925 142.840 ;
        RECT 87.160 142.640 87.480 142.700 ;
        RECT 87.635 142.655 87.925 142.700 ;
        RECT 88.540 142.640 88.860 142.900 ;
        RECT 89.000 142.840 89.320 142.900 ;
        RECT 90.930 142.885 91.070 143.380 ;
        RECT 91.760 143.320 92.080 143.380 ;
        RECT 95.440 143.320 95.760 143.580 ;
        RECT 96.360 143.520 96.680 143.580 ;
        RECT 98.675 143.520 98.965 143.565 ;
        RECT 96.360 143.380 98.965 143.520 ;
        RECT 96.360 143.320 96.680 143.380 ;
        RECT 98.675 143.335 98.965 143.380 ;
        RECT 107.875 143.520 108.165 143.565 ;
        RECT 108.320 143.520 108.640 143.580 ;
        RECT 107.875 143.380 108.640 143.520 ;
        RECT 107.875 143.335 108.165 143.380 ;
        RECT 95.530 143.180 95.670 143.320 ;
        RECT 92.310 143.040 96.590 143.180 ;
        RECT 92.310 142.885 92.450 143.040 ;
        RECT 90.855 142.840 91.145 142.885 ;
        RECT 89.000 142.700 91.145 142.840 ;
        RECT 89.000 142.640 89.320 142.700 ;
        RECT 90.855 142.655 91.145 142.700 ;
        RECT 91.775 142.655 92.065 142.885 ;
        RECT 92.235 142.655 92.525 142.885 ;
        RECT 93.155 142.840 93.445 142.885 ;
        RECT 95.900 142.840 96.220 142.900 ;
        RECT 96.450 142.885 96.590 143.040 ;
        RECT 93.155 142.700 96.220 142.840 ;
        RECT 93.155 142.655 93.445 142.700 ;
        RECT 81.665 142.500 81.955 142.545 ;
        RECT 84.185 142.500 84.475 142.545 ;
        RECT 85.375 142.500 85.665 142.545 ;
        RECT 81.665 142.360 85.665 142.500 ;
        RECT 81.665 142.315 81.955 142.360 ;
        RECT 84.185 142.315 84.475 142.360 ;
        RECT 85.375 142.315 85.665 142.360 ;
        RECT 88.080 142.500 88.400 142.560 ;
        RECT 89.935 142.500 90.225 142.545 ;
        RECT 88.080 142.360 90.225 142.500 ;
        RECT 88.080 142.300 88.400 142.360 ;
        RECT 89.935 142.315 90.225 142.360 ;
        RECT 82.100 142.160 82.390 142.205 ;
        RECT 83.670 142.160 83.960 142.205 ;
        RECT 85.770 142.160 86.060 142.205 ;
        RECT 91.850 142.160 91.990 142.655 ;
        RECT 95.900 142.640 96.220 142.700 ;
        RECT 96.375 142.840 96.665 142.885 ;
        RECT 96.835 142.840 97.125 142.885 ;
        RECT 96.375 142.700 97.125 142.840 ;
        RECT 98.750 142.840 98.890 143.335 ;
        RECT 108.320 143.320 108.640 143.380 ;
        RECT 110.620 143.520 110.940 143.580 ;
        RECT 111.555 143.520 111.845 143.565 ;
        RECT 110.620 143.380 111.845 143.520 ;
        RECT 110.620 143.320 110.940 143.380 ;
        RECT 111.555 143.335 111.845 143.380 ;
        RECT 135.475 143.520 135.765 143.565 ;
        RECT 135.920 143.520 136.240 143.580 ;
        RECT 147.055 143.520 147.345 143.565 ;
        RECT 135.475 143.380 136.240 143.520 ;
        RECT 135.475 143.335 135.765 143.380 ;
        RECT 135.920 143.320 136.240 143.380 ;
        RECT 141.070 143.380 145.810 143.520 ;
        RECT 103.735 143.180 104.025 143.225 ;
        RECT 110.160 143.180 110.480 143.240 ;
        RECT 120.280 143.180 120.600 143.240 ;
        RECT 103.735 143.040 110.480 143.180 ;
        RECT 103.735 142.995 104.025 143.040 ;
        RECT 110.160 142.980 110.480 143.040 ;
        RECT 112.550 143.040 120.600 143.180 ;
        RECT 101.895 142.840 102.185 142.885 ;
        RECT 98.750 142.700 102.185 142.840 ;
        RECT 96.375 142.655 96.665 142.700 ;
        RECT 96.835 142.655 97.125 142.700 ;
        RECT 101.895 142.655 102.185 142.700 ;
        RECT 104.180 142.640 104.500 142.900 ;
        RECT 105.575 142.840 105.865 142.885 ;
        RECT 107.860 142.840 108.180 142.900 ;
        RECT 105.575 142.700 108.180 142.840 ;
        RECT 105.575 142.655 105.865 142.700 ;
        RECT 92.695 142.160 92.985 142.205 ;
        RECT 82.100 142.020 86.060 142.160 ;
        RECT 82.100 141.975 82.390 142.020 ;
        RECT 83.670 141.975 83.960 142.020 ;
        RECT 85.770 141.975 86.060 142.020 ;
        RECT 88.710 142.020 92.985 142.160 ;
        RECT 88.710 141.820 88.850 142.020 ;
        RECT 92.695 141.975 92.985 142.020 ;
        RECT 76.210 141.680 88.850 141.820 ;
        RECT 89.460 141.620 89.780 141.880 ;
        RECT 93.600 141.820 93.920 141.880 ;
        RECT 95.990 141.865 96.130 142.640 ;
        RECT 102.800 142.500 103.120 142.560 ;
        RECT 105.650 142.500 105.790 142.655 ;
        RECT 107.860 142.640 108.180 142.700 ;
        RECT 108.780 142.640 109.100 142.900 ;
        RECT 112.550 142.885 112.690 143.040 ;
        RECT 120.280 142.980 120.600 143.040 ;
        RECT 137.760 143.180 138.080 143.240 ;
        RECT 141.070 143.225 141.210 143.380 ;
        RECT 140.995 143.180 141.285 143.225 ;
        RECT 137.760 143.040 141.285 143.180 ;
        RECT 137.760 142.980 138.080 143.040 ;
        RECT 140.995 142.995 141.285 143.040 ;
        RECT 141.440 143.180 141.760 143.240 ;
        RECT 141.995 143.180 142.285 143.225 ;
        RECT 141.440 143.040 142.285 143.180 ;
        RECT 141.440 142.980 141.760 143.040 ;
        RECT 141.995 142.995 142.285 143.040 ;
        RECT 143.755 143.180 144.045 143.225 ;
        RECT 144.200 143.180 144.520 143.240 ;
        RECT 143.755 143.040 144.520 143.180 ;
        RECT 143.755 142.995 144.045 143.040 ;
        RECT 112.475 142.840 112.765 142.885 ;
        RECT 109.330 142.700 112.765 142.840 ;
        RECT 102.800 142.360 105.790 142.500 ;
        RECT 102.800 142.300 103.120 142.360 ;
        RECT 96.360 142.160 96.680 142.220 ;
        RECT 109.330 142.160 109.470 142.700 ;
        RECT 112.475 142.655 112.765 142.700 ;
        RECT 113.380 142.640 113.700 142.900 ;
        RECT 115.220 142.640 115.540 142.900 ;
        RECT 118.915 142.840 119.205 142.885 ;
        RECT 122.120 142.840 122.440 142.900 ;
        RECT 124.420 142.840 124.740 142.900 ;
        RECT 127.195 142.840 127.485 142.885 ;
        RECT 131.795 142.840 132.085 142.885 ;
        RECT 118.915 142.700 127.485 142.840 ;
        RECT 118.915 142.655 119.205 142.700 ;
        RECT 109.700 142.500 110.020 142.560 ;
        RECT 111.540 142.500 111.860 142.560 ;
        RECT 118.990 142.500 119.130 142.655 ;
        RECT 122.120 142.640 122.440 142.700 ;
        RECT 124.420 142.640 124.740 142.700 ;
        RECT 127.195 142.655 127.485 142.700 ;
        RECT 130.260 142.700 132.085 142.840 ;
        RECT 109.700 142.360 119.130 142.500 ;
        RECT 109.700 142.300 110.020 142.360 ;
        RECT 111.540 142.300 111.860 142.360 ;
        RECT 119.835 142.315 120.125 142.545 ;
        RECT 126.275 142.500 126.565 142.545 ;
        RECT 129.020 142.500 129.340 142.560 ;
        RECT 130.260 142.500 130.400 142.700 ;
        RECT 131.795 142.655 132.085 142.700 ;
        RECT 132.240 142.640 132.560 142.900 ;
        RECT 133.620 142.640 133.940 142.900 ;
        RECT 135.935 142.840 136.225 142.885 ;
        RECT 139.615 142.840 139.905 142.885 ;
        RECT 135.935 142.700 139.905 142.840 ;
        RECT 135.935 142.655 136.225 142.700 ;
        RECT 139.615 142.655 139.905 142.700 ;
        RECT 140.535 142.840 140.825 142.885 ;
        RECT 143.280 142.840 143.600 142.900 ;
        RECT 143.830 142.840 143.970 142.995 ;
        RECT 144.200 142.980 144.520 143.040 ;
        RECT 144.675 143.180 144.965 143.225 ;
        RECT 145.120 143.180 145.440 143.240 ;
        RECT 144.675 143.040 145.440 143.180 ;
        RECT 145.670 143.180 145.810 143.380 ;
        RECT 146.590 143.380 147.345 143.520 ;
        RECT 146.040 143.180 146.360 143.240 ;
        RECT 145.670 143.040 146.360 143.180 ;
        RECT 144.675 142.995 144.965 143.040 ;
        RECT 140.535 142.700 143.970 142.840 ;
        RECT 140.535 142.655 140.825 142.700 ;
        RECT 126.275 142.360 130.400 142.500 ;
        RECT 139.690 142.500 139.830 142.655 ;
        RECT 143.280 142.640 143.600 142.700 ;
        RECT 142.360 142.500 142.680 142.560 ;
        RECT 144.750 142.500 144.890 142.995 ;
        RECT 145.120 142.980 145.440 143.040 ;
        RECT 146.040 142.980 146.360 143.040 ;
        RECT 145.595 142.840 145.885 142.885 ;
        RECT 146.590 142.840 146.730 143.380 ;
        RECT 147.055 143.335 147.345 143.380 ;
        RECT 147.895 143.335 148.185 143.565 ;
        RECT 149.275 143.520 149.565 143.565 ;
        RECT 149.720 143.520 150.040 143.580 ;
        RECT 149.275 143.380 150.040 143.520 ;
        RECT 149.275 143.335 149.565 143.380 ;
        RECT 145.595 142.700 146.730 142.840 ;
        RECT 147.970 142.840 148.110 143.335 ;
        RECT 149.720 143.320 150.040 143.380 ;
        RECT 148.355 142.840 148.645 142.885 ;
        RECT 147.970 142.700 148.645 142.840 ;
        RECT 145.595 142.655 145.885 142.700 ;
        RECT 148.355 142.655 148.645 142.700 ;
        RECT 139.690 142.360 144.890 142.500 ;
        RECT 126.275 142.315 126.565 142.360 ;
        RECT 96.360 142.020 109.470 142.160 ;
        RECT 110.160 142.160 110.480 142.220 ;
        RECT 119.360 142.160 119.680 142.220 ;
        RECT 110.160 142.020 119.680 142.160 ;
        RECT 119.910 142.160 120.050 142.315 ;
        RECT 129.020 142.300 129.340 142.360 ;
        RECT 142.360 142.300 142.680 142.360 ;
        RECT 121.200 142.160 121.520 142.220 ;
        RECT 144.200 142.160 144.520 142.220 ;
        RECT 119.910 142.020 133.390 142.160 ;
        RECT 96.360 141.960 96.680 142.020 ;
        RECT 110.160 141.960 110.480 142.020 ;
        RECT 119.360 141.960 119.680 142.020 ;
        RECT 121.200 141.960 121.520 142.020 ;
        RECT 94.075 141.820 94.365 141.865 ;
        RECT 93.600 141.680 94.365 141.820 ;
        RECT 93.600 141.620 93.920 141.680 ;
        RECT 94.075 141.635 94.365 141.680 ;
        RECT 95.915 141.820 96.205 141.865 ;
        RECT 98.675 141.820 98.965 141.865 ;
        RECT 95.915 141.680 98.965 141.820 ;
        RECT 95.915 141.635 96.205 141.680 ;
        RECT 98.675 141.635 98.965 141.680 ;
        RECT 99.580 141.620 99.900 141.880 ;
        RECT 101.420 141.820 101.740 141.880 ;
        RECT 106.035 141.820 106.325 141.865 ;
        RECT 112.000 141.820 112.320 141.880 ;
        RECT 101.420 141.680 112.320 141.820 ;
        RECT 101.420 141.620 101.740 141.680 ;
        RECT 106.035 141.635 106.325 141.680 ;
        RECT 112.000 141.620 112.320 141.680 ;
        RECT 116.140 141.620 116.460 141.880 ;
        RECT 117.980 141.620 118.300 141.880 ;
        RECT 128.100 141.620 128.420 141.880 ;
        RECT 130.875 141.820 131.165 141.865 ;
        RECT 132.700 141.820 133.020 141.880 ;
        RECT 133.250 141.865 133.390 142.020 ;
        RECT 140.150 142.020 147.190 142.160 ;
        RECT 130.875 141.680 133.020 141.820 ;
        RECT 130.875 141.635 131.165 141.680 ;
        RECT 132.700 141.620 133.020 141.680 ;
        RECT 133.175 141.820 133.465 141.865 ;
        RECT 136.380 141.820 136.700 141.880 ;
        RECT 133.175 141.680 136.700 141.820 ;
        RECT 133.175 141.635 133.465 141.680 ;
        RECT 136.380 141.620 136.700 141.680 ;
        RECT 138.680 141.820 139.000 141.880 ;
        RECT 140.150 141.865 140.290 142.020 ;
        RECT 144.200 141.960 144.520 142.020 ;
        RECT 140.075 141.820 140.365 141.865 ;
        RECT 138.680 141.680 140.365 141.820 ;
        RECT 138.680 141.620 139.000 141.680 ;
        RECT 140.075 141.635 140.365 141.680 ;
        RECT 141.900 141.620 142.220 141.880 ;
        RECT 142.835 141.820 143.125 141.865 ;
        RECT 145.580 141.820 145.900 141.880 ;
        RECT 147.050 141.865 147.190 142.020 ;
        RECT 142.835 141.680 145.900 141.820 ;
        RECT 142.835 141.635 143.125 141.680 ;
        RECT 145.580 141.620 145.900 141.680 ;
        RECT 146.975 141.635 147.265 141.865 ;
        RECT 22.690 141.000 157.010 141.480 ;
        RECT 26.900 140.600 27.220 140.860 ;
        RECT 28.740 140.600 29.060 140.860 ;
        RECT 33.800 140.600 34.120 140.860 ;
        RECT 40.700 140.600 41.020 140.860 ;
        RECT 41.160 140.800 41.480 140.860 ;
        RECT 41.635 140.800 41.925 140.845 ;
        RECT 41.160 140.660 41.925 140.800 ;
        RECT 41.160 140.600 41.480 140.660 ;
        RECT 41.635 140.615 41.925 140.660 ;
        RECT 42.555 140.800 42.845 140.845 ;
        RECT 43.000 140.800 43.320 140.860 ;
        RECT 42.555 140.660 43.320 140.800 ;
        RECT 42.555 140.615 42.845 140.660 ;
        RECT 43.000 140.600 43.320 140.660 ;
        RECT 49.915 140.800 50.205 140.845 ;
        RECT 50.835 140.800 51.125 140.845 ;
        RECT 49.915 140.660 51.125 140.800 ;
        RECT 49.915 140.615 50.205 140.660 ;
        RECT 50.835 140.615 51.125 140.660 ;
        RECT 53.120 140.800 53.440 140.860 ;
        RECT 54.055 140.800 54.345 140.845 ;
        RECT 65.080 140.800 65.400 140.860 ;
        RECT 53.120 140.660 54.345 140.800 ;
        RECT 53.120 140.600 53.440 140.660 ;
        RECT 54.055 140.615 54.345 140.660 ;
        RECT 61.950 140.660 65.400 140.800 ;
        RECT 28.830 140.120 28.970 140.600 ;
        RECT 32.895 140.460 33.185 140.505 ;
        RECT 34.720 140.460 35.040 140.520 ;
        RECT 39.795 140.460 40.085 140.505 ;
        RECT 32.895 140.320 40.085 140.460 ;
        RECT 32.895 140.275 33.185 140.320 ;
        RECT 34.720 140.260 35.040 140.320 ;
        RECT 39.795 140.275 40.085 140.320 ;
        RECT 29.215 140.120 29.505 140.165 ;
        RECT 28.830 139.980 29.505 140.120 ;
        RECT 29.215 139.935 29.505 139.980 ;
        RECT 29.660 140.120 29.980 140.180 ;
        RECT 32.420 140.120 32.740 140.180 ;
        RECT 29.660 139.980 32.740 140.120 ;
        RECT 29.660 139.920 29.980 139.980 ;
        RECT 32.420 139.920 32.740 139.980 ;
        RECT 27.835 139.780 28.125 139.825 ;
        RECT 28.280 139.780 28.600 139.840 ;
        RECT 27.835 139.640 28.600 139.780 ;
        RECT 27.835 139.595 28.125 139.640 ;
        RECT 28.280 139.580 28.600 139.640 ;
        RECT 28.755 139.780 29.045 139.825 ;
        RECT 29.750 139.780 29.890 139.920 ;
        RECT 37.480 139.780 37.800 139.840 ;
        RECT 38.875 139.780 39.165 139.825 ;
        RECT 28.755 139.640 29.890 139.780 ;
        RECT 32.050 139.640 39.165 139.780 ;
        RECT 28.755 139.595 29.045 139.640 ;
        RECT 32.050 139.160 32.190 139.640 ;
        RECT 37.480 139.580 37.800 139.640 ;
        RECT 38.875 139.595 39.165 139.640 ;
        RECT 34.735 139.440 35.025 139.485 ;
        RECT 36.560 139.440 36.880 139.500 ;
        RECT 34.735 139.300 36.880 139.440 ;
        RECT 40.790 139.440 40.930 140.600 ;
        RECT 43.500 140.460 43.790 140.505 ;
        RECT 45.600 140.460 45.890 140.505 ;
        RECT 47.170 140.460 47.460 140.505 ;
        RECT 61.950 140.460 62.090 140.660 ;
        RECT 65.080 140.600 65.400 140.660 ;
        RECT 65.540 140.800 65.860 140.860 ;
        RECT 68.300 140.800 68.620 140.860 ;
        RECT 65.540 140.660 68.620 140.800 ;
        RECT 65.540 140.600 65.860 140.660 ;
        RECT 68.300 140.600 68.620 140.660 ;
        RECT 72.900 140.800 73.220 140.860 ;
        RECT 74.740 140.800 75.060 140.860 ;
        RECT 89.935 140.800 90.225 140.845 ;
        RECT 90.840 140.800 91.160 140.860 ;
        RECT 72.900 140.660 89.690 140.800 ;
        RECT 72.900 140.600 73.220 140.660 ;
        RECT 74.740 140.600 75.060 140.660 ;
        RECT 43.500 140.320 47.460 140.460 ;
        RECT 43.500 140.275 43.790 140.320 ;
        RECT 45.600 140.275 45.890 140.320 ;
        RECT 47.170 140.275 47.460 140.320 ;
        RECT 52.750 140.320 62.090 140.460 ;
        RECT 62.360 140.460 62.650 140.505 ;
        RECT 64.460 140.460 64.750 140.505 ;
        RECT 66.030 140.460 66.320 140.505 ;
        RECT 62.360 140.320 66.320 140.460 ;
        RECT 43.895 140.120 44.185 140.165 ;
        RECT 45.085 140.120 45.375 140.165 ;
        RECT 47.605 140.120 47.895 140.165 ;
        RECT 51.280 140.120 51.600 140.180 ;
        RECT 52.750 140.165 52.890 140.320 ;
        RECT 62.360 140.275 62.650 140.320 ;
        RECT 64.460 140.275 64.750 140.320 ;
        RECT 66.030 140.275 66.320 140.320 ;
        RECT 68.775 140.460 69.065 140.505 ;
        RECT 73.835 140.460 74.125 140.505 ;
        RECT 68.775 140.320 70.370 140.460 ;
        RECT 68.775 140.275 69.065 140.320 ;
        RECT 43.895 139.980 47.895 140.120 ;
        RECT 43.895 139.935 44.185 139.980 ;
        RECT 45.085 139.935 45.375 139.980 ;
        RECT 47.605 139.935 47.895 139.980 ;
        RECT 49.990 139.980 51.600 140.120 ;
        RECT 43.015 139.780 43.305 139.825 ;
        RECT 49.990 139.780 50.130 139.980 ;
        RECT 51.280 139.920 51.600 139.980 ;
        RECT 52.675 139.935 52.965 140.165 ;
        RECT 59.560 140.120 59.880 140.180 ;
        RECT 62.755 140.120 63.045 140.165 ;
        RECT 63.945 140.120 64.235 140.165 ;
        RECT 66.465 140.120 66.755 140.165 ;
        RECT 59.560 139.980 60.710 140.120 ;
        RECT 59.560 139.920 59.880 139.980 ;
        RECT 43.015 139.640 50.130 139.780 ;
        RECT 43.015 139.595 43.305 139.640 ;
        RECT 50.360 139.580 50.680 139.840 ;
        RECT 54.960 139.580 55.280 139.840 ;
        RECT 58.655 139.780 58.945 139.825 ;
        RECT 60.020 139.780 60.340 139.840 ;
        RECT 60.570 139.825 60.710 139.980 ;
        RECT 62.755 139.980 66.755 140.120 ;
        RECT 62.755 139.935 63.045 139.980 ;
        RECT 63.945 139.935 64.235 139.980 ;
        RECT 66.465 139.935 66.755 139.980 ;
        RECT 70.230 139.840 70.370 140.320 ;
        RECT 71.150 140.320 74.125 140.460 ;
        RECT 71.150 140.180 71.290 140.320 ;
        RECT 73.835 140.275 74.125 140.320 ;
        RECT 79.815 140.275 80.105 140.505 ;
        RECT 82.560 140.460 82.850 140.505 ;
        RECT 84.130 140.460 84.420 140.505 ;
        RECT 86.230 140.460 86.520 140.505 ;
        RECT 82.560 140.320 86.520 140.460 ;
        RECT 89.550 140.460 89.690 140.660 ;
        RECT 89.935 140.660 91.160 140.800 ;
        RECT 89.935 140.615 90.225 140.660 ;
        RECT 90.840 140.600 91.160 140.660 ;
        RECT 94.980 140.800 95.300 140.860 ;
        RECT 101.420 140.800 101.740 140.860 ;
        RECT 106.495 140.800 106.785 140.845 ;
        RECT 94.980 140.660 101.740 140.800 ;
        RECT 94.980 140.600 95.300 140.660 ;
        RECT 101.420 140.600 101.740 140.660 ;
        RECT 101.970 140.660 106.785 140.800 ;
        RECT 101.970 140.460 102.110 140.660 ;
        RECT 106.495 140.615 106.785 140.660 ;
        RECT 107.415 140.800 107.705 140.845 ;
        RECT 108.780 140.800 109.100 140.860 ;
        RECT 107.415 140.660 109.100 140.800 ;
        RECT 107.415 140.615 107.705 140.660 ;
        RECT 89.550 140.320 102.110 140.460 ;
        RECT 102.340 140.460 102.660 140.520 ;
        RECT 106.570 140.460 106.710 140.615 ;
        RECT 108.780 140.600 109.100 140.660 ;
        RECT 110.710 140.660 119.590 140.800 ;
        RECT 109.700 140.460 110.020 140.520 ;
        RECT 102.340 140.320 104.870 140.460 ;
        RECT 106.570 140.320 110.020 140.460 ;
        RECT 82.560 140.275 82.850 140.320 ;
        RECT 84.130 140.275 84.420 140.320 ;
        RECT 86.230 140.275 86.520 140.320 ;
        RECT 71.060 139.920 71.380 140.180 ;
        RECT 71.520 139.920 71.840 140.180 ;
        RECT 76.135 140.120 76.425 140.165 ;
        RECT 74.370 139.980 76.425 140.120 ;
        RECT 57.350 139.640 60.340 139.780 ;
        RECT 44.380 139.485 44.700 139.500 ;
        RECT 41.635 139.440 41.925 139.485 ;
        RECT 44.350 139.440 44.700 139.485 ;
        RECT 40.790 139.300 41.925 139.440 ;
        RECT 44.185 139.300 44.700 139.440 ;
        RECT 34.735 139.255 35.025 139.300 ;
        RECT 36.560 139.240 36.880 139.300 ;
        RECT 41.635 139.255 41.925 139.300 ;
        RECT 44.350 139.255 44.700 139.300 ;
        RECT 44.380 139.240 44.700 139.255 ;
        RECT 54.500 139.440 54.820 139.500 ;
        RECT 57.350 139.440 57.490 139.640 ;
        RECT 58.655 139.595 58.945 139.640 ;
        RECT 60.020 139.580 60.340 139.640 ;
        RECT 60.495 139.595 60.785 139.825 ;
        RECT 60.955 139.780 61.245 139.825 ;
        RECT 61.875 139.780 62.165 139.825 ;
        RECT 69.680 139.780 70.000 139.840 ;
        RECT 60.955 139.640 61.630 139.780 ;
        RECT 60.955 139.595 61.245 139.640 ;
        RECT 61.490 139.500 61.630 139.640 ;
        RECT 61.875 139.640 70.000 139.780 ;
        RECT 61.875 139.595 62.165 139.640 ;
        RECT 69.680 139.580 70.000 139.640 ;
        RECT 70.140 139.580 70.460 139.840 ;
        RECT 71.980 139.825 72.300 139.840 ;
        RECT 71.975 139.780 72.300 139.825 ;
        RECT 71.785 139.640 72.300 139.780 ;
        RECT 71.975 139.595 72.300 139.640 ;
        RECT 71.980 139.580 72.300 139.595 ;
        RECT 72.440 139.780 72.760 139.840 ;
        RECT 74.370 139.825 74.510 139.980 ;
        RECT 76.135 139.935 76.425 139.980 ;
        RECT 72.915 139.780 73.205 139.825 ;
        RECT 72.440 139.640 73.205 139.780 ;
        RECT 72.440 139.580 72.760 139.640 ;
        RECT 72.915 139.595 73.205 139.640 ;
        RECT 74.295 139.780 74.585 139.825 ;
        RECT 74.740 139.780 75.060 139.840 ;
        RECT 74.295 139.640 75.060 139.780 ;
        RECT 74.295 139.595 74.585 139.640 ;
        RECT 74.740 139.580 75.060 139.640 ;
        RECT 75.660 139.780 75.980 139.840 ;
        RECT 79.890 139.780 80.030 140.275 ;
        RECT 102.340 140.260 102.660 140.320 ;
        RECT 82.125 140.120 82.415 140.165 ;
        RECT 84.645 140.120 84.935 140.165 ;
        RECT 85.835 140.120 86.125 140.165 ;
        RECT 82.125 139.980 86.125 140.120 ;
        RECT 82.125 139.935 82.415 139.980 ;
        RECT 84.645 139.935 84.935 139.980 ;
        RECT 85.835 139.935 86.125 139.980 ;
        RECT 89.460 139.920 89.780 140.180 ;
        RECT 89.920 140.120 90.240 140.180 ;
        RECT 94.980 140.120 95.300 140.180 ;
        RECT 104.730 140.120 104.870 140.320 ;
        RECT 109.700 140.260 110.020 140.320 ;
        RECT 110.160 140.120 110.480 140.180 ;
        RECT 89.920 139.980 95.300 140.120 ;
        RECT 89.920 139.920 90.240 139.980 ;
        RECT 94.980 139.920 95.300 139.980 ;
        RECT 101.510 139.980 104.410 140.120 ;
        RECT 104.730 139.980 110.480 140.120 ;
        RECT 86.715 139.780 87.005 139.825 ;
        RECT 89.550 139.780 89.690 139.920 ;
        RECT 75.660 139.640 80.030 139.780 ;
        RECT 82.190 139.640 87.005 139.780 ;
        RECT 75.660 139.580 75.980 139.640 ;
        RECT 82.190 139.500 82.330 139.640 ;
        RECT 86.715 139.595 87.005 139.640 ;
        RECT 87.250 139.640 89.690 139.780 ;
        RECT 90.855 139.780 91.145 139.825 ;
        RECT 91.300 139.780 91.620 139.840 ;
        RECT 101.510 139.825 101.650 139.980 ;
        RECT 101.435 139.780 101.725 139.825 ;
        RECT 90.855 139.640 91.620 139.780 ;
        RECT 54.500 139.300 57.490 139.440 ;
        RECT 57.720 139.440 58.040 139.500 ;
        RECT 57.720 139.300 60.710 139.440 ;
        RECT 54.500 139.240 54.820 139.300 ;
        RECT 57.720 139.240 58.040 139.300 ;
        RECT 31.960 138.900 32.280 139.160 ;
        RECT 32.420 139.100 32.740 139.160 ;
        RECT 33.685 139.100 33.975 139.145 ;
        RECT 32.420 138.960 33.975 139.100 ;
        RECT 32.420 138.900 32.740 138.960 ;
        RECT 33.685 138.915 33.975 138.960 ;
        RECT 36.100 138.900 36.420 139.160 ;
        RECT 60.020 138.900 60.340 139.160 ;
        RECT 60.570 139.100 60.710 139.300 ;
        RECT 61.400 139.240 61.720 139.500 ;
        RECT 63.210 139.440 63.500 139.485 ;
        RECT 65.080 139.440 65.400 139.500 ;
        RECT 63.210 139.300 65.400 139.440 ;
        RECT 63.210 139.255 63.500 139.300 ;
        RECT 65.080 139.240 65.400 139.300 ;
        RECT 82.100 139.240 82.420 139.500 ;
        RECT 85.490 139.440 85.780 139.485 ;
        RECT 87.250 139.440 87.390 139.640 ;
        RECT 90.855 139.595 91.145 139.640 ;
        RECT 91.300 139.580 91.620 139.640 ;
        RECT 93.690 139.640 101.725 139.780 ;
        RECT 93.690 139.500 93.830 139.640 ;
        RECT 101.435 139.595 101.725 139.640 ;
        RECT 102.815 139.780 103.105 139.825 ;
        RECT 103.260 139.780 103.580 139.840 ;
        RECT 102.815 139.640 103.580 139.780 ;
        RECT 102.815 139.595 103.105 139.640 ;
        RECT 103.260 139.580 103.580 139.640 ;
        RECT 103.720 139.580 104.040 139.840 ;
        RECT 104.270 139.825 104.410 139.980 ;
        RECT 110.160 139.920 110.480 139.980 ;
        RECT 104.195 139.595 104.485 139.825 ;
        RECT 104.640 139.580 104.960 139.840 ;
        RECT 105.560 139.780 105.880 139.840 ;
        RECT 110.710 139.780 110.850 140.660 ;
        RECT 114.800 140.460 115.090 140.505 ;
        RECT 116.900 140.460 117.190 140.505 ;
        RECT 118.470 140.460 118.760 140.505 ;
        RECT 114.800 140.320 118.760 140.460 ;
        RECT 114.800 140.275 115.090 140.320 ;
        RECT 116.900 140.275 117.190 140.320 ;
        RECT 118.470 140.275 118.760 140.320 ;
        RECT 115.195 140.120 115.485 140.165 ;
        RECT 116.385 140.120 116.675 140.165 ;
        RECT 118.905 140.120 119.195 140.165 ;
        RECT 115.195 139.980 119.195 140.120 ;
        RECT 119.450 140.120 119.590 140.660 ;
        RECT 121.200 140.600 121.520 140.860 ;
        RECT 129.020 140.600 129.340 140.860 ;
        RECT 141.900 140.800 142.220 140.860 ;
        RECT 145.595 140.800 145.885 140.845 ;
        RECT 141.900 140.660 147.190 140.800 ;
        RECT 141.900 140.600 142.220 140.660 ;
        RECT 145.595 140.615 145.885 140.660 ;
        RECT 122.620 140.460 122.910 140.505 ;
        RECT 124.720 140.460 125.010 140.505 ;
        RECT 126.290 140.460 126.580 140.505 ;
        RECT 122.620 140.320 126.580 140.460 ;
        RECT 122.620 140.275 122.910 140.320 ;
        RECT 124.720 140.275 125.010 140.320 ;
        RECT 126.290 140.275 126.580 140.320 ;
        RECT 123.015 140.120 123.305 140.165 ;
        RECT 124.205 140.120 124.495 140.165 ;
        RECT 126.725 140.120 127.015 140.165 ;
        RECT 119.450 139.980 122.810 140.120 ;
        RECT 115.195 139.935 115.485 139.980 ;
        RECT 116.385 139.935 116.675 139.980 ;
        RECT 118.905 139.935 119.195 139.980 ;
        RECT 105.560 139.640 110.850 139.780 ;
        RECT 114.300 139.780 114.620 139.840 ;
        RECT 117.060 139.780 117.380 139.840 ;
        RECT 122.135 139.780 122.425 139.825 ;
        RECT 114.300 139.640 122.425 139.780 ;
        RECT 122.670 139.780 122.810 139.980 ;
        RECT 123.015 139.980 127.015 140.120 ;
        RECT 123.015 139.935 123.305 139.980 ;
        RECT 124.205 139.935 124.495 139.980 ;
        RECT 126.725 139.935 127.015 139.980 ;
        RECT 129.110 139.780 129.250 140.600 ;
        RECT 132.240 140.260 132.560 140.520 ;
        RECT 133.620 140.460 133.940 140.520 ;
        RECT 139.600 140.460 139.920 140.520 ;
        RECT 133.620 140.320 139.920 140.460 ;
        RECT 133.620 140.260 133.940 140.320 ;
        RECT 132.330 140.120 132.470 140.260 ;
        RECT 137.390 140.165 137.530 140.320 ;
        RECT 139.600 140.260 139.920 140.320 ;
        RECT 132.330 139.980 133.390 140.120 ;
        RECT 133.250 139.825 133.390 139.980 ;
        RECT 134.630 139.980 136.150 140.120 ;
        RECT 132.485 139.780 132.775 139.825 ;
        RECT 122.670 139.640 126.950 139.780 ;
        RECT 129.110 139.640 132.775 139.780 ;
        RECT 105.560 139.580 105.880 139.640 ;
        RECT 114.300 139.580 114.620 139.640 ;
        RECT 117.060 139.580 117.380 139.640 ;
        RECT 122.135 139.595 122.425 139.640 ;
        RECT 85.490 139.300 87.390 139.440 ;
        RECT 85.490 139.255 85.780 139.300 ;
        RECT 87.620 139.240 87.940 139.500 ;
        RECT 88.555 139.440 88.845 139.485 ;
        RECT 89.000 139.440 89.320 139.500 ;
        RECT 88.555 139.300 89.320 139.440 ;
        RECT 88.555 139.255 88.845 139.300 ;
        RECT 89.000 139.240 89.320 139.300 ;
        RECT 89.475 139.440 89.765 139.485 ;
        RECT 93.600 139.440 93.920 139.500 ;
        RECT 89.475 139.300 93.920 139.440 ;
        RECT 89.475 139.255 89.765 139.300 ;
        RECT 93.600 139.240 93.920 139.300 ;
        RECT 100.500 139.240 100.820 139.500 ;
        RECT 104.730 139.440 104.870 139.580 ;
        RECT 109.715 139.440 110.005 139.485 ;
        RECT 114.760 139.440 115.080 139.500 ;
        RECT 104.730 139.300 115.080 139.440 ;
        RECT 109.715 139.255 110.005 139.300 ;
        RECT 114.760 139.240 115.080 139.300 ;
        RECT 115.650 139.440 115.940 139.485 ;
        RECT 116.140 139.440 116.460 139.500 ;
        RECT 115.650 139.300 116.460 139.440 ;
        RECT 115.650 139.255 115.940 139.300 ;
        RECT 116.140 139.240 116.460 139.300 ;
        RECT 121.660 139.440 121.980 139.500 ;
        RECT 123.360 139.440 123.650 139.485 ;
        RECT 121.660 139.300 123.650 139.440 ;
        RECT 121.660 139.240 121.980 139.300 ;
        RECT 123.360 139.255 123.650 139.300 ;
        RECT 126.810 139.160 126.950 139.640 ;
        RECT 132.485 139.595 132.775 139.640 ;
        RECT 133.175 139.595 133.465 139.825 ;
        RECT 133.635 139.780 133.925 139.825 ;
        RECT 134.080 139.780 134.400 139.840 ;
        RECT 134.630 139.825 134.770 139.980 ;
        RECT 136.010 139.840 136.150 139.980 ;
        RECT 137.315 139.935 137.605 140.165 ;
        RECT 144.200 140.120 144.520 140.180 ;
        RECT 143.830 139.980 144.520 140.120 ;
        RECT 133.635 139.640 134.400 139.780 ;
        RECT 133.635 139.595 133.925 139.640 ;
        RECT 69.235 139.100 69.525 139.145 ;
        RECT 60.570 138.960 69.525 139.100 ;
        RECT 69.235 138.915 69.525 138.960 ;
        RECT 70.600 139.100 70.920 139.160 ;
        RECT 75.215 139.100 75.505 139.145 ;
        RECT 70.600 138.960 75.505 139.100 ;
        RECT 70.600 138.900 70.920 138.960 ;
        RECT 75.215 138.915 75.505 138.960 ;
        RECT 79.340 138.900 79.660 139.160 ;
        RECT 94.060 138.900 94.380 139.160 ;
        RECT 101.420 138.900 101.740 139.160 ;
        RECT 104.640 138.900 104.960 139.160 ;
        RECT 109.240 138.900 109.560 139.160 ;
        RECT 126.720 138.900 127.040 139.160 ;
        RECT 131.780 138.900 132.100 139.160 ;
        RECT 133.250 139.100 133.390 139.595 ;
        RECT 134.080 139.580 134.400 139.640 ;
        RECT 134.550 139.595 134.840 139.825 ;
        RECT 135.015 139.780 135.305 139.825 ;
        RECT 135.015 139.640 135.690 139.780 ;
        RECT 135.015 139.595 135.305 139.640 ;
        RECT 135.550 139.160 135.690 139.640 ;
        RECT 135.920 139.580 136.240 139.840 ;
        RECT 136.380 139.580 136.700 139.840 ;
        RECT 143.830 139.825 143.970 139.980 ;
        RECT 144.200 139.920 144.520 139.980 ;
        RECT 144.750 139.980 146.730 140.120 ;
        RECT 140.075 139.780 140.365 139.825 ;
        RECT 140.075 139.640 143.510 139.780 ;
        RECT 140.075 139.595 140.365 139.640 ;
        RECT 143.370 139.485 143.510 139.640 ;
        RECT 143.755 139.595 144.045 139.825 ;
        RECT 144.750 139.780 144.890 139.980 ;
        RECT 146.590 139.840 146.730 139.980 ;
        RECT 144.290 139.640 144.890 139.780 ;
        RECT 145.120 139.780 145.440 139.840 ;
        RECT 146.055 139.780 146.345 139.825 ;
        RECT 145.120 139.640 146.345 139.780 ;
        RECT 143.295 139.440 143.585 139.485 ;
        RECT 144.290 139.440 144.430 139.640 ;
        RECT 145.120 139.580 145.440 139.640 ;
        RECT 146.055 139.595 146.345 139.640 ;
        RECT 146.500 139.580 146.820 139.840 ;
        RECT 147.050 139.825 147.190 140.660 ;
        RECT 147.920 140.460 148.210 140.505 ;
        RECT 150.020 140.460 150.310 140.505 ;
        RECT 151.590 140.460 151.880 140.505 ;
        RECT 147.920 140.320 151.880 140.460 ;
        RECT 147.920 140.275 148.210 140.320 ;
        RECT 150.020 140.275 150.310 140.320 ;
        RECT 151.590 140.275 151.880 140.320 ;
        RECT 147.420 139.920 147.740 140.180 ;
        RECT 148.315 140.120 148.605 140.165 ;
        RECT 149.505 140.120 149.795 140.165 ;
        RECT 152.025 140.120 152.315 140.165 ;
        RECT 148.315 139.980 152.315 140.120 ;
        RECT 148.315 139.935 148.605 139.980 ;
        RECT 149.505 139.935 149.795 139.980 ;
        RECT 152.025 139.935 152.315 139.980 ;
        RECT 146.975 139.595 147.265 139.825 ;
        RECT 143.295 139.300 144.430 139.440 ;
        RECT 143.295 139.255 143.585 139.300 ;
        RECT 144.660 139.240 144.980 139.500 ;
        RECT 148.800 139.485 149.120 139.500 ;
        RECT 145.210 139.300 146.730 139.440 ;
        RECT 145.210 139.160 145.350 139.300 ;
        RECT 135.000 139.100 135.320 139.160 ;
        RECT 133.250 138.960 135.320 139.100 ;
        RECT 135.000 138.900 135.320 138.960 ;
        RECT 135.460 138.900 135.780 139.160 ;
        RECT 140.520 138.900 140.840 139.160 ;
        RECT 140.980 139.100 141.300 139.160 ;
        RECT 141.455 139.100 141.745 139.145 ;
        RECT 140.980 138.960 141.745 139.100 ;
        RECT 140.980 138.900 141.300 138.960 ;
        RECT 141.455 138.915 141.745 138.960 ;
        RECT 141.900 138.900 142.220 139.160 ;
        RECT 142.375 139.100 142.665 139.145 ;
        RECT 145.120 139.100 145.440 139.160 ;
        RECT 142.375 138.960 145.440 139.100 ;
        RECT 142.375 138.915 142.665 138.960 ;
        RECT 145.120 138.900 145.440 138.960 ;
        RECT 146.040 138.900 146.360 139.160 ;
        RECT 146.590 139.100 146.730 139.300 ;
        RECT 148.770 139.255 149.120 139.485 ;
        RECT 148.800 139.240 149.120 139.255 ;
        RECT 154.335 139.100 154.625 139.145 ;
        RECT 146.590 138.960 154.625 139.100 ;
        RECT 154.335 138.915 154.625 138.960 ;
        RECT 22.690 138.280 157.810 138.760 ;
        RECT 31.960 137.880 32.280 138.140 ;
        RECT 36.115 138.080 36.405 138.125 ;
        RECT 36.560 138.080 36.880 138.140 ;
        RECT 36.115 137.940 36.880 138.080 ;
        RECT 36.115 137.895 36.405 137.940 ;
        RECT 36.560 137.880 36.880 137.940 ;
        RECT 42.080 137.880 42.400 138.140 ;
        RECT 54.975 138.080 55.265 138.125 ;
        RECT 54.590 137.940 55.265 138.080 ;
        RECT 25.060 137.200 25.380 137.460 ;
        RECT 26.410 137.400 26.700 137.445 ;
        RECT 26.410 137.260 30.350 137.400 ;
        RECT 26.410 137.215 26.700 137.260 ;
        RECT 25.955 137.060 26.245 137.105 ;
        RECT 27.145 137.060 27.435 137.105 ;
        RECT 29.665 137.060 29.955 137.105 ;
        RECT 25.955 136.920 29.955 137.060 ;
        RECT 30.210 137.060 30.350 137.260 ;
        RECT 33.340 137.200 33.660 137.460 ;
        RECT 34.260 137.400 34.580 137.460 ;
        RECT 34.735 137.400 35.025 137.445 ;
        RECT 36.100 137.400 36.420 137.460 ;
        RECT 34.260 137.260 36.420 137.400 ;
        RECT 34.260 137.200 34.580 137.260 ;
        RECT 34.735 137.215 35.025 137.260 ;
        RECT 36.100 137.200 36.420 137.260 ;
        RECT 41.735 137.400 42.025 137.445 ;
        RECT 42.170 137.400 42.310 137.880 ;
        RECT 54.590 137.460 54.730 137.940 ;
        RECT 54.975 137.895 55.265 137.940 ;
        RECT 59.100 137.880 59.420 138.140 ;
        RECT 60.020 137.880 60.340 138.140 ;
        RECT 62.320 138.080 62.640 138.140 ;
        RECT 62.320 137.940 64.850 138.080 ;
        RECT 62.320 137.880 62.640 137.940 ;
        RECT 59.190 137.740 59.330 137.880 ;
        RECT 59.575 137.740 59.865 137.785 ;
        RECT 55.050 137.600 57.950 137.740 ;
        RECT 55.050 137.460 55.190 137.600 ;
        RECT 57.810 137.460 57.950 137.600 ;
        RECT 58.270 137.600 59.865 137.740 ;
        RECT 60.110 137.740 60.250 137.880 ;
        RECT 64.710 137.740 64.850 137.940 ;
        RECT 65.080 137.880 65.400 138.140 ;
        RECT 71.060 138.080 71.380 138.140 ;
        RECT 70.690 137.940 71.380 138.080 ;
        RECT 70.690 137.785 70.830 137.940 ;
        RECT 71.060 137.880 71.380 137.940 ;
        RECT 71.520 138.080 71.840 138.140 ;
        RECT 72.455 138.080 72.745 138.125 ;
        RECT 71.520 137.940 72.745 138.080 ;
        RECT 71.520 137.880 71.840 137.940 ;
        RECT 72.455 137.895 72.745 137.940 ;
        RECT 74.280 137.880 74.600 138.140 ;
        RECT 74.740 137.880 75.060 138.140 ;
        RECT 85.320 138.080 85.640 138.140 ;
        RECT 86.255 138.080 86.545 138.125 ;
        RECT 95.440 138.080 95.760 138.140 ;
        RECT 85.320 137.940 95.760 138.080 ;
        RECT 85.320 137.880 85.640 137.940 ;
        RECT 86.255 137.895 86.545 137.940 ;
        RECT 95.440 137.880 95.760 137.940 ;
        RECT 95.915 138.080 96.205 138.125 ;
        RECT 95.915 137.940 97.050 138.080 ;
        RECT 95.915 137.895 96.205 137.940 ;
        RECT 65.555 137.740 65.845 137.785 ;
        RECT 60.110 137.600 62.550 137.740 ;
        RECT 64.710 137.600 65.845 137.740 ;
        RECT 41.735 137.260 42.310 137.400 ;
        RECT 41.735 137.215 42.025 137.260 ;
        RECT 54.040 137.200 54.360 137.460 ;
        RECT 54.500 137.200 54.820 137.460 ;
        RECT 54.960 137.200 55.280 137.460 ;
        RECT 57.720 137.200 58.040 137.460 ;
        RECT 58.270 137.445 58.410 137.600 ;
        RECT 59.575 137.555 59.865 137.600 ;
        RECT 58.195 137.215 58.485 137.445 ;
        RECT 59.115 137.400 59.405 137.445 ;
        RECT 60.495 137.400 60.785 137.445 ;
        RECT 60.940 137.400 61.260 137.460 ;
        RECT 59.115 137.260 61.260 137.400 ;
        RECT 59.115 137.215 59.405 137.260 ;
        RECT 60.495 137.215 60.785 137.260 ;
        RECT 60.940 137.200 61.260 137.260 ;
        RECT 61.415 137.390 61.705 137.445 ;
        RECT 61.860 137.390 62.180 137.460 ;
        RECT 62.410 137.445 62.550 137.600 ;
        RECT 65.555 137.555 65.845 137.600 ;
        RECT 66.705 137.570 66.995 137.615 ;
        RECT 61.415 137.250 62.180 137.390 ;
        RECT 61.415 137.215 61.705 137.250 ;
        RECT 61.860 137.200 62.180 137.250 ;
        RECT 62.335 137.215 62.625 137.445 ;
        RECT 62.780 137.400 63.100 137.460 ;
        RECT 66.630 137.400 66.995 137.570 ;
        RECT 70.615 137.555 70.905 137.785 ;
        RECT 74.370 137.740 74.510 137.880 ;
        RECT 71.150 137.600 74.510 137.740 ;
        RECT 82.190 137.600 89.230 137.740 ;
        RECT 62.780 137.385 66.995 137.400 ;
        RECT 69.695 137.400 69.985 137.445 ;
        RECT 70.140 137.400 70.460 137.460 ;
        RECT 71.150 137.445 71.290 137.600 ;
        RECT 82.190 137.460 82.330 137.600 ;
        RECT 71.075 137.400 71.365 137.445 ;
        RECT 62.780 137.260 66.770 137.385 ;
        RECT 69.695 137.260 70.460 137.400 ;
        RECT 62.780 137.200 63.100 137.260 ;
        RECT 69.695 137.215 69.985 137.260 ;
        RECT 70.140 137.200 70.460 137.260 ;
        RECT 70.690 137.260 71.365 137.400 ;
        RECT 32.435 137.060 32.725 137.105 ;
        RECT 30.210 136.920 32.725 137.060 ;
        RECT 25.955 136.875 26.245 136.920 ;
        RECT 27.145 136.875 27.435 136.920 ;
        RECT 29.665 136.875 29.955 136.920 ;
        RECT 32.435 136.875 32.725 136.920 ;
        RECT 38.425 137.060 38.715 137.105 ;
        RECT 40.945 137.060 41.235 137.105 ;
        RECT 42.135 137.060 42.425 137.105 ;
        RECT 38.425 136.920 42.425 137.060 ;
        RECT 38.425 136.875 38.715 136.920 ;
        RECT 40.945 136.875 41.235 136.920 ;
        RECT 42.135 136.875 42.425 136.920 ;
        RECT 43.015 136.875 43.305 137.105 ;
        RECT 25.560 136.720 25.850 136.765 ;
        RECT 27.660 136.720 27.950 136.765 ;
        RECT 29.230 136.720 29.520 136.765 ;
        RECT 25.560 136.580 29.520 136.720 ;
        RECT 25.560 136.535 25.850 136.580 ;
        RECT 27.660 136.535 27.950 136.580 ;
        RECT 29.230 136.535 29.520 136.580 ;
        RECT 34.275 136.720 34.565 136.765 ;
        RECT 34.720 136.720 35.040 136.780 ;
        RECT 34.275 136.580 35.040 136.720 ;
        RECT 34.275 136.535 34.565 136.580 ;
        RECT 34.720 136.520 35.040 136.580 ;
        RECT 38.860 136.720 39.150 136.765 ;
        RECT 40.430 136.720 40.720 136.765 ;
        RECT 42.530 136.720 42.820 136.765 ;
        RECT 38.860 136.580 42.820 136.720 ;
        RECT 38.860 136.535 39.150 136.580 ;
        RECT 40.430 136.535 40.720 136.580 ;
        RECT 42.530 136.535 42.820 136.580 ;
        RECT 42.080 136.380 42.400 136.440 ;
        RECT 43.090 136.380 43.230 136.875 ;
        RECT 52.660 136.860 52.980 137.120 ;
        RECT 53.120 137.060 53.440 137.120 ;
        RECT 57.275 137.060 57.565 137.105 ;
        RECT 53.120 136.920 57.565 137.060 ;
        RECT 53.120 136.860 53.440 136.920 ;
        RECT 57.275 136.875 57.565 136.920 ;
        RECT 65.080 137.060 65.400 137.120 ;
        RECT 70.690 137.060 70.830 137.260 ;
        RECT 71.075 137.215 71.365 137.260 ;
        RECT 71.520 137.200 71.840 137.460 ;
        RECT 75.200 137.400 75.520 137.460 ;
        RECT 80.320 137.400 80.610 137.445 ;
        RECT 75.200 137.260 80.610 137.400 ;
        RECT 75.200 137.200 75.520 137.260 ;
        RECT 80.320 137.215 80.610 137.260 ;
        RECT 81.655 137.400 81.945 137.445 ;
        RECT 82.100 137.400 82.420 137.460 ;
        RECT 81.655 137.260 82.420 137.400 ;
        RECT 81.655 137.215 81.945 137.260 ;
        RECT 82.100 137.200 82.420 137.260 ;
        RECT 83.020 137.400 83.340 137.460 ;
        RECT 89.090 137.445 89.230 137.600 ;
        RECT 90.010 137.600 96.590 137.740 ;
        RECT 85.335 137.400 85.625 137.445 ;
        RECT 83.020 137.260 88.850 137.400 ;
        RECT 83.020 137.200 83.340 137.260 ;
        RECT 85.335 137.215 85.625 137.260 ;
        RECT 65.080 136.920 70.830 137.060 ;
        RECT 77.065 137.060 77.355 137.105 ;
        RECT 79.585 137.060 79.875 137.105 ;
        RECT 80.775 137.060 81.065 137.105 ;
        RECT 77.065 136.920 81.065 137.060 ;
        RECT 88.710 137.060 88.850 137.260 ;
        RECT 89.015 137.215 89.305 137.445 ;
        RECT 90.010 137.400 90.150 137.600 ;
        RECT 90.380 137.445 90.700 137.460 ;
        RECT 89.550 137.260 90.150 137.400 ;
        RECT 89.550 137.060 89.690 137.260 ;
        RECT 90.350 137.215 90.700 137.445 ;
        RECT 90.380 137.200 90.700 137.215 ;
        RECT 88.710 136.920 89.690 137.060 ;
        RECT 89.895 137.060 90.185 137.105 ;
        RECT 91.085 137.060 91.375 137.105 ;
        RECT 93.605 137.060 93.895 137.105 ;
        RECT 89.895 136.920 93.895 137.060 ;
        RECT 52.750 136.720 52.890 136.860 ;
        RECT 57.350 136.720 57.490 136.875 ;
        RECT 65.080 136.860 65.400 136.920 ;
        RECT 77.065 136.875 77.355 136.920 ;
        RECT 79.585 136.875 79.875 136.920 ;
        RECT 80.775 136.875 81.065 136.920 ;
        RECT 89.895 136.875 90.185 136.920 ;
        RECT 91.085 136.875 91.375 136.920 ;
        RECT 93.605 136.875 93.895 136.920 ;
        RECT 72.900 136.720 73.220 136.780 ;
        RECT 52.750 136.580 57.030 136.720 ;
        RECT 57.350 136.580 73.220 136.720 ;
        RECT 42.080 136.240 43.230 136.380 ;
        RECT 52.200 136.380 52.520 136.440 ;
        RECT 53.135 136.380 53.425 136.425 ;
        RECT 52.200 136.240 53.425 136.380 ;
        RECT 56.890 136.380 57.030 136.580 ;
        RECT 72.900 136.520 73.220 136.580 ;
        RECT 77.500 136.720 77.790 136.765 ;
        RECT 79.070 136.720 79.360 136.765 ;
        RECT 81.170 136.720 81.460 136.765 ;
        RECT 77.500 136.580 81.460 136.720 ;
        RECT 77.500 136.535 77.790 136.580 ;
        RECT 79.070 136.535 79.360 136.580 ;
        RECT 81.170 136.535 81.460 136.580 ;
        RECT 89.500 136.720 89.790 136.765 ;
        RECT 91.600 136.720 91.890 136.765 ;
        RECT 93.170 136.720 93.460 136.765 ;
        RECT 89.500 136.580 93.460 136.720 ;
        RECT 96.450 136.720 96.590 137.600 ;
        RECT 96.910 137.460 97.050 137.940 ;
        RECT 99.580 137.880 99.900 138.140 ;
        RECT 101.435 138.080 101.725 138.125 ;
        RECT 102.340 138.080 102.660 138.140 ;
        RECT 101.435 137.940 102.660 138.080 ;
        RECT 101.435 137.895 101.725 137.940 ;
        RECT 102.340 137.880 102.660 137.940 ;
        RECT 102.815 138.080 103.105 138.125 ;
        RECT 108.320 138.080 108.640 138.140 ;
        RECT 102.815 137.940 108.640 138.080 ;
        RECT 102.815 137.895 103.105 137.940 ;
        RECT 96.820 137.400 97.140 137.460 ;
        RECT 97.295 137.400 97.585 137.445 ;
        RECT 96.820 137.260 97.585 137.400 ;
        RECT 96.820 137.200 97.140 137.260 ;
        RECT 97.295 137.215 97.585 137.260 ;
        RECT 98.215 137.400 98.505 137.445 ;
        RECT 99.670 137.400 99.810 137.880 ;
        RECT 100.515 137.400 100.805 137.445 ;
        RECT 102.890 137.400 103.030 137.895 ;
        RECT 104.270 137.460 104.410 137.940 ;
        RECT 108.320 137.880 108.640 137.940 ;
        RECT 109.240 138.080 109.560 138.140 ;
        RECT 112.475 138.080 112.765 138.125 ;
        RECT 109.240 137.940 112.765 138.080 ;
        RECT 109.240 137.880 109.560 137.940 ;
        RECT 112.475 137.895 112.765 137.940 ;
        RECT 114.300 137.880 114.620 138.140 ;
        RECT 114.760 137.880 115.080 138.140 ;
        RECT 115.220 137.880 115.540 138.140 ;
        RECT 117.075 138.080 117.365 138.125 ;
        RECT 117.980 138.080 118.300 138.140 ;
        RECT 117.075 137.940 118.300 138.080 ;
        RECT 117.075 137.895 117.365 137.940 ;
        RECT 117.980 137.880 118.300 137.940 ;
        RECT 121.660 138.080 121.980 138.140 ;
        RECT 122.595 138.080 122.885 138.125 ;
        RECT 121.660 137.940 122.885 138.080 ;
        RECT 121.660 137.880 121.980 137.940 ;
        RECT 122.595 137.895 122.885 137.940 ;
        RECT 126.275 137.895 126.565 138.125 ;
        RECT 114.390 137.740 114.530 137.880 ;
        RECT 105.190 137.600 114.530 137.740 ;
        RECT 114.850 137.740 114.990 137.880 ;
        RECT 117.535 137.740 117.825 137.785 ;
        RECT 114.850 137.600 117.825 137.740 ;
        RECT 98.215 137.260 99.350 137.400 ;
        RECT 99.670 137.260 100.805 137.400 ;
        RECT 98.215 137.215 98.505 137.260 ;
        RECT 99.210 137.060 99.350 137.260 ;
        RECT 100.515 137.215 100.805 137.260 ;
        RECT 101.050 137.260 103.030 137.400 ;
        RECT 101.050 137.060 101.190 137.260 ;
        RECT 103.735 137.215 104.025 137.445 ;
        RECT 99.210 136.920 101.190 137.060 ;
        RECT 103.810 137.060 103.950 137.215 ;
        RECT 104.180 137.200 104.500 137.460 ;
        RECT 105.190 137.445 105.330 137.600 ;
        RECT 117.535 137.555 117.825 137.600 ;
        RECT 105.115 137.215 105.405 137.445 ;
        RECT 105.560 137.200 105.880 137.460 ;
        RECT 106.450 137.400 106.740 137.445 ;
        RECT 107.860 137.400 108.180 137.460 ;
        RECT 106.450 137.260 108.180 137.400 ;
        RECT 106.450 137.215 106.740 137.260 ;
        RECT 107.860 137.200 108.180 137.260 ;
        RECT 108.320 137.400 108.640 137.460 ;
        RECT 113.395 137.400 113.685 137.445 ;
        RECT 117.060 137.400 117.380 137.460 ;
        RECT 108.320 137.260 113.150 137.400 ;
        RECT 108.320 137.200 108.640 137.260 ;
        RECT 105.650 137.060 105.790 137.200 ;
        RECT 103.810 136.920 105.790 137.060 ;
        RECT 105.995 137.060 106.285 137.105 ;
        RECT 107.185 137.060 107.475 137.105 ;
        RECT 109.705 137.060 109.995 137.105 ;
        RECT 105.995 136.920 109.995 137.060 ;
        RECT 113.010 137.060 113.150 137.260 ;
        RECT 113.395 137.260 117.380 137.400 ;
        RECT 113.395 137.215 113.685 137.260 ;
        RECT 114.315 137.060 114.605 137.105 ;
        RECT 113.010 136.920 114.605 137.060 ;
        RECT 103.810 136.720 103.950 136.920 ;
        RECT 105.995 136.875 106.285 136.920 ;
        RECT 107.185 136.875 107.475 136.920 ;
        RECT 109.705 136.875 109.995 136.920 ;
        RECT 114.315 136.875 114.605 136.920 ;
        RECT 96.450 136.580 103.950 136.720 ;
        RECT 105.600 136.720 105.890 136.765 ;
        RECT 107.700 136.720 107.990 136.765 ;
        RECT 109.270 136.720 109.560 136.765 ;
        RECT 105.600 136.580 109.560 136.720 ;
        RECT 89.500 136.535 89.790 136.580 ;
        RECT 91.600 136.535 91.890 136.580 ;
        RECT 93.170 136.535 93.460 136.580 ;
        RECT 105.600 136.535 105.890 136.580 ;
        RECT 107.700 136.535 107.990 136.580 ;
        RECT 109.270 136.535 109.560 136.580 ;
        RECT 112.015 136.720 112.305 136.765 ;
        RECT 114.850 136.720 114.990 137.260 ;
        RECT 117.060 137.200 117.380 137.260 ;
        RECT 123.515 137.400 123.805 137.445 ;
        RECT 126.350 137.400 126.490 137.895 ;
        RECT 128.100 137.880 128.420 138.140 ;
        RECT 128.575 138.080 128.865 138.125 ;
        RECT 129.940 138.080 130.260 138.140 ;
        RECT 128.575 137.940 130.260 138.080 ;
        RECT 128.575 137.895 128.865 137.940 ;
        RECT 129.940 137.880 130.260 137.940 ;
        RECT 130.400 137.880 130.720 138.140 ;
        RECT 131.780 137.880 132.100 138.140 ;
        RECT 132.700 138.080 133.020 138.140 ;
        RECT 135.000 138.080 135.320 138.140 ;
        RECT 140.995 138.080 141.285 138.125 ;
        RECT 141.440 138.080 141.760 138.140 ;
        RECT 132.700 137.940 134.770 138.080 ;
        RECT 132.700 137.880 133.020 137.940 ;
        RECT 130.490 137.740 130.630 137.880 ;
        RECT 131.870 137.740 132.010 137.880 ;
        RECT 134.630 137.785 134.770 137.940 ;
        RECT 135.000 137.940 140.750 138.080 ;
        RECT 135.000 137.880 135.320 137.940 ;
        RECT 134.555 137.740 134.845 137.785 ;
        RECT 138.680 137.740 139.000 137.800 ;
        RECT 140.610 137.740 140.750 137.940 ;
        RECT 140.995 137.940 141.760 138.080 ;
        RECT 140.995 137.895 141.285 137.940 ;
        RECT 141.440 137.880 141.760 137.940 ;
        RECT 143.295 138.080 143.585 138.125 ;
        RECT 143.740 138.080 144.060 138.140 ;
        RECT 143.295 137.940 144.060 138.080 ;
        RECT 143.295 137.895 143.585 137.940 ;
        RECT 143.740 137.880 144.060 137.940 ;
        RECT 144.215 137.895 144.505 138.125 ;
        RECT 144.660 138.080 144.980 138.140 ;
        RECT 145.135 138.080 145.425 138.125 ;
        RECT 144.660 137.940 145.425 138.080 ;
        RECT 144.290 137.740 144.430 137.895 ;
        RECT 144.660 137.880 144.980 137.940 ;
        RECT 145.135 137.895 145.425 137.940 ;
        RECT 145.580 138.080 145.900 138.140 ;
        RECT 145.580 137.940 147.190 138.080 ;
        RECT 145.580 137.880 145.900 137.940 ;
        RECT 130.490 137.600 131.550 137.740 ;
        RECT 131.870 137.600 132.930 137.740 ;
        RECT 123.515 137.260 126.490 137.400 ;
        RECT 126.720 137.400 127.040 137.460 ;
        RECT 131.410 137.400 131.550 137.600 ;
        RECT 132.790 137.445 132.930 137.600 ;
        RECT 134.555 137.600 135.690 137.740 ;
        RECT 134.555 137.555 134.845 137.600 ;
        RECT 132.255 137.400 132.545 137.445 ;
        RECT 126.720 137.260 131.090 137.400 ;
        RECT 131.410 137.260 132.545 137.400 ;
        RECT 123.515 137.215 123.805 137.260 ;
        RECT 126.720 137.200 127.040 137.260 ;
        RECT 118.440 137.060 118.760 137.120 ;
        RECT 129.035 137.060 129.325 137.105 ;
        RECT 118.440 136.920 129.325 137.060 ;
        RECT 130.950 137.060 131.090 137.260 ;
        RECT 132.255 137.215 132.545 137.260 ;
        RECT 132.715 137.215 133.005 137.445 ;
        RECT 135.000 137.200 135.320 137.460 ;
        RECT 135.550 137.445 135.690 137.600 ;
        RECT 138.680 137.600 140.290 137.740 ;
        RECT 140.610 137.600 141.210 137.740 ;
        RECT 144.290 137.600 146.730 137.740 ;
        RECT 138.680 137.540 139.000 137.600 ;
        RECT 140.150 137.445 140.290 137.600 ;
        RECT 135.475 137.215 135.765 137.445 ;
        RECT 140.075 137.215 140.365 137.445 ;
        RECT 140.520 137.200 140.840 137.460 ;
        RECT 141.070 137.445 141.210 137.600 ;
        RECT 140.995 137.400 141.285 137.445 ;
        RECT 144.660 137.400 144.980 137.460 ;
        RECT 140.995 137.260 144.980 137.400 ;
        RECT 140.995 137.215 141.285 137.260 ;
        RECT 144.660 137.200 144.980 137.260 ;
        RECT 145.120 137.400 145.440 137.460 ;
        RECT 146.590 137.445 146.730 137.600 ;
        RECT 145.595 137.400 145.885 137.445 ;
        RECT 145.120 137.260 145.885 137.400 ;
        RECT 145.120 137.200 145.440 137.260 ;
        RECT 145.595 137.215 145.885 137.260 ;
        RECT 146.515 137.215 146.805 137.445 ;
        RECT 147.050 137.400 147.190 137.940 ;
        RECT 147.435 137.895 147.725 138.125 ;
        RECT 147.510 137.740 147.650 137.895 ;
        RECT 148.800 137.880 149.120 138.140 ;
        RECT 151.100 137.740 151.420 137.800 ;
        RECT 147.510 137.600 151.420 137.740 ;
        RECT 151.100 137.540 151.420 137.600 ;
        RECT 147.895 137.400 148.185 137.445 ;
        RECT 147.050 137.260 148.185 137.400 ;
        RECT 147.895 137.215 148.185 137.260 ;
        RECT 140.610 137.060 140.750 137.200 ;
        RECT 141.440 137.060 141.760 137.120 ;
        RECT 130.950 136.920 137.530 137.060 ;
        RECT 140.610 136.920 141.760 137.060 ;
        RECT 118.440 136.860 118.760 136.920 ;
        RECT 129.035 136.875 129.325 136.920 ;
        RECT 135.000 136.720 135.320 136.780 ;
        RECT 137.390 136.720 137.530 136.920 ;
        RECT 141.440 136.860 141.760 136.920 ;
        RECT 142.820 136.860 143.140 137.120 ;
        RECT 142.910 136.720 143.050 136.860 ;
        RECT 112.015 136.580 114.990 136.720 ;
        RECT 134.170 136.580 136.610 136.720 ;
        RECT 137.390 136.580 143.050 136.720 ;
        RECT 143.370 136.580 146.270 136.720 ;
        RECT 112.015 136.535 112.305 136.580 ;
        RECT 57.720 136.380 58.040 136.440 ;
        RECT 56.890 136.240 58.040 136.380 ;
        RECT 42.080 136.180 42.400 136.240 ;
        RECT 52.200 136.180 52.520 136.240 ;
        RECT 53.135 136.195 53.425 136.240 ;
        RECT 57.720 136.180 58.040 136.240 ;
        RECT 58.655 136.380 58.945 136.425 ;
        RECT 61.400 136.380 61.720 136.440 ;
        RECT 66.475 136.380 66.765 136.425 ;
        RECT 58.655 136.240 66.765 136.380 ;
        RECT 58.655 136.195 58.945 136.240 ;
        RECT 61.400 136.180 61.720 136.240 ;
        RECT 66.475 136.195 66.765 136.240 ;
        RECT 67.395 136.380 67.685 136.425 ;
        RECT 74.280 136.380 74.600 136.440 ;
        RECT 67.395 136.240 74.600 136.380 ;
        RECT 67.395 136.195 67.685 136.240 ;
        RECT 74.280 136.180 74.600 136.240 ;
        RECT 76.120 136.380 76.440 136.440 ;
        RECT 88.540 136.380 88.860 136.440 ;
        RECT 76.120 136.240 88.860 136.380 ;
        RECT 76.120 136.180 76.440 136.240 ;
        RECT 88.540 136.180 88.860 136.240 ;
        RECT 96.360 136.180 96.680 136.440 ;
        RECT 131.335 136.380 131.625 136.425 ;
        RECT 131.780 136.380 132.100 136.440 ;
        RECT 134.170 136.425 134.310 136.580 ;
        RECT 135.000 136.520 135.320 136.580 ;
        RECT 136.470 136.440 136.610 136.580 ;
        RECT 131.335 136.240 132.100 136.380 ;
        RECT 131.335 136.195 131.625 136.240 ;
        RECT 131.780 136.180 132.100 136.240 ;
        RECT 134.095 136.195 134.385 136.425 ;
        RECT 135.460 136.180 135.780 136.440 ;
        RECT 136.380 136.180 136.700 136.440 ;
        RECT 136.840 136.180 137.160 136.440 ;
        RECT 143.370 136.425 143.510 136.580 ;
        RECT 146.130 136.440 146.270 136.580 ;
        RECT 143.295 136.195 143.585 136.425 ;
        RECT 146.040 136.180 146.360 136.440 ;
        RECT 22.690 135.560 157.010 136.040 ;
        RECT 33.340 135.160 33.660 135.420 ;
        RECT 49.455 135.360 49.745 135.405 ;
        RECT 50.820 135.360 51.140 135.420 ;
        RECT 49.455 135.220 51.140 135.360 ;
        RECT 49.455 135.175 49.745 135.220 ;
        RECT 50.820 135.160 51.140 135.220 ;
        RECT 64.160 135.160 64.480 135.420 ;
        RECT 66.920 135.160 67.240 135.420 ;
        RECT 75.200 135.160 75.520 135.420 ;
        RECT 75.660 135.360 75.980 135.420 ;
        RECT 77.040 135.360 77.360 135.420 ;
        RECT 80.735 135.360 81.025 135.405 ;
        RECT 75.660 135.220 81.025 135.360 ;
        RECT 75.660 135.160 75.980 135.220 ;
        RECT 77.040 135.160 77.360 135.220 ;
        RECT 80.735 135.175 81.025 135.220 ;
        RECT 90.380 135.360 90.700 135.420 ;
        RECT 91.315 135.360 91.605 135.405 ;
        RECT 97.740 135.360 98.060 135.420 ;
        RECT 102.340 135.360 102.660 135.420 ;
        RECT 118.440 135.360 118.760 135.420 ;
        RECT 90.380 135.220 91.605 135.360 ;
        RECT 90.380 135.160 90.700 135.220 ;
        RECT 91.315 135.175 91.605 135.220 ;
        RECT 96.450 135.220 102.660 135.360 ;
        RECT 43.040 135.020 43.330 135.065 ;
        RECT 45.140 135.020 45.430 135.065 ;
        RECT 46.710 135.020 47.000 135.065 ;
        RECT 43.040 134.880 47.000 135.020 ;
        RECT 43.040 134.835 43.330 134.880 ;
        RECT 45.140 134.835 45.430 134.880 ;
        RECT 46.710 134.835 47.000 134.880 ;
        RECT 50.400 135.020 50.690 135.065 ;
        RECT 52.500 135.020 52.790 135.065 ;
        RECT 54.070 135.020 54.360 135.065 ;
        RECT 50.400 134.880 54.360 135.020 ;
        RECT 50.400 134.835 50.690 134.880 ;
        RECT 52.500 134.835 52.790 134.880 ;
        RECT 54.070 134.835 54.360 134.880 ;
        RECT 56.815 134.835 57.105 135.065 ;
        RECT 67.010 135.020 67.150 135.160 ;
        RECT 76.580 135.020 76.900 135.080 ;
        RECT 84.400 135.020 84.720 135.080 ;
        RECT 67.010 134.880 84.720 135.020 ;
        RECT 32.880 134.680 33.200 134.740 ;
        RECT 43.435 134.680 43.725 134.725 ;
        RECT 44.625 134.680 44.915 134.725 ;
        RECT 47.145 134.680 47.435 134.725 ;
        RECT 30.210 134.540 37.250 134.680 ;
        RECT 30.210 134.385 30.350 134.540 ;
        RECT 32.880 134.480 33.200 134.540 ;
        RECT 30.135 134.155 30.425 134.385 ;
        RECT 30.580 134.140 30.900 134.400 ;
        RECT 31.055 134.155 31.345 134.385 ;
        RECT 28.280 134.000 28.600 134.060 ;
        RECT 29.660 134.000 29.980 134.060 ;
        RECT 31.130 134.000 31.270 134.155 ;
        RECT 31.960 134.140 32.280 134.400 ;
        RECT 32.435 134.155 32.725 134.385 ;
        RECT 28.280 133.860 29.430 134.000 ;
        RECT 28.280 133.800 28.600 133.860 ;
        RECT 28.740 133.460 29.060 133.720 ;
        RECT 29.290 133.660 29.430 133.860 ;
        RECT 29.660 133.860 31.270 134.000 ;
        RECT 31.500 134.000 31.820 134.060 ;
        RECT 32.510 134.000 32.650 134.155 ;
        RECT 34.260 134.140 34.580 134.400 ;
        RECT 34.720 134.140 35.040 134.400 ;
        RECT 37.110 134.385 37.250 134.540 ;
        RECT 43.435 134.540 47.435 134.680 ;
        RECT 43.435 134.495 43.725 134.540 ;
        RECT 44.625 134.495 44.915 134.540 ;
        RECT 47.145 134.495 47.435 134.540 ;
        RECT 50.795 134.680 51.085 134.725 ;
        RECT 51.985 134.680 52.275 134.725 ;
        RECT 54.505 134.680 54.795 134.725 ;
        RECT 50.795 134.540 54.795 134.680 ;
        RECT 56.890 134.680 57.030 134.835 ;
        RECT 76.580 134.820 76.900 134.880 ;
        RECT 84.400 134.820 84.720 134.880 ;
        RECT 60.035 134.680 60.325 134.725 ;
        RECT 56.890 134.540 60.325 134.680 ;
        RECT 50.795 134.495 51.085 134.540 ;
        RECT 51.985 134.495 52.275 134.540 ;
        RECT 54.505 134.495 54.795 134.540 ;
        RECT 60.035 134.495 60.325 134.540 ;
        RECT 60.940 134.680 61.260 134.740 ;
        RECT 65.080 134.680 65.400 134.740 ;
        RECT 94.520 134.680 94.840 134.740 ;
        RECT 95.455 134.680 95.745 134.725 ;
        RECT 60.940 134.540 65.400 134.680 ;
        RECT 60.940 134.480 61.260 134.540 ;
        RECT 65.080 134.480 65.400 134.540 ;
        RECT 70.690 134.540 94.290 134.680 ;
        RECT 37.035 134.155 37.325 134.385 ;
        RECT 42.080 134.340 42.400 134.400 ;
        RECT 42.555 134.340 42.845 134.385 ;
        RECT 49.915 134.340 50.205 134.385 ;
        RECT 42.080 134.200 50.205 134.340 ;
        RECT 42.080 134.140 42.400 134.200 ;
        RECT 42.555 134.155 42.845 134.200 ;
        RECT 49.915 134.155 50.205 134.200 ;
        RECT 50.360 134.340 50.680 134.400 ;
        RECT 70.690 134.385 70.830 134.540 ;
        RECT 50.360 134.200 57.950 134.340 ;
        RECT 50.360 134.140 50.680 134.200 ;
        RECT 36.560 134.000 36.880 134.060 ;
        RECT 37.955 134.000 38.245 134.045 ;
        RECT 31.500 133.860 32.650 134.000 ;
        RECT 33.660 133.860 36.330 134.000 ;
        RECT 29.660 133.800 29.980 133.860 ;
        RECT 31.500 133.800 31.820 133.860 ;
        RECT 33.660 133.660 33.800 133.860 ;
        RECT 36.190 133.705 36.330 133.860 ;
        RECT 36.560 133.860 38.245 134.000 ;
        RECT 36.560 133.800 36.880 133.860 ;
        RECT 37.955 133.815 38.245 133.860 ;
        RECT 43.890 134.000 44.180 134.045 ;
        RECT 51.250 134.000 51.540 134.045 ;
        RECT 52.660 134.000 52.980 134.060 ;
        RECT 43.890 133.860 50.130 134.000 ;
        RECT 43.890 133.815 44.180 133.860 ;
        RECT 29.290 133.520 33.800 133.660 ;
        RECT 36.115 133.475 36.405 133.705 ;
        RECT 49.990 133.660 50.130 133.860 ;
        RECT 51.250 133.860 52.980 134.000 ;
        RECT 51.250 133.815 51.540 133.860 ;
        RECT 52.660 133.800 52.980 133.860 ;
        RECT 52.200 133.660 52.520 133.720 ;
        RECT 49.990 133.520 52.520 133.660 ;
        RECT 52.200 133.460 52.520 133.520 ;
        RECT 57.260 133.460 57.580 133.720 ;
        RECT 57.810 133.660 57.950 134.200 ;
        RECT 70.615 134.155 70.905 134.385 ;
        RECT 74.755 134.340 75.045 134.385 ;
        RECT 74.755 134.200 75.890 134.340 ;
        RECT 74.755 134.155 75.045 134.200 ;
        RECT 58.180 134.000 58.500 134.060 ;
        RECT 69.680 134.000 70.000 134.060 ;
        RECT 73.360 134.000 73.680 134.060 ;
        RECT 58.180 133.860 73.680 134.000 ;
        RECT 58.180 133.800 58.500 133.860 ;
        RECT 69.680 133.800 70.000 133.860 ;
        RECT 73.360 133.800 73.680 133.860 ;
        RECT 75.200 133.800 75.520 134.060 ;
        RECT 75.290 133.660 75.430 133.800 ;
        RECT 57.810 133.520 75.430 133.660 ;
        RECT 75.750 133.660 75.890 134.200 ;
        RECT 76.120 134.140 76.440 134.400 ;
        RECT 76.580 134.140 76.900 134.400 ;
        RECT 77.975 134.340 78.265 134.385 ;
        RECT 79.340 134.340 79.660 134.400 ;
        RECT 87.160 134.340 87.480 134.400 ;
        RECT 77.975 134.200 79.660 134.340 ;
        RECT 77.975 134.155 78.265 134.200 ;
        RECT 79.340 134.140 79.660 134.200 ;
        RECT 79.890 134.200 87.480 134.340 ;
        RECT 77.055 134.000 77.345 134.045 ;
        RECT 79.890 134.000 80.030 134.200 ;
        RECT 87.160 134.140 87.480 134.200 ;
        RECT 92.235 134.340 92.525 134.385 ;
        RECT 92.235 134.200 93.370 134.340 ;
        RECT 92.235 134.155 92.525 134.200 ;
        RECT 77.055 133.860 80.030 134.000 ;
        RECT 77.055 133.815 77.345 133.860 ;
        RECT 80.275 133.815 80.565 134.045 ;
        RECT 78.420 133.660 78.740 133.720 ;
        RECT 80.350 133.660 80.490 133.815 ;
        RECT 93.230 133.705 93.370 134.200 ;
        RECT 94.150 134.060 94.290 134.540 ;
        RECT 94.520 134.540 95.745 134.680 ;
        RECT 94.520 134.480 94.840 134.540 ;
        RECT 95.455 134.495 95.745 134.540 ;
        RECT 95.915 134.680 96.205 134.725 ;
        RECT 96.450 134.680 96.590 135.220 ;
        RECT 97.740 135.160 98.060 135.220 ;
        RECT 102.340 135.160 102.660 135.220 ;
        RECT 102.890 135.220 118.760 135.360 ;
        RECT 102.890 135.020 103.030 135.220 ;
        RECT 118.440 135.160 118.760 135.220 ;
        RECT 119.820 135.160 120.140 135.420 ;
        RECT 146.500 135.360 146.820 135.420 ;
        RECT 146.975 135.360 147.265 135.405 ;
        RECT 146.500 135.220 147.265 135.360 ;
        RECT 146.500 135.160 146.820 135.220 ;
        RECT 146.975 135.175 147.265 135.220 ;
        RECT 123.515 135.020 123.805 135.065 ;
        RECT 95.915 134.540 96.590 134.680 ;
        RECT 97.370 134.880 103.030 135.020 ;
        RECT 112.090 134.880 123.805 135.020 ;
        RECT 95.915 134.495 96.205 134.540 ;
        RECT 97.370 134.400 97.510 134.880 ;
        RECT 98.660 134.480 98.980 134.740 ;
        RECT 112.090 134.400 112.230 134.880 ;
        RECT 123.515 134.835 123.805 134.880 ;
        RECT 149.720 135.020 150.010 135.065 ;
        RECT 151.290 135.020 151.580 135.065 ;
        RECT 153.390 135.020 153.680 135.065 ;
        RECT 149.720 134.880 153.680 135.020 ;
        RECT 149.720 134.835 150.010 134.880 ;
        RECT 151.290 134.835 151.580 134.880 ;
        RECT 153.390 134.835 153.680 134.880 ;
        RECT 149.285 134.680 149.575 134.725 ;
        RECT 151.805 134.680 152.095 134.725 ;
        RECT 152.995 134.680 153.285 134.725 ;
        RECT 149.285 134.540 153.285 134.680 ;
        RECT 149.285 134.495 149.575 134.540 ;
        RECT 151.805 134.495 152.095 134.540 ;
        RECT 152.995 134.495 153.285 134.540 ;
        RECT 94.995 134.340 95.285 134.385 ;
        RECT 96.360 134.340 96.680 134.400 ;
        RECT 94.995 134.200 96.680 134.340 ;
        RECT 94.995 134.155 95.285 134.200 ;
        RECT 96.360 134.140 96.680 134.200 ;
        RECT 97.280 134.140 97.600 134.400 ;
        RECT 99.135 134.340 99.425 134.385 ;
        RECT 100.515 134.340 100.805 134.385 ;
        RECT 99.135 134.200 100.805 134.340 ;
        RECT 99.135 134.155 99.425 134.200 ;
        RECT 100.515 134.155 100.805 134.200 ;
        RECT 100.960 134.340 101.280 134.400 ;
        RECT 103.275 134.340 103.565 134.385 ;
        RECT 100.960 134.200 103.565 134.340 ;
        RECT 100.960 134.140 101.280 134.200 ;
        RECT 103.275 134.155 103.565 134.200 ;
        RECT 107.415 134.340 107.705 134.385 ;
        RECT 108.780 134.340 109.100 134.400 ;
        RECT 107.415 134.200 109.100 134.340 ;
        RECT 107.415 134.155 107.705 134.200 ;
        RECT 108.780 134.140 109.100 134.200 ;
        RECT 111.540 134.140 111.860 134.400 ;
        RECT 112.000 134.140 112.320 134.400 ;
        RECT 122.120 134.340 122.440 134.400 ;
        RECT 122.595 134.340 122.885 134.385 ;
        RECT 122.120 134.200 122.885 134.340 ;
        RECT 122.120 134.140 122.440 134.200 ;
        RECT 122.595 134.155 122.885 134.200 ;
        RECT 124.435 134.155 124.725 134.385 ;
        RECT 94.060 134.000 94.380 134.060 ;
        RECT 113.395 134.000 113.685 134.045 ;
        RECT 94.060 133.860 113.685 134.000 ;
        RECT 94.060 133.800 94.380 133.860 ;
        RECT 113.395 133.815 113.685 133.860 ;
        RECT 113.840 134.000 114.160 134.060 ;
        RECT 124.510 134.000 124.650 134.155 ;
        RECT 125.340 134.140 125.660 134.400 ;
        RECT 133.160 134.340 133.480 134.400 ;
        RECT 138.680 134.340 139.000 134.400 ;
        RECT 133.160 134.200 139.000 134.340 ;
        RECT 133.160 134.140 133.480 134.200 ;
        RECT 138.680 134.140 139.000 134.200 ;
        RECT 140.520 134.340 140.840 134.400 ;
        RECT 143.740 134.340 144.060 134.400 ;
        RECT 140.520 134.200 144.060 134.340 ;
        RECT 140.520 134.140 140.840 134.200 ;
        RECT 143.740 134.140 144.060 134.200 ;
        RECT 151.100 134.340 151.420 134.400 ;
        RECT 152.540 134.340 152.830 134.385 ;
        RECT 151.100 134.200 152.830 134.340 ;
        RECT 151.100 134.140 151.420 134.200 ;
        RECT 152.540 134.155 152.830 134.200 ;
        RECT 153.875 134.340 154.165 134.385 ;
        RECT 154.320 134.340 154.640 134.400 ;
        RECT 153.875 134.200 154.640 134.340 ;
        RECT 153.875 134.155 154.165 134.200 ;
        RECT 154.320 134.140 154.640 134.200 ;
        RECT 113.840 133.860 127.410 134.000 ;
        RECT 113.840 133.800 114.160 133.860 ;
        RECT 127.270 133.720 127.410 133.860 ;
        RECT 75.750 133.520 80.490 133.660 ;
        RECT 78.420 133.460 78.740 133.520 ;
        RECT 93.155 133.475 93.445 133.705 ;
        RECT 97.280 133.460 97.600 133.720 ;
        RECT 108.320 133.460 108.640 133.720 ;
        RECT 109.700 133.660 110.020 133.720 ;
        RECT 110.635 133.660 110.925 133.705 ;
        RECT 109.700 133.520 110.925 133.660 ;
        RECT 109.700 133.460 110.020 133.520 ;
        RECT 110.635 133.475 110.925 133.520 ;
        RECT 124.420 133.460 124.740 133.720 ;
        RECT 127.180 133.460 127.500 133.720 ;
        RECT 137.760 133.660 138.080 133.720 ;
        RECT 140.995 133.660 141.285 133.705 ;
        RECT 143.280 133.660 143.600 133.720 ;
        RECT 137.760 133.520 143.600 133.660 ;
        RECT 137.760 133.460 138.080 133.520 ;
        RECT 140.995 133.475 141.285 133.520 ;
        RECT 143.280 133.460 143.600 133.520 ;
        RECT 22.690 132.840 157.810 133.320 ;
        RECT 28.280 132.440 28.600 132.700 ;
        RECT 28.740 132.440 29.060 132.700 ;
        RECT 32.435 132.640 32.725 132.685 ;
        RECT 32.880 132.640 33.200 132.700 ;
        RECT 32.435 132.500 33.200 132.640 ;
        RECT 32.435 132.455 32.725 132.500 ;
        RECT 32.880 132.440 33.200 132.500 ;
        RECT 53.595 132.640 53.885 132.685 ;
        RECT 54.040 132.640 54.360 132.700 ;
        RECT 53.595 132.500 54.360 132.640 ;
        RECT 53.595 132.455 53.885 132.500 ;
        RECT 54.040 132.440 54.360 132.500 ;
        RECT 57.260 132.440 57.580 132.700 ;
        RECT 57.720 132.640 58.040 132.700 ;
        RECT 62.320 132.640 62.640 132.700 ;
        RECT 57.720 132.500 62.640 132.640 ;
        RECT 57.720 132.440 58.040 132.500 ;
        RECT 28.370 132.300 28.510 132.440 ;
        RECT 26.990 132.160 28.510 132.300 ;
        RECT 24.600 131.960 24.920 132.020 ;
        RECT 26.990 132.005 27.130 132.160 ;
        RECT 28.830 132.005 28.970 132.440 ;
        RECT 42.080 132.300 42.400 132.360 ;
        RECT 57.350 132.300 57.490 132.440 ;
        RECT 59.190 132.345 59.330 132.500 ;
        RECT 62.320 132.440 62.640 132.500 ;
        RECT 65.080 132.440 65.400 132.700 ;
        RECT 72.455 132.455 72.745 132.685 ;
        RECT 60.020 132.345 60.340 132.360 ;
        RECT 36.190 132.160 42.400 132.300 ;
        RECT 25.995 131.960 26.285 132.005 ;
        RECT 24.600 131.820 26.285 131.960 ;
        RECT 24.600 131.760 24.920 131.820 ;
        RECT 25.995 131.775 26.285 131.820 ;
        RECT 26.455 131.775 26.745 132.005 ;
        RECT 26.915 131.775 27.205 132.005 ;
        RECT 27.835 131.775 28.125 132.005 ;
        RECT 28.755 131.775 29.045 132.005 ;
        RECT 26.530 131.280 26.670 131.775 ;
        RECT 27.910 131.620 28.050 131.775 ;
        RECT 31.960 131.760 32.280 132.020 ;
        RECT 32.050 131.620 32.190 131.760 ;
        RECT 27.910 131.480 32.190 131.620 ;
        RECT 35.640 131.420 35.960 131.680 ;
        RECT 36.190 131.665 36.330 132.160 ;
        RECT 42.080 132.100 42.400 132.160 ;
        RECT 48.150 132.160 57.490 132.300 ;
        RECT 37.480 132.005 37.800 132.020 ;
        RECT 37.450 131.775 37.800 132.005 ;
        RECT 37.480 131.760 37.800 131.775 ;
        RECT 41.160 131.960 41.480 132.020 ;
        RECT 48.150 132.005 48.290 132.160 ;
        RECT 41.160 131.820 46.910 131.960 ;
        RECT 41.160 131.760 41.480 131.820 ;
        RECT 36.115 131.435 36.405 131.665 ;
        RECT 36.995 131.620 37.285 131.665 ;
        RECT 38.185 131.620 38.475 131.665 ;
        RECT 40.705 131.620 40.995 131.665 ;
        RECT 36.995 131.480 40.995 131.620 ;
        RECT 36.995 131.435 37.285 131.480 ;
        RECT 38.185 131.435 38.475 131.480 ;
        RECT 40.705 131.435 40.995 131.480 ;
        RECT 46.235 131.435 46.525 131.665 ;
        RECT 46.770 131.620 46.910 131.820 ;
        RECT 48.075 131.775 48.365 132.005 ;
        RECT 49.455 131.960 49.745 132.005 ;
        RECT 50.360 131.960 50.680 132.020 ;
        RECT 49.455 131.820 50.680 131.960 ;
        RECT 49.455 131.775 49.745 131.820 ;
        RECT 49.530 131.620 49.670 131.775 ;
        RECT 50.360 131.760 50.680 131.820 ;
        RECT 50.820 131.760 51.140 132.020 ;
        RECT 52.290 132.005 52.430 132.160 ;
        RECT 59.115 132.115 59.405 132.345 ;
        RECT 60.020 132.115 60.405 132.345 ;
        RECT 70.770 132.300 71.060 132.345 ;
        RECT 72.530 132.300 72.670 132.455 ;
        RECT 74.280 132.440 74.600 132.700 ;
        RECT 96.375 132.640 96.665 132.685 ;
        RECT 98.200 132.640 98.520 132.700 ;
        RECT 99.580 132.640 99.900 132.700 ;
        RECT 96.375 132.500 99.900 132.640 ;
        RECT 96.375 132.455 96.665 132.500 ;
        RECT 98.200 132.440 98.520 132.500 ;
        RECT 99.580 132.440 99.900 132.500 ;
        RECT 100.515 132.640 100.805 132.685 ;
        RECT 100.960 132.640 101.280 132.700 ;
        RECT 100.515 132.500 101.280 132.640 ;
        RECT 100.515 132.455 100.805 132.500 ;
        RECT 100.960 132.440 101.280 132.500 ;
        RECT 108.320 132.440 108.640 132.700 ;
        RECT 111.540 132.640 111.860 132.700 ;
        RECT 114.775 132.640 115.065 132.685 ;
        RECT 111.540 132.500 115.065 132.640 ;
        RECT 111.540 132.440 111.860 132.500 ;
        RECT 114.775 132.455 115.065 132.500 ;
        RECT 124.895 132.640 125.185 132.685 ;
        RECT 126.260 132.640 126.580 132.700 ;
        RECT 124.895 132.500 126.580 132.640 ;
        RECT 124.895 132.455 125.185 132.500 ;
        RECT 70.770 132.160 72.670 132.300 ;
        RECT 70.770 132.115 71.060 132.160 ;
        RECT 60.020 132.100 60.340 132.115 ;
        RECT 52.215 131.775 52.505 132.005 ;
        RECT 52.675 131.960 52.965 132.005 ;
        RECT 53.120 131.960 53.440 132.020 ;
        RECT 52.675 131.820 53.440 131.960 ;
        RECT 52.675 131.775 52.965 131.820 ;
        RECT 53.120 131.760 53.440 131.820 ;
        RECT 53.580 131.960 53.900 132.020 ;
        RECT 54.055 131.960 54.345 132.005 ;
        RECT 53.580 131.820 54.345 131.960 ;
        RECT 53.580 131.760 53.900 131.820 ;
        RECT 54.055 131.775 54.345 131.820 ;
        RECT 56.355 131.775 56.645 132.005 ;
        RECT 71.520 131.960 71.840 132.020 ;
        RECT 71.995 131.960 72.285 132.005 ;
        RECT 56.890 131.820 64.850 131.960 ;
        RECT 46.770 131.480 49.670 131.620 ;
        RECT 50.910 131.620 51.050 131.760 ;
        RECT 56.430 131.620 56.570 131.775 ;
        RECT 50.910 131.480 56.570 131.620 ;
        RECT 30.580 131.280 30.900 131.340 ;
        RECT 36.190 131.280 36.330 131.435 ;
        RECT 26.530 131.140 30.900 131.280 ;
        RECT 30.580 131.080 30.900 131.140 ;
        RECT 33.890 131.140 36.330 131.280 ;
        RECT 36.600 131.280 36.890 131.325 ;
        RECT 38.700 131.280 38.990 131.325 ;
        RECT 40.270 131.280 40.560 131.325 ;
        RECT 36.600 131.140 40.560 131.280 ;
        RECT 33.890 131.000 34.030 131.140 ;
        RECT 36.600 131.095 36.890 131.140 ;
        RECT 38.700 131.095 38.990 131.140 ;
        RECT 40.270 131.095 40.560 131.140 ;
        RECT 43.015 131.280 43.305 131.325 ;
        RECT 46.310 131.280 46.450 131.435 ;
        RECT 43.015 131.140 46.450 131.280 ;
        RECT 48.520 131.280 48.840 131.340 ;
        RECT 50.835 131.280 51.125 131.325 ;
        RECT 56.890 131.280 57.030 131.820 ;
        RECT 57.260 131.420 57.580 131.680 ;
        RECT 61.860 131.620 62.180 131.680 ;
        RECT 64.175 131.620 64.465 131.665 ;
        RECT 61.860 131.480 64.465 131.620 ;
        RECT 61.860 131.420 62.180 131.480 ;
        RECT 64.175 131.435 64.465 131.480 ;
        RECT 61.415 131.280 61.705 131.325 ;
        RECT 48.520 131.140 57.030 131.280 ;
        RECT 60.110 131.140 61.705 131.280 ;
        RECT 43.015 131.095 43.305 131.140 ;
        RECT 24.615 130.940 24.905 130.985 ;
        RECT 25.520 130.940 25.840 131.000 ;
        RECT 24.615 130.800 25.840 130.940 ;
        RECT 24.615 130.755 24.905 130.800 ;
        RECT 25.520 130.740 25.840 130.800 ;
        RECT 27.820 130.940 28.140 131.000 ;
        RECT 31.500 130.940 31.820 131.000 ;
        RECT 27.820 130.800 31.820 130.940 ;
        RECT 27.820 130.740 28.140 130.800 ;
        RECT 31.500 130.740 31.820 130.800 ;
        RECT 31.960 130.740 32.280 131.000 ;
        RECT 33.800 130.740 34.120 131.000 ;
        RECT 40.700 130.940 41.020 131.000 ;
        RECT 43.090 130.940 43.230 131.095 ;
        RECT 48.520 131.080 48.840 131.140 ;
        RECT 50.835 131.095 51.125 131.140 ;
        RECT 40.700 130.800 43.230 130.940 ;
        RECT 40.700 130.740 41.020 130.800 ;
        RECT 43.460 130.740 43.780 131.000 ;
        RECT 47.600 130.740 47.920 131.000 ;
        RECT 60.110 130.985 60.250 131.140 ;
        RECT 61.415 131.095 61.705 131.140 ;
        RECT 60.035 130.755 60.325 130.985 ;
        RECT 60.955 130.940 61.245 130.985 ;
        RECT 63.240 130.940 63.560 131.000 ;
        RECT 60.955 130.800 63.560 130.940 ;
        RECT 64.710 130.940 64.850 131.820 ;
        RECT 71.520 131.820 72.285 131.960 ;
        RECT 71.520 131.760 71.840 131.820 ;
        RECT 71.995 131.775 72.285 131.820 ;
        RECT 73.375 131.960 73.665 132.005 ;
        RECT 74.370 131.960 74.510 132.440 ;
        RECT 87.620 132.300 87.940 132.360 ;
        RECT 87.620 132.160 92.450 132.300 ;
        RECT 87.620 132.100 87.940 132.160 ;
        RECT 76.120 132.005 76.440 132.020 ;
        RECT 76.090 131.960 76.440 132.005 ;
        RECT 73.375 131.820 74.510 131.960 ;
        RECT 75.925 131.820 76.440 131.960 ;
        RECT 73.375 131.775 73.665 131.820 ;
        RECT 76.090 131.775 76.440 131.820 ;
        RECT 67.405 131.620 67.695 131.665 ;
        RECT 69.925 131.620 70.215 131.665 ;
        RECT 71.115 131.620 71.405 131.665 ;
        RECT 67.405 131.480 71.405 131.620 ;
        RECT 72.070 131.620 72.210 131.775 ;
        RECT 76.120 131.760 76.440 131.775 ;
        RECT 82.100 131.760 82.420 132.020 ;
        RECT 83.480 132.005 83.800 132.020 ;
        RECT 83.450 131.775 83.800 132.005 ;
        RECT 83.480 131.760 83.800 131.775 ;
        RECT 84.860 131.960 85.180 132.020 ;
        RECT 91.300 131.960 91.620 132.020 ;
        RECT 84.860 131.820 91.620 131.960 ;
        RECT 84.860 131.760 85.180 131.820 ;
        RECT 91.300 131.760 91.620 131.820 ;
        RECT 74.755 131.620 75.045 131.665 ;
        RECT 72.070 131.480 75.045 131.620 ;
        RECT 67.405 131.435 67.695 131.480 ;
        RECT 69.925 131.435 70.215 131.480 ;
        RECT 71.115 131.435 71.405 131.480 ;
        RECT 74.755 131.435 75.045 131.480 ;
        RECT 75.635 131.620 75.925 131.665 ;
        RECT 76.825 131.620 77.115 131.665 ;
        RECT 79.345 131.620 79.635 131.665 ;
        RECT 75.635 131.480 79.635 131.620 ;
        RECT 75.635 131.435 75.925 131.480 ;
        RECT 76.825 131.435 77.115 131.480 ;
        RECT 79.345 131.435 79.635 131.480 ;
        RECT 82.995 131.620 83.285 131.665 ;
        RECT 84.185 131.620 84.475 131.665 ;
        RECT 86.705 131.620 86.995 131.665 ;
        RECT 82.995 131.480 86.995 131.620 ;
        RECT 82.995 131.435 83.285 131.480 ;
        RECT 84.185 131.435 84.475 131.480 ;
        RECT 86.705 131.435 86.995 131.480 ;
        RECT 89.000 131.620 89.320 131.680 ;
        RECT 92.310 131.665 92.450 132.160 ;
        RECT 97.280 132.100 97.600 132.360 ;
        RECT 99.135 132.300 99.425 132.345 ;
        RECT 106.080 132.300 106.370 132.345 ;
        RECT 99.135 132.160 106.370 132.300 ;
        RECT 108.410 132.300 108.550 132.440 ;
        RECT 109.100 132.300 109.390 132.345 ;
        RECT 108.410 132.160 109.390 132.300 ;
        RECT 99.135 132.115 99.425 132.160 ;
        RECT 106.080 132.115 106.370 132.160 ;
        RECT 109.100 132.115 109.390 132.160 ;
        RECT 113.840 132.100 114.160 132.360 ;
        RECT 114.850 132.300 114.990 132.455 ;
        RECT 126.260 132.440 126.580 132.500 ;
        RECT 134.095 132.640 134.385 132.685 ;
        RECT 135.935 132.640 136.225 132.685 ;
        RECT 136.380 132.640 136.700 132.700 ;
        RECT 134.095 132.500 135.230 132.640 ;
        RECT 134.095 132.455 134.385 132.500 ;
        RECT 130.875 132.300 131.165 132.345 ;
        RECT 135.090 132.300 135.230 132.500 ;
        RECT 135.935 132.500 136.700 132.640 ;
        RECT 135.935 132.455 136.225 132.500 ;
        RECT 136.380 132.440 136.700 132.500 ;
        RECT 137.850 132.500 143.050 132.640 ;
        RECT 137.850 132.300 137.990 132.500 ;
        RECT 142.910 132.360 143.050 132.500 ;
        RECT 140.075 132.300 140.365 132.345 ;
        RECT 140.520 132.300 140.840 132.360 ;
        RECT 114.850 132.160 119.590 132.300 ;
        RECT 95.900 131.760 96.220 132.020 ;
        RECT 97.370 131.960 97.510 132.100 ;
        RECT 98.675 131.960 98.965 132.005 ;
        RECT 97.370 131.820 98.965 131.960 ;
        RECT 98.675 131.775 98.965 131.820 ;
        RECT 99.595 131.960 99.885 132.005 ;
        RECT 113.930 131.960 114.070 132.100 ;
        RECT 99.595 131.820 114.070 131.960 ;
        RECT 116.615 131.960 116.905 132.005 ;
        RECT 117.980 131.960 118.300 132.020 ;
        RECT 119.450 132.005 119.590 132.160 ;
        RECT 130.875 132.160 134.770 132.300 ;
        RECT 135.090 132.160 137.990 132.300 ;
        RECT 130.875 132.115 131.165 132.160 ;
        RECT 116.615 131.820 118.300 131.960 ;
        RECT 99.595 131.775 99.885 131.820 ;
        RECT 116.615 131.775 116.905 131.820 ;
        RECT 91.775 131.620 92.065 131.665 ;
        RECT 89.000 131.480 92.065 131.620 ;
        RECT 89.000 131.420 89.320 131.480 ;
        RECT 91.775 131.435 92.065 131.480 ;
        RECT 92.235 131.435 92.525 131.665 ;
        RECT 97.295 131.620 97.585 131.665 ;
        RECT 97.740 131.620 98.060 131.680 ;
        RECT 97.295 131.480 98.060 131.620 ;
        RECT 97.295 131.435 97.585 131.480 ;
        RECT 97.740 131.420 98.060 131.480 ;
        RECT 67.840 131.280 68.130 131.325 ;
        RECT 69.410 131.280 69.700 131.325 ;
        RECT 71.510 131.280 71.800 131.325 ;
        RECT 67.840 131.140 71.800 131.280 ;
        RECT 67.840 131.095 68.130 131.140 ;
        RECT 69.410 131.095 69.700 131.140 ;
        RECT 71.510 131.095 71.800 131.140 ;
        RECT 75.240 131.280 75.530 131.325 ;
        RECT 77.340 131.280 77.630 131.325 ;
        RECT 78.910 131.280 79.200 131.325 ;
        RECT 82.600 131.280 82.890 131.325 ;
        RECT 84.700 131.280 84.990 131.325 ;
        RECT 86.270 131.280 86.560 131.325 ;
        RECT 99.670 131.280 99.810 131.775 ;
        RECT 117.980 131.760 118.300 131.820 ;
        RECT 119.375 131.775 119.665 132.005 ;
        RECT 123.515 131.960 123.805 132.005 ;
        RECT 124.880 131.960 125.200 132.020 ;
        RECT 123.515 131.820 125.200 131.960 ;
        RECT 123.515 131.775 123.805 131.820 ;
        RECT 124.880 131.760 125.200 131.820 ;
        RECT 130.415 131.775 130.705 132.005 ;
        RECT 131.335 131.960 131.625 132.005 ;
        RECT 133.160 131.960 133.480 132.020 ;
        RECT 134.110 131.960 134.400 132.005 ;
        RECT 131.335 131.820 132.010 131.960 ;
        RECT 131.335 131.775 131.625 131.820 ;
        RECT 102.825 131.620 103.115 131.665 ;
        RECT 105.345 131.620 105.635 131.665 ;
        RECT 106.535 131.620 106.825 131.665 ;
        RECT 102.825 131.480 106.825 131.620 ;
        RECT 102.825 131.435 103.115 131.480 ;
        RECT 105.345 131.435 105.635 131.480 ;
        RECT 106.535 131.435 106.825 131.480 ;
        RECT 107.415 131.620 107.705 131.665 ;
        RECT 107.860 131.620 108.180 131.680 ;
        RECT 107.415 131.480 108.180 131.620 ;
        RECT 107.415 131.435 107.705 131.480 ;
        RECT 107.860 131.420 108.180 131.480 ;
        RECT 108.755 131.620 109.045 131.665 ;
        RECT 109.945 131.620 110.235 131.665 ;
        RECT 112.465 131.620 112.755 131.665 ;
        RECT 108.755 131.480 112.755 131.620 ;
        RECT 108.755 131.435 109.045 131.480 ;
        RECT 109.945 131.435 110.235 131.480 ;
        RECT 112.465 131.435 112.755 131.480 ;
        RECT 117.060 131.420 117.380 131.680 ;
        RECT 121.200 131.620 121.520 131.680 ;
        RECT 126.275 131.620 126.565 131.665 ;
        RECT 121.200 131.480 126.565 131.620 ;
        RECT 121.200 131.420 121.520 131.480 ;
        RECT 126.275 131.435 126.565 131.480 ;
        RECT 75.240 131.140 79.200 131.280 ;
        RECT 75.240 131.095 75.530 131.140 ;
        RECT 77.340 131.095 77.630 131.140 ;
        RECT 78.910 131.095 79.200 131.140 ;
        RECT 79.430 131.140 82.330 131.280 ;
        RECT 79.430 130.940 79.570 131.140 ;
        RECT 64.710 130.800 79.570 130.940 ;
        RECT 60.955 130.755 61.245 130.800 ;
        RECT 63.240 130.740 63.560 130.800 ;
        RECT 81.640 130.740 81.960 131.000 ;
        RECT 82.190 130.940 82.330 131.140 ;
        RECT 82.600 131.140 86.560 131.280 ;
        RECT 82.600 131.095 82.890 131.140 ;
        RECT 84.700 131.095 84.990 131.140 ;
        RECT 86.270 131.095 86.560 131.140 ;
        RECT 86.790 131.140 99.810 131.280 ;
        RECT 103.260 131.280 103.550 131.325 ;
        RECT 104.830 131.280 105.120 131.325 ;
        RECT 106.930 131.280 107.220 131.325 ;
        RECT 103.260 131.140 107.220 131.280 ;
        RECT 86.790 130.940 86.930 131.140 ;
        RECT 103.260 131.095 103.550 131.140 ;
        RECT 104.830 131.095 105.120 131.140 ;
        RECT 106.930 131.095 107.220 131.140 ;
        RECT 108.360 131.280 108.650 131.325 ;
        RECT 110.460 131.280 110.750 131.325 ;
        RECT 112.030 131.280 112.320 131.325 ;
        RECT 108.360 131.140 112.320 131.280 ;
        RECT 108.360 131.095 108.650 131.140 ;
        RECT 110.460 131.095 110.750 131.140 ;
        RECT 112.030 131.095 112.320 131.140 ;
        RECT 116.600 131.080 116.920 131.340 ;
        RECT 130.490 131.280 130.630 131.775 ;
        RECT 131.870 131.665 132.010 131.820 ;
        RECT 133.160 131.820 134.400 131.960 ;
        RECT 134.630 131.960 134.770 132.160 ;
        RECT 135.935 131.960 136.225 132.005 ;
        RECT 137.300 131.960 137.620 132.020 ;
        RECT 137.850 132.005 137.990 132.160 ;
        RECT 138.310 132.160 139.830 132.300 ;
        RECT 138.310 132.005 138.450 132.160 ;
        RECT 134.630 131.820 137.620 131.960 ;
        RECT 133.160 131.760 133.480 131.820 ;
        RECT 134.110 131.775 134.400 131.820 ;
        RECT 135.935 131.775 136.225 131.820 ;
        RECT 137.300 131.760 137.620 131.820 ;
        RECT 137.775 131.775 138.065 132.005 ;
        RECT 138.235 131.775 138.525 132.005 ;
        RECT 138.680 131.760 139.000 132.020 ;
        RECT 139.155 131.775 139.445 132.005 ;
        RECT 139.690 131.960 139.830 132.160 ;
        RECT 140.075 132.160 140.840 132.300 ;
        RECT 140.075 132.115 140.365 132.160 ;
        RECT 140.520 132.100 140.840 132.160 ;
        RECT 141.440 132.300 141.760 132.360 ;
        RECT 141.915 132.300 142.205 132.345 ;
        RECT 141.440 132.160 142.205 132.300 ;
        RECT 141.440 132.100 141.760 132.160 ;
        RECT 141.915 132.115 142.205 132.160 ;
        RECT 142.820 132.100 143.140 132.360 ;
        RECT 142.360 131.960 142.680 132.020 ;
        RECT 139.690 131.820 142.680 131.960 ;
        RECT 131.795 131.620 132.085 131.665 ;
        RECT 134.540 131.620 134.860 131.680 ;
        RECT 136.380 131.620 136.700 131.680 ;
        RECT 131.795 131.480 134.860 131.620 ;
        RECT 131.795 131.435 132.085 131.480 ;
        RECT 134.540 131.420 134.860 131.480 ;
        RECT 135.090 131.480 136.700 131.620 ;
        RECT 131.320 131.280 131.640 131.340 ;
        RECT 132.255 131.280 132.545 131.325 ;
        RECT 130.490 131.140 132.545 131.280 ;
        RECT 131.320 131.080 131.640 131.140 ;
        RECT 132.255 131.095 132.545 131.140 ;
        RECT 82.190 130.800 86.930 130.940 ;
        RECT 87.160 130.940 87.480 131.000 ;
        RECT 89.015 130.940 89.305 130.985 ;
        RECT 87.160 130.800 89.305 130.940 ;
        RECT 87.160 130.740 87.480 130.800 ;
        RECT 89.015 130.755 89.305 130.800 ;
        RECT 89.460 130.740 89.780 131.000 ;
        RECT 94.060 130.740 94.380 131.000 ;
        RECT 129.480 130.740 129.800 131.000 ;
        RECT 135.090 130.985 135.230 131.480 ;
        RECT 136.380 131.420 136.700 131.480 ;
        RECT 137.315 131.280 137.605 131.325 ;
        RECT 138.770 131.280 138.910 131.760 ;
        RECT 137.315 131.140 138.910 131.280 ;
        RECT 137.315 131.095 137.605 131.140 ;
        RECT 135.015 130.755 135.305 130.985 ;
        RECT 137.760 130.940 138.080 131.000 ;
        RECT 139.230 130.940 139.370 131.775 ;
        RECT 142.360 131.760 142.680 131.820 ;
        RECT 146.960 131.760 147.280 132.020 ;
        RECT 137.760 130.800 139.370 130.940 ;
        RECT 137.760 130.740 138.080 130.800 ;
        RECT 143.740 130.740 144.060 131.000 ;
        RECT 147.895 130.940 148.185 130.985 ;
        RECT 151.100 130.940 151.420 131.000 ;
        RECT 147.895 130.800 151.420 130.940 ;
        RECT 147.895 130.755 148.185 130.800 ;
        RECT 151.100 130.740 151.420 130.800 ;
        RECT 22.690 130.120 157.010 130.600 ;
        RECT 24.600 129.720 24.920 129.980 ;
        RECT 30.120 129.920 30.440 129.980 ;
        RECT 33.340 129.920 33.660 129.980 ;
        RECT 28.370 129.780 33.660 129.920 ;
        RECT 25.060 129.240 25.380 129.300 ;
        RECT 28.370 129.285 28.510 129.780 ;
        RECT 30.120 129.720 30.440 129.780 ;
        RECT 33.340 129.720 33.660 129.780 ;
        RECT 37.480 129.920 37.800 129.980 ;
        RECT 39.335 129.920 39.625 129.965 ;
        RECT 37.480 129.780 39.625 129.920 ;
        RECT 37.480 129.720 37.800 129.780 ;
        RECT 39.335 129.735 39.625 129.780 ;
        RECT 42.080 129.920 42.400 129.980 ;
        RECT 46.695 129.920 46.985 129.965 ;
        RECT 42.080 129.780 46.985 129.920 ;
        RECT 42.080 129.720 42.400 129.780 ;
        RECT 46.695 129.735 46.985 129.780 ;
        RECT 28.780 129.580 29.070 129.625 ;
        RECT 30.880 129.580 31.170 129.625 ;
        RECT 32.450 129.580 32.740 129.625 ;
        RECT 42.540 129.580 42.860 129.640 ;
        RECT 28.780 129.440 32.740 129.580 ;
        RECT 28.780 129.395 29.070 129.440 ;
        RECT 30.880 129.395 31.170 129.440 ;
        RECT 32.450 129.395 32.740 129.440 ;
        RECT 37.570 129.440 42.860 129.580 ;
        RECT 28.295 129.240 28.585 129.285 ;
        RECT 25.060 129.100 28.585 129.240 ;
        RECT 25.060 129.040 25.380 129.100 ;
        RECT 28.295 129.055 28.585 129.100 ;
        RECT 29.175 129.240 29.465 129.285 ;
        RECT 30.365 129.240 30.655 129.285 ;
        RECT 32.885 129.240 33.175 129.285 ;
        RECT 29.175 129.100 33.175 129.240 ;
        RECT 29.175 129.055 29.465 129.100 ;
        RECT 30.365 129.055 30.655 129.100 ;
        RECT 32.885 129.055 33.175 129.100 ;
        RECT 27.835 128.715 28.125 128.945 ;
        RECT 29.630 128.900 29.920 128.945 ;
        RECT 31.960 128.900 32.280 128.960 ;
        RECT 29.630 128.760 32.280 128.900 ;
        RECT 29.630 128.715 29.920 128.760 ;
        RECT 27.910 128.560 28.050 128.715 ;
        RECT 31.960 128.700 32.280 128.760 ;
        RECT 32.420 128.900 32.740 128.960 ;
        RECT 37.570 128.945 37.710 129.440 ;
        RECT 42.540 129.380 42.860 129.440 ;
        RECT 43.460 129.380 43.780 129.640 ;
        RECT 46.770 129.580 46.910 129.735 ;
        RECT 52.660 129.720 52.980 129.980 ;
        RECT 53.135 129.920 53.425 129.965 ;
        RECT 54.960 129.920 55.280 129.980 ;
        RECT 53.135 129.780 55.280 129.920 ;
        RECT 53.135 129.735 53.425 129.780 ;
        RECT 54.960 129.720 55.280 129.780 ;
        RECT 60.955 129.920 61.245 129.965 ;
        RECT 61.860 129.920 62.180 129.980 ;
        RECT 60.955 129.780 62.180 129.920 ;
        RECT 60.955 129.735 61.245 129.780 ;
        RECT 61.860 129.720 62.180 129.780 ;
        RECT 71.060 129.920 71.380 129.980 ;
        RECT 84.860 129.920 85.180 129.980 ;
        RECT 71.060 129.780 85.180 129.920 ;
        RECT 71.060 129.720 71.380 129.780 ;
        RECT 84.860 129.720 85.180 129.780 ;
        RECT 86.715 129.920 87.005 129.965 ;
        RECT 89.000 129.920 89.320 129.980 ;
        RECT 86.715 129.780 89.320 129.920 ;
        RECT 86.715 129.735 87.005 129.780 ;
        RECT 89.000 129.720 89.320 129.780 ;
        RECT 93.600 129.920 93.920 129.980 ;
        RECT 95.900 129.920 96.220 129.980 ;
        RECT 93.600 129.780 96.220 129.920 ;
        RECT 93.600 129.720 93.920 129.780 ;
        RECT 95.900 129.720 96.220 129.780 ;
        RECT 107.875 129.920 108.165 129.965 ;
        RECT 108.780 129.920 109.100 129.980 ;
        RECT 107.875 129.780 109.100 129.920 ;
        RECT 107.875 129.735 108.165 129.780 ;
        RECT 108.780 129.720 109.100 129.780 ;
        RECT 117.995 129.920 118.285 129.965 ;
        RECT 121.200 129.920 121.520 129.980 ;
        RECT 117.995 129.780 121.520 129.920 ;
        RECT 117.995 129.735 118.285 129.780 ;
        RECT 121.200 129.720 121.520 129.780 ;
        RECT 125.340 129.920 125.660 129.980 ;
        RECT 126.735 129.920 127.025 129.965 ;
        RECT 125.340 129.780 127.025 129.920 ;
        RECT 125.340 129.720 125.660 129.780 ;
        RECT 126.735 129.735 127.025 129.780 ;
        RECT 136.380 129.720 136.700 129.980 ;
        RECT 143.740 129.920 144.060 129.980 ;
        RECT 144.215 129.920 144.505 129.965 ;
        RECT 143.740 129.780 144.505 129.920 ;
        RECT 143.740 129.720 144.060 129.780 ;
        RECT 144.215 129.735 144.505 129.780 ;
        RECT 145.135 129.920 145.425 129.965 ;
        RECT 146.960 129.920 147.280 129.980 ;
        RECT 145.135 129.780 147.280 129.920 ;
        RECT 145.135 129.735 145.425 129.780 ;
        RECT 146.960 129.720 147.280 129.780 ;
        RECT 54.540 129.580 54.830 129.625 ;
        RECT 56.640 129.580 56.930 129.625 ;
        RECT 58.210 129.580 58.500 129.625 ;
        RECT 46.770 129.440 54.270 129.580 ;
        RECT 43.550 129.240 43.690 129.380 ;
        RECT 54.130 129.300 54.270 129.440 ;
        RECT 54.540 129.440 58.500 129.580 ;
        RECT 54.540 129.395 54.830 129.440 ;
        RECT 56.640 129.395 56.930 129.440 ;
        RECT 58.210 129.395 58.500 129.440 ;
        RECT 65.580 129.580 65.870 129.625 ;
        RECT 67.680 129.580 67.970 129.625 ;
        RECT 69.250 129.580 69.540 129.625 ;
        RECT 65.580 129.440 69.540 129.580 ;
        RECT 65.580 129.395 65.870 129.440 ;
        RECT 67.680 129.395 67.970 129.440 ;
        RECT 69.250 129.395 69.540 129.440 ;
        RECT 71.995 129.580 72.285 129.625 ;
        RECT 81.195 129.580 81.485 129.625 ;
        RECT 83.020 129.580 83.340 129.640 ;
        RECT 71.995 129.440 74.510 129.580 ;
        RECT 71.995 129.395 72.285 129.440 ;
        RECT 38.030 129.100 43.690 129.240 ;
        RECT 49.455 129.240 49.745 129.285 ;
        RECT 51.280 129.240 51.600 129.300 ;
        RECT 49.455 129.100 51.600 129.240 ;
        RECT 38.030 128.945 38.170 129.100 ;
        RECT 49.455 129.055 49.745 129.100 ;
        RECT 51.280 129.040 51.600 129.100 ;
        RECT 52.200 129.240 52.520 129.300 ;
        RECT 52.675 129.240 52.965 129.285 ;
        RECT 52.200 129.100 52.965 129.240 ;
        RECT 52.200 129.040 52.520 129.100 ;
        RECT 52.675 129.055 52.965 129.100 ;
        RECT 54.040 129.040 54.360 129.300 ;
        RECT 54.935 129.240 55.225 129.285 ;
        RECT 56.125 129.240 56.415 129.285 ;
        RECT 58.645 129.240 58.935 129.285 ;
        RECT 65.975 129.240 66.265 129.285 ;
        RECT 67.165 129.240 67.455 129.285 ;
        RECT 69.685 129.240 69.975 129.285 ;
        RECT 54.935 129.100 58.935 129.240 ;
        RECT 54.935 129.055 55.225 129.100 ;
        RECT 56.125 129.055 56.415 129.100 ;
        RECT 58.645 129.055 58.935 129.100 ;
        RECT 59.190 129.100 64.390 129.240 ;
        RECT 36.115 128.900 36.405 128.945 ;
        RECT 32.420 128.760 36.405 128.900 ;
        RECT 32.420 128.700 32.740 128.760 ;
        RECT 36.115 128.715 36.405 128.760 ;
        RECT 37.035 128.715 37.325 128.945 ;
        RECT 37.495 128.715 37.785 128.945 ;
        RECT 37.955 128.715 38.245 128.945 ;
        RECT 38.400 128.900 38.720 128.960 ;
        RECT 40.255 128.900 40.545 128.945 ;
        RECT 38.400 128.760 53.350 128.900 ;
        RECT 37.110 128.560 37.250 128.715 ;
        RECT 38.400 128.700 38.720 128.760 ;
        RECT 40.255 128.715 40.545 128.760 ;
        RECT 45.300 128.560 45.620 128.620 ;
        RECT 27.910 128.420 31.730 128.560 ;
        RECT 37.110 128.420 45.620 128.560 ;
        RECT 31.590 128.280 31.730 128.420 ;
        RECT 45.300 128.360 45.620 128.420 ;
        RECT 47.600 128.360 47.920 128.620 ;
        RECT 50.375 128.375 50.665 128.605 ;
        RECT 50.820 128.560 51.140 128.620 ;
        RECT 51.295 128.560 51.585 128.605 ;
        RECT 50.820 128.420 51.585 128.560 ;
        RECT 31.500 128.020 31.820 128.280 ;
        RECT 35.195 128.220 35.485 128.265 ;
        RECT 35.640 128.220 35.960 128.280 ;
        RECT 37.020 128.220 37.340 128.280 ;
        RECT 35.195 128.080 37.340 128.220 ;
        RECT 47.690 128.220 47.830 128.360 ;
        RECT 50.450 128.220 50.590 128.375 ;
        RECT 50.820 128.360 51.140 128.420 ;
        RECT 51.295 128.375 51.585 128.420 ;
        RECT 51.740 128.360 52.060 128.620 ;
        RECT 53.210 128.560 53.350 128.760 ;
        RECT 53.580 128.700 53.900 128.960 ;
        RECT 59.190 128.900 59.330 129.100 ;
        RECT 64.250 128.960 64.390 129.100 ;
        RECT 64.710 129.100 65.770 129.240 ;
        RECT 62.335 128.900 62.625 128.945 ;
        RECT 55.050 128.760 59.330 128.900 ;
        RECT 59.650 128.760 62.625 128.900 ;
        RECT 55.050 128.560 55.190 128.760 ;
        RECT 53.210 128.420 55.190 128.560 ;
        RECT 55.390 128.560 55.680 128.605 ;
        RECT 59.650 128.560 59.790 128.760 ;
        RECT 62.335 128.715 62.625 128.760 ;
        RECT 63.240 128.700 63.560 128.960 ;
        RECT 64.160 128.700 64.480 128.960 ;
        RECT 64.710 128.945 64.850 129.100 ;
        RECT 64.635 128.715 64.925 128.945 ;
        RECT 65.095 128.715 65.385 128.945 ;
        RECT 65.170 128.560 65.310 128.715 ;
        RECT 65.630 128.620 65.770 129.100 ;
        RECT 65.975 129.100 69.975 129.240 ;
        RECT 65.975 129.055 66.265 129.100 ;
        RECT 67.165 129.055 67.455 129.100 ;
        RECT 69.685 129.055 69.975 129.100 ;
        RECT 74.370 129.240 74.510 129.440 ;
        RECT 81.195 129.440 83.340 129.580 ;
        RECT 81.195 129.395 81.485 129.440 ;
        RECT 83.020 129.380 83.340 129.440 ;
        RECT 83.480 129.380 83.800 129.640 ;
        RECT 90.380 129.580 90.700 129.640 ;
        RECT 92.680 129.580 93.000 129.640 ;
        RECT 90.380 129.440 93.000 129.580 ;
        RECT 90.380 129.380 90.700 129.440 ;
        RECT 92.680 129.380 93.000 129.440 ;
        RECT 97.740 129.380 98.060 129.640 ;
        RECT 120.740 129.580 121.030 129.625 ;
        RECT 122.310 129.580 122.600 129.625 ;
        RECT 124.410 129.580 124.700 129.625 ;
        RECT 120.740 129.440 124.700 129.580 ;
        RECT 120.740 129.395 121.030 129.440 ;
        RECT 122.310 129.395 122.600 129.440 ;
        RECT 124.410 129.395 124.700 129.440 ;
        RECT 134.540 129.580 134.860 129.640 ;
        RECT 139.615 129.580 139.905 129.625 ;
        RECT 150.640 129.580 150.930 129.625 ;
        RECT 152.210 129.580 152.500 129.625 ;
        RECT 154.310 129.580 154.600 129.625 ;
        RECT 134.540 129.440 146.730 129.580 ;
        RECT 134.540 129.380 134.860 129.440 ;
        RECT 139.615 129.395 139.905 129.440 ;
        RECT 75.215 129.240 75.505 129.285 ;
        RECT 89.460 129.240 89.780 129.300 ;
        RECT 95.915 129.240 96.205 129.285 ;
        RECT 96.820 129.240 97.140 129.300 ;
        RECT 74.370 129.100 75.505 129.240 ;
        RECT 74.370 128.960 74.510 129.100 ;
        RECT 75.215 129.055 75.505 129.100 ;
        RECT 84.490 129.100 89.780 129.240 ;
        RECT 68.300 128.900 68.620 128.960 ;
        RECT 68.300 128.760 72.210 128.900 ;
        RECT 68.300 128.700 68.620 128.760 ;
        RECT 55.390 128.420 59.790 128.560 ;
        RECT 61.490 128.420 65.310 128.560 ;
        RECT 55.390 128.375 55.680 128.420 ;
        RECT 61.490 128.280 61.630 128.420 ;
        RECT 65.540 128.360 65.860 128.620 ;
        RECT 66.430 128.560 66.720 128.605 ;
        RECT 66.920 128.560 67.240 128.620 ;
        RECT 66.430 128.420 67.240 128.560 ;
        RECT 72.070 128.560 72.210 128.760 ;
        RECT 74.280 128.700 74.600 128.960 ;
        RECT 78.895 128.900 79.185 128.945 ;
        RECT 81.640 128.900 81.960 128.960 ;
        RECT 84.490 128.945 84.630 129.100 ;
        RECT 89.460 129.040 89.780 129.100 ;
        RECT 91.850 129.100 94.750 129.240 ;
        RECT 91.850 128.960 91.990 129.100 ;
        RECT 94.610 128.960 94.750 129.100 ;
        RECT 95.915 129.100 97.140 129.240 ;
        RECT 95.915 129.055 96.205 129.100 ;
        RECT 96.820 129.040 97.140 129.100 ;
        RECT 99.595 129.240 99.885 129.285 ;
        RECT 100.960 129.240 101.280 129.300 ;
        RECT 99.595 129.100 101.280 129.240 ;
        RECT 99.595 129.055 99.885 129.100 ;
        RECT 100.960 129.040 101.280 129.100 ;
        RECT 110.160 129.240 110.480 129.300 ;
        RECT 110.635 129.240 110.925 129.285 ;
        RECT 110.160 129.100 110.925 129.240 ;
        RECT 110.160 129.040 110.480 129.100 ;
        RECT 110.635 129.055 110.925 129.100 ;
        RECT 120.305 129.240 120.595 129.285 ;
        RECT 122.825 129.240 123.115 129.285 ;
        RECT 124.015 129.240 124.305 129.285 ;
        RECT 120.305 129.100 124.305 129.240 ;
        RECT 120.305 129.055 120.595 129.100 ;
        RECT 122.825 129.055 123.115 129.100 ;
        RECT 124.015 129.055 124.305 129.100 ;
        RECT 128.575 129.240 128.865 129.285 ;
        RECT 138.220 129.240 138.540 129.300 ;
        RECT 128.575 129.100 138.540 129.240 ;
        RECT 128.575 129.055 128.865 129.100 ;
        RECT 138.220 129.040 138.540 129.100 ;
        RECT 78.895 128.760 81.960 128.900 ;
        RECT 78.895 128.715 79.185 128.760 ;
        RECT 81.640 128.700 81.960 128.760 ;
        RECT 84.415 128.715 84.705 128.945 ;
        RECT 85.320 128.700 85.640 128.960 ;
        RECT 85.780 128.900 86.100 128.960 ;
        RECT 87.160 128.900 87.480 128.960 ;
        RECT 91.315 128.900 91.605 128.945 ;
        RECT 85.780 128.760 87.480 128.900 ;
        RECT 85.780 128.700 86.100 128.760 ;
        RECT 87.160 128.700 87.480 128.760 ;
        RECT 88.170 128.760 91.605 128.900 ;
        RECT 78.420 128.560 78.740 128.620 ;
        RECT 88.170 128.605 88.310 128.760 ;
        RECT 91.315 128.715 91.605 128.760 ;
        RECT 88.095 128.560 88.385 128.605 ;
        RECT 72.070 128.420 73.130 128.560 ;
        RECT 66.430 128.375 66.720 128.420 ;
        RECT 66.920 128.360 67.240 128.420 ;
        RECT 53.580 128.220 53.900 128.280 ;
        RECT 47.690 128.080 53.900 128.220 ;
        RECT 35.195 128.035 35.485 128.080 ;
        RECT 35.640 128.020 35.960 128.080 ;
        RECT 37.020 128.020 37.340 128.080 ;
        RECT 53.580 128.020 53.900 128.080 ;
        RECT 61.400 128.020 61.720 128.280 ;
        RECT 64.175 128.220 64.465 128.265 ;
        RECT 71.060 128.220 71.380 128.280 ;
        RECT 64.175 128.080 71.380 128.220 ;
        RECT 64.175 128.035 64.465 128.080 ;
        RECT 71.060 128.020 71.380 128.080 ;
        RECT 72.440 128.020 72.760 128.280 ;
        RECT 72.990 128.220 73.130 128.420 ;
        RECT 78.420 128.420 88.385 128.560 ;
        RECT 78.420 128.360 78.740 128.420 ;
        RECT 88.095 128.375 88.385 128.420 ;
        RECT 89.935 128.560 90.225 128.605 ;
        RECT 90.380 128.560 90.700 128.620 ;
        RECT 89.935 128.420 90.700 128.560 ;
        RECT 89.935 128.375 90.225 128.420 ;
        RECT 90.380 128.360 90.700 128.420 ;
        RECT 78.895 128.220 79.185 128.265 ;
        RECT 72.990 128.080 79.185 128.220 ;
        RECT 78.895 128.035 79.185 128.080 ;
        RECT 80.260 128.220 80.580 128.280 ;
        RECT 87.620 128.220 87.940 128.280 ;
        RECT 80.260 128.080 87.940 128.220 ;
        RECT 91.390 128.220 91.530 128.715 ;
        RECT 91.760 128.700 92.080 128.960 ;
        RECT 92.235 128.715 92.525 128.945 ;
        RECT 93.155 128.900 93.445 128.945 ;
        RECT 93.600 128.900 93.920 128.960 ;
        RECT 93.155 128.760 93.920 128.900 ;
        RECT 93.155 128.715 93.445 128.760 ;
        RECT 92.310 128.560 92.450 128.715 ;
        RECT 93.600 128.700 93.920 128.760 ;
        RECT 94.520 128.700 94.840 128.960 ;
        RECT 97.755 128.715 98.045 128.945 ;
        RECT 96.360 128.560 96.680 128.620 ;
        RECT 97.830 128.560 97.970 128.715 ;
        RECT 109.700 128.700 110.020 128.960 ;
        RECT 123.615 128.900 123.905 128.945 ;
        RECT 124.420 128.900 124.740 128.960 ;
        RECT 124.895 128.900 125.185 128.945 ;
        RECT 123.615 128.760 124.190 128.900 ;
        RECT 123.615 128.715 123.905 128.760 ;
        RECT 112.000 128.560 112.320 128.620 ;
        RECT 116.140 128.560 116.460 128.620 ;
        RECT 117.075 128.560 117.365 128.605 ;
        RECT 92.310 128.420 97.970 128.560 ;
        RECT 108.870 128.420 117.365 128.560 ;
        RECT 96.360 128.360 96.680 128.420 ;
        RECT 108.870 128.220 109.010 128.420 ;
        RECT 112.000 128.360 112.320 128.420 ;
        RECT 116.140 128.360 116.460 128.420 ;
        RECT 117.075 128.375 117.365 128.420 ;
        RECT 124.050 128.280 124.190 128.760 ;
        RECT 124.420 128.760 125.185 128.900 ;
        RECT 124.420 128.700 124.740 128.760 ;
        RECT 124.895 128.715 125.185 128.760 ;
        RECT 128.115 128.900 128.405 128.945 ;
        RECT 129.480 128.900 129.800 128.960 ;
        RECT 128.115 128.760 129.800 128.900 ;
        RECT 128.115 128.715 128.405 128.760 ;
        RECT 129.480 128.700 129.800 128.760 ;
        RECT 134.080 128.700 134.400 128.960 ;
        RECT 137.300 128.700 137.620 128.960 ;
        RECT 140.075 128.715 140.365 128.945 ;
        RECT 140.535 128.900 140.825 128.945 ;
        RECT 141.070 128.900 141.210 129.440 ;
        RECT 140.535 128.760 141.210 128.900 ;
        RECT 140.535 128.715 140.825 128.760 ;
        RECT 141.455 128.715 141.745 128.945 ;
        RECT 140.150 128.560 140.290 128.715 ;
        RECT 141.530 128.560 141.670 128.715 ;
        RECT 141.900 128.700 142.220 128.960 ;
        RECT 142.820 128.900 143.140 128.960 ;
        RECT 146.590 128.945 146.730 129.440 ;
        RECT 150.640 129.440 154.600 129.580 ;
        RECT 150.640 129.395 150.930 129.440 ;
        RECT 152.210 129.395 152.500 129.440 ;
        RECT 154.310 129.395 154.600 129.440 ;
        RECT 150.205 129.240 150.495 129.285 ;
        RECT 152.725 129.240 153.015 129.285 ;
        RECT 153.915 129.240 154.205 129.285 ;
        RECT 150.205 129.100 154.205 129.240 ;
        RECT 150.205 129.055 150.495 129.100 ;
        RECT 152.725 129.055 153.015 129.100 ;
        RECT 153.915 129.055 154.205 129.100 ;
        RECT 142.820 128.760 146.270 128.900 ;
        RECT 142.820 128.700 143.140 128.760 ;
        RECT 140.150 128.420 141.210 128.560 ;
        RECT 141.530 128.420 143.050 128.560 ;
        RECT 91.390 128.080 109.010 128.220 ;
        RECT 110.175 128.220 110.465 128.265 ;
        RECT 111.080 128.220 111.400 128.280 ;
        RECT 110.175 128.080 111.400 128.220 ;
        RECT 80.260 128.020 80.580 128.080 ;
        RECT 87.620 128.020 87.940 128.080 ;
        RECT 110.175 128.035 110.465 128.080 ;
        RECT 111.080 128.020 111.400 128.080 ;
        RECT 111.540 128.220 111.860 128.280 ;
        RECT 115.695 128.220 115.985 128.265 ;
        RECT 111.540 128.080 115.985 128.220 ;
        RECT 111.540 128.020 111.860 128.080 ;
        RECT 115.695 128.035 115.985 128.080 ;
        RECT 123.960 128.020 124.280 128.280 ;
        RECT 131.320 128.020 131.640 128.280 ;
        RECT 135.000 128.020 135.320 128.280 ;
        RECT 140.520 128.020 140.840 128.280 ;
        RECT 141.070 128.220 141.210 128.420 ;
        RECT 141.900 128.220 142.220 128.280 ;
        RECT 142.910 128.265 143.050 128.420 ;
        RECT 143.280 128.360 143.600 128.620 ;
        RECT 144.375 128.560 144.665 128.605 ;
        RECT 145.595 128.560 145.885 128.605 ;
        RECT 143.830 128.420 145.885 128.560 ;
        RECT 146.130 128.560 146.270 128.760 ;
        RECT 146.515 128.715 146.805 128.945 ;
        RECT 151.100 128.900 151.420 128.960 ;
        RECT 153.460 128.900 153.750 128.945 ;
        RECT 151.100 128.760 153.750 128.900 ;
        RECT 151.100 128.700 151.420 128.760 ;
        RECT 153.460 128.715 153.750 128.760 ;
        RECT 154.320 128.900 154.640 128.960 ;
        RECT 154.795 128.900 155.085 128.945 ;
        RECT 154.320 128.760 155.085 128.900 ;
        RECT 154.320 128.700 154.640 128.760 ;
        RECT 154.795 128.715 155.085 128.760 ;
        RECT 146.130 128.420 148.110 128.560 ;
        RECT 141.070 128.080 142.220 128.220 ;
        RECT 141.900 128.020 142.220 128.080 ;
        RECT 142.835 128.220 143.125 128.265 ;
        RECT 143.830 128.220 143.970 128.420 ;
        RECT 144.375 128.375 144.665 128.420 ;
        RECT 145.595 128.375 145.885 128.420 ;
        RECT 142.835 128.080 143.970 128.220 ;
        RECT 146.040 128.220 146.360 128.280 ;
        RECT 147.970 128.265 148.110 128.420 ;
        RECT 147.435 128.220 147.725 128.265 ;
        RECT 146.040 128.080 147.725 128.220 ;
        RECT 142.835 128.035 143.125 128.080 ;
        RECT 146.040 128.020 146.360 128.080 ;
        RECT 147.435 128.035 147.725 128.080 ;
        RECT 147.895 128.035 148.185 128.265 ;
        RECT 22.690 127.400 157.810 127.880 ;
        RECT 25.060 127.000 25.380 127.260 ;
        RECT 42.540 127.200 42.860 127.260 ;
        RECT 33.660 127.060 42.860 127.200 ;
        RECT 24.155 126.520 24.445 126.565 ;
        RECT 25.150 126.520 25.290 127.000 ;
        RECT 33.660 126.920 33.800 127.060 ;
        RECT 42.540 127.000 42.860 127.060 ;
        RECT 51.740 127.200 52.060 127.260 ;
        RECT 54.500 127.200 54.820 127.260 ;
        RECT 51.740 127.060 54.820 127.200 ;
        RECT 51.740 127.000 52.060 127.060 ;
        RECT 54.500 127.000 54.820 127.060 ;
        RECT 57.260 127.000 57.580 127.260 ;
        RECT 60.020 127.000 60.340 127.260 ;
        RECT 60.480 127.200 60.800 127.260 ;
        RECT 60.480 127.060 65.770 127.200 ;
        RECT 60.480 127.000 60.800 127.060 ;
        RECT 25.520 126.905 25.840 126.920 ;
        RECT 25.490 126.860 25.840 126.905 ;
        RECT 28.740 126.860 29.060 126.920 ;
        RECT 30.580 126.860 30.900 126.920 ;
        RECT 33.340 126.860 33.800 126.920 ;
        RECT 36.560 126.860 36.880 126.920 ;
        RECT 51.280 126.860 51.600 126.920 ;
        RECT 57.350 126.860 57.490 127.000 ;
        RECT 25.490 126.720 25.990 126.860 ;
        RECT 28.740 126.720 34.490 126.860 ;
        RECT 25.490 126.675 25.840 126.720 ;
        RECT 25.520 126.660 25.840 126.675 ;
        RECT 28.740 126.660 29.060 126.720 ;
        RECT 30.580 126.660 30.900 126.720 ;
        RECT 33.340 126.660 33.660 126.720 ;
        RECT 24.155 126.380 25.290 126.520 ;
        RECT 32.420 126.520 32.740 126.580 ;
        RECT 32.895 126.520 33.185 126.565 ;
        RECT 32.420 126.380 33.185 126.520 ;
        RECT 24.155 126.335 24.445 126.380 ;
        RECT 32.420 126.320 32.740 126.380 ;
        RECT 32.895 126.335 33.185 126.380 ;
        RECT 33.800 126.320 34.120 126.580 ;
        RECT 34.350 126.565 34.490 126.720 ;
        RECT 36.560 126.720 51.600 126.860 ;
        RECT 36.560 126.660 36.880 126.720 ;
        RECT 51.280 126.660 51.600 126.720 ;
        RECT 51.830 126.720 57.490 126.860 ;
        RECT 60.110 126.860 60.250 127.000 ;
        RECT 65.080 126.905 65.400 126.920 ;
        RECT 64.935 126.860 65.400 126.905 ;
        RECT 60.110 126.720 65.400 126.860 ;
        RECT 65.630 126.860 65.770 127.060 ;
        RECT 66.920 127.000 67.240 127.260 ;
        RECT 67.380 127.200 67.700 127.260 ;
        RECT 70.535 127.200 70.825 127.245 ;
        RECT 79.340 127.200 79.660 127.260 ;
        RECT 88.080 127.200 88.400 127.260 ;
        RECT 67.380 127.060 88.400 127.200 ;
        RECT 67.380 127.000 67.700 127.060 ;
        RECT 70.535 127.015 70.825 127.060 ;
        RECT 66.015 126.860 66.305 126.905 ;
        RECT 71.060 126.860 71.380 126.920 ;
        RECT 71.535 126.860 71.825 126.905 ;
        RECT 65.630 126.720 66.305 126.860 ;
        RECT 34.275 126.335 34.565 126.565 ;
        RECT 34.735 126.520 35.025 126.565 ;
        RECT 40.255 126.520 40.545 126.565 ;
        RECT 34.735 126.380 40.545 126.520 ;
        RECT 34.735 126.335 35.025 126.380 ;
        RECT 40.255 126.335 40.545 126.380 ;
        RECT 42.540 126.520 42.860 126.580 ;
        RECT 51.830 126.520 51.970 126.720 ;
        RECT 64.935 126.675 65.400 126.720 ;
        RECT 66.015 126.675 66.305 126.720 ;
        RECT 66.505 126.720 69.450 126.860 ;
        RECT 65.080 126.660 65.400 126.675 ;
        RECT 42.540 126.380 51.970 126.520 ;
        RECT 53.595 126.520 53.885 126.565 ;
        RECT 54.040 126.520 54.360 126.580 ;
        RECT 53.595 126.380 54.360 126.520 ;
        RECT 42.540 126.320 42.860 126.380 ;
        RECT 53.595 126.335 53.885 126.380 ;
        RECT 54.040 126.320 54.360 126.380 ;
        RECT 54.930 126.520 55.220 126.565 ;
        RECT 61.415 126.520 61.705 126.565 ;
        RECT 54.930 126.380 61.705 126.520 ;
        RECT 54.930 126.335 55.220 126.380 ;
        RECT 61.415 126.335 61.705 126.380 ;
        RECT 62.335 126.335 62.625 126.565 ;
        RECT 25.035 126.180 25.325 126.225 ;
        RECT 26.225 126.180 26.515 126.225 ;
        RECT 28.745 126.180 29.035 126.225 ;
        RECT 25.035 126.040 29.035 126.180 ;
        RECT 25.035 125.995 25.325 126.040 ;
        RECT 26.225 125.995 26.515 126.040 ;
        RECT 28.745 125.995 29.035 126.040 ;
        RECT 36.115 126.180 36.405 126.225 ;
        RECT 36.575 126.180 36.865 126.225 ;
        RECT 36.115 126.040 36.865 126.180 ;
        RECT 36.115 125.995 36.405 126.040 ;
        RECT 36.575 125.995 36.865 126.040 ;
        RECT 37.480 126.180 37.800 126.240 ;
        RECT 43.015 126.180 43.305 126.225 ;
        RECT 37.480 126.040 43.305 126.180 ;
        RECT 37.480 125.980 37.800 126.040 ;
        RECT 43.015 125.995 43.305 126.040 ;
        RECT 43.920 126.180 44.240 126.240 ;
        RECT 44.855 126.180 45.145 126.225 ;
        RECT 43.920 126.040 45.145 126.180 ;
        RECT 43.920 125.980 44.240 126.040 ;
        RECT 44.855 125.995 45.145 126.040 ;
        RECT 52.675 125.995 52.965 126.225 ;
        RECT 54.475 126.180 54.765 126.225 ;
        RECT 55.665 126.180 55.955 126.225 ;
        RECT 58.185 126.180 58.475 126.225 ;
        RECT 54.475 126.040 58.475 126.180 ;
        RECT 62.410 126.180 62.550 126.335 ;
        RECT 63.240 126.320 63.560 126.580 ;
        RECT 63.715 126.520 64.005 126.565 ;
        RECT 63.715 126.380 64.850 126.520 ;
        RECT 63.715 126.335 64.005 126.380 ;
        RECT 64.710 126.180 64.850 126.380 ;
        RECT 65.540 126.180 65.860 126.240 ;
        RECT 66.505 126.180 66.645 126.720 ;
        RECT 67.840 126.320 68.160 126.580 ;
        RECT 68.760 126.320 69.080 126.580 ;
        RECT 69.310 126.565 69.450 126.720 ;
        RECT 71.060 126.720 71.825 126.860 ;
        RECT 71.060 126.660 71.380 126.720 ;
        RECT 71.535 126.675 71.825 126.720 ;
        RECT 72.070 126.565 72.210 127.060 ;
        RECT 79.340 127.000 79.660 127.060 ;
        RECT 88.080 127.000 88.400 127.060 ;
        RECT 89.015 127.015 89.305 127.245 ;
        RECT 75.200 126.860 75.520 126.920 ;
        RECT 79.800 126.860 80.120 126.920 ;
        RECT 81.195 126.860 81.485 126.905 ;
        RECT 75.200 126.720 81.485 126.860 ;
        RECT 89.090 126.860 89.230 127.015 ;
        RECT 94.060 127.000 94.380 127.260 ;
        RECT 96.360 127.000 96.680 127.260 ;
        RECT 116.140 127.200 116.460 127.260 ;
        RECT 131.320 127.200 131.640 127.260 ;
        RECT 116.140 127.060 128.790 127.200 ;
        RECT 116.140 127.000 116.460 127.060 ;
        RECT 90.700 126.860 90.990 126.905 ;
        RECT 89.090 126.720 90.990 126.860 ;
        RECT 75.200 126.660 75.520 126.720 ;
        RECT 79.800 126.660 80.120 126.720 ;
        RECT 81.195 126.675 81.485 126.720 ;
        RECT 90.700 126.675 90.990 126.720 ;
        RECT 69.235 126.520 69.525 126.565 ;
        RECT 69.235 126.380 70.830 126.520 ;
        RECT 69.235 126.335 69.525 126.380 ;
        RECT 62.410 126.040 64.390 126.180 ;
        RECT 64.710 126.040 66.645 126.180 ;
        RECT 70.690 126.180 70.830 126.380 ;
        RECT 71.995 126.335 72.285 126.565 ;
        RECT 88.095 126.520 88.385 126.565 ;
        RECT 94.150 126.520 94.290 127.000 ;
        RECT 117.980 126.860 118.300 126.920 ;
        RECT 94.610 126.720 118.300 126.860 ;
        RECT 94.610 126.580 94.750 126.720 ;
        RECT 88.095 126.380 94.290 126.520 ;
        RECT 88.095 126.335 88.385 126.380 ;
        RECT 94.520 126.320 94.840 126.580 ;
        RECT 108.410 126.565 108.550 126.720 ;
        RECT 117.980 126.660 118.300 126.720 ;
        RECT 119.360 126.860 119.680 126.920 ;
        RECT 122.210 126.905 122.350 127.060 ;
        RECT 119.360 126.720 121.890 126.860 ;
        RECT 119.360 126.660 119.680 126.720 ;
        RECT 121.750 126.580 121.890 126.720 ;
        RECT 122.135 126.675 122.425 126.905 ;
        RECT 126.260 126.860 126.580 126.920 ;
        RECT 127.655 126.860 127.945 126.905 ;
        RECT 126.260 126.720 127.945 126.860 ;
        RECT 126.260 126.660 126.580 126.720 ;
        RECT 127.655 126.675 127.945 126.720 ;
        RECT 103.275 126.520 103.565 126.565 ;
        RECT 103.275 126.380 104.870 126.520 ;
        RECT 103.275 126.335 103.565 126.380 ;
        RECT 72.455 126.180 72.745 126.225 ;
        RECT 70.690 126.040 72.745 126.180 ;
        RECT 54.475 125.995 54.765 126.040 ;
        RECT 55.665 125.995 55.955 126.040 ;
        RECT 58.185 125.995 58.475 126.040 ;
        RECT 24.640 125.840 24.930 125.885 ;
        RECT 26.740 125.840 27.030 125.885 ;
        RECT 28.310 125.840 28.600 125.885 ;
        RECT 24.640 125.700 28.600 125.840 ;
        RECT 24.640 125.655 24.930 125.700 ;
        RECT 26.740 125.655 27.030 125.700 ;
        RECT 28.310 125.655 28.600 125.700 ;
        RECT 39.795 125.840 40.085 125.885 ;
        RECT 41.620 125.840 41.940 125.900 ;
        RECT 39.795 125.700 41.940 125.840 ;
        RECT 39.795 125.655 40.085 125.700 ;
        RECT 41.620 125.640 41.940 125.700 ;
        RECT 48.075 125.840 48.365 125.885 ;
        RECT 51.740 125.840 52.060 125.900 ;
        RECT 48.075 125.700 52.060 125.840 ;
        RECT 48.075 125.655 48.365 125.700 ;
        RECT 51.740 125.640 52.060 125.700 ;
        RECT 31.055 125.500 31.345 125.545 ;
        RECT 31.500 125.500 31.820 125.560 ;
        RECT 31.055 125.360 31.820 125.500 ;
        RECT 31.055 125.315 31.345 125.360 ;
        RECT 31.500 125.300 31.820 125.360 ;
        RECT 49.440 125.300 49.760 125.560 ;
        RECT 52.750 125.500 52.890 125.995 ;
        RECT 64.250 125.885 64.390 126.040 ;
        RECT 65.540 125.980 65.860 126.040 ;
        RECT 72.455 125.995 72.745 126.040 ;
        RECT 54.080 125.840 54.370 125.885 ;
        RECT 56.180 125.840 56.470 125.885 ;
        RECT 57.750 125.840 58.040 125.885 ;
        RECT 54.080 125.700 58.040 125.840 ;
        RECT 54.080 125.655 54.370 125.700 ;
        RECT 56.180 125.655 56.470 125.700 ;
        RECT 57.750 125.655 58.040 125.700 ;
        RECT 64.175 125.655 64.465 125.885 ;
        RECT 67.840 125.840 68.160 125.900 ;
        RECT 69.695 125.840 69.985 125.885 ;
        RECT 71.980 125.840 72.300 125.900 ;
        RECT 67.840 125.700 69.985 125.840 ;
        RECT 67.840 125.640 68.160 125.700 ;
        RECT 69.695 125.655 69.985 125.700 ;
        RECT 70.690 125.700 72.300 125.840 ;
        RECT 72.530 125.840 72.670 125.995 ;
        RECT 74.740 125.980 75.060 126.240 ;
        RECT 80.260 125.980 80.580 126.240 ;
        RECT 80.720 125.980 81.040 126.240 ;
        RECT 89.475 125.995 89.765 126.225 ;
        RECT 90.355 126.180 90.645 126.225 ;
        RECT 91.545 126.180 91.835 126.225 ;
        RECT 94.065 126.180 94.355 126.225 ;
        RECT 90.355 126.040 94.355 126.180 ;
        RECT 90.355 125.995 90.645 126.040 ;
        RECT 91.545 125.995 91.835 126.040 ;
        RECT 94.065 125.995 94.355 126.040 ;
        RECT 76.120 125.840 76.440 125.900 ;
        RECT 72.530 125.700 79.110 125.840 ;
        RECT 54.960 125.500 55.280 125.560 ;
        RECT 52.750 125.360 55.280 125.500 ;
        RECT 54.960 125.300 55.280 125.360 ;
        RECT 62.320 125.500 62.640 125.560 ;
        RECT 65.095 125.500 65.385 125.545 ;
        RECT 69.220 125.500 69.540 125.560 ;
        RECT 70.690 125.545 70.830 125.700 ;
        RECT 71.980 125.640 72.300 125.700 ;
        RECT 76.120 125.640 76.440 125.700 ;
        RECT 78.970 125.560 79.110 125.700 ;
        RECT 62.320 125.360 69.540 125.500 ;
        RECT 62.320 125.300 62.640 125.360 ;
        RECT 65.095 125.315 65.385 125.360 ;
        RECT 69.220 125.300 69.540 125.360 ;
        RECT 70.615 125.315 70.905 125.545 ;
        RECT 77.960 125.300 78.280 125.560 ;
        RECT 78.880 125.300 79.200 125.560 ;
        RECT 83.020 125.300 83.340 125.560 ;
        RECT 89.550 125.500 89.690 125.995 ;
        RECT 104.180 125.980 104.500 126.240 ;
        RECT 104.730 126.180 104.870 126.380 ;
        RECT 108.335 126.335 108.625 126.565 ;
        RECT 112.000 126.320 112.320 126.580 ;
        RECT 112.920 126.520 113.240 126.580 ;
        RECT 114.300 126.520 114.620 126.580 ;
        RECT 117.535 126.520 117.825 126.565 ;
        RECT 119.835 126.520 120.125 126.565 ;
        RECT 112.920 126.380 114.070 126.520 ;
        RECT 112.920 126.320 113.240 126.380 ;
        RECT 105.100 126.180 105.420 126.240 ;
        RECT 107.875 126.180 108.165 126.225 ;
        RECT 104.730 126.040 108.165 126.180 ;
        RECT 105.100 125.980 105.420 126.040 ;
        RECT 107.875 125.995 108.165 126.040 ;
        RECT 110.620 125.980 110.940 126.240 ;
        RECT 113.380 125.980 113.700 126.240 ;
        RECT 113.930 126.180 114.070 126.380 ;
        RECT 114.300 126.380 117.825 126.520 ;
        RECT 114.300 126.320 114.620 126.380 ;
        RECT 117.535 126.335 117.825 126.380 ;
        RECT 118.070 126.380 120.125 126.520 ;
        RECT 118.070 126.180 118.210 126.380 ;
        RECT 119.835 126.335 120.125 126.380 ;
        RECT 121.660 126.520 121.980 126.580 ;
        RECT 123.055 126.520 123.345 126.565 ;
        RECT 127.195 126.520 127.485 126.565 ;
        RECT 121.660 126.380 127.485 126.520 ;
        RECT 121.660 126.320 121.980 126.380 ;
        RECT 123.055 126.335 123.345 126.380 ;
        RECT 127.195 126.335 127.485 126.380 ;
        RECT 128.115 126.335 128.405 126.565 ;
        RECT 113.930 126.040 118.210 126.180 ;
        RECT 118.440 126.180 118.760 126.240 ;
        RECT 118.915 126.180 119.205 126.225 ;
        RECT 119.360 126.180 119.680 126.240 ;
        RECT 118.440 126.040 119.680 126.180 ;
        RECT 118.440 125.980 118.760 126.040 ;
        RECT 118.915 125.995 119.205 126.040 ;
        RECT 119.360 125.980 119.680 126.040 ;
        RECT 89.960 125.840 90.250 125.885 ;
        RECT 92.060 125.840 92.350 125.885 ;
        RECT 93.630 125.840 93.920 125.885 ;
        RECT 89.960 125.700 93.920 125.840 ;
        RECT 104.270 125.840 104.410 125.980 ;
        RECT 113.470 125.840 113.610 125.980 ;
        RECT 128.190 125.840 128.330 126.335 ;
        RECT 128.650 126.180 128.790 127.060 ;
        RECT 130.260 127.060 131.640 127.200 ;
        RECT 130.260 126.860 130.400 127.060 ;
        RECT 131.320 127.000 131.640 127.060 ;
        RECT 131.780 127.000 132.100 127.260 ;
        RECT 135.000 127.200 135.320 127.260 ;
        RECT 134.170 127.060 135.320 127.200 ;
        RECT 129.110 126.720 130.400 126.860 ;
        RECT 129.110 126.565 129.250 126.720 ;
        RECT 129.035 126.335 129.325 126.565 ;
        RECT 129.955 126.335 130.245 126.565 ;
        RECT 131.870 126.520 132.010 127.000 ;
        RECT 134.170 126.905 134.310 127.060 ;
        RECT 135.000 127.000 135.320 127.060 ;
        RECT 135.550 127.060 137.070 127.200 ;
        RECT 134.095 126.675 134.385 126.905 ;
        RECT 135.550 126.860 135.690 127.060 ;
        RECT 136.930 126.920 137.070 127.060 ;
        RECT 140.520 127.000 140.840 127.260 ;
        RECT 141.440 127.200 141.760 127.260 ;
        RECT 142.375 127.200 142.665 127.245 ;
        RECT 141.440 127.060 142.665 127.200 ;
        RECT 141.440 127.000 141.760 127.060 ;
        RECT 142.375 127.015 142.665 127.060 ;
        RECT 142.820 127.000 143.140 127.260 ;
        RECT 143.280 127.200 143.600 127.260 ;
        RECT 146.040 127.200 146.360 127.260 ;
        RECT 148.895 127.200 149.185 127.245 ;
        RECT 143.280 127.060 145.810 127.200 ;
        RECT 143.280 127.000 143.600 127.060 ;
        RECT 134.630 126.720 135.690 126.860 ;
        RECT 133.175 126.520 133.465 126.565 ;
        RECT 131.870 126.380 133.465 126.520 ;
        RECT 133.175 126.335 133.465 126.380 ;
        RECT 133.635 126.520 133.925 126.565 ;
        RECT 134.630 126.520 134.770 126.720 ;
        RECT 136.840 126.660 137.160 126.920 ;
        RECT 133.635 126.380 134.770 126.520 ;
        RECT 133.635 126.335 133.925 126.380 ;
        RECT 130.030 126.180 130.170 126.335 ;
        RECT 135.000 126.320 135.320 126.580 ;
        RECT 135.920 126.565 136.240 126.580 ;
        RECT 135.465 126.285 135.755 126.515 ;
        RECT 135.920 126.335 136.345 126.565 ;
        RECT 135.920 126.320 136.240 126.335 ;
        RECT 128.650 126.040 130.170 126.180 ;
        RECT 104.270 125.700 113.610 125.840 ;
        RECT 124.970 125.700 128.330 125.840 ;
        RECT 135.550 125.840 135.690 126.285 ;
        RECT 140.610 126.180 140.750 127.000 ;
        RECT 141.900 126.860 142.220 126.920 ;
        RECT 141.900 126.720 143.510 126.860 ;
        RECT 141.900 126.660 142.220 126.720 ;
        RECT 143.370 126.565 143.510 126.720 ;
        RECT 143.295 126.520 143.585 126.565 ;
        RECT 145.120 126.520 145.440 126.580 ;
        RECT 143.295 126.380 145.440 126.520 ;
        RECT 145.670 126.520 145.810 127.060 ;
        RECT 146.040 127.060 149.185 127.200 ;
        RECT 146.040 127.000 146.360 127.060 ;
        RECT 148.895 127.015 149.185 127.060 ;
        RECT 149.735 127.015 150.025 127.245 ;
        RECT 146.515 126.860 146.805 126.905 ;
        RECT 147.420 126.860 147.740 126.920 ;
        RECT 146.515 126.720 147.740 126.860 ;
        RECT 146.515 126.675 146.805 126.720 ;
        RECT 147.420 126.660 147.740 126.720 ;
        RECT 147.895 126.675 148.185 126.905 ;
        RECT 146.960 126.520 147.280 126.580 ;
        RECT 147.970 126.520 148.110 126.675 ;
        RECT 145.670 126.380 148.110 126.520 ;
        RECT 149.810 126.520 149.950 127.015 ;
        RECT 150.195 126.520 150.485 126.565 ;
        RECT 149.810 126.380 150.485 126.520 ;
        RECT 143.295 126.335 143.585 126.380 ;
        RECT 145.120 126.320 145.440 126.380 ;
        RECT 146.960 126.320 147.280 126.380 ;
        RECT 150.195 126.335 150.485 126.380 ;
        RECT 152.955 126.335 153.245 126.565 ;
        RECT 153.030 126.180 153.170 126.335 ;
        RECT 140.610 126.040 147.190 126.180 ;
        RECT 143.740 125.840 144.060 125.900 ;
        RECT 135.550 125.700 144.060 125.840 ;
        RECT 89.960 125.655 90.250 125.700 ;
        RECT 92.060 125.655 92.350 125.700 ;
        RECT 93.630 125.655 93.920 125.700 ;
        RECT 124.970 125.560 125.110 125.700 ;
        RECT 143.740 125.640 144.060 125.700 ;
        RECT 144.200 125.640 144.520 125.900 ;
        RECT 144.675 125.840 144.965 125.885 ;
        RECT 145.580 125.840 145.900 125.900 ;
        RECT 144.675 125.700 145.900 125.840 ;
        RECT 144.675 125.655 144.965 125.700 ;
        RECT 93.140 125.500 93.460 125.560 ;
        RECT 89.550 125.360 93.460 125.500 ;
        RECT 93.140 125.300 93.460 125.360 ;
        RECT 102.340 125.300 102.660 125.560 ;
        RECT 117.520 125.500 117.840 125.560 ;
        RECT 117.995 125.500 118.285 125.545 ;
        RECT 117.520 125.360 118.285 125.500 ;
        RECT 117.520 125.300 117.840 125.360 ;
        RECT 117.995 125.315 118.285 125.360 ;
        RECT 118.440 125.300 118.760 125.560 ;
        RECT 118.900 125.500 119.220 125.560 ;
        RECT 120.295 125.500 120.585 125.545 ;
        RECT 121.200 125.500 121.520 125.560 ;
        RECT 118.900 125.360 121.520 125.500 ;
        RECT 118.900 125.300 119.220 125.360 ;
        RECT 120.295 125.315 120.585 125.360 ;
        RECT 121.200 125.300 121.520 125.360 ;
        RECT 123.975 125.500 124.265 125.545 ;
        RECT 124.880 125.500 125.200 125.560 ;
        RECT 123.975 125.360 125.200 125.500 ;
        RECT 123.975 125.315 124.265 125.360 ;
        RECT 124.880 125.300 125.200 125.360 ;
        RECT 126.275 125.500 126.565 125.545 ;
        RECT 127.640 125.500 127.960 125.560 ;
        RECT 126.275 125.360 127.960 125.500 ;
        RECT 126.275 125.315 126.565 125.360 ;
        RECT 127.640 125.300 127.960 125.360 ;
        RECT 131.320 125.300 131.640 125.560 ;
        RECT 132.240 125.300 132.560 125.560 ;
        RECT 136.395 125.500 136.685 125.545 ;
        RECT 138.680 125.500 139.000 125.560 ;
        RECT 136.395 125.360 139.000 125.500 ;
        RECT 136.395 125.315 136.685 125.360 ;
        RECT 138.680 125.300 139.000 125.360 ;
        RECT 141.455 125.500 141.745 125.545 ;
        RECT 144.750 125.500 144.890 125.655 ;
        RECT 145.580 125.640 145.900 125.700 ;
        RECT 141.455 125.360 144.890 125.500 ;
        RECT 141.455 125.315 141.745 125.360 ;
        RECT 146.500 125.300 146.820 125.560 ;
        RECT 147.050 125.500 147.190 126.040 ;
        RECT 147.510 126.040 153.170 126.180 ;
        RECT 147.510 125.885 147.650 126.040 ;
        RECT 147.435 125.655 147.725 125.885 ;
        RECT 150.640 125.840 150.960 125.900 ;
        RECT 152.035 125.840 152.325 125.885 ;
        RECT 150.640 125.700 152.325 125.840 ;
        RECT 150.640 125.640 150.960 125.700 ;
        RECT 152.035 125.655 152.325 125.700 ;
        RECT 148.815 125.500 149.105 125.545 ;
        RECT 147.050 125.360 149.105 125.500 ;
        RECT 148.815 125.315 149.105 125.360 ;
        RECT 151.100 125.300 151.420 125.560 ;
        RECT 22.690 124.680 157.010 125.160 ;
        RECT 26.915 124.480 27.205 124.525 ;
        RECT 33.800 124.480 34.120 124.540 ;
        RECT 26.915 124.340 34.120 124.480 ;
        RECT 26.915 124.295 27.205 124.340 ;
        RECT 33.800 124.280 34.120 124.340 ;
        RECT 36.115 124.480 36.405 124.525 ;
        RECT 37.480 124.480 37.800 124.540 ;
        RECT 36.115 124.340 37.800 124.480 ;
        RECT 36.115 124.295 36.405 124.340 ;
        RECT 37.480 124.280 37.800 124.340 ;
        RECT 42.080 124.480 42.400 124.540 ;
        RECT 45.300 124.480 45.620 124.540 ;
        RECT 53.135 124.480 53.425 124.525 ;
        RECT 42.080 124.340 43.230 124.480 ;
        RECT 42.080 124.280 42.400 124.340 ;
        RECT 38.860 124.140 39.150 124.185 ;
        RECT 40.430 124.140 40.720 124.185 ;
        RECT 42.530 124.140 42.820 124.185 ;
        RECT 38.860 124.000 42.820 124.140 ;
        RECT 38.860 123.955 39.150 124.000 ;
        RECT 40.430 123.955 40.720 124.000 ;
        RECT 42.530 123.955 42.820 124.000 ;
        RECT 43.090 123.845 43.230 124.340 ;
        RECT 45.300 124.340 53.425 124.480 ;
        RECT 45.300 124.280 45.620 124.340 ;
        RECT 53.135 124.295 53.425 124.340 ;
        RECT 54.040 124.280 54.360 124.540 ;
        RECT 54.960 124.280 55.280 124.540 ;
        RECT 55.895 124.480 56.185 124.525 ;
        RECT 57.260 124.480 57.580 124.540 ;
        RECT 55.895 124.340 57.580 124.480 ;
        RECT 55.895 124.295 56.185 124.340 ;
        RECT 46.680 124.140 46.970 124.185 ;
        RECT 48.250 124.140 48.540 124.185 ;
        RECT 50.350 124.140 50.640 124.185 ;
        RECT 46.680 124.000 50.640 124.140 ;
        RECT 46.680 123.955 46.970 124.000 ;
        RECT 48.250 123.955 48.540 124.000 ;
        RECT 50.350 123.955 50.640 124.000 ;
        RECT 38.425 123.800 38.715 123.845 ;
        RECT 40.945 123.800 41.235 123.845 ;
        RECT 42.135 123.800 42.425 123.845 ;
        RECT 26.070 123.660 33.110 123.800 ;
        RECT 26.070 123.505 26.210 123.660 ;
        RECT 25.995 123.275 26.285 123.505 ;
        RECT 27.375 123.275 27.665 123.505 ;
        RECT 32.970 123.460 33.110 123.660 ;
        RECT 33.660 123.660 34.950 123.800 ;
        RECT 33.660 123.460 33.800 123.660 ;
        RECT 32.970 123.320 33.800 123.460 ;
        RECT 25.075 122.935 25.365 123.165 ;
        RECT 26.440 123.120 26.760 123.180 ;
        RECT 27.450 123.120 27.590 123.275 ;
        RECT 34.260 123.260 34.580 123.520 ;
        RECT 34.810 123.460 34.950 123.660 ;
        RECT 38.425 123.660 42.425 123.800 ;
        RECT 38.425 123.615 38.715 123.660 ;
        RECT 40.945 123.615 41.235 123.660 ;
        RECT 42.135 123.615 42.425 123.660 ;
        RECT 43.015 123.615 43.305 123.845 ;
        RECT 46.245 123.800 46.535 123.845 ;
        RECT 48.765 123.800 49.055 123.845 ;
        RECT 49.955 123.800 50.245 123.845 ;
        RECT 46.245 123.660 50.245 123.800 ;
        RECT 46.245 123.615 46.535 123.660 ;
        RECT 48.765 123.615 49.055 123.660 ;
        RECT 49.955 123.615 50.245 123.660 ;
        RECT 50.820 123.800 51.140 123.860 ;
        RECT 54.130 123.800 54.270 124.280 ;
        RECT 55.970 124.140 56.110 124.295 ;
        RECT 57.260 124.280 57.580 124.340 ;
        RECT 63.240 124.480 63.560 124.540 ;
        RECT 75.200 124.480 75.520 124.540 ;
        RECT 63.240 124.340 75.520 124.480 ;
        RECT 63.240 124.280 63.560 124.340 ;
        RECT 75.200 124.280 75.520 124.340 ;
        RECT 80.720 124.480 81.040 124.540 ;
        RECT 83.495 124.480 83.785 124.525 ;
        RECT 80.720 124.340 83.785 124.480 ;
        RECT 80.720 124.280 81.040 124.340 ;
        RECT 83.495 124.295 83.785 124.340 ;
        RECT 105.100 124.480 105.420 124.540 ;
        RECT 105.575 124.480 105.865 124.525 ;
        RECT 105.100 124.340 105.865 124.480 ;
        RECT 105.100 124.280 105.420 124.340 ;
        RECT 105.575 124.295 105.865 124.340 ;
        RECT 119.360 124.480 119.680 124.540 ;
        RECT 133.620 124.480 133.940 124.540 ;
        RECT 119.360 124.340 133.940 124.480 ;
        RECT 119.360 124.280 119.680 124.340 ;
        RECT 133.620 124.280 133.940 124.340 ;
        RECT 140.980 124.480 141.300 124.540 ;
        RECT 140.980 124.340 144.430 124.480 ;
        RECT 140.980 124.280 141.300 124.340 ;
        RECT 50.820 123.660 54.270 123.800 ;
        RECT 54.590 124.000 56.110 124.140 ;
        RECT 50.820 123.600 51.140 123.660 ;
        RECT 40.240 123.460 40.560 123.520 ;
        RECT 34.810 123.320 40.560 123.460 ;
        RECT 40.240 123.260 40.560 123.320 ;
        RECT 41.620 123.505 41.940 123.520 ;
        RECT 49.440 123.505 49.760 123.520 ;
        RECT 41.620 123.460 41.970 123.505 ;
        RECT 49.440 123.460 49.790 123.505 ;
        RECT 50.360 123.460 50.680 123.520 ;
        RECT 53.595 123.460 53.885 123.505 ;
        RECT 41.620 123.320 42.135 123.460 ;
        RECT 49.440 123.320 49.955 123.460 ;
        RECT 50.360 123.320 53.885 123.460 ;
        RECT 41.620 123.275 41.970 123.320 ;
        RECT 49.440 123.275 49.790 123.320 ;
        RECT 41.620 123.260 41.940 123.275 ;
        RECT 49.440 123.260 49.760 123.275 ;
        RECT 50.360 123.260 50.680 123.320 ;
        RECT 53.595 123.275 53.885 123.320 ;
        RECT 54.055 123.460 54.345 123.505 ;
        RECT 54.590 123.460 54.730 124.000 ;
        RECT 56.355 123.955 56.645 124.185 ;
        RECT 76.620 124.140 76.910 124.185 ;
        RECT 78.720 124.140 79.010 124.185 ;
        RECT 80.290 124.140 80.580 124.185 ;
        RECT 94.060 124.140 94.380 124.200 ;
        RECT 76.620 124.000 80.580 124.140 ;
        RECT 76.620 123.955 76.910 124.000 ;
        RECT 78.720 123.955 79.010 124.000 ;
        RECT 80.290 123.955 80.580 124.000 ;
        RECT 85.410 124.000 94.380 124.140 ;
        RECT 56.430 123.800 56.570 123.955 ;
        RECT 85.410 123.860 85.550 124.000 ;
        RECT 55.050 123.660 56.570 123.800 ;
        RECT 56.815 123.800 57.105 123.845 ;
        RECT 58.180 123.800 58.500 123.860 ;
        RECT 77.015 123.800 77.305 123.845 ;
        RECT 78.205 123.800 78.495 123.845 ;
        RECT 80.725 123.800 81.015 123.845 ;
        RECT 56.815 123.660 58.500 123.800 ;
        RECT 55.050 123.505 55.190 123.660 ;
        RECT 56.815 123.615 57.105 123.660 ;
        RECT 54.055 123.320 54.730 123.460 ;
        RECT 54.055 123.275 54.345 123.320 ;
        RECT 54.975 123.275 55.265 123.505 ;
        RECT 55.435 123.275 55.725 123.505 ;
        RECT 56.890 123.460 57.030 123.615 ;
        RECT 58.180 123.600 58.500 123.660 ;
        RECT 65.170 123.660 76.810 123.800 ;
        RECT 56.475 123.320 57.030 123.460 ;
        RECT 64.160 123.460 64.480 123.520 ;
        RECT 65.170 123.505 65.310 123.660 ;
        RECT 76.670 123.520 76.810 123.660 ;
        RECT 77.015 123.660 81.015 123.800 ;
        RECT 77.015 123.615 77.305 123.660 ;
        RECT 78.205 123.615 78.495 123.660 ;
        RECT 80.725 123.615 81.015 123.660 ;
        RECT 85.320 123.600 85.640 123.860 ;
        RECT 91.760 123.800 92.080 123.860 ;
        RECT 93.230 123.845 93.370 124.000 ;
        RECT 94.060 123.940 94.380 124.000 ;
        RECT 99.160 124.140 99.450 124.185 ;
        RECT 101.260 124.140 101.550 124.185 ;
        RECT 102.830 124.140 103.120 124.185 ;
        RECT 99.160 124.000 103.120 124.140 ;
        RECT 99.160 123.955 99.450 124.000 ;
        RECT 101.260 123.955 101.550 124.000 ;
        RECT 102.830 123.955 103.120 124.000 ;
        RECT 107.415 123.955 107.705 124.185 ;
        RECT 127.680 124.140 127.970 124.185 ;
        RECT 129.780 124.140 130.070 124.185 ;
        RECT 131.350 124.140 131.640 124.185 ;
        RECT 127.680 124.000 131.640 124.140 ;
        RECT 127.680 123.955 127.970 124.000 ;
        RECT 129.780 123.955 130.070 124.000 ;
        RECT 131.350 123.955 131.640 124.000 ;
        RECT 134.095 124.140 134.385 124.185 ;
        RECT 135.920 124.140 136.240 124.200 ;
        RECT 139.140 124.140 139.460 124.200 ;
        RECT 144.290 124.140 144.430 124.340 ;
        RECT 144.660 124.280 144.980 124.540 ;
        RECT 145.120 124.480 145.440 124.540 ;
        RECT 147.895 124.480 148.185 124.525 ;
        RECT 145.120 124.340 148.185 124.480 ;
        RECT 145.120 124.280 145.440 124.340 ;
        RECT 147.895 124.295 148.185 124.340 ;
        RECT 146.515 124.140 146.805 124.185 ;
        RECT 134.095 124.000 137.530 124.140 ;
        RECT 134.095 123.955 134.385 124.000 ;
        RECT 87.250 123.660 92.080 123.800 ;
        RECT 65.095 123.460 65.385 123.505 ;
        RECT 76.135 123.460 76.425 123.505 ;
        RECT 64.160 123.320 65.385 123.460 ;
        RECT 36.560 123.120 36.880 123.180 ;
        RECT 26.440 122.980 27.590 123.120 ;
        RECT 27.910 122.980 36.880 123.120 ;
        RECT 25.150 122.780 25.290 122.935 ;
        RECT 26.440 122.920 26.760 122.980 ;
        RECT 25.520 122.780 25.840 122.840 ;
        RECT 27.910 122.780 28.050 122.980 ;
        RECT 36.560 122.920 36.880 122.980 ;
        RECT 43.550 122.980 51.050 123.120 ;
        RECT 25.150 122.640 28.050 122.780 ;
        RECT 25.520 122.580 25.840 122.640 ;
        RECT 30.580 122.580 30.900 122.840 ;
        RECT 31.040 122.580 31.360 122.840 ;
        RECT 35.180 122.780 35.500 122.840 ;
        RECT 43.550 122.780 43.690 122.980 ;
        RECT 35.180 122.640 43.690 122.780 ;
        RECT 35.180 122.580 35.500 122.640 ;
        RECT 43.920 122.580 44.240 122.840 ;
        RECT 50.910 122.780 51.050 122.980 ;
        RECT 51.280 122.920 51.600 123.180 ;
        RECT 51.740 123.120 52.060 123.180 ;
        RECT 52.215 123.120 52.505 123.165 ;
        RECT 55.510 123.120 55.650 123.275 ;
        RECT 51.740 122.980 55.650 123.120 ;
        RECT 51.740 122.920 52.060 122.980 ;
        RECT 52.215 122.935 52.505 122.980 ;
        RECT 56.475 122.780 56.615 123.320 ;
        RECT 64.160 123.260 64.480 123.320 ;
        RECT 65.095 123.275 65.385 123.320 ;
        RECT 73.910 123.320 76.425 123.460 ;
        RECT 60.940 122.920 61.260 123.180 ;
        RECT 50.910 122.640 56.615 122.780 ;
        RECT 61.030 122.780 61.170 122.920 ;
        RECT 73.910 122.840 74.050 123.320 ;
        RECT 76.135 123.275 76.425 123.320 ;
        RECT 76.580 123.260 76.900 123.520 ;
        RECT 83.480 123.460 83.800 123.520 ;
        RECT 84.415 123.460 84.705 123.505 ;
        RECT 83.480 123.320 84.705 123.460 ;
        RECT 83.480 123.260 83.800 123.320 ;
        RECT 84.415 123.275 84.705 123.320 ;
        RECT 77.470 123.120 77.760 123.165 ;
        RECT 81.180 123.120 81.500 123.180 ;
        RECT 87.250 123.120 87.390 123.660 ;
        RECT 91.760 123.600 92.080 123.660 ;
        RECT 93.155 123.615 93.445 123.845 ;
        RECT 93.600 123.800 93.920 123.860 ;
        RECT 98.675 123.800 98.965 123.845 ;
        RECT 93.600 123.660 98.965 123.800 ;
        RECT 93.600 123.600 93.920 123.660 ;
        RECT 98.675 123.615 98.965 123.660 ;
        RECT 99.555 123.800 99.845 123.845 ;
        RECT 100.745 123.800 101.035 123.845 ;
        RECT 103.265 123.800 103.555 123.845 ;
        RECT 99.555 123.660 103.555 123.800 ;
        RECT 99.555 123.615 99.845 123.660 ;
        RECT 100.745 123.615 101.035 123.660 ;
        RECT 103.265 123.615 103.555 123.660 ;
        RECT 87.635 123.275 87.925 123.505 ;
        RECT 88.555 123.460 88.845 123.505 ;
        RECT 88.170 123.320 88.845 123.460 ;
        RECT 77.470 122.980 81.500 123.120 ;
        RECT 77.470 122.935 77.760 122.980 ;
        RECT 81.180 122.920 81.500 122.980 ;
        RECT 81.960 122.980 87.390 123.120 ;
        RECT 71.520 122.780 71.840 122.840 ;
        RECT 73.820 122.780 74.140 122.840 ;
        RECT 61.030 122.640 74.140 122.780 ;
        RECT 71.520 122.580 71.840 122.640 ;
        RECT 73.820 122.580 74.140 122.640 ;
        RECT 75.200 122.780 75.520 122.840 ;
        RECT 81.960 122.780 82.100 122.980 ;
        RECT 75.200 122.640 82.100 122.780 ;
        RECT 83.035 122.780 83.325 122.825 ;
        RECT 83.480 122.780 83.800 122.840 ;
        RECT 83.035 122.640 83.800 122.780 ;
        RECT 75.200 122.580 75.520 122.640 ;
        RECT 83.035 122.595 83.325 122.640 ;
        RECT 83.480 122.580 83.800 122.640 ;
        RECT 85.320 122.780 85.640 122.840 ;
        RECT 87.710 122.780 87.850 123.275 ;
        RECT 88.170 122.840 88.310 123.320 ;
        RECT 88.555 123.275 88.845 123.320 ;
        RECT 92.680 123.260 93.000 123.520 ;
        RECT 94.075 123.275 94.365 123.505 ;
        RECT 94.150 123.120 94.290 123.275 ;
        RECT 97.280 123.260 97.600 123.520 ;
        RECT 99.955 123.460 100.245 123.505 ;
        RECT 98.290 123.320 100.245 123.460 ;
        RECT 92.310 122.980 94.290 123.120 ;
        RECT 92.310 122.840 92.450 122.980 ;
        RECT 85.320 122.640 87.850 122.780 ;
        RECT 85.320 122.580 85.640 122.640 ;
        RECT 88.080 122.580 88.400 122.840 ;
        RECT 89.475 122.780 89.765 122.825 ;
        RECT 90.840 122.780 91.160 122.840 ;
        RECT 89.475 122.640 91.160 122.780 ;
        RECT 89.475 122.595 89.765 122.640 ;
        RECT 90.840 122.580 91.160 122.640 ;
        RECT 91.300 122.780 91.620 122.840 ;
        RECT 91.775 122.780 92.065 122.825 ;
        RECT 91.300 122.640 92.065 122.780 ;
        RECT 91.300 122.580 91.620 122.640 ;
        RECT 91.775 122.595 92.065 122.640 ;
        RECT 92.220 122.580 92.540 122.840 ;
        RECT 94.980 122.580 95.300 122.840 ;
        RECT 98.290 122.825 98.430 123.320 ;
        RECT 99.955 123.275 100.245 123.320 ;
        RECT 106.955 123.460 107.245 123.505 ;
        RECT 107.490 123.460 107.630 123.955 ;
        RECT 135.920 123.940 136.240 124.000 ;
        RECT 110.160 123.800 110.480 123.860 ;
        RECT 106.955 123.320 107.630 123.460 ;
        RECT 107.850 123.660 110.480 123.800 ;
        RECT 106.955 123.275 107.245 123.320 ;
        RECT 103.260 123.120 103.580 123.180 ;
        RECT 107.850 123.120 107.990 123.660 ;
        RECT 110.160 123.600 110.480 123.660 ;
        RECT 112.920 123.600 113.240 123.860 ;
        RECT 137.390 123.845 137.530 124.000 ;
        RECT 139.140 124.000 143.050 124.140 ;
        RECT 144.290 124.000 146.805 124.140 ;
        RECT 139.140 123.940 139.460 124.000 ;
        RECT 128.075 123.800 128.365 123.845 ;
        RECT 129.265 123.800 129.555 123.845 ;
        RECT 131.785 123.800 132.075 123.845 ;
        RECT 128.075 123.660 132.075 123.800 ;
        RECT 128.075 123.615 128.365 123.660 ;
        RECT 129.265 123.615 129.555 123.660 ;
        RECT 131.785 123.615 132.075 123.660 ;
        RECT 137.315 123.615 137.605 123.845 ;
        RECT 138.680 123.800 139.000 123.860 ;
        RECT 141.915 123.800 142.205 123.845 ;
        RECT 138.680 123.660 142.205 123.800 ;
        RECT 138.680 123.600 139.000 123.660 ;
        RECT 141.915 123.615 142.205 123.660 ;
        RECT 108.780 123.460 109.100 123.520 ;
        RECT 109.715 123.460 110.005 123.505 ;
        RECT 113.010 123.460 113.150 123.600 ;
        RECT 108.780 123.320 113.150 123.460 ;
        RECT 117.995 123.460 118.285 123.505 ;
        RECT 119.820 123.460 120.140 123.520 ;
        RECT 122.120 123.460 122.440 123.520 ;
        RECT 127.195 123.460 127.485 123.505 ;
        RECT 117.995 123.320 122.440 123.460 ;
        RECT 108.780 123.260 109.100 123.320 ;
        RECT 109.715 123.275 110.005 123.320 ;
        RECT 117.995 123.275 118.285 123.320 ;
        RECT 119.820 123.260 120.140 123.320 ;
        RECT 122.120 123.260 122.440 123.320 ;
        RECT 124.510 123.320 127.485 123.460 ;
        RECT 103.260 122.980 107.990 123.120 ;
        RECT 103.260 122.920 103.580 122.980 ;
        RECT 124.510 122.840 124.650 123.320 ;
        RECT 127.195 123.275 127.485 123.320 ;
        RECT 134.080 123.460 134.400 123.520 ;
        RECT 140.075 123.460 140.365 123.505 ;
        RECT 134.080 123.320 140.365 123.460 ;
        RECT 134.080 123.260 134.400 123.320 ;
        RECT 140.075 123.275 140.365 123.320 ;
        RECT 140.535 123.460 140.825 123.505 ;
        RECT 140.980 123.460 141.300 123.520 ;
        RECT 140.535 123.320 141.300 123.460 ;
        RECT 140.535 123.275 140.825 123.320 ;
        RECT 125.340 123.120 125.660 123.180 ;
        RECT 128.420 123.120 128.710 123.165 ;
        RECT 125.340 122.980 128.710 123.120 ;
        RECT 125.340 122.920 125.660 122.980 ;
        RECT 128.420 122.935 128.710 122.980 ;
        RECT 138.220 123.120 138.540 123.180 ;
        RECT 140.610 123.120 140.750 123.275 ;
        RECT 140.980 123.260 141.300 123.320 ;
        RECT 138.220 122.980 140.750 123.120 ;
        RECT 141.900 123.120 142.220 123.180 ;
        RECT 142.375 123.120 142.665 123.165 ;
        RECT 141.900 122.980 142.665 123.120 ;
        RECT 142.910 123.120 143.050 124.000 ;
        RECT 146.515 123.955 146.805 124.000 ;
        RECT 150.640 124.140 150.930 124.185 ;
        RECT 152.210 124.140 152.500 124.185 ;
        RECT 154.310 124.140 154.600 124.185 ;
        RECT 150.640 124.000 154.600 124.140 ;
        RECT 150.640 123.955 150.930 124.000 ;
        RECT 152.210 123.955 152.500 124.000 ;
        RECT 154.310 123.955 154.600 124.000 ;
        RECT 143.740 123.800 144.060 123.860 ;
        RECT 144.215 123.800 144.505 123.845 ;
        RECT 143.740 123.660 144.505 123.800 ;
        RECT 143.740 123.600 144.060 123.660 ;
        RECT 144.215 123.615 144.505 123.660 ;
        RECT 150.205 123.800 150.495 123.845 ;
        RECT 152.725 123.800 153.015 123.845 ;
        RECT 153.915 123.800 154.205 123.845 ;
        RECT 150.205 123.660 154.205 123.800 ;
        RECT 150.205 123.615 150.495 123.660 ;
        RECT 152.725 123.615 153.015 123.660 ;
        RECT 153.915 123.615 154.205 123.660 ;
        RECT 145.595 123.460 145.885 123.505 ;
        RECT 144.750 123.320 145.885 123.460 ;
        RECT 144.750 123.120 144.890 123.320 ;
        RECT 145.595 123.275 145.885 123.320 ;
        RECT 146.055 123.275 146.345 123.505 ;
        RECT 151.100 123.460 151.420 123.520 ;
        RECT 153.460 123.460 153.750 123.505 ;
        RECT 151.100 123.320 153.750 123.460 ;
        RECT 146.130 123.120 146.270 123.275 ;
        RECT 151.100 123.260 151.420 123.320 ;
        RECT 153.460 123.275 153.750 123.320 ;
        RECT 154.320 123.460 154.640 123.520 ;
        RECT 154.795 123.460 155.085 123.505 ;
        RECT 154.320 123.320 155.085 123.460 ;
        RECT 154.320 123.260 154.640 123.320 ;
        RECT 154.795 123.275 155.085 123.320 ;
        RECT 142.910 122.980 144.890 123.120 ;
        RECT 145.670 122.980 146.270 123.120 ;
        RECT 138.220 122.920 138.540 122.980 ;
        RECT 141.900 122.920 142.220 122.980 ;
        RECT 142.375 122.935 142.665 122.980 ;
        RECT 98.215 122.595 98.505 122.825 ;
        RECT 106.035 122.780 106.325 122.825 ;
        RECT 106.480 122.780 106.800 122.840 ;
        RECT 106.035 122.640 106.800 122.780 ;
        RECT 106.035 122.595 106.325 122.640 ;
        RECT 106.480 122.580 106.800 122.640 ;
        RECT 109.240 122.580 109.560 122.840 ;
        RECT 124.420 122.580 124.740 122.840 ;
        RECT 134.540 122.580 134.860 122.840 ;
        RECT 137.300 122.780 137.620 122.840 ;
        RECT 142.835 122.780 143.125 122.825 ;
        RECT 137.300 122.640 143.125 122.780 ;
        RECT 137.300 122.580 137.620 122.640 ;
        RECT 142.835 122.595 143.125 122.640 ;
        RECT 144.200 122.780 144.520 122.840 ;
        RECT 145.670 122.780 145.810 122.980 ;
        RECT 144.200 122.640 145.810 122.780 ;
        RECT 144.200 122.580 144.520 122.640 ;
        RECT 22.690 121.960 157.810 122.440 ;
        RECT 31.040 121.760 31.360 121.820 ;
        RECT 30.670 121.620 31.360 121.760 ;
        RECT 29.830 121.420 30.120 121.465 ;
        RECT 30.670 121.420 30.810 121.620 ;
        RECT 31.040 121.560 31.360 121.620 ;
        RECT 32.420 121.560 32.740 121.820 ;
        RECT 33.340 121.560 33.660 121.820 ;
        RECT 34.260 121.760 34.580 121.820 ;
        RECT 34.735 121.760 35.025 121.805 ;
        RECT 43.920 121.760 44.240 121.820 ;
        RECT 34.260 121.620 35.025 121.760 ;
        RECT 34.260 121.560 34.580 121.620 ;
        RECT 34.735 121.575 35.025 121.620 ;
        RECT 38.490 121.620 44.240 121.760 ;
        RECT 32.510 121.420 32.650 121.560 ;
        RECT 33.430 121.420 33.570 121.560 ;
        RECT 29.830 121.280 30.810 121.420 ;
        RECT 31.590 121.280 32.650 121.420 ;
        RECT 32.970 121.280 33.570 121.420 ;
        RECT 36.115 121.420 36.405 121.465 ;
        RECT 36.560 121.420 36.880 121.480 ;
        RECT 36.115 121.280 36.880 121.420 ;
        RECT 29.830 121.235 30.120 121.280 ;
        RECT 30.580 120.880 30.900 121.140 ;
        RECT 31.040 120.880 31.360 121.140 ;
        RECT 31.590 121.125 31.730 121.280 ;
        RECT 31.515 120.895 31.805 121.125 ;
        RECT 31.960 121.080 32.280 121.140 ;
        RECT 32.970 121.125 33.110 121.280 ;
        RECT 36.115 121.235 36.405 121.280 ;
        RECT 36.560 121.220 36.880 121.280 ;
        RECT 37.020 121.220 37.340 121.480 ;
        RECT 32.435 121.080 32.725 121.125 ;
        RECT 31.960 120.940 32.725 121.080 ;
        RECT 31.960 120.880 32.280 120.940 ;
        RECT 32.435 120.895 32.725 120.940 ;
        RECT 32.895 120.895 33.185 121.125 ;
        RECT 33.355 120.895 33.645 121.125 ;
        RECT 37.480 121.080 37.800 121.140 ;
        RECT 38.490 121.125 38.630 121.620 ;
        RECT 43.920 121.560 44.240 121.620 ;
        RECT 46.695 121.760 46.985 121.805 ;
        RECT 50.360 121.760 50.680 121.820 ;
        RECT 46.695 121.620 50.680 121.760 ;
        RECT 46.695 121.575 46.985 121.620 ;
        RECT 50.360 121.560 50.680 121.620 ;
        RECT 66.935 121.760 67.225 121.805 ;
        RECT 68.760 121.760 69.080 121.820 ;
        RECT 74.740 121.760 75.060 121.820 ;
        RECT 66.935 121.620 75.060 121.760 ;
        RECT 66.935 121.575 67.225 121.620 ;
        RECT 68.760 121.560 69.080 121.620 ;
        RECT 74.740 121.560 75.060 121.620 ;
        RECT 81.180 121.560 81.500 121.820 ;
        RECT 83.020 121.760 83.340 121.820 ;
        RECT 82.190 121.620 83.340 121.760 ;
        RECT 39.795 121.420 40.085 121.465 ;
        RECT 44.855 121.420 45.145 121.465 ;
        RECT 49.900 121.420 50.220 121.480 ;
        RECT 39.795 121.280 45.145 121.420 ;
        RECT 39.795 121.235 40.085 121.280 ;
        RECT 44.855 121.235 45.145 121.280 ;
        RECT 49.530 121.280 50.220 121.420 ;
        RECT 37.955 121.080 38.245 121.125 ;
        RECT 37.480 120.940 38.245 121.080 ;
        RECT 26.465 120.740 26.755 120.785 ;
        RECT 28.985 120.740 29.275 120.785 ;
        RECT 30.175 120.740 30.465 120.785 ;
        RECT 26.465 120.600 30.465 120.740 ;
        RECT 30.670 120.740 30.810 120.880 ;
        RECT 33.430 120.740 33.570 120.895 ;
        RECT 37.480 120.880 37.800 120.940 ;
        RECT 37.955 120.895 38.245 120.940 ;
        RECT 38.415 120.895 38.705 121.125 ;
        RECT 40.700 120.880 41.020 121.140 ;
        RECT 49.530 121.125 49.670 121.280 ;
        RECT 49.900 121.220 50.220 121.280 ;
        RECT 50.790 121.420 51.080 121.465 ;
        RECT 51.280 121.420 51.600 121.480 ;
        RECT 50.790 121.280 51.600 121.420 ;
        RECT 50.790 121.235 51.080 121.280 ;
        RECT 51.280 121.220 51.600 121.280 ;
        RECT 72.610 121.420 72.900 121.465 ;
        RECT 78.435 121.420 78.725 121.465 ;
        RECT 72.610 121.280 78.725 121.420 ;
        RECT 72.610 121.235 72.900 121.280 ;
        RECT 78.435 121.235 78.725 121.280 ;
        RECT 78.880 121.420 79.200 121.480 ;
        RECT 78.880 121.280 80.950 121.420 ;
        RECT 78.880 121.220 79.200 121.280 ;
        RECT 42.095 120.895 42.385 121.125 ;
        RECT 49.455 120.895 49.745 121.125 ;
        RECT 60.480 121.080 60.800 121.140 ;
        RECT 61.415 121.080 61.705 121.125 ;
        RECT 75.200 121.080 75.520 121.140 ;
        RECT 49.990 120.940 56.570 121.080 ;
        RECT 30.670 120.600 33.570 120.740 ;
        RECT 26.465 120.555 26.755 120.600 ;
        RECT 28.985 120.555 29.275 120.600 ;
        RECT 30.175 120.555 30.465 120.600 ;
        RECT 26.900 120.400 27.190 120.445 ;
        RECT 28.470 120.400 28.760 120.445 ;
        RECT 30.570 120.400 30.860 120.445 ;
        RECT 26.900 120.260 30.860 120.400 ;
        RECT 26.900 120.215 27.190 120.260 ;
        RECT 28.470 120.215 28.760 120.260 ;
        RECT 30.570 120.215 30.860 120.260 ;
        RECT 39.335 120.400 39.625 120.445 ;
        RECT 41.175 120.400 41.465 120.445 ;
        RECT 39.335 120.260 41.465 120.400 ;
        RECT 39.335 120.215 39.625 120.260 ;
        RECT 41.175 120.215 41.465 120.260 ;
        RECT 41.635 120.215 41.925 120.445 ;
        RECT 42.170 120.400 42.310 120.895 ;
        RECT 43.920 120.540 44.240 120.800 ;
        RECT 44.395 120.740 44.685 120.785 ;
        RECT 49.990 120.740 50.130 120.940 ;
        RECT 44.395 120.600 50.130 120.740 ;
        RECT 50.335 120.740 50.625 120.785 ;
        RECT 51.525 120.740 51.815 120.785 ;
        RECT 54.045 120.740 54.335 120.785 ;
        RECT 50.335 120.600 54.335 120.740 ;
        RECT 44.395 120.555 44.685 120.600 ;
        RECT 50.335 120.555 50.625 120.600 ;
        RECT 51.525 120.555 51.815 120.600 ;
        RECT 54.045 120.555 54.335 120.600 ;
        RECT 56.430 120.740 56.570 120.940 ;
        RECT 60.480 120.940 61.705 121.080 ;
        RECT 60.480 120.880 60.800 120.940 ;
        RECT 61.415 120.895 61.705 120.940 ;
        RECT 62.410 120.940 75.520 121.080 ;
        RECT 58.180 120.740 58.500 120.800 ;
        RECT 59.575 120.740 59.865 120.785 ;
        RECT 56.430 120.600 59.865 120.740 ;
        RECT 49.440 120.400 49.760 120.460 ;
        RECT 56.430 120.445 56.570 120.600 ;
        RECT 58.180 120.540 58.500 120.600 ;
        RECT 59.575 120.555 59.865 120.600 ;
        RECT 61.860 120.540 62.180 120.800 ;
        RECT 42.170 120.260 49.760 120.400 ;
        RECT 24.155 120.060 24.445 120.105 ;
        RECT 25.980 120.060 26.300 120.120 ;
        RECT 24.155 119.920 26.300 120.060 ;
        RECT 24.155 119.875 24.445 119.920 ;
        RECT 25.980 119.860 26.300 119.920 ;
        RECT 35.640 119.860 35.960 120.120 ;
        RECT 38.415 120.060 38.705 120.105 ;
        RECT 40.240 120.060 40.560 120.120 ;
        RECT 38.415 119.920 40.560 120.060 ;
        RECT 41.710 120.060 41.850 120.215 ;
        RECT 49.440 120.200 49.760 120.260 ;
        RECT 49.940 120.400 50.230 120.445 ;
        RECT 52.040 120.400 52.330 120.445 ;
        RECT 53.610 120.400 53.900 120.445 ;
        RECT 49.940 120.260 53.900 120.400 ;
        RECT 49.940 120.215 50.230 120.260 ;
        RECT 52.040 120.215 52.330 120.260 ;
        RECT 53.610 120.215 53.900 120.260 ;
        RECT 56.355 120.215 56.645 120.445 ;
        RECT 58.640 120.400 58.960 120.460 ;
        RECT 62.410 120.400 62.550 120.940 ;
        RECT 75.200 120.880 75.520 120.940 ;
        RECT 79.340 120.880 79.660 121.140 ;
        RECT 80.810 121.125 80.950 121.280 ;
        RECT 82.190 121.125 82.330 121.620 ;
        RECT 83.020 121.560 83.340 121.620 ;
        RECT 92.220 121.760 92.540 121.820 ;
        RECT 96.835 121.760 97.125 121.805 ;
        RECT 92.220 121.620 97.125 121.760 ;
        RECT 92.220 121.560 92.540 121.620 ;
        RECT 96.835 121.575 97.125 121.620 ;
        RECT 97.280 121.760 97.600 121.820 ;
        RECT 100.515 121.760 100.805 121.805 ;
        RECT 97.280 121.620 100.805 121.760 ;
        RECT 97.280 121.560 97.600 121.620 ;
        RECT 100.515 121.575 100.805 121.620 ;
        RECT 102.340 121.560 102.660 121.820 ;
        RECT 112.000 121.560 112.320 121.820 ;
        RECT 113.855 121.760 114.145 121.805 ;
        RECT 114.300 121.760 114.620 121.820 ;
        RECT 113.855 121.620 114.620 121.760 ;
        RECT 113.855 121.575 114.145 121.620 ;
        RECT 114.300 121.560 114.620 121.620 ;
        RECT 122.135 121.760 122.425 121.805 ;
        RECT 125.340 121.760 125.660 121.820 ;
        RECT 122.135 121.620 125.660 121.760 ;
        RECT 122.135 121.575 122.425 121.620 ;
        RECT 125.340 121.560 125.660 121.620 ;
        RECT 133.175 121.760 133.465 121.805 ;
        RECT 134.080 121.760 134.400 121.820 ;
        RECT 133.175 121.620 134.400 121.760 ;
        RECT 133.175 121.575 133.465 121.620 ;
        RECT 134.080 121.560 134.400 121.620 ;
        RECT 135.000 121.760 135.320 121.820 ;
        RECT 136.855 121.760 137.145 121.805 ;
        RECT 140.535 121.760 140.825 121.805 ;
        RECT 135.000 121.620 137.145 121.760 ;
        RECT 135.000 121.560 135.320 121.620 ;
        RECT 136.855 121.575 137.145 121.620 ;
        RECT 139.690 121.620 143.510 121.760 ;
        RECT 102.815 121.420 103.105 121.465 ;
        RECT 124.420 121.420 124.740 121.480 ;
        RECT 134.540 121.420 134.860 121.480 ;
        RECT 82.650 121.280 93.830 121.420 ;
        RECT 82.650 121.125 82.790 121.280 ;
        RECT 83.940 121.125 84.260 121.140 ;
        RECT 90.010 121.125 90.150 121.280 ;
        RECT 93.690 121.140 93.830 121.280 ;
        RECT 95.990 121.280 103.950 121.420 ;
        RECT 91.300 121.125 91.620 121.140 ;
        RECT 80.275 120.895 80.565 121.125 ;
        RECT 80.735 120.895 81.025 121.125 ;
        RECT 82.115 120.895 82.405 121.125 ;
        RECT 82.575 120.895 82.865 121.125 ;
        RECT 83.910 120.895 84.260 121.125 ;
        RECT 89.935 120.895 90.225 121.125 ;
        RECT 91.270 121.080 91.620 121.125 ;
        RECT 91.105 120.940 91.620 121.080 ;
        RECT 91.270 120.895 91.620 120.940 ;
        RECT 69.245 120.740 69.535 120.785 ;
        RECT 71.765 120.740 72.055 120.785 ;
        RECT 72.955 120.740 73.245 120.785 ;
        RECT 69.245 120.600 73.245 120.740 ;
        RECT 69.245 120.555 69.535 120.600 ;
        RECT 71.765 120.555 72.055 120.600 ;
        RECT 72.955 120.555 73.245 120.600 ;
        RECT 73.820 120.540 74.140 120.800 ;
        RECT 74.280 120.740 74.600 120.800 ;
        RECT 77.515 120.740 77.805 120.785 ;
        RECT 74.280 120.600 77.805 120.740 ;
        RECT 74.280 120.540 74.600 120.600 ;
        RECT 77.515 120.555 77.805 120.600 ;
        RECT 58.640 120.260 62.550 120.400 ;
        RECT 69.680 120.400 69.970 120.445 ;
        RECT 71.250 120.400 71.540 120.445 ;
        RECT 73.350 120.400 73.640 120.445 ;
        RECT 69.680 120.260 73.640 120.400 ;
        RECT 80.350 120.400 80.490 120.895 ;
        RECT 83.940 120.880 84.260 120.895 ;
        RECT 91.300 120.880 91.620 120.895 ;
        RECT 93.600 120.880 93.920 121.140 ;
        RECT 95.990 120.800 96.130 121.280 ;
        RECT 102.815 121.235 103.105 121.280 ;
        RECT 83.455 120.740 83.745 120.785 ;
        RECT 84.645 120.740 84.935 120.785 ;
        RECT 87.165 120.740 87.455 120.785 ;
        RECT 83.455 120.600 87.455 120.740 ;
        RECT 83.455 120.555 83.745 120.600 ;
        RECT 84.645 120.555 84.935 120.600 ;
        RECT 87.165 120.555 87.455 120.600 ;
        RECT 89.460 120.540 89.780 120.800 ;
        RECT 90.815 120.740 91.105 120.785 ;
        RECT 92.005 120.740 92.295 120.785 ;
        RECT 94.525 120.740 94.815 120.785 ;
        RECT 90.815 120.600 94.815 120.740 ;
        RECT 90.815 120.555 91.105 120.600 ;
        RECT 92.005 120.555 92.295 120.600 ;
        RECT 94.525 120.555 94.815 120.600 ;
        RECT 95.900 120.540 96.220 120.800 ;
        RECT 103.260 120.540 103.580 120.800 ;
        RECT 83.060 120.400 83.350 120.445 ;
        RECT 85.160 120.400 85.450 120.445 ;
        RECT 86.730 120.400 87.020 120.445 ;
        RECT 89.550 120.400 89.690 120.540 ;
        RECT 80.350 120.260 82.100 120.400 ;
        RECT 58.640 120.200 58.960 120.260 ;
        RECT 69.680 120.215 69.970 120.260 ;
        RECT 71.250 120.215 71.540 120.260 ;
        RECT 73.350 120.215 73.640 120.260 ;
        RECT 54.500 120.060 54.820 120.120 ;
        RECT 41.710 119.920 54.820 120.060 ;
        RECT 38.415 119.875 38.705 119.920 ;
        RECT 40.240 119.860 40.560 119.920 ;
        RECT 54.500 119.860 54.820 119.920 ;
        RECT 56.800 119.860 57.120 120.120 ;
        RECT 62.780 119.860 63.100 120.120 ;
        RECT 74.740 119.860 75.060 120.120 ;
        RECT 81.960 120.060 82.100 120.260 ;
        RECT 83.060 120.260 87.020 120.400 ;
        RECT 83.060 120.215 83.350 120.260 ;
        RECT 85.160 120.215 85.450 120.260 ;
        RECT 86.730 120.215 87.020 120.260 ;
        RECT 87.710 120.260 89.690 120.400 ;
        RECT 90.420 120.400 90.710 120.445 ;
        RECT 92.520 120.400 92.810 120.445 ;
        RECT 94.090 120.400 94.380 120.445 ;
        RECT 90.420 120.260 94.380 120.400 ;
        RECT 87.710 120.060 87.850 120.260 ;
        RECT 90.420 120.215 90.710 120.260 ;
        RECT 92.520 120.215 92.810 120.260 ;
        RECT 94.090 120.215 94.380 120.260 ;
        RECT 81.960 119.920 87.850 120.060 ;
        RECT 88.080 120.060 88.400 120.120 ;
        RECT 89.475 120.060 89.765 120.105 ;
        RECT 88.080 119.920 89.765 120.060 ;
        RECT 103.810 120.060 103.950 121.280 ;
        RECT 105.190 121.280 126.490 121.420 ;
        RECT 105.190 121.125 105.330 121.280 ;
        RECT 107.950 121.140 108.090 121.280 ;
        RECT 106.480 121.125 106.800 121.140 ;
        RECT 105.115 120.895 105.405 121.125 ;
        RECT 106.450 121.080 106.800 121.125 ;
        RECT 106.285 120.940 106.800 121.080 ;
        RECT 106.450 120.895 106.800 120.940 ;
        RECT 106.480 120.880 106.800 120.895 ;
        RECT 107.860 120.880 108.180 121.140 ;
        RECT 119.360 121.125 119.680 121.140 ;
        RECT 120.830 121.125 120.970 121.280 ;
        RECT 124.420 121.220 124.740 121.280 ;
        RECT 126.350 121.140 126.490 121.280 ;
        RECT 126.810 121.280 134.860 121.420 ;
        RECT 119.360 120.895 119.710 121.125 ;
        RECT 120.755 120.895 121.045 121.125 ;
        RECT 119.360 120.880 119.680 120.895 ;
        RECT 121.200 120.880 121.520 121.140 ;
        RECT 121.660 121.080 121.980 121.140 ;
        RECT 122.580 121.080 122.900 121.140 ;
        RECT 123.055 121.080 123.345 121.125 ;
        RECT 121.660 120.940 123.345 121.080 ;
        RECT 121.660 120.880 121.980 120.940 ;
        RECT 122.580 120.880 122.900 120.940 ;
        RECT 123.055 120.895 123.345 120.940 ;
        RECT 123.515 120.895 123.805 121.125 ;
        RECT 123.975 120.895 124.265 121.125 ;
        RECT 124.895 120.895 125.185 121.125 ;
        RECT 105.995 120.740 106.285 120.785 ;
        RECT 107.185 120.740 107.475 120.785 ;
        RECT 109.705 120.740 109.995 120.785 ;
        RECT 105.995 120.600 109.995 120.740 ;
        RECT 105.995 120.555 106.285 120.600 ;
        RECT 107.185 120.555 107.475 120.600 ;
        RECT 109.705 120.555 109.995 120.600 ;
        RECT 116.165 120.740 116.455 120.785 ;
        RECT 118.685 120.740 118.975 120.785 ;
        RECT 119.875 120.740 120.165 120.785 ;
        RECT 116.165 120.600 120.165 120.740 ;
        RECT 121.290 120.740 121.430 120.880 ;
        RECT 123.590 120.740 123.730 120.895 ;
        RECT 121.290 120.600 123.730 120.740 ;
        RECT 116.165 120.555 116.455 120.600 ;
        RECT 118.685 120.555 118.975 120.600 ;
        RECT 119.875 120.555 120.165 120.600 ;
        RECT 105.600 120.400 105.890 120.445 ;
        RECT 107.700 120.400 107.990 120.445 ;
        RECT 109.270 120.400 109.560 120.445 ;
        RECT 105.600 120.260 109.560 120.400 ;
        RECT 105.600 120.215 105.890 120.260 ;
        RECT 107.700 120.215 107.990 120.260 ;
        RECT 109.270 120.215 109.560 120.260 ;
        RECT 116.600 120.400 116.890 120.445 ;
        RECT 118.170 120.400 118.460 120.445 ;
        RECT 120.270 120.400 120.560 120.445 ;
        RECT 116.600 120.260 120.560 120.400 ;
        RECT 124.050 120.400 124.190 120.895 ;
        RECT 124.970 120.740 125.110 120.895 ;
        RECT 126.260 120.880 126.580 121.140 ;
        RECT 126.810 120.740 126.950 121.280 ;
        RECT 134.540 121.220 134.860 121.280 ;
        RECT 135.090 121.280 137.530 121.420 ;
        RECT 127.640 121.125 127.960 121.140 ;
        RECT 127.610 121.080 127.960 121.125 ;
        RECT 127.445 120.940 127.960 121.080 ;
        RECT 127.610 120.895 127.960 120.940 ;
        RECT 127.640 120.880 127.960 120.895 ;
        RECT 132.240 120.880 132.560 121.140 ;
        RECT 135.090 121.125 135.230 121.280 ;
        RECT 137.390 121.140 137.530 121.280 ;
        RECT 135.015 120.895 135.305 121.125 ;
        RECT 135.935 121.080 136.225 121.125 ;
        RECT 136.380 121.080 136.700 121.140 ;
        RECT 135.935 120.940 136.700 121.080 ;
        RECT 135.935 120.895 136.225 120.940 ;
        RECT 136.380 120.880 136.700 120.940 ;
        RECT 137.300 120.880 137.620 121.140 ;
        RECT 137.775 120.895 138.065 121.125 ;
        RECT 124.970 120.600 126.950 120.740 ;
        RECT 127.155 120.740 127.445 120.785 ;
        RECT 128.345 120.740 128.635 120.785 ;
        RECT 130.865 120.740 131.155 120.785 ;
        RECT 127.155 120.600 131.155 120.740 ;
        RECT 132.330 120.740 132.470 120.880 ;
        RECT 134.555 120.740 134.845 120.785 ;
        RECT 132.330 120.600 134.845 120.740 ;
        RECT 127.155 120.555 127.445 120.600 ;
        RECT 128.345 120.555 128.635 120.600 ;
        RECT 130.865 120.555 131.155 120.600 ;
        RECT 134.555 120.555 134.845 120.600 ;
        RECT 135.460 120.540 135.780 120.800 ;
        RECT 125.340 120.400 125.660 120.460 ;
        RECT 124.050 120.260 125.660 120.400 ;
        RECT 116.600 120.215 116.890 120.260 ;
        RECT 118.170 120.215 118.460 120.260 ;
        RECT 120.270 120.215 120.560 120.260 ;
        RECT 125.340 120.200 125.660 120.260 ;
        RECT 126.760 120.400 127.050 120.445 ;
        RECT 128.860 120.400 129.150 120.445 ;
        RECT 130.430 120.400 130.720 120.445 ;
        RECT 126.760 120.260 130.720 120.400 ;
        RECT 126.760 120.215 127.050 120.260 ;
        RECT 128.860 120.215 129.150 120.260 ;
        RECT 130.430 120.215 130.720 120.260 ;
        RECT 134.080 120.400 134.400 120.460 ;
        RECT 137.850 120.400 137.990 120.895 ;
        RECT 138.220 120.880 138.540 121.140 ;
        RECT 138.680 120.880 139.000 121.140 ;
        RECT 139.140 120.880 139.460 121.140 ;
        RECT 139.690 121.125 139.830 121.620 ;
        RECT 140.535 121.575 140.825 121.620 ;
        RECT 143.370 121.420 143.510 121.620 ;
        RECT 144.200 121.560 144.520 121.820 ;
        RECT 144.660 121.560 144.980 121.820 ;
        RECT 144.750 121.420 144.890 121.560 ;
        RECT 143.370 121.280 144.890 121.420 ;
        RECT 149.890 121.420 150.180 121.465 ;
        RECT 150.640 121.420 150.960 121.480 ;
        RECT 149.890 121.280 150.960 121.420 ;
        RECT 149.890 121.235 150.180 121.280 ;
        RECT 150.640 121.220 150.960 121.280 ;
        RECT 139.615 120.895 139.905 121.125 ;
        RECT 140.075 120.895 140.365 121.125 ;
        RECT 140.995 120.895 141.285 121.125 ;
        RECT 142.375 121.080 142.665 121.125 ;
        RECT 151.115 121.080 151.405 121.125 ;
        RECT 154.320 121.080 154.640 121.140 ;
        RECT 142.375 120.940 145.810 121.080 ;
        RECT 142.375 120.895 142.665 120.940 ;
        RECT 138.770 120.740 138.910 120.880 ;
        RECT 140.150 120.740 140.290 120.895 ;
        RECT 138.770 120.600 140.290 120.740 ;
        RECT 134.080 120.260 137.990 120.400 ;
        RECT 141.070 120.400 141.210 120.895 ;
        RECT 145.670 120.800 145.810 120.940 ;
        RECT 151.115 120.940 154.640 121.080 ;
        RECT 151.115 120.895 151.405 120.940 ;
        RECT 154.320 120.880 154.640 120.940 ;
        RECT 143.295 120.740 143.585 120.785 ;
        RECT 145.120 120.740 145.440 120.800 ;
        RECT 143.295 120.600 145.440 120.740 ;
        RECT 143.295 120.555 143.585 120.600 ;
        RECT 141.900 120.400 142.220 120.460 ;
        RECT 143.370 120.400 143.510 120.555 ;
        RECT 145.120 120.540 145.440 120.600 ;
        RECT 145.580 120.540 145.900 120.800 ;
        RECT 146.525 120.740 146.815 120.785 ;
        RECT 149.045 120.740 149.335 120.785 ;
        RECT 150.235 120.740 150.525 120.785 ;
        RECT 146.525 120.600 150.525 120.740 ;
        RECT 146.525 120.555 146.815 120.600 ;
        RECT 149.045 120.555 149.335 120.600 ;
        RECT 150.235 120.555 150.525 120.600 ;
        RECT 141.070 120.260 143.510 120.400 ;
        RECT 146.960 120.400 147.250 120.445 ;
        RECT 148.530 120.400 148.820 120.445 ;
        RECT 150.630 120.400 150.920 120.445 ;
        RECT 146.960 120.260 150.920 120.400 ;
        RECT 134.080 120.200 134.400 120.260 ;
        RECT 141.900 120.200 142.220 120.260 ;
        RECT 146.960 120.215 147.250 120.260 ;
        RECT 148.530 120.215 148.820 120.260 ;
        RECT 150.630 120.215 150.920 120.260 ;
        RECT 121.200 120.060 121.520 120.120 ;
        RECT 103.810 119.920 121.520 120.060 ;
        RECT 88.080 119.860 88.400 119.920 ;
        RECT 89.475 119.875 89.765 119.920 ;
        RECT 121.200 119.860 121.520 119.920 ;
        RECT 123.040 120.060 123.360 120.120 ;
        RECT 133.635 120.060 133.925 120.105 ;
        RECT 137.760 120.060 138.080 120.120 ;
        RECT 123.040 119.920 138.080 120.060 ;
        RECT 123.040 119.860 123.360 119.920 ;
        RECT 133.635 119.875 133.925 119.920 ;
        RECT 137.760 119.860 138.080 119.920 ;
        RECT 141.440 119.860 141.760 120.120 ;
        RECT 22.690 119.240 157.010 119.720 ;
        RECT 27.835 119.040 28.125 119.085 ;
        RECT 31.960 119.040 32.280 119.100 ;
        RECT 27.835 118.900 32.280 119.040 ;
        RECT 27.835 118.855 28.125 118.900 ;
        RECT 31.960 118.840 32.280 118.900 ;
        RECT 51.280 118.840 51.600 119.100 ;
        RECT 56.800 118.840 57.120 119.100 ;
        RECT 59.575 119.040 59.865 119.085 ;
        RECT 60.480 119.040 60.800 119.100 ;
        RECT 59.575 118.900 60.800 119.040 ;
        RECT 59.575 118.855 59.865 118.900 ;
        RECT 60.480 118.840 60.800 118.900 ;
        RECT 62.780 118.840 63.100 119.100 ;
        RECT 74.740 118.840 75.060 119.100 ;
        RECT 78.420 118.840 78.740 119.100 ;
        RECT 79.340 118.840 79.660 119.100 ;
        RECT 83.940 118.840 84.260 119.100 ;
        RECT 87.250 118.900 90.150 119.040 ;
        RECT 31.040 118.700 31.330 118.745 ;
        RECT 32.610 118.700 32.900 118.745 ;
        RECT 34.710 118.700 35.000 118.745 ;
        RECT 45.300 118.700 45.620 118.760 ;
        RECT 55.435 118.700 55.725 118.745 ;
        RECT 31.040 118.560 35.000 118.700 ;
        RECT 31.040 118.515 31.330 118.560 ;
        RECT 32.610 118.515 32.900 118.560 ;
        RECT 34.710 118.515 35.000 118.560 ;
        RECT 41.710 118.560 45.620 118.700 ;
        RECT 30.605 118.360 30.895 118.405 ;
        RECT 33.125 118.360 33.415 118.405 ;
        RECT 34.315 118.360 34.605 118.405 ;
        RECT 30.605 118.220 34.605 118.360 ;
        RECT 30.605 118.175 30.895 118.220 ;
        RECT 33.125 118.175 33.415 118.220 ;
        RECT 34.315 118.175 34.605 118.220 ;
        RECT 25.520 118.020 25.840 118.080 ;
        RECT 25.995 118.020 26.285 118.065 ;
        RECT 25.520 117.880 26.285 118.020 ;
        RECT 25.520 117.820 25.840 117.880 ;
        RECT 25.995 117.835 26.285 117.880 ;
        RECT 31.040 118.020 31.360 118.080 ;
        RECT 41.710 118.065 41.850 118.560 ;
        RECT 45.300 118.500 45.620 118.560 ;
        RECT 49.070 118.560 55.725 118.700 ;
        RECT 43.090 118.220 46.910 118.360 ;
        RECT 35.195 118.020 35.485 118.065 ;
        RECT 31.040 117.880 35.485 118.020 ;
        RECT 31.040 117.820 31.360 117.880 ;
        RECT 35.195 117.835 35.485 117.880 ;
        RECT 38.875 117.835 39.165 118.065 ;
        RECT 41.175 117.835 41.465 118.065 ;
        RECT 41.635 117.835 41.925 118.065 ;
        RECT 26.915 117.680 27.205 117.725 ;
        RECT 31.500 117.680 31.820 117.740 ;
        RECT 33.340 117.680 33.660 117.740 ;
        RECT 26.915 117.540 33.660 117.680 ;
        RECT 26.915 117.495 27.205 117.540 ;
        RECT 31.500 117.480 31.820 117.540 ;
        RECT 33.340 117.480 33.660 117.540 ;
        RECT 33.800 117.725 34.120 117.740 ;
        RECT 33.800 117.495 34.150 117.725 ;
        RECT 38.950 117.680 39.090 117.835 ;
        RECT 35.730 117.540 39.090 117.680 ;
        RECT 41.250 117.680 41.390 117.835 ;
        RECT 42.080 117.820 42.400 118.080 ;
        RECT 43.090 118.065 43.230 118.220 ;
        RECT 43.015 117.835 43.305 118.065 ;
        RECT 43.920 118.020 44.240 118.080 ;
        RECT 46.235 118.020 46.525 118.065 ;
        RECT 43.920 117.880 46.525 118.020 ;
        RECT 43.920 117.820 44.240 117.880 ;
        RECT 46.235 117.835 46.525 117.880 ;
        RECT 46.770 118.020 46.910 118.220 ;
        RECT 48.075 118.020 48.365 118.065 ;
        RECT 48.520 118.020 48.840 118.080 ;
        RECT 49.070 118.065 49.210 118.560 ;
        RECT 55.435 118.515 55.725 118.560 ;
        RECT 56.890 118.360 57.030 118.840 ;
        RECT 49.990 118.220 57.030 118.360 ;
        RECT 49.990 118.065 50.130 118.220 ;
        RECT 58.640 118.160 58.960 118.420 ;
        RECT 62.870 118.360 63.010 118.840 ;
        RECT 68.315 118.360 68.605 118.405 ;
        RECT 62.870 118.220 68.605 118.360 ;
        RECT 68.315 118.175 68.605 118.220 ;
        RECT 68.760 118.160 69.080 118.420 ;
        RECT 46.770 117.880 48.840 118.020 ;
        RECT 43.475 117.680 43.765 117.725 ;
        RECT 41.250 117.540 43.765 117.680 ;
        RECT 33.800 117.480 34.120 117.495 ;
        RECT 35.730 117.400 35.870 117.540 ;
        RECT 43.475 117.495 43.765 117.540 ;
        RECT 44.840 117.680 45.160 117.740 ;
        RECT 46.770 117.680 46.910 117.880 ;
        RECT 48.075 117.835 48.365 117.880 ;
        RECT 48.520 117.820 48.840 117.880 ;
        RECT 48.995 117.835 49.285 118.065 ;
        RECT 49.455 117.835 49.745 118.065 ;
        RECT 49.915 117.835 50.205 118.065 ;
        RECT 49.530 117.680 49.670 117.835 ;
        RECT 52.200 117.820 52.520 118.080 ;
        RECT 58.730 118.020 58.870 118.160 ;
        RECT 52.750 117.880 58.870 118.020 ;
        RECT 60.035 118.020 60.325 118.065 ;
        RECT 68.850 118.020 68.990 118.160 ;
        RECT 60.035 117.880 68.990 118.020 ;
        RECT 71.075 118.020 71.365 118.065 ;
        RECT 74.830 118.020 74.970 118.840 ;
        RECT 80.260 118.700 80.580 118.760 ;
        RECT 87.250 118.700 87.390 118.900 ;
        RECT 80.260 118.560 87.390 118.700 ;
        RECT 80.260 118.500 80.580 118.560 ;
        RECT 87.635 118.515 87.925 118.745 ;
        RECT 90.010 118.700 90.150 118.900 ;
        RECT 92.680 118.840 93.000 119.100 ;
        RECT 109.240 119.040 109.560 119.100 ;
        RECT 110.635 119.040 110.925 119.085 ;
        RECT 109.240 118.900 110.925 119.040 ;
        RECT 109.240 118.840 109.560 118.900 ;
        RECT 110.635 118.855 110.925 118.900 ;
        RECT 119.360 119.040 119.680 119.100 ;
        RECT 119.835 119.040 120.125 119.085 ;
        RECT 135.460 119.040 135.780 119.100 ;
        RECT 135.935 119.040 136.225 119.085 ;
        RECT 119.360 118.900 120.125 119.040 ;
        RECT 119.360 118.840 119.680 118.900 ;
        RECT 119.835 118.855 120.125 118.900 ;
        RECT 121.290 118.900 134.310 119.040 ;
        RECT 113.840 118.700 114.160 118.760 ;
        RECT 115.680 118.700 116.000 118.760 ;
        RECT 121.290 118.700 121.430 118.900 ;
        RECT 90.010 118.560 121.430 118.700 ;
        RECT 121.660 118.700 121.980 118.760 ;
        RECT 122.595 118.700 122.885 118.745 ;
        RECT 121.660 118.560 122.885 118.700 ;
        RECT 83.495 118.360 83.785 118.405 ;
        RECT 85.320 118.360 85.640 118.420 ;
        RECT 83.495 118.220 85.640 118.360 ;
        RECT 83.495 118.175 83.785 118.220 ;
        RECT 85.320 118.160 85.640 118.220 ;
        RECT 79.800 118.020 80.120 118.080 ;
        RECT 71.075 117.880 74.970 118.020 ;
        RECT 78.670 117.895 80.120 118.020 ;
        RECT 78.665 117.880 80.120 117.895 ;
        RECT 44.840 117.540 46.910 117.680 ;
        RECT 49.070 117.540 49.670 117.680 ;
        RECT 44.840 117.480 45.160 117.540 ;
        RECT 26.440 117.340 26.760 117.400 ;
        RECT 28.295 117.340 28.585 117.385 ;
        RECT 35.640 117.340 35.960 117.400 ;
        RECT 26.440 117.200 35.960 117.340 ;
        RECT 26.440 117.140 26.760 117.200 ;
        RECT 28.295 117.155 28.585 117.200 ;
        RECT 35.640 117.140 35.960 117.200 ;
        RECT 36.100 117.140 36.420 117.400 ;
        RECT 39.780 117.140 40.100 117.400 ;
        RECT 45.300 117.340 45.620 117.400 ;
        RECT 49.070 117.340 49.210 117.540 ;
        RECT 45.300 117.200 49.210 117.340 ;
        RECT 49.440 117.340 49.760 117.400 ;
        RECT 52.750 117.340 52.890 117.880 ;
        RECT 60.035 117.835 60.325 117.880 ;
        RECT 71.075 117.835 71.365 117.880 ;
        RECT 54.960 117.680 55.280 117.740 ;
        RECT 56.355 117.680 56.645 117.725 ;
        RECT 54.960 117.540 56.645 117.680 ;
        RECT 54.960 117.480 55.280 117.540 ;
        RECT 56.355 117.495 56.645 117.540 ;
        RECT 57.260 117.480 57.580 117.740 ;
        RECT 67.855 117.680 68.145 117.725 ;
        RECT 74.280 117.680 74.600 117.740 ;
        RECT 67.855 117.540 74.600 117.680 ;
        RECT 67.855 117.495 68.145 117.540 ;
        RECT 74.280 117.480 74.600 117.540 ;
        RECT 77.515 117.680 77.805 117.725 ;
        RECT 77.960 117.680 78.280 117.740 ;
        RECT 77.515 117.540 78.280 117.680 ;
        RECT 78.665 117.665 78.955 117.880 ;
        RECT 79.800 117.820 80.120 117.880 ;
        RECT 80.735 118.020 81.025 118.065 ;
        RECT 82.100 118.020 82.420 118.080 ;
        RECT 80.735 117.880 82.420 118.020 ;
        RECT 80.735 117.835 81.025 117.880 ;
        RECT 82.100 117.820 82.420 117.880 ;
        RECT 82.575 117.835 82.865 118.065 ;
        RECT 84.875 118.020 85.165 118.065 ;
        RECT 87.710 118.020 87.850 118.515 ;
        RECT 113.840 118.500 114.160 118.560 ;
        RECT 115.680 118.500 116.000 118.560 ;
        RECT 121.660 118.500 121.980 118.560 ;
        RECT 122.595 118.515 122.885 118.560 ;
        RECT 89.000 118.360 89.320 118.420 ;
        RECT 90.395 118.360 90.685 118.405 ;
        RECT 89.000 118.220 90.685 118.360 ;
        RECT 89.000 118.160 89.320 118.220 ;
        RECT 90.395 118.175 90.685 118.220 ;
        RECT 90.840 118.160 91.160 118.420 ;
        RECT 95.915 118.360 96.205 118.405 ;
        RECT 98.660 118.360 98.980 118.420 ;
        RECT 101.420 118.360 101.740 118.420 ;
        RECT 101.895 118.360 102.185 118.405 ;
        RECT 95.915 118.220 102.185 118.360 ;
        RECT 95.915 118.175 96.205 118.220 ;
        RECT 98.660 118.160 98.980 118.220 ;
        RECT 101.420 118.160 101.740 118.220 ;
        RECT 101.895 118.175 102.185 118.220 ;
        RECT 112.460 118.160 112.780 118.420 ;
        RECT 114.300 118.360 114.620 118.420 ;
        RECT 116.155 118.360 116.445 118.405 ;
        RECT 114.300 118.220 116.445 118.360 ;
        RECT 114.300 118.160 114.620 118.220 ;
        RECT 116.155 118.175 116.445 118.220 ;
        RECT 117.520 118.360 117.840 118.420 ;
        RECT 123.040 118.360 123.360 118.420 ;
        RECT 129.035 118.360 129.325 118.405 ;
        RECT 117.520 118.220 123.360 118.360 ;
        RECT 117.520 118.160 117.840 118.220 ;
        RECT 84.875 117.880 87.850 118.020 ;
        RECT 89.935 118.020 90.225 118.065 ;
        RECT 90.930 118.020 91.070 118.160 ;
        RECT 89.935 117.880 91.070 118.020 ;
        RECT 94.535 118.020 94.825 118.065 ;
        RECT 94.980 118.020 95.300 118.080 ;
        RECT 94.535 117.880 95.300 118.020 ;
        RECT 84.875 117.835 85.165 117.880 ;
        RECT 89.935 117.835 90.225 117.880 ;
        RECT 94.535 117.835 94.825 117.880 ;
        RECT 77.515 117.495 77.805 117.540 ;
        RECT 77.960 117.480 78.280 117.540 ;
        RECT 82.650 117.400 82.790 117.835 ;
        RECT 94.980 117.820 95.300 117.880 ;
        RECT 100.960 117.820 101.280 118.080 ;
        RECT 111.080 117.820 111.400 118.080 ;
        RECT 111.555 118.020 111.845 118.065 ;
        RECT 112.000 118.020 112.320 118.080 ;
        RECT 111.555 117.880 112.320 118.020 ;
        RECT 111.555 117.835 111.845 117.880 ;
        RECT 112.000 117.820 112.320 117.880 ;
        RECT 113.395 118.020 113.685 118.065 ;
        RECT 117.980 118.020 118.300 118.080 ;
        RECT 113.395 117.880 118.300 118.020 ;
        RECT 113.395 117.835 113.685 117.880 ;
        RECT 89.460 117.680 89.780 117.740 ;
        RECT 95.440 117.680 95.760 117.740 ;
        RECT 101.435 117.680 101.725 117.725 ;
        RECT 111.170 117.680 111.310 117.820 ;
        RECT 113.470 117.680 113.610 117.835 ;
        RECT 117.980 117.820 118.300 117.880 ;
        RECT 118.440 118.020 118.760 118.080 ;
        RECT 122.210 118.065 122.350 118.220 ;
        RECT 123.040 118.160 123.360 118.220 ;
        RECT 124.510 118.220 129.325 118.360 ;
        RECT 120.755 118.020 121.045 118.065 ;
        RECT 118.440 117.880 121.045 118.020 ;
        RECT 118.440 117.820 118.760 117.880 ;
        RECT 120.755 117.835 121.045 117.880 ;
        RECT 122.135 117.835 122.425 118.065 ;
        RECT 122.580 117.820 122.900 118.080 ;
        RECT 123.500 117.820 123.820 118.080 ;
        RECT 124.510 118.065 124.650 118.220 ;
        RECT 129.035 118.175 129.325 118.220 ;
        RECT 130.260 118.220 133.850 118.360 ;
        RECT 124.435 117.835 124.725 118.065 ;
        RECT 126.275 118.020 126.565 118.065 ;
        RECT 130.260 118.020 130.400 118.220 ;
        RECT 124.970 117.880 130.400 118.020 ;
        RECT 89.460 117.540 101.190 117.680 ;
        RECT 89.460 117.480 89.780 117.540 ;
        RECT 95.440 117.480 95.760 117.540 ;
        RECT 49.440 117.200 52.890 117.340 ;
        RECT 57.735 117.340 58.025 117.385 ;
        RECT 61.400 117.340 61.720 117.400 ;
        RECT 57.735 117.200 61.720 117.340 ;
        RECT 45.300 117.140 45.620 117.200 ;
        RECT 49.440 117.140 49.760 117.200 ;
        RECT 57.735 117.155 58.025 117.200 ;
        RECT 61.400 117.140 61.720 117.200 ;
        RECT 66.000 117.140 66.320 117.400 ;
        RECT 70.600 117.140 70.920 117.400 ;
        RECT 79.800 117.140 80.120 117.400 ;
        RECT 81.640 117.140 81.960 117.400 ;
        RECT 82.560 117.140 82.880 117.400 ;
        RECT 84.400 117.340 84.720 117.400 ;
        RECT 94.995 117.340 95.285 117.385 ;
        RECT 95.900 117.340 96.220 117.400 ;
        RECT 84.400 117.200 96.220 117.340 ;
        RECT 84.400 117.140 84.720 117.200 ;
        RECT 94.995 117.155 95.285 117.200 ;
        RECT 95.900 117.140 96.220 117.200 ;
        RECT 99.120 117.140 99.440 117.400 ;
        RECT 101.050 117.340 101.190 117.540 ;
        RECT 101.435 117.540 113.610 117.680 ;
        RECT 113.840 117.680 114.160 117.740 ;
        RECT 114.775 117.680 115.065 117.725 ;
        RECT 122.670 117.680 122.810 117.820 ;
        RECT 124.970 117.680 125.110 117.880 ;
        RECT 126.275 117.835 126.565 117.880 ;
        RECT 132.240 117.820 132.560 118.080 ;
        RECT 133.710 118.065 133.850 118.220 ;
        RECT 134.170 118.065 134.310 118.900 ;
        RECT 135.460 118.900 136.225 119.040 ;
        RECT 135.460 118.840 135.780 118.900 ;
        RECT 135.935 118.855 136.225 118.900 ;
        RECT 139.140 119.040 139.460 119.100 ;
        RECT 142.375 119.040 142.665 119.085 ;
        RECT 139.140 118.900 142.665 119.040 ;
        RECT 139.140 118.840 139.460 118.900 ;
        RECT 142.375 118.855 142.665 118.900 ;
        RECT 143.280 119.040 143.600 119.100 ;
        RECT 151.100 119.040 151.420 119.100 ;
        RECT 143.280 118.900 151.420 119.040 ;
        RECT 140.535 118.700 140.825 118.745 ;
        RECT 141.440 118.700 141.760 118.760 ;
        RECT 140.535 118.560 141.760 118.700 ;
        RECT 142.450 118.700 142.590 118.855 ;
        RECT 143.280 118.840 143.600 118.900 ;
        RECT 151.100 118.840 151.420 118.900 ;
        RECT 146.500 118.700 146.820 118.760 ;
        RECT 142.450 118.560 146.820 118.700 ;
        RECT 140.535 118.515 140.825 118.560 ;
        RECT 141.440 118.500 141.760 118.560 ;
        RECT 146.500 118.500 146.820 118.560 ;
        RECT 150.180 118.700 150.470 118.745 ;
        RECT 151.750 118.700 152.040 118.745 ;
        RECT 153.850 118.700 154.140 118.745 ;
        RECT 150.180 118.560 154.140 118.700 ;
        RECT 150.180 118.515 150.470 118.560 ;
        RECT 151.750 118.515 152.040 118.560 ;
        RECT 153.850 118.515 154.140 118.560 ;
        RECT 139.615 118.360 139.905 118.405 ;
        RECT 147.420 118.360 147.740 118.420 ;
        RECT 139.615 118.220 147.740 118.360 ;
        RECT 139.615 118.175 139.905 118.220 ;
        RECT 147.420 118.160 147.740 118.220 ;
        RECT 149.745 118.360 150.035 118.405 ;
        RECT 152.265 118.360 152.555 118.405 ;
        RECT 153.455 118.360 153.745 118.405 ;
        RECT 149.745 118.220 153.745 118.360 ;
        RECT 149.745 118.175 150.035 118.220 ;
        RECT 152.265 118.175 152.555 118.220 ;
        RECT 153.455 118.175 153.745 118.220 ;
        RECT 154.320 118.160 154.640 118.420 ;
        RECT 133.635 117.835 133.925 118.065 ;
        RECT 134.095 117.835 134.385 118.065 ;
        RECT 135.460 117.820 135.780 118.080 ;
        RECT 138.220 118.020 138.540 118.080 ;
        RECT 139.155 118.020 139.445 118.065 ;
        RECT 138.220 117.880 139.445 118.020 ;
        RECT 138.220 117.820 138.540 117.880 ;
        RECT 139.155 117.835 139.445 117.880 ;
        RECT 140.075 118.020 140.365 118.065 ;
        RECT 146.040 118.020 146.360 118.080 ;
        RECT 140.075 117.880 146.360 118.020 ;
        RECT 140.075 117.835 140.365 117.880 ;
        RECT 146.040 117.820 146.360 117.880 ;
        RECT 146.500 117.820 146.820 118.080 ;
        RECT 113.840 117.540 115.065 117.680 ;
        RECT 101.435 117.495 101.725 117.540 ;
        RECT 113.840 117.480 114.160 117.540 ;
        RECT 114.775 117.495 115.065 117.540 ;
        RECT 118.990 117.540 122.350 117.680 ;
        RECT 122.670 117.540 125.110 117.680 ;
        RECT 118.990 117.340 119.130 117.540 ;
        RECT 101.050 117.200 119.130 117.340 ;
        RECT 119.375 117.340 119.665 117.385 ;
        RECT 121.675 117.340 121.965 117.385 ;
        RECT 119.375 117.200 121.965 117.340 ;
        RECT 122.210 117.340 122.350 117.540 ;
        RECT 125.340 117.480 125.660 117.740 ;
        RECT 125.800 117.480 126.120 117.740 ;
        RECT 126.350 117.540 133.390 117.680 ;
        RECT 124.880 117.340 125.200 117.400 ;
        RECT 122.210 117.200 125.200 117.340 ;
        RECT 125.430 117.340 125.570 117.480 ;
        RECT 126.350 117.340 126.490 117.540 ;
        RECT 125.430 117.200 126.490 117.340 ;
        RECT 119.375 117.155 119.665 117.200 ;
        RECT 121.675 117.155 121.965 117.200 ;
        RECT 124.880 117.140 125.200 117.200 ;
        RECT 127.180 117.140 127.500 117.400 ;
        RECT 132.700 117.140 133.020 117.400 ;
        RECT 133.250 117.340 133.390 117.540 ;
        RECT 134.555 117.495 134.845 117.725 ;
        RECT 134.630 117.340 134.770 117.495 ;
        RECT 136.840 117.480 137.160 117.740 ;
        RECT 137.760 117.480 138.080 117.740 ;
        RECT 144.660 117.680 144.980 117.740 ;
        RECT 142.450 117.540 144.980 117.680 ;
        RECT 142.450 117.385 142.590 117.540 ;
        RECT 144.660 117.480 144.980 117.540 ;
        RECT 152.940 117.725 153.260 117.740 ;
        RECT 152.940 117.495 153.290 117.725 ;
        RECT 152.940 117.480 153.260 117.495 ;
        RECT 133.250 117.200 134.770 117.340 ;
        RECT 142.375 117.155 142.665 117.385 ;
        RECT 143.280 117.140 143.600 117.400 ;
        RECT 143.740 117.140 144.060 117.400 ;
        RECT 145.120 117.340 145.440 117.400 ;
        RECT 147.435 117.340 147.725 117.385 ;
        RECT 145.120 117.200 147.725 117.340 ;
        RECT 145.120 117.140 145.440 117.200 ;
        RECT 147.435 117.155 147.725 117.200 ;
        RECT 22.690 116.520 157.810 117.000 ;
        RECT 26.915 116.320 27.205 116.365 ;
        RECT 29.660 116.320 29.980 116.380 ;
        RECT 26.915 116.180 29.980 116.320 ;
        RECT 26.915 116.135 27.205 116.180 ;
        RECT 29.660 116.120 29.980 116.180 ;
        RECT 33.800 116.320 34.120 116.380 ;
        RECT 34.275 116.320 34.565 116.365 ;
        RECT 33.800 116.180 34.565 116.320 ;
        RECT 33.800 116.120 34.120 116.180 ;
        RECT 34.275 116.135 34.565 116.180 ;
        RECT 36.100 116.120 36.420 116.380 ;
        RECT 37.035 116.320 37.325 116.365 ;
        RECT 40.700 116.320 41.020 116.380 ;
        RECT 37.035 116.180 41.020 116.320 ;
        RECT 37.035 116.135 37.325 116.180 ;
        RECT 40.700 116.120 41.020 116.180 ;
        RECT 58.640 116.120 58.960 116.380 ;
        RECT 70.600 116.120 70.920 116.380 ;
        RECT 79.800 116.320 80.120 116.380 ;
        RECT 77.130 116.180 80.120 116.320 ;
        RECT 36.190 115.980 36.330 116.120 ;
        RECT 29.290 115.840 36.330 115.980 ;
        RECT 25.060 115.440 25.380 115.700 ;
        RECT 25.995 115.455 26.285 115.685 ;
        RECT 27.375 115.455 27.665 115.685 ;
        RECT 26.070 114.960 26.210 115.455 ;
        RECT 27.450 115.300 27.590 115.455 ;
        RECT 28.280 115.440 28.600 115.700 ;
        RECT 28.740 115.440 29.060 115.700 ;
        RECT 29.290 115.685 29.430 115.840 ;
        RECT 37.480 115.780 37.800 116.040 ;
        RECT 38.830 115.980 39.120 116.025 ;
        RECT 39.780 115.980 40.100 116.040 ;
        RECT 48.075 115.980 48.365 116.025 ;
        RECT 56.400 115.980 56.690 116.025 ;
        RECT 38.830 115.840 40.100 115.980 ;
        RECT 38.830 115.795 39.120 115.840 ;
        RECT 39.780 115.780 40.100 115.840 ;
        RECT 45.390 115.840 46.450 115.980 ;
        RECT 29.215 115.455 29.505 115.685 ;
        RECT 32.420 115.640 32.740 115.700 ;
        RECT 29.750 115.500 32.740 115.640 ;
        RECT 29.750 115.300 29.890 115.500 ;
        RECT 32.420 115.440 32.740 115.500 ;
        RECT 34.720 115.440 35.040 115.700 ;
        RECT 35.640 115.440 35.960 115.700 ;
        RECT 36.115 115.455 36.405 115.685 ;
        RECT 37.570 115.640 37.710 115.780 ;
        RECT 45.390 115.700 45.530 115.840 ;
        RECT 36.650 115.500 37.710 115.640 ;
        RECT 27.450 115.160 29.890 115.300 ;
        RECT 30.595 115.300 30.885 115.345 ;
        RECT 31.055 115.300 31.345 115.345 ;
        RECT 30.595 115.160 31.345 115.300 ;
        RECT 30.595 115.115 30.885 115.160 ;
        RECT 31.055 115.115 31.345 115.160 ;
        RECT 33.800 115.300 34.120 115.360 ;
        RECT 36.190 115.300 36.330 115.455 ;
        RECT 33.800 115.160 36.330 115.300 ;
        RECT 33.800 115.100 34.120 115.160 ;
        RECT 36.650 114.960 36.790 115.500 ;
        RECT 44.840 115.440 45.160 115.700 ;
        RECT 45.300 115.440 45.620 115.700 ;
        RECT 46.310 115.685 46.450 115.840 ;
        RECT 48.075 115.840 56.690 115.980 ;
        RECT 48.075 115.795 48.365 115.840 ;
        RECT 56.400 115.795 56.690 115.840 ;
        RECT 63.715 115.980 64.005 116.025 ;
        RECT 64.620 115.980 64.940 116.040 ;
        RECT 68.300 115.980 68.620 116.040 ;
        RECT 63.715 115.840 64.940 115.980 ;
        RECT 63.715 115.795 64.005 115.840 ;
        RECT 64.620 115.780 64.940 115.840 ;
        RECT 65.630 115.840 68.620 115.980 ;
        RECT 65.630 115.700 65.770 115.840 ;
        RECT 68.300 115.780 68.620 115.840 ;
        RECT 76.550 115.980 76.840 116.025 ;
        RECT 77.130 115.980 77.270 116.180 ;
        RECT 79.800 116.120 80.120 116.180 ;
        RECT 93.600 116.120 93.920 116.380 ;
        RECT 97.295 116.135 97.585 116.365 ;
        RECT 98.200 116.320 98.520 116.380 ;
        RECT 99.120 116.320 99.440 116.380 ;
        RECT 98.200 116.180 99.440 116.320 ;
        RECT 76.550 115.840 77.270 115.980 ;
        RECT 77.500 115.980 77.820 116.040 ;
        RECT 83.495 115.980 83.785 116.025 ;
        RECT 77.500 115.840 83.785 115.980 ;
        RECT 76.550 115.795 76.840 115.840 ;
        RECT 77.500 115.780 77.820 115.840 ;
        RECT 83.495 115.795 83.785 115.840 ;
        RECT 92.235 115.980 92.525 116.025 ;
        RECT 93.690 115.980 93.830 116.120 ;
        RECT 92.235 115.840 93.830 115.980 ;
        RECT 97.370 115.980 97.510 116.135 ;
        RECT 98.200 116.120 98.520 116.180 ;
        RECT 99.120 116.120 99.440 116.180 ;
        RECT 99.595 116.320 99.885 116.365 ;
        RECT 100.960 116.320 101.280 116.380 ;
        RECT 99.595 116.180 101.280 116.320 ;
        RECT 99.595 116.135 99.885 116.180 ;
        RECT 100.960 116.120 101.280 116.180 ;
        RECT 117.980 116.120 118.300 116.380 ;
        RECT 123.515 116.320 123.805 116.365 ;
        RECT 124.420 116.320 124.740 116.380 ;
        RECT 129.940 116.320 130.260 116.380 ;
        RECT 123.515 116.180 124.740 116.320 ;
        RECT 123.515 116.135 123.805 116.180 ;
        RECT 124.420 116.120 124.740 116.180 ;
        RECT 124.970 116.180 130.260 116.320 ;
        RECT 106.080 115.980 106.370 116.025 ;
        RECT 97.370 115.840 106.370 115.980 ;
        RECT 92.235 115.795 92.525 115.840 ;
        RECT 106.080 115.795 106.370 115.840 ;
        RECT 121.200 115.980 121.520 116.040 ;
        RECT 124.970 115.980 125.110 116.180 ;
        RECT 129.940 116.120 130.260 116.180 ;
        RECT 132.240 116.320 132.560 116.380 ;
        RECT 133.175 116.320 133.465 116.365 ;
        RECT 134.540 116.320 134.860 116.380 ;
        RECT 132.240 116.180 134.860 116.320 ;
        RECT 132.240 116.120 132.560 116.180 ;
        RECT 133.175 116.135 133.465 116.180 ;
        RECT 134.540 116.120 134.860 116.180 ;
        RECT 135.460 116.320 135.780 116.380 ;
        RECT 136.855 116.320 137.145 116.365 ;
        RECT 139.155 116.320 139.445 116.365 ;
        RECT 135.460 116.180 137.145 116.320 ;
        RECT 135.460 116.120 135.780 116.180 ;
        RECT 136.855 116.135 137.145 116.180 ;
        RECT 137.850 116.180 139.445 116.320 ;
        RECT 127.640 116.025 127.960 116.040 ;
        RECT 121.200 115.840 125.110 115.980 ;
        RECT 45.775 115.455 46.065 115.685 ;
        RECT 46.235 115.455 46.525 115.685 ;
        RECT 46.695 115.640 46.985 115.685 ;
        RECT 54.960 115.640 55.280 115.700 ;
        RECT 46.695 115.500 55.280 115.640 ;
        RECT 46.695 115.455 46.985 115.500 ;
        RECT 37.495 115.115 37.785 115.345 ;
        RECT 38.375 115.300 38.665 115.345 ;
        RECT 39.565 115.300 39.855 115.345 ;
        RECT 42.085 115.300 42.375 115.345 ;
        RECT 38.375 115.160 42.375 115.300 ;
        RECT 38.375 115.115 38.665 115.160 ;
        RECT 39.565 115.115 39.855 115.160 ;
        RECT 42.085 115.115 42.375 115.160 ;
        RECT 26.070 114.820 36.790 114.960 ;
        RECT 25.520 114.620 25.840 114.680 ;
        RECT 34.735 114.620 35.025 114.665 ;
        RECT 25.520 114.480 35.025 114.620 ;
        RECT 37.570 114.620 37.710 115.115 ;
        RECT 37.980 114.960 38.270 115.005 ;
        RECT 40.080 114.960 40.370 115.005 ;
        RECT 41.650 114.960 41.940 115.005 ;
        RECT 37.980 114.820 41.940 114.960 ;
        RECT 44.930 114.960 45.070 115.440 ;
        RECT 45.850 115.300 45.990 115.455 ;
        RECT 54.960 115.440 55.280 115.500 ;
        RECT 58.180 115.440 58.500 115.700 ;
        RECT 60.940 115.440 61.260 115.700 ;
        RECT 61.400 115.440 61.720 115.700 ;
        RECT 62.320 115.440 62.640 115.700 ;
        RECT 63.240 115.640 63.560 115.700 ;
        RECT 64.175 115.640 64.465 115.685 ;
        RECT 63.240 115.500 64.465 115.640 ;
        RECT 63.240 115.440 63.560 115.500 ;
        RECT 64.175 115.455 64.465 115.500 ;
        RECT 65.095 115.455 65.385 115.685 ;
        RECT 52.660 115.300 52.980 115.360 ;
        RECT 45.850 115.160 52.980 115.300 ;
        RECT 52.660 115.100 52.980 115.160 ;
        RECT 53.145 115.300 53.435 115.345 ;
        RECT 55.665 115.300 55.955 115.345 ;
        RECT 56.855 115.300 57.145 115.345 ;
        RECT 53.145 115.160 57.145 115.300 ;
        RECT 53.145 115.115 53.435 115.160 ;
        RECT 55.665 115.115 55.955 115.160 ;
        RECT 56.855 115.115 57.145 115.160 ;
        RECT 57.720 115.300 58.040 115.360 ;
        RECT 61.030 115.300 61.170 115.440 ;
        RECT 57.720 115.160 61.170 115.300 ;
        RECT 57.720 115.100 58.040 115.160 ;
        RECT 53.580 114.960 53.870 115.005 ;
        RECT 55.150 114.960 55.440 115.005 ;
        RECT 57.250 114.960 57.540 115.005 ;
        RECT 44.930 114.820 47.370 114.960 ;
        RECT 37.980 114.775 38.270 114.820 ;
        RECT 40.080 114.775 40.370 114.820 ;
        RECT 41.650 114.775 41.940 114.820 ;
        RECT 47.230 114.680 47.370 114.820 ;
        RECT 53.580 114.820 57.540 114.960 ;
        RECT 53.580 114.775 53.870 114.820 ;
        RECT 55.150 114.775 55.440 114.820 ;
        RECT 57.250 114.775 57.540 114.820 ;
        RECT 42.080 114.620 42.400 114.680 ;
        RECT 37.570 114.480 42.400 114.620 ;
        RECT 25.520 114.420 25.840 114.480 ;
        RECT 34.735 114.435 35.025 114.480 ;
        RECT 42.080 114.420 42.400 114.480 ;
        RECT 43.920 114.620 44.240 114.680 ;
        RECT 44.395 114.620 44.685 114.665 ;
        RECT 43.920 114.480 44.685 114.620 ;
        RECT 43.920 114.420 44.240 114.480 ;
        RECT 44.395 114.435 44.685 114.480 ;
        RECT 47.140 114.420 47.460 114.680 ;
        RECT 50.835 114.620 51.125 114.665 ;
        RECT 52.200 114.620 52.520 114.680 ;
        RECT 54.040 114.620 54.360 114.680 ;
        RECT 50.835 114.480 54.360 114.620 ;
        RECT 64.250 114.620 64.390 115.455 ;
        RECT 65.170 115.300 65.310 115.455 ;
        RECT 65.540 115.440 65.860 115.700 ;
        RECT 66.460 115.440 66.780 115.700 ;
        RECT 68.390 115.300 68.530 115.780 ;
        RECT 73.835 115.640 74.125 115.685 ;
        RECT 72.530 115.500 74.125 115.640 ;
        RECT 69.235 115.300 69.525 115.345 ;
        RECT 65.170 115.160 66.690 115.300 ;
        RECT 68.390 115.160 69.525 115.300 ;
        RECT 66.550 114.680 66.690 115.160 ;
        RECT 69.235 115.115 69.525 115.160 ;
        RECT 70.140 115.100 70.460 115.360 ;
        RECT 72.530 115.005 72.670 115.500 ;
        RECT 73.835 115.455 74.125 115.500 ;
        RECT 75.200 115.640 75.520 115.700 ;
        RECT 79.340 115.640 79.660 115.700 ;
        RECT 92.310 115.640 92.450 115.795 ;
        RECT 121.200 115.780 121.520 115.840 ;
        RECT 127.500 115.795 127.960 116.025 ;
        RECT 137.850 115.980 137.990 116.180 ;
        RECT 139.155 116.135 139.445 116.180 ;
        RECT 146.500 116.320 146.820 116.380 ;
        RECT 151.115 116.320 151.405 116.365 ;
        RECT 146.500 116.180 151.405 116.320 ;
        RECT 146.500 116.120 146.820 116.180 ;
        RECT 151.115 116.135 151.405 116.180 ;
        RECT 152.940 116.120 153.260 116.380 ;
        RECT 127.640 115.780 127.960 115.795 ;
        RECT 136.930 115.840 137.990 115.980 ;
        RECT 138.220 115.980 138.540 116.040 ;
        RECT 149.720 115.980 150.040 116.040 ;
        RECT 154.320 115.980 154.640 116.040 ;
        RECT 138.220 115.840 154.640 115.980 ;
        RECT 75.200 115.500 92.450 115.640 ;
        RECT 75.200 115.440 75.520 115.500 ;
        RECT 79.340 115.440 79.660 115.500 ;
        RECT 92.680 115.440 93.000 115.700 ;
        RECT 93.615 115.455 93.905 115.685 ;
        RECT 76.095 115.300 76.385 115.345 ;
        RECT 77.285 115.300 77.575 115.345 ;
        RECT 79.805 115.300 80.095 115.345 ;
        RECT 76.095 115.160 80.095 115.300 ;
        RECT 76.095 115.115 76.385 115.160 ;
        RECT 77.285 115.115 77.575 115.160 ;
        RECT 79.805 115.115 80.095 115.160 ;
        RECT 72.455 114.775 72.745 115.005 ;
        RECT 75.700 114.960 75.990 115.005 ;
        RECT 77.800 114.960 78.090 115.005 ;
        RECT 79.370 114.960 79.660 115.005 ;
        RECT 75.700 114.820 79.660 114.960 ;
        RECT 93.690 114.960 93.830 115.455 ;
        RECT 94.060 115.440 94.380 115.700 ;
        RECT 96.375 115.640 96.665 115.685 ;
        RECT 98.200 115.640 98.520 115.700 ;
        RECT 96.375 115.500 98.520 115.640 ;
        RECT 96.375 115.455 96.665 115.500 ;
        RECT 98.200 115.440 98.520 115.500 ;
        RECT 98.675 115.455 98.965 115.685 ;
        RECT 103.260 115.640 103.580 115.700 ;
        RECT 109.700 115.685 110.020 115.700 ;
        RECT 103.260 115.500 107.630 115.640 ;
        RECT 94.150 115.300 94.290 115.440 ;
        RECT 97.755 115.300 98.045 115.345 ;
        RECT 94.150 115.160 98.045 115.300 ;
        RECT 97.755 115.115 98.045 115.160 ;
        RECT 98.750 114.960 98.890 115.455 ;
        RECT 103.260 115.440 103.580 115.500 ;
        RECT 107.490 115.345 107.630 115.500 ;
        RECT 109.670 115.455 110.020 115.685 ;
        RECT 109.700 115.440 110.020 115.455 ;
        RECT 117.520 115.440 117.840 115.700 ;
        RECT 118.900 115.640 119.220 115.700 ;
        RECT 121.675 115.640 121.965 115.685 ;
        RECT 118.900 115.500 121.965 115.640 ;
        RECT 118.900 115.440 119.220 115.500 ;
        RECT 121.675 115.455 121.965 115.500 ;
        RECT 126.260 115.440 126.580 115.700 ;
        RECT 102.825 115.300 103.115 115.345 ;
        RECT 105.345 115.300 105.635 115.345 ;
        RECT 106.535 115.300 106.825 115.345 ;
        RECT 102.825 115.160 106.825 115.300 ;
        RECT 102.825 115.115 103.115 115.160 ;
        RECT 105.345 115.115 105.635 115.160 ;
        RECT 106.535 115.115 106.825 115.160 ;
        RECT 107.415 115.300 107.705 115.345 ;
        RECT 108.335 115.300 108.625 115.345 ;
        RECT 107.415 115.160 108.625 115.300 ;
        RECT 107.415 115.115 107.705 115.160 ;
        RECT 108.335 115.115 108.625 115.160 ;
        RECT 109.215 115.300 109.505 115.345 ;
        RECT 110.405 115.300 110.695 115.345 ;
        RECT 112.925 115.300 113.215 115.345 ;
        RECT 118.455 115.300 118.745 115.345 ;
        RECT 119.820 115.300 120.140 115.360 ;
        RECT 120.295 115.300 120.585 115.345 ;
        RECT 109.215 115.160 113.215 115.300 ;
        RECT 109.215 115.115 109.505 115.160 ;
        RECT 110.405 115.115 110.695 115.160 ;
        RECT 112.925 115.115 113.215 115.160 ;
        RECT 113.470 115.160 120.585 115.300 ;
        RECT 100.515 114.960 100.805 115.005 ;
        RECT 93.690 114.820 100.805 114.960 ;
        RECT 75.700 114.775 75.990 114.820 ;
        RECT 77.800 114.775 78.090 114.820 ;
        RECT 79.370 114.775 79.660 114.820 ;
        RECT 100.515 114.775 100.805 114.820 ;
        RECT 103.260 114.960 103.550 115.005 ;
        RECT 104.830 114.960 105.120 115.005 ;
        RECT 106.930 114.960 107.220 115.005 ;
        RECT 103.260 114.820 107.220 114.960 ;
        RECT 103.260 114.775 103.550 114.820 ;
        RECT 104.830 114.775 105.120 114.820 ;
        RECT 106.930 114.775 107.220 114.820 ;
        RECT 108.820 114.960 109.110 115.005 ;
        RECT 110.920 114.960 111.210 115.005 ;
        RECT 112.490 114.960 112.780 115.005 ;
        RECT 108.820 114.820 112.780 114.960 ;
        RECT 108.820 114.775 109.110 114.820 ;
        RECT 110.920 114.775 111.210 114.820 ;
        RECT 112.490 114.775 112.780 114.820 ;
        RECT 65.555 114.620 65.845 114.665 ;
        RECT 64.250 114.480 65.845 114.620 ;
        RECT 50.835 114.435 51.125 114.480 ;
        RECT 52.200 114.420 52.520 114.480 ;
        RECT 54.040 114.420 54.360 114.480 ;
        RECT 65.555 114.435 65.845 114.480 ;
        RECT 66.460 114.420 66.780 114.680 ;
        RECT 67.840 114.420 68.160 114.680 ;
        RECT 71.520 114.620 71.840 114.680 ;
        RECT 72.915 114.620 73.205 114.665 ;
        RECT 71.520 114.480 73.205 114.620 ;
        RECT 71.520 114.420 71.840 114.480 ;
        RECT 72.915 114.435 73.205 114.480 ;
        RECT 82.115 114.620 82.405 114.665 ;
        RECT 82.560 114.620 82.880 114.680 ;
        RECT 86.700 114.620 87.020 114.680 ;
        RECT 82.115 114.480 87.020 114.620 ;
        RECT 82.115 114.435 82.405 114.480 ;
        RECT 82.560 114.420 82.880 114.480 ;
        RECT 86.700 114.420 87.020 114.480 ;
        RECT 91.760 114.620 92.080 114.680 ;
        RECT 92.695 114.620 92.985 114.665 ;
        RECT 91.760 114.480 92.985 114.620 ;
        RECT 91.760 114.420 92.080 114.480 ;
        RECT 92.695 114.435 92.985 114.480 ;
        RECT 108.320 114.620 108.640 114.680 ;
        RECT 113.470 114.620 113.610 115.160 ;
        RECT 118.455 115.115 118.745 115.160 ;
        RECT 119.820 115.100 120.140 115.160 ;
        RECT 120.295 115.115 120.585 115.160 ;
        RECT 127.155 115.300 127.445 115.345 ;
        RECT 128.345 115.300 128.635 115.345 ;
        RECT 130.865 115.300 131.155 115.345 ;
        RECT 127.155 115.160 131.155 115.300 ;
        RECT 127.155 115.115 127.445 115.160 ;
        RECT 128.345 115.115 128.635 115.160 ;
        RECT 130.865 115.115 131.155 115.160 ;
        RECT 134.080 115.100 134.400 115.360 ;
        RECT 126.760 114.960 127.050 115.005 ;
        RECT 128.860 114.960 129.150 115.005 ;
        RECT 130.430 114.960 130.720 115.005 ;
        RECT 126.760 114.820 130.720 114.960 ;
        RECT 126.760 114.775 127.050 114.820 ;
        RECT 128.860 114.775 129.150 114.820 ;
        RECT 130.430 114.775 130.720 114.820 ;
        RECT 136.930 114.680 137.070 115.840 ;
        RECT 138.220 115.780 138.540 115.840 ;
        RECT 139.140 115.640 139.460 115.700 ;
        RECT 144.290 115.685 144.430 115.840 ;
        RECT 149.720 115.780 150.040 115.840 ;
        RECT 154.320 115.780 154.640 115.840 ;
        RECT 137.850 115.500 139.460 115.640 ;
        RECT 137.850 115.360 137.990 115.500 ;
        RECT 139.140 115.440 139.460 115.500 ;
        RECT 139.615 115.640 139.905 115.685 ;
        RECT 139.615 115.500 143.510 115.640 ;
        RECT 139.615 115.455 139.905 115.500 ;
        RECT 137.315 115.300 137.605 115.345 ;
        RECT 137.760 115.300 138.080 115.360 ;
        RECT 137.315 115.160 138.080 115.300 ;
        RECT 137.315 115.115 137.605 115.160 ;
        RECT 137.760 115.100 138.080 115.160 ;
        RECT 138.235 115.300 138.525 115.345 ;
        RECT 142.835 115.300 143.125 115.345 ;
        RECT 138.235 115.160 143.125 115.300 ;
        RECT 138.235 115.115 138.525 115.160 ;
        RECT 142.835 115.115 143.125 115.160 ;
        RECT 143.370 114.960 143.510 115.500 ;
        RECT 144.215 115.455 144.505 115.685 ;
        RECT 145.495 115.640 145.785 115.685 ;
        RECT 144.750 115.500 145.785 115.640 ;
        RECT 143.740 115.300 144.060 115.360 ;
        RECT 144.750 115.300 144.890 115.500 ;
        RECT 145.495 115.455 145.785 115.500 ;
        RECT 152.020 115.440 152.340 115.700 ;
        RECT 143.740 115.160 144.890 115.300 ;
        RECT 145.095 115.300 145.385 115.345 ;
        RECT 146.285 115.300 146.575 115.345 ;
        RECT 148.805 115.300 149.095 115.345 ;
        RECT 145.095 115.160 149.095 115.300 ;
        RECT 143.740 115.100 144.060 115.160 ;
        RECT 145.095 115.115 145.385 115.160 ;
        RECT 146.285 115.115 146.575 115.160 ;
        RECT 148.805 115.115 149.095 115.160 ;
        RECT 144.700 114.960 144.990 115.005 ;
        RECT 146.800 114.960 147.090 115.005 ;
        RECT 148.370 114.960 148.660 115.005 ;
        RECT 143.370 114.820 144.430 114.960 ;
        RECT 144.290 114.680 144.430 114.820 ;
        RECT 144.700 114.820 148.660 114.960 ;
        RECT 144.700 114.775 144.990 114.820 ;
        RECT 146.800 114.775 147.090 114.820 ;
        RECT 148.370 114.775 148.660 114.820 ;
        RECT 108.320 114.480 113.610 114.620 ;
        RECT 108.320 114.420 108.640 114.480 ;
        RECT 115.220 114.420 115.540 114.680 ;
        RECT 115.680 114.420 116.000 114.680 ;
        RECT 136.840 114.420 137.160 114.680 ;
        RECT 138.680 114.620 139.000 114.680 ;
        RECT 140.075 114.620 140.365 114.665 ;
        RECT 138.680 114.480 140.365 114.620 ;
        RECT 138.680 114.420 139.000 114.480 ;
        RECT 140.075 114.435 140.365 114.480 ;
        RECT 144.200 114.420 144.520 114.680 ;
        RECT 22.690 113.800 157.010 114.280 ;
        RECT 36.560 113.600 36.880 113.660 ;
        RECT 40.240 113.600 40.560 113.660 ;
        RECT 57.260 113.600 57.580 113.660 ;
        RECT 26.990 113.460 57.580 113.600 ;
        RECT 25.980 112.380 26.300 112.640 ;
        RECT 26.990 112.625 27.130 113.460 ;
        RECT 36.560 113.400 36.880 113.460 ;
        RECT 40.240 113.400 40.560 113.460 ;
        RECT 57.260 113.400 57.580 113.460 ;
        RECT 62.320 113.600 62.640 113.660 ;
        RECT 65.555 113.600 65.845 113.645 ;
        RECT 62.320 113.460 65.845 113.600 ;
        RECT 62.320 113.400 62.640 113.460 ;
        RECT 65.555 113.415 65.845 113.460 ;
        RECT 82.100 113.400 82.420 113.660 ;
        RECT 88.540 113.400 88.860 113.660 ;
        RECT 109.700 113.400 110.020 113.660 ;
        RECT 115.235 113.600 115.525 113.645 ;
        RECT 117.520 113.600 117.840 113.660 ;
        RECT 126.260 113.600 126.580 113.660 ;
        RECT 115.235 113.460 117.840 113.600 ;
        RECT 115.235 113.415 115.525 113.460 ;
        RECT 117.520 113.400 117.840 113.460 ;
        RECT 125.430 113.460 126.580 113.600 ;
        RECT 33.340 113.260 33.660 113.320 ;
        RECT 29.290 113.120 33.660 113.260 ;
        RECT 26.915 112.395 27.205 112.625 ;
        RECT 28.740 112.380 29.060 112.640 ;
        RECT 29.290 112.625 29.430 113.120 ;
        RECT 33.340 113.060 33.660 113.120 ;
        RECT 34.720 113.060 35.040 113.320 ;
        RECT 41.635 113.260 41.925 113.305 ;
        RECT 44.840 113.260 45.160 113.320 ;
        RECT 40.330 113.120 45.160 113.260 ;
        RECT 34.275 112.920 34.565 112.965 ;
        RECT 34.810 112.920 34.950 113.060 ;
        RECT 34.275 112.780 34.950 112.920 ;
        RECT 34.275 112.735 34.565 112.780 ;
        RECT 29.215 112.395 29.505 112.625 ;
        RECT 29.675 112.580 29.965 112.625 ;
        RECT 30.595 112.580 30.885 112.625 ;
        RECT 32.420 112.580 32.740 112.640 ;
        RECT 29.675 112.440 30.350 112.580 ;
        RECT 29.675 112.395 29.965 112.440 ;
        RECT 25.075 112.240 25.365 112.285 ;
        RECT 25.075 112.100 29.430 112.240 ;
        RECT 25.075 112.055 25.365 112.100 ;
        RECT 27.360 111.700 27.680 111.960 ;
        RECT 29.290 111.900 29.430 112.100 ;
        RECT 30.210 111.900 30.350 112.440 ;
        RECT 30.595 112.440 32.740 112.580 ;
        RECT 30.595 112.395 30.885 112.440 ;
        RECT 32.420 112.380 32.740 112.440 ;
        RECT 33.340 112.580 33.660 112.640 ;
        RECT 40.330 112.580 40.470 113.120 ;
        RECT 41.635 113.075 41.925 113.120 ;
        RECT 44.840 113.060 45.160 113.120 ;
        RECT 47.180 113.260 47.470 113.305 ;
        RECT 49.280 113.260 49.570 113.305 ;
        RECT 50.850 113.260 51.140 113.305 ;
        RECT 47.180 113.120 51.140 113.260 ;
        RECT 47.180 113.075 47.470 113.120 ;
        RECT 49.280 113.075 49.570 113.120 ;
        RECT 50.850 113.075 51.140 113.120 ;
        RECT 54.540 113.260 54.830 113.305 ;
        RECT 56.640 113.260 56.930 113.305 ;
        RECT 58.210 113.260 58.500 113.305 ;
        RECT 54.540 113.120 58.500 113.260 ;
        RECT 54.540 113.075 54.830 113.120 ;
        RECT 56.640 113.075 56.930 113.120 ;
        RECT 58.210 113.075 58.500 113.120 ;
        RECT 60.955 113.260 61.245 113.305 ;
        RECT 70.180 113.260 70.470 113.305 ;
        RECT 72.280 113.260 72.570 113.305 ;
        RECT 73.850 113.260 74.140 113.305 ;
        RECT 60.955 113.120 68.530 113.260 ;
        RECT 60.955 113.075 61.245 113.120 ;
        RECT 42.080 112.920 42.400 112.980 ;
        RECT 44.380 112.920 44.700 112.980 ;
        RECT 68.390 112.965 68.530 113.120 ;
        RECT 70.180 113.120 74.140 113.260 ;
        RECT 70.180 113.075 70.470 113.120 ;
        RECT 72.280 113.075 72.570 113.120 ;
        RECT 73.850 113.075 74.140 113.120 ;
        RECT 79.430 113.120 86.010 113.260 ;
        RECT 46.695 112.920 46.985 112.965 ;
        RECT 42.080 112.780 46.985 112.920 ;
        RECT 42.080 112.720 42.400 112.780 ;
        RECT 44.380 112.720 44.700 112.780 ;
        RECT 46.695 112.735 46.985 112.780 ;
        RECT 47.575 112.920 47.865 112.965 ;
        RECT 48.765 112.920 49.055 112.965 ;
        RECT 51.285 112.920 51.575 112.965 ;
        RECT 47.575 112.780 51.575 112.920 ;
        RECT 47.575 112.735 47.865 112.780 ;
        RECT 48.765 112.735 49.055 112.780 ;
        RECT 51.285 112.735 51.575 112.780 ;
        RECT 54.935 112.920 55.225 112.965 ;
        RECT 56.125 112.920 56.415 112.965 ;
        RECT 58.645 112.920 58.935 112.965 ;
        RECT 54.935 112.780 58.935 112.920 ;
        RECT 54.935 112.735 55.225 112.780 ;
        RECT 56.125 112.735 56.415 112.780 ;
        RECT 58.645 112.735 58.935 112.780 ;
        RECT 68.315 112.735 68.605 112.965 ;
        RECT 70.575 112.920 70.865 112.965 ;
        RECT 71.765 112.920 72.055 112.965 ;
        RECT 74.285 112.920 74.575 112.965 ;
        RECT 70.575 112.780 74.575 112.920 ;
        RECT 70.575 112.735 70.865 112.780 ;
        RECT 71.765 112.735 72.055 112.780 ;
        RECT 74.285 112.735 74.575 112.780 ;
        RECT 75.200 112.720 75.520 112.980 ;
        RECT 79.430 112.965 79.570 113.120 ;
        RECT 79.355 112.735 79.645 112.965 ;
        RECT 79.815 112.920 80.105 112.965 ;
        RECT 81.640 112.920 81.960 112.980 ;
        RECT 85.870 112.965 86.010 113.120 ;
        RECT 79.815 112.780 81.960 112.920 ;
        RECT 79.815 112.735 80.105 112.780 ;
        RECT 81.640 112.720 81.960 112.780 ;
        RECT 85.795 112.920 86.085 112.965 ;
        RECT 88.630 112.920 88.770 113.400 ;
        RECT 89.040 113.260 89.330 113.305 ;
        RECT 91.140 113.260 91.430 113.305 ;
        RECT 92.710 113.260 93.000 113.305 ;
        RECT 89.040 113.120 93.000 113.260 ;
        RECT 89.040 113.075 89.330 113.120 ;
        RECT 91.140 113.075 91.430 113.120 ;
        RECT 92.710 113.075 93.000 113.120 ;
        RECT 95.915 113.075 96.205 113.305 ;
        RECT 115.680 113.260 116.000 113.320 ;
        RECT 110.710 113.120 116.000 113.260 ;
        RECT 85.795 112.780 88.770 112.920 ;
        RECT 89.435 112.920 89.725 112.965 ;
        RECT 90.625 112.920 90.915 112.965 ;
        RECT 93.145 112.920 93.435 112.965 ;
        RECT 89.435 112.780 93.435 112.920 ;
        RECT 85.795 112.735 86.085 112.780 ;
        RECT 89.435 112.735 89.725 112.780 ;
        RECT 90.625 112.735 90.915 112.780 ;
        RECT 93.145 112.735 93.435 112.780 ;
        RECT 93.600 112.720 93.920 112.980 ;
        RECT 33.340 112.440 40.470 112.580 ;
        RECT 33.340 112.380 33.660 112.440 ;
        RECT 40.715 112.395 41.005 112.625 ;
        RECT 40.790 111.960 40.930 112.395 ;
        RECT 42.540 112.380 42.860 112.640 ;
        RECT 43.000 112.380 43.320 112.640 ;
        RECT 54.055 112.580 54.345 112.625 ;
        RECT 57.720 112.580 58.040 112.640 ;
        RECT 54.055 112.440 58.040 112.580 ;
        RECT 54.055 112.395 54.345 112.440 ;
        RECT 57.720 112.380 58.040 112.440 ;
        RECT 63.255 112.395 63.545 112.625 ;
        RECT 46.235 112.240 46.525 112.285 ;
        RECT 47.920 112.240 48.210 112.285 ;
        RECT 46.235 112.100 48.210 112.240 ;
        RECT 46.235 112.055 46.525 112.100 ;
        RECT 47.920 112.055 48.210 112.100 ;
        RECT 55.390 112.240 55.680 112.285 ;
        RECT 58.640 112.240 58.960 112.300 ;
        RECT 55.390 112.100 58.960 112.240 ;
        RECT 63.330 112.240 63.470 112.395 ;
        RECT 63.700 112.380 64.020 112.640 ;
        RECT 64.160 112.380 64.480 112.640 ;
        RECT 65.095 112.580 65.385 112.625 ;
        RECT 65.540 112.580 65.860 112.640 ;
        RECT 65.095 112.440 65.860 112.580 ;
        RECT 65.095 112.395 65.385 112.440 ;
        RECT 65.540 112.380 65.860 112.440 ;
        RECT 66.460 112.380 66.780 112.640 ;
        RECT 69.695 112.580 69.985 112.625 ;
        RECT 75.290 112.580 75.430 112.720 ;
        RECT 69.695 112.440 75.430 112.580 ;
        RECT 69.695 112.395 69.985 112.440 ;
        RECT 77.055 112.395 77.345 112.625 ;
        RECT 66.550 112.240 66.690 112.380 ;
        RECT 63.330 112.100 66.690 112.240 ;
        RECT 71.030 112.240 71.320 112.285 ;
        RECT 71.520 112.240 71.840 112.300 ;
        RECT 71.030 112.100 71.840 112.240 ;
        RECT 77.130 112.240 77.270 112.395 ;
        RECT 80.260 112.380 80.580 112.640 ;
        RECT 84.400 112.380 84.720 112.640 ;
        RECT 88.555 112.580 88.845 112.625 ;
        RECT 92.220 112.580 92.540 112.640 ;
        RECT 93.690 112.580 93.830 112.720 ;
        RECT 95.990 112.580 96.130 113.075 ;
        RECT 98.660 112.720 98.980 112.980 ;
        RECT 104.640 112.920 104.960 112.980 ;
        RECT 107.875 112.920 108.165 112.965 ;
        RECT 108.320 112.920 108.640 112.980 ;
        RECT 104.640 112.780 108.640 112.920 ;
        RECT 104.640 112.720 104.960 112.780 ;
        RECT 107.875 112.735 108.165 112.780 ;
        RECT 108.320 112.720 108.640 112.780 ;
        RECT 88.555 112.440 93.830 112.580 ;
        RECT 94.150 112.440 96.130 112.580 ;
        RECT 98.215 112.580 98.505 112.625 ;
        RECT 102.800 112.580 103.120 112.640 ;
        RECT 110.710 112.625 110.850 113.120 ;
        RECT 115.680 113.060 116.000 113.120 ;
        RECT 118.900 113.260 119.190 113.305 ;
        RECT 120.470 113.260 120.760 113.305 ;
        RECT 122.570 113.260 122.860 113.305 ;
        RECT 118.900 113.120 122.860 113.260 ;
        RECT 118.900 113.075 119.190 113.120 ;
        RECT 120.470 113.075 120.760 113.120 ;
        RECT 122.570 113.075 122.860 113.120 ;
        RECT 115.220 112.720 115.540 112.980 ;
        RECT 125.430 112.965 125.570 113.460 ;
        RECT 126.260 113.400 126.580 113.460 ;
        RECT 134.080 113.400 134.400 113.660 ;
        RECT 134.540 113.600 134.860 113.660 ;
        RECT 135.475 113.600 135.765 113.645 ;
        RECT 134.540 113.460 135.765 113.600 ;
        RECT 134.540 113.400 134.860 113.460 ;
        RECT 135.475 113.415 135.765 113.460 ;
        RECT 136.395 113.600 136.685 113.645 ;
        RECT 137.300 113.600 137.620 113.660 ;
        RECT 136.395 113.460 137.620 113.600 ;
        RECT 136.395 113.415 136.685 113.460 ;
        RECT 125.840 113.260 126.130 113.305 ;
        RECT 127.940 113.260 128.230 113.305 ;
        RECT 129.510 113.260 129.800 113.305 ;
        RECT 125.840 113.120 129.800 113.260 ;
        RECT 125.840 113.075 126.130 113.120 ;
        RECT 127.940 113.075 128.230 113.120 ;
        RECT 129.510 113.075 129.800 113.120 ;
        RECT 132.255 113.260 132.545 113.305 ;
        RECT 134.170 113.260 134.310 113.400 ;
        RECT 132.255 113.120 134.310 113.260 ;
        RECT 132.255 113.075 132.545 113.120 ;
        RECT 118.465 112.920 118.755 112.965 ;
        RECT 120.985 112.920 121.275 112.965 ;
        RECT 122.175 112.920 122.465 112.965 ;
        RECT 118.465 112.780 122.465 112.920 ;
        RECT 118.465 112.735 118.755 112.780 ;
        RECT 120.985 112.735 121.275 112.780 ;
        RECT 122.175 112.735 122.465 112.780 ;
        RECT 123.055 112.920 123.345 112.965 ;
        RECT 125.355 112.920 125.645 112.965 ;
        RECT 123.055 112.780 125.645 112.920 ;
        RECT 123.055 112.735 123.345 112.780 ;
        RECT 125.355 112.735 125.645 112.780 ;
        RECT 126.235 112.920 126.525 112.965 ;
        RECT 127.425 112.920 127.715 112.965 ;
        RECT 129.945 112.920 130.235 112.965 ;
        RECT 126.235 112.780 130.235 112.920 ;
        RECT 126.235 112.735 126.525 112.780 ;
        RECT 127.425 112.735 127.715 112.780 ;
        RECT 129.945 112.735 130.235 112.780 ;
        RECT 107.415 112.580 107.705 112.625 ;
        RECT 98.215 112.440 107.705 112.580 ;
        RECT 88.555 112.395 88.845 112.440 ;
        RECT 92.220 112.380 92.540 112.440 ;
        RECT 89.890 112.240 90.180 112.285 ;
        RECT 90.840 112.240 91.160 112.300 ;
        RECT 77.130 112.100 82.100 112.240 ;
        RECT 55.390 112.055 55.680 112.100 ;
        RECT 58.640 112.040 58.960 112.100 ;
        RECT 71.030 112.055 71.320 112.100 ;
        RECT 71.520 112.040 71.840 112.100 ;
        RECT 29.290 111.760 30.350 111.900 ;
        RECT 30.580 111.900 30.900 111.960 ;
        RECT 31.055 111.900 31.345 111.945 ;
        RECT 33.800 111.900 34.120 111.960 ;
        RECT 30.580 111.760 34.120 111.900 ;
        RECT 30.580 111.700 30.900 111.760 ;
        RECT 31.055 111.715 31.345 111.760 ;
        RECT 33.800 111.700 34.120 111.760 ;
        RECT 36.100 111.900 36.420 111.960 ;
        RECT 37.495 111.900 37.785 111.945 ;
        RECT 36.100 111.760 37.785 111.900 ;
        RECT 36.100 111.700 36.420 111.760 ;
        RECT 37.495 111.715 37.785 111.760 ;
        RECT 40.700 111.700 41.020 111.960 ;
        RECT 52.660 111.900 52.980 111.960 ;
        RECT 53.595 111.900 53.885 111.945 ;
        RECT 52.660 111.760 53.885 111.900 ;
        RECT 52.660 111.700 52.980 111.760 ;
        RECT 53.595 111.715 53.885 111.760 ;
        RECT 61.860 111.700 62.180 111.960 ;
        RECT 76.120 111.900 76.440 111.960 ;
        RECT 76.595 111.900 76.885 111.945 ;
        RECT 76.120 111.760 76.885 111.900 ;
        RECT 76.120 111.700 76.440 111.760 ;
        RECT 76.595 111.715 76.885 111.760 ;
        RECT 77.960 111.700 78.280 111.960 ;
        RECT 81.960 111.900 82.100 112.100 ;
        RECT 89.890 112.100 91.160 112.240 ;
        RECT 89.890 112.055 90.180 112.100 ;
        RECT 90.840 112.040 91.160 112.100 ;
        RECT 91.300 112.240 91.620 112.300 ;
        RECT 94.150 112.240 94.290 112.440 ;
        RECT 98.215 112.395 98.505 112.440 ;
        RECT 102.800 112.380 103.120 112.440 ;
        RECT 107.415 112.395 107.705 112.440 ;
        RECT 110.635 112.395 110.925 112.625 ;
        RECT 111.080 112.580 111.400 112.640 ;
        RECT 113.380 112.580 113.700 112.640 ;
        RECT 111.080 112.440 113.700 112.580 ;
        RECT 111.080 112.380 111.400 112.440 ;
        RECT 113.380 112.380 113.700 112.440 ;
        RECT 114.315 112.580 114.605 112.625 ;
        RECT 115.310 112.580 115.450 112.720 ;
        RECT 114.315 112.440 115.450 112.580 ;
        RECT 121.660 112.625 121.980 112.640 ;
        RECT 114.315 112.395 114.605 112.440 ;
        RECT 121.660 112.395 122.010 112.625 ;
        RECT 126.690 112.580 126.980 112.625 ;
        RECT 132.700 112.580 133.020 112.640 ;
        RECT 134.170 112.625 134.310 113.120 ;
        RECT 126.690 112.440 133.020 112.580 ;
        RECT 126.690 112.395 126.980 112.440 ;
        RECT 121.660 112.380 121.980 112.395 ;
        RECT 132.700 112.380 133.020 112.440 ;
        RECT 134.095 112.395 134.385 112.625 ;
        RECT 134.555 112.580 134.845 112.625 ;
        RECT 134.555 112.440 135.230 112.580 ;
        RECT 134.555 112.395 134.845 112.440 ;
        RECT 135.090 112.300 135.230 112.440 ;
        RECT 91.300 112.100 94.290 112.240 ;
        RECT 94.980 112.240 95.300 112.300 ;
        RECT 97.755 112.240 98.045 112.285 ;
        RECT 94.980 112.100 98.045 112.240 ;
        RECT 91.300 112.040 91.620 112.100 ;
        RECT 94.980 112.040 95.300 112.100 ;
        RECT 97.755 112.055 98.045 112.100 ;
        RECT 135.000 112.040 135.320 112.300 ;
        RECT 135.550 112.240 135.690 113.415 ;
        RECT 137.300 113.400 137.620 113.460 ;
        RECT 139.615 113.600 139.905 113.645 ;
        RECT 142.820 113.600 143.140 113.660 ;
        RECT 139.615 113.460 143.140 113.600 ;
        RECT 139.615 113.415 139.905 113.460 ;
        RECT 142.820 113.400 143.140 113.460 ;
        RECT 143.740 113.400 144.060 113.660 ;
        RECT 144.215 113.600 144.505 113.645 ;
        RECT 144.660 113.600 144.980 113.660 ;
        RECT 144.215 113.460 144.980 113.600 ;
        RECT 144.215 113.415 144.505 113.460 ;
        RECT 144.660 113.400 144.980 113.460 ;
        RECT 153.875 113.600 154.165 113.645 ;
        RECT 154.320 113.600 154.640 113.660 ;
        RECT 153.875 113.460 154.640 113.600 ;
        RECT 153.875 113.415 154.165 113.460 ;
        RECT 154.320 113.400 154.640 113.460 ;
        RECT 137.760 113.260 138.080 113.320 ;
        RECT 137.760 113.120 138.450 113.260 ;
        RECT 137.760 113.060 138.080 113.120 ;
        RECT 136.840 112.920 137.160 112.980 ;
        RECT 138.310 112.920 138.450 113.120 ;
        RECT 144.660 112.920 144.980 112.980 ;
        RECT 136.010 112.780 137.990 112.920 ;
        RECT 138.310 112.780 140.750 112.920 ;
        RECT 136.010 112.625 136.150 112.780 ;
        RECT 136.840 112.720 137.160 112.780 ;
        RECT 137.850 112.640 137.990 112.780 ;
        RECT 135.935 112.395 136.225 112.625 ;
        RECT 137.315 112.580 137.605 112.625 ;
        RECT 136.470 112.440 137.605 112.580 ;
        RECT 136.470 112.240 136.610 112.440 ;
        RECT 137.315 112.395 137.605 112.440 ;
        RECT 137.760 112.380 138.080 112.640 ;
        RECT 140.610 112.625 140.750 112.780 ;
        RECT 141.530 112.780 144.980 112.920 ;
        RECT 141.530 112.625 141.670 112.780 ;
        RECT 144.660 112.720 144.980 112.780 ;
        RECT 139.155 112.395 139.445 112.625 ;
        RECT 140.075 112.580 140.365 112.625 ;
        RECT 139.690 112.440 140.365 112.580 ;
        RECT 135.550 112.100 136.610 112.240 ;
        RECT 136.840 112.240 137.160 112.300 ;
        RECT 139.230 112.240 139.370 112.395 ;
        RECT 136.840 112.100 139.370 112.240 ;
        RECT 136.840 112.040 137.160 112.100 ;
        RECT 82.575 111.900 82.865 111.945 ;
        RECT 81.960 111.760 82.865 111.900 ;
        RECT 82.575 111.715 82.865 111.760 ;
        RECT 84.860 111.700 85.180 111.960 ;
        RECT 95.440 111.700 95.760 111.960 ;
        RECT 102.800 111.900 103.120 111.960 ;
        RECT 105.115 111.900 105.405 111.945 ;
        RECT 102.800 111.760 105.405 111.900 ;
        RECT 102.800 111.700 103.120 111.760 ;
        RECT 105.115 111.715 105.405 111.760 ;
        RECT 106.940 111.700 107.260 111.960 ;
        RECT 116.140 111.700 116.460 111.960 ;
        RECT 133.175 111.900 133.465 111.945 ;
        RECT 136.380 111.900 136.700 111.960 ;
        RECT 139.690 111.900 139.830 112.440 ;
        RECT 140.075 112.395 140.365 112.440 ;
        RECT 140.535 112.395 140.825 112.625 ;
        RECT 141.455 112.395 141.745 112.625 ;
        RECT 141.915 112.395 142.205 112.625 ;
        RECT 142.375 112.395 142.665 112.625 ;
        RECT 145.580 112.580 145.900 112.640 ;
        RECT 146.055 112.580 146.345 112.625 ;
        RECT 145.580 112.440 146.345 112.580 ;
        RECT 133.175 111.760 139.830 111.900 ;
        RECT 141.990 111.900 142.130 112.395 ;
        RECT 142.450 112.240 142.590 112.395 ;
        RECT 145.580 112.380 145.900 112.440 ;
        RECT 146.055 112.395 146.345 112.440 ;
        RECT 142.450 112.100 143.510 112.240 ;
        RECT 143.370 111.960 143.510 112.100 ;
        RECT 145.120 112.040 145.440 112.300 ;
        RECT 146.515 112.055 146.805 112.285 ;
        RECT 142.360 111.900 142.680 111.960 ;
        RECT 141.990 111.760 142.680 111.900 ;
        RECT 133.175 111.715 133.465 111.760 ;
        RECT 136.380 111.700 136.700 111.760 ;
        RECT 142.360 111.700 142.680 111.760 ;
        RECT 143.280 111.700 143.600 111.960 ;
        RECT 143.740 111.900 144.060 111.960 ;
        RECT 146.590 111.900 146.730 112.055 ;
        RECT 143.740 111.760 146.730 111.900 ;
        RECT 143.740 111.700 144.060 111.760 ;
        RECT 22.690 111.080 157.810 111.560 ;
        RECT 28.740 110.880 29.060 110.940 ;
        RECT 30.580 110.880 30.900 110.940 ;
        RECT 28.740 110.740 30.900 110.880 ;
        RECT 28.740 110.680 29.060 110.740 ;
        RECT 30.580 110.680 30.900 110.740 ;
        RECT 31.055 110.880 31.345 110.925 ;
        RECT 34.720 110.880 35.040 110.940 ;
        RECT 31.055 110.740 35.040 110.880 ;
        RECT 31.055 110.695 31.345 110.740 ;
        RECT 34.720 110.680 35.040 110.740 ;
        RECT 43.000 110.680 43.320 110.940 ;
        RECT 54.500 110.880 54.820 110.940 ;
        RECT 55.435 110.880 55.725 110.925 ;
        RECT 54.500 110.740 55.725 110.880 ;
        RECT 54.500 110.680 54.820 110.740 ;
        RECT 55.435 110.695 55.725 110.740 ;
        RECT 58.640 110.680 58.960 110.940 ;
        RECT 61.860 110.680 62.180 110.940 ;
        RECT 63.700 110.680 64.020 110.940 ;
        RECT 64.160 110.880 64.480 110.940 ;
        RECT 64.635 110.880 64.925 110.925 ;
        RECT 64.160 110.740 64.925 110.880 ;
        RECT 64.160 110.680 64.480 110.740 ;
        RECT 64.635 110.695 64.925 110.740 ;
        RECT 67.840 110.680 68.160 110.940 ;
        RECT 69.235 110.880 69.525 110.925 ;
        RECT 70.140 110.880 70.460 110.940 ;
        RECT 69.235 110.740 70.460 110.880 ;
        RECT 69.235 110.695 69.525 110.740 ;
        RECT 70.140 110.680 70.460 110.740 ;
        RECT 84.860 110.880 85.180 110.940 ;
        RECT 87.175 110.880 87.465 110.925 ;
        RECT 84.860 110.740 87.465 110.880 ;
        RECT 84.860 110.680 85.180 110.740 ;
        RECT 87.175 110.695 87.465 110.740 ;
        RECT 90.395 110.880 90.685 110.925 ;
        RECT 90.840 110.880 91.160 110.940 ;
        RECT 92.680 110.880 93.000 110.940 ;
        RECT 90.395 110.740 91.160 110.880 ;
        RECT 90.395 110.695 90.685 110.740 ;
        RECT 90.840 110.680 91.160 110.740 ;
        RECT 92.310 110.740 93.000 110.880 ;
        RECT 41.635 110.540 41.925 110.585 ;
        RECT 43.920 110.540 44.240 110.600 ;
        RECT 49.455 110.540 49.745 110.585 ;
        RECT 56.815 110.540 57.105 110.585 ;
        RECT 33.660 110.400 41.390 110.540 ;
        RECT 25.520 110.245 25.840 110.260 ;
        RECT 25.490 110.015 25.840 110.245 ;
        RECT 32.895 110.200 33.185 110.245 ;
        RECT 33.660 110.200 33.800 110.400 ;
        RECT 41.250 110.260 41.390 110.400 ;
        RECT 41.635 110.400 44.240 110.540 ;
        RECT 41.635 110.355 41.925 110.400 ;
        RECT 43.920 110.340 44.240 110.400 ;
        RECT 44.470 110.400 57.105 110.540 ;
        RECT 34.720 110.245 35.040 110.260 ;
        RECT 32.895 110.060 33.800 110.200 ;
        RECT 32.895 110.015 33.185 110.060 ;
        RECT 34.690 110.015 35.040 110.245 ;
        RECT 25.520 110.000 25.840 110.015 ;
        RECT 34.720 110.000 35.040 110.015 ;
        RECT 40.240 110.200 40.560 110.260 ;
        RECT 40.715 110.200 41.005 110.245 ;
        RECT 40.240 110.060 41.005 110.200 ;
        RECT 40.240 110.000 40.560 110.060 ;
        RECT 40.715 110.015 41.005 110.060 ;
        RECT 41.160 110.000 41.480 110.260 ;
        RECT 44.470 110.245 44.610 110.400 ;
        RECT 49.455 110.355 49.745 110.400 ;
        RECT 56.815 110.355 57.105 110.400 ;
        RECT 57.260 110.540 57.580 110.600 ;
        RECT 57.735 110.540 58.025 110.585 ;
        RECT 57.260 110.400 58.025 110.540 ;
        RECT 57.260 110.340 57.580 110.400 ;
        RECT 57.735 110.355 58.025 110.400 ;
        RECT 44.395 110.015 44.685 110.245 ;
        RECT 44.840 110.000 45.160 110.260 ;
        RECT 45.315 110.015 45.605 110.245 ;
        RECT 46.235 110.200 46.525 110.245 ;
        RECT 47.140 110.200 47.460 110.260 ;
        RECT 46.235 110.060 47.460 110.200 ;
        RECT 46.235 110.015 46.525 110.060 ;
        RECT 24.155 109.675 24.445 109.905 ;
        RECT 25.035 109.860 25.325 109.905 ;
        RECT 26.225 109.860 26.515 109.905 ;
        RECT 28.745 109.860 29.035 109.905 ;
        RECT 33.355 109.860 33.645 109.905 ;
        RECT 25.035 109.720 29.035 109.860 ;
        RECT 25.035 109.675 25.325 109.720 ;
        RECT 26.225 109.675 26.515 109.720 ;
        RECT 28.745 109.675 29.035 109.720 ;
        RECT 30.670 109.720 33.645 109.860 ;
        RECT 24.230 109.180 24.370 109.675 ;
        RECT 24.640 109.520 24.930 109.565 ;
        RECT 26.740 109.520 27.030 109.565 ;
        RECT 28.310 109.520 28.600 109.565 ;
        RECT 24.640 109.380 28.600 109.520 ;
        RECT 24.640 109.335 24.930 109.380 ;
        RECT 26.740 109.335 27.030 109.380 ;
        RECT 28.310 109.335 28.600 109.380 ;
        RECT 30.670 109.240 30.810 109.720 ;
        RECT 33.355 109.675 33.645 109.720 ;
        RECT 34.235 109.860 34.525 109.905 ;
        RECT 35.425 109.860 35.715 109.905 ;
        RECT 37.945 109.860 38.235 109.905 ;
        RECT 34.235 109.720 38.235 109.860 ;
        RECT 34.235 109.675 34.525 109.720 ;
        RECT 35.425 109.675 35.715 109.720 ;
        RECT 37.945 109.675 38.235 109.720 ;
        RECT 42.555 109.860 42.845 109.905 ;
        RECT 45.390 109.860 45.530 110.015 ;
        RECT 47.140 110.000 47.460 110.060 ;
        RECT 52.660 110.000 52.980 110.260 ;
        RECT 53.120 110.000 53.440 110.260 ;
        RECT 53.580 110.000 53.900 110.260 ;
        RECT 54.040 110.000 54.360 110.260 ;
        RECT 54.500 110.000 54.820 110.260 ;
        RECT 61.950 110.245 62.090 110.680 ;
        RECT 63.790 110.540 63.930 110.680 ;
        RECT 65.555 110.540 65.845 110.585 ;
        RECT 63.790 110.400 65.845 110.540 ;
        RECT 65.555 110.355 65.845 110.400 ;
        RECT 61.875 110.015 62.165 110.245 ;
        RECT 62.335 110.200 62.625 110.245 ;
        RECT 63.240 110.200 63.560 110.260 ;
        RECT 62.335 110.060 63.560 110.200 ;
        RECT 62.335 110.015 62.625 110.060 ;
        RECT 63.240 110.000 63.560 110.060 ;
        RECT 64.620 110.200 64.940 110.260 ;
        RECT 65.095 110.200 65.385 110.245 ;
        RECT 64.620 110.060 65.385 110.200 ;
        RECT 64.620 110.000 64.940 110.060 ;
        RECT 65.095 110.015 65.385 110.060 ;
        RECT 67.395 110.015 67.685 110.245 ;
        RECT 42.555 109.720 45.530 109.860 ;
        RECT 42.555 109.675 42.845 109.720 ;
        RECT 31.975 109.520 32.265 109.565 ;
        RECT 32.420 109.520 32.740 109.580 ;
        RECT 31.975 109.380 32.740 109.520 ;
        RECT 31.975 109.335 32.265 109.380 ;
        RECT 32.420 109.320 32.740 109.380 ;
        RECT 33.840 109.520 34.130 109.565 ;
        RECT 35.940 109.520 36.230 109.565 ;
        RECT 37.510 109.520 37.800 109.565 ;
        RECT 33.840 109.380 37.800 109.520 ;
        RECT 33.840 109.335 34.130 109.380 ;
        RECT 35.940 109.335 36.230 109.380 ;
        RECT 37.510 109.335 37.800 109.380 ;
        RECT 40.255 109.520 40.545 109.565 ;
        RECT 40.700 109.520 41.020 109.580 ;
        RECT 40.255 109.380 50.590 109.520 ;
        RECT 40.255 109.335 40.545 109.380 ;
        RECT 40.700 109.320 41.020 109.380 ;
        RECT 50.450 109.240 50.590 109.380 ;
        RECT 30.580 109.180 30.900 109.240 ;
        RECT 24.230 109.040 30.900 109.180 ;
        RECT 30.580 108.980 30.900 109.040 ;
        RECT 50.360 108.980 50.680 109.240 ;
        RECT 52.750 109.180 52.890 110.000 ;
        RECT 53.670 109.860 53.810 110.000 ;
        RECT 55.895 109.860 56.185 109.905 ;
        RECT 53.670 109.720 56.185 109.860 ;
        RECT 55.895 109.675 56.185 109.720 ;
        RECT 67.470 109.520 67.610 110.015 ;
        RECT 67.930 109.905 68.070 110.680 ;
        RECT 68.300 110.540 68.620 110.600 ;
        RECT 71.075 110.540 71.365 110.585 ;
        RECT 68.300 110.400 71.365 110.540 ;
        RECT 68.300 110.340 68.620 110.400 ;
        RECT 71.075 110.355 71.365 110.400 ;
        RECT 77.960 110.540 78.280 110.600 ;
        RECT 80.580 110.540 80.870 110.585 ;
        RECT 92.310 110.540 92.450 110.740 ;
        RECT 92.680 110.680 93.000 110.740 ;
        RECT 94.980 110.680 95.300 110.940 ;
        RECT 95.440 110.680 95.760 110.940 ;
        RECT 102.800 110.680 103.120 110.940 ;
        RECT 103.275 110.695 103.565 110.925 ;
        RECT 106.940 110.880 107.260 110.940 ;
        RECT 111.095 110.880 111.385 110.925 ;
        RECT 106.940 110.740 111.385 110.880 ;
        RECT 77.960 110.400 80.870 110.540 ;
        RECT 77.960 110.340 78.280 110.400 ;
        RECT 80.580 110.355 80.870 110.400 ;
        RECT 90.930 110.400 92.450 110.540 ;
        RECT 90.930 110.260 91.070 110.400 ;
        RECT 68.760 110.200 69.080 110.260 ;
        RECT 69.695 110.200 69.985 110.245 ;
        RECT 68.760 110.060 69.985 110.200 ;
        RECT 68.760 110.000 69.080 110.060 ;
        RECT 69.695 110.015 69.985 110.060 ;
        RECT 70.140 110.000 70.460 110.260 ;
        RECT 75.675 110.200 75.965 110.245 ;
        RECT 76.120 110.200 76.440 110.260 ;
        RECT 75.675 110.060 76.440 110.200 ;
        RECT 75.675 110.015 75.965 110.060 ;
        RECT 76.120 110.000 76.440 110.060 ;
        RECT 79.340 110.245 79.660 110.260 ;
        RECT 79.340 110.200 79.680 110.245 ;
        RECT 88.095 110.200 88.385 110.245 ;
        RECT 79.340 110.060 79.855 110.200 ;
        RECT 86.330 110.060 88.385 110.200 ;
        RECT 79.340 110.015 79.680 110.060 ;
        RECT 79.340 110.000 79.660 110.015 ;
        RECT 67.855 109.675 68.145 109.905 ;
        RECT 76.595 109.675 76.885 109.905 ;
        RECT 80.235 109.860 80.525 109.905 ;
        RECT 81.425 109.860 81.715 109.905 ;
        RECT 83.945 109.860 84.235 109.905 ;
        RECT 80.235 109.720 84.235 109.860 ;
        RECT 80.235 109.675 80.525 109.720 ;
        RECT 81.425 109.675 81.715 109.720 ;
        RECT 83.945 109.675 84.235 109.720 ;
        RECT 75.200 109.520 75.520 109.580 ;
        RECT 76.670 109.520 76.810 109.675 ;
        RECT 67.470 109.380 76.810 109.520 ;
        RECT 79.840 109.520 80.130 109.565 ;
        RECT 81.940 109.520 82.230 109.565 ;
        RECT 83.510 109.520 83.800 109.565 ;
        RECT 79.840 109.380 83.800 109.520 ;
        RECT 75.200 109.320 75.520 109.380 ;
        RECT 79.840 109.335 80.130 109.380 ;
        RECT 81.940 109.335 82.230 109.380 ;
        RECT 83.510 109.335 83.800 109.380 ;
        RECT 53.135 109.180 53.425 109.225 ;
        RECT 52.750 109.040 53.425 109.180 ;
        RECT 53.135 108.995 53.425 109.040 ;
        RECT 62.320 109.180 62.640 109.240 ;
        RECT 62.795 109.180 63.085 109.225 ;
        RECT 62.320 109.040 63.085 109.180 ;
        RECT 62.320 108.980 62.640 109.040 ;
        RECT 62.795 108.995 63.085 109.040 ;
        RECT 66.920 109.180 67.240 109.240 ;
        RECT 68.760 109.180 69.080 109.240 ;
        RECT 66.920 109.040 69.080 109.180 ;
        RECT 66.920 108.980 67.240 109.040 ;
        RECT 68.760 108.980 69.080 109.040 ;
        RECT 71.060 108.980 71.380 109.240 ;
        RECT 84.860 109.180 85.180 109.240 ;
        RECT 86.330 109.225 86.470 110.060 ;
        RECT 88.095 110.015 88.385 110.060 ;
        RECT 89.015 110.015 89.305 110.245 ;
        RECT 89.090 109.520 89.230 110.015 ;
        RECT 90.840 110.000 91.160 110.260 ;
        RECT 91.300 110.000 91.620 110.260 ;
        RECT 91.775 110.200 92.065 110.245 ;
        RECT 92.310 110.200 92.450 110.400 ;
        RECT 91.775 110.060 92.450 110.200 ;
        RECT 92.695 110.200 92.985 110.245 ;
        RECT 94.075 110.200 94.365 110.245 ;
        RECT 95.530 110.200 95.670 110.680 ;
        RECT 92.695 110.060 95.670 110.200 ;
        RECT 102.355 110.200 102.645 110.245 ;
        RECT 102.890 110.200 103.030 110.680 ;
        RECT 103.350 110.540 103.490 110.695 ;
        RECT 106.940 110.680 107.260 110.740 ;
        RECT 111.095 110.695 111.385 110.740 ;
        RECT 118.900 110.680 119.220 110.940 ;
        RECT 134.080 110.680 134.400 110.940 ;
        RECT 137.760 110.880 138.080 110.940 ;
        RECT 149.735 110.880 150.025 110.925 ;
        RECT 137.760 110.740 150.025 110.880 ;
        RECT 137.760 110.680 138.080 110.740 ;
        RECT 149.735 110.695 150.025 110.740 ;
        RECT 104.960 110.540 105.250 110.585 ;
        RECT 103.350 110.400 105.250 110.540 ;
        RECT 104.960 110.355 105.250 110.400 ;
        RECT 116.140 110.540 116.460 110.600 ;
        RECT 134.170 110.540 134.310 110.680 ;
        RECT 116.140 110.400 118.210 110.540 ;
        RECT 116.140 110.340 116.460 110.400 ;
        RECT 112.000 110.200 112.320 110.260 ;
        RECT 118.070 110.245 118.210 110.400 ;
        RECT 133.250 110.400 134.310 110.540 ;
        RECT 134.555 110.540 134.845 110.585 ;
        RECT 137.300 110.540 137.620 110.600 ;
        RECT 134.555 110.400 137.620 110.540 ;
        RECT 133.250 110.245 133.390 110.400 ;
        RECT 134.555 110.355 134.845 110.400 ;
        RECT 137.300 110.340 137.620 110.400 ;
        RECT 138.680 110.540 139.000 110.600 ;
        RECT 139.460 110.540 139.750 110.585 ;
        RECT 138.680 110.400 139.750 110.540 ;
        RECT 138.680 110.340 139.000 110.400 ;
        RECT 139.460 110.355 139.750 110.400 ;
        RECT 102.355 110.060 103.030 110.200 ;
        RECT 110.710 110.060 112.320 110.200 ;
        RECT 91.775 110.015 92.065 110.060 ;
        RECT 92.695 110.015 92.985 110.060 ;
        RECT 94.075 110.015 94.365 110.060 ;
        RECT 102.355 110.015 102.645 110.060 ;
        RECT 93.155 109.860 93.445 109.905 ;
        RECT 103.260 109.860 103.580 109.920 ;
        RECT 103.735 109.860 104.025 109.905 ;
        RECT 93.155 109.720 94.290 109.860 ;
        RECT 93.155 109.675 93.445 109.720 ;
        RECT 94.150 109.580 94.290 109.720 ;
        RECT 103.260 109.720 104.025 109.860 ;
        RECT 103.260 109.660 103.580 109.720 ;
        RECT 103.735 109.675 104.025 109.720 ;
        RECT 104.615 109.860 104.905 109.905 ;
        RECT 105.805 109.860 106.095 109.905 ;
        RECT 108.325 109.860 108.615 109.905 ;
        RECT 104.615 109.720 108.615 109.860 ;
        RECT 104.615 109.675 104.905 109.720 ;
        RECT 105.805 109.675 106.095 109.720 ;
        RECT 108.325 109.675 108.615 109.720 ;
        RECT 94.060 109.520 94.380 109.580 ;
        RECT 110.710 109.565 110.850 110.060 ;
        RECT 112.000 110.000 112.320 110.060 ;
        RECT 117.995 110.015 118.285 110.245 ;
        RECT 133.175 110.015 133.465 110.245 ;
        RECT 133.635 110.200 133.925 110.245 ;
        RECT 135.000 110.200 135.320 110.260 ;
        RECT 137.775 110.200 138.065 110.245 ;
        RECT 146.500 110.200 146.820 110.260 ;
        RECT 133.635 110.060 137.530 110.200 ;
        RECT 133.635 110.015 133.925 110.060 ;
        RECT 135.000 110.000 135.320 110.060 ;
        RECT 111.080 109.860 111.400 109.920 ;
        RECT 112.935 109.860 113.225 109.905 ;
        RECT 117.060 109.860 117.380 109.920 ;
        RECT 137.390 109.905 137.530 110.060 ;
        RECT 137.775 110.060 146.820 110.200 ;
        RECT 137.775 110.015 138.065 110.060 ;
        RECT 146.500 110.000 146.820 110.060 ;
        RECT 148.815 110.200 149.105 110.245 ;
        RECT 149.275 110.200 149.565 110.245 ;
        RECT 148.815 110.060 149.565 110.200 ;
        RECT 148.815 110.015 149.105 110.060 ;
        RECT 149.275 110.015 149.565 110.060 ;
        RECT 111.080 109.720 117.380 109.860 ;
        RECT 111.080 109.660 111.400 109.720 ;
        RECT 112.935 109.675 113.225 109.720 ;
        RECT 117.060 109.660 117.380 109.720 ;
        RECT 137.315 109.675 137.605 109.905 ;
        RECT 138.220 109.660 138.540 109.920 ;
        RECT 139.115 109.860 139.405 109.905 ;
        RECT 140.305 109.860 140.595 109.905 ;
        RECT 142.825 109.860 143.115 109.905 ;
        RECT 139.115 109.720 143.115 109.860 ;
        RECT 139.115 109.675 139.405 109.720 ;
        RECT 140.305 109.675 140.595 109.720 ;
        RECT 142.825 109.675 143.115 109.720 ;
        RECT 145.595 109.675 145.885 109.905 ;
        RECT 89.090 109.380 94.380 109.520 ;
        RECT 94.060 109.320 94.380 109.380 ;
        RECT 104.220 109.520 104.510 109.565 ;
        RECT 106.320 109.520 106.610 109.565 ;
        RECT 107.890 109.520 108.180 109.565 ;
        RECT 104.220 109.380 108.180 109.520 ;
        RECT 104.220 109.335 104.510 109.380 ;
        RECT 106.320 109.335 106.610 109.380 ;
        RECT 107.890 109.335 108.180 109.380 ;
        RECT 110.635 109.335 110.925 109.565 ;
        RECT 134.555 109.520 134.845 109.565 ;
        RECT 136.840 109.520 137.160 109.580 ;
        RECT 134.555 109.380 137.160 109.520 ;
        RECT 134.555 109.335 134.845 109.380 ;
        RECT 136.840 109.320 137.160 109.380 ;
        RECT 138.720 109.520 139.010 109.565 ;
        RECT 140.820 109.520 141.110 109.565 ;
        RECT 142.390 109.520 142.680 109.565 ;
        RECT 138.720 109.380 142.680 109.520 ;
        RECT 138.720 109.335 139.010 109.380 ;
        RECT 140.820 109.335 141.110 109.380 ;
        RECT 142.390 109.335 142.680 109.380 ;
        RECT 145.135 109.520 145.425 109.565 ;
        RECT 145.670 109.520 145.810 109.675 ;
        RECT 145.135 109.380 145.810 109.520 ;
        RECT 145.135 109.335 145.425 109.380 ;
        RECT 86.255 109.180 86.545 109.225 ;
        RECT 84.860 109.040 86.545 109.180 ;
        RECT 84.860 108.980 85.180 109.040 ;
        RECT 86.255 108.995 86.545 109.040 ;
        RECT 91.300 109.180 91.620 109.240 ;
        RECT 92.695 109.180 92.985 109.225 ;
        RECT 91.300 109.040 92.985 109.180 ;
        RECT 91.300 108.980 91.620 109.040 ;
        RECT 92.695 108.995 92.985 109.040 ;
        RECT 22.690 108.360 157.010 108.840 ;
        RECT 25.520 108.160 25.840 108.220 ;
        RECT 27.375 108.160 27.665 108.205 ;
        RECT 25.520 108.020 27.665 108.160 ;
        RECT 25.520 107.960 25.840 108.020 ;
        RECT 27.375 107.975 27.665 108.020 ;
        RECT 28.280 107.960 28.600 108.220 ;
        RECT 44.840 108.160 45.160 108.220 ;
        RECT 53.580 108.160 53.900 108.220 ;
        RECT 44.840 108.020 53.900 108.160 ;
        RECT 44.840 107.960 45.160 108.020 ;
        RECT 53.580 107.960 53.900 108.020 ;
        RECT 54.040 108.160 54.360 108.220 ;
        RECT 59.575 108.160 59.865 108.205 ;
        RECT 54.040 108.020 59.865 108.160 ;
        RECT 54.040 107.960 54.360 108.020 ;
        RECT 59.575 107.975 59.865 108.020 ;
        RECT 67.855 108.160 68.145 108.205 ;
        RECT 70.140 108.160 70.460 108.220 ;
        RECT 67.855 108.020 70.460 108.160 ;
        RECT 67.855 107.975 68.145 108.020 ;
        RECT 26.915 107.820 27.205 107.865 ;
        RECT 28.370 107.820 28.510 107.960 ;
        RECT 47.600 107.820 47.920 107.880 ;
        RECT 48.980 107.820 49.300 107.880 ;
        RECT 26.915 107.680 28.510 107.820 ;
        RECT 36.190 107.680 47.920 107.820 ;
        RECT 26.915 107.635 27.205 107.680 ;
        RECT 27.360 107.480 27.680 107.540 ;
        RECT 30.135 107.480 30.425 107.525 ;
        RECT 27.360 107.340 30.425 107.480 ;
        RECT 27.360 107.280 27.680 107.340 ;
        RECT 30.135 107.295 30.425 107.340 ;
        RECT 25.060 106.940 25.380 107.200 ;
        RECT 25.980 106.940 26.300 107.200 ;
        RECT 35.195 106.955 35.485 107.185 ;
        RECT 36.190 107.140 36.330 107.680 ;
        RECT 47.600 107.620 47.920 107.680 ;
        RECT 48.610 107.680 49.300 107.820 ;
        RECT 36.560 107.480 36.880 107.540 ;
        RECT 48.610 107.525 48.750 107.680 ;
        RECT 48.980 107.620 49.300 107.680 ;
        RECT 51.280 107.820 51.600 107.880 ;
        RECT 51.280 107.680 58.870 107.820 ;
        RECT 51.280 107.620 51.600 107.680 ;
        RECT 41.175 107.480 41.465 107.525 ;
        RECT 44.395 107.480 44.685 107.525 ;
        RECT 36.560 107.340 38.170 107.480 ;
        RECT 36.560 107.280 36.880 107.340 ;
        RECT 38.030 107.185 38.170 107.340 ;
        RECT 41.175 107.340 44.685 107.480 ;
        RECT 41.175 107.295 41.465 107.340 ;
        RECT 44.395 107.295 44.685 107.340 ;
        RECT 48.535 107.295 48.825 107.525 ;
        RECT 53.670 107.480 55.190 107.520 ;
        RECT 51.830 107.380 55.190 107.480 ;
        RECT 51.830 107.340 53.810 107.380 ;
        RECT 37.035 107.140 37.325 107.185 ;
        RECT 36.190 107.000 37.325 107.140 ;
        RECT 37.035 106.955 37.325 107.000 ;
        RECT 37.955 106.955 38.245 107.185 ;
        RECT 35.270 106.520 35.410 106.955 ;
        RECT 38.400 106.940 38.720 107.200 ;
        RECT 38.875 106.955 39.165 107.185 ;
        RECT 37.480 106.800 37.800 106.860 ;
        RECT 38.950 106.800 39.090 106.955 ;
        RECT 44.840 106.940 45.160 107.200 ;
        RECT 45.760 106.940 46.080 107.200 ;
        RECT 46.235 106.955 46.525 107.185 ;
        RECT 46.695 106.955 46.985 107.185 ;
        RECT 47.600 107.140 47.920 107.200 ;
        RECT 51.830 107.140 51.970 107.340 ;
        RECT 47.600 107.000 51.970 107.140 ;
        RECT 52.660 107.140 52.980 107.200 ;
        RECT 53.135 107.140 53.425 107.185 ;
        RECT 52.660 107.000 53.425 107.140 ;
        RECT 37.480 106.660 39.090 106.800 ;
        RECT 44.930 106.800 45.070 106.940 ;
        RECT 46.310 106.800 46.450 106.955 ;
        RECT 44.930 106.660 46.450 106.800 ;
        RECT 46.770 106.800 46.910 106.955 ;
        RECT 47.600 106.940 47.920 107.000 ;
        RECT 52.660 106.940 52.980 107.000 ;
        RECT 53.135 106.955 53.425 107.000 ;
        RECT 53.580 106.940 53.900 107.200 ;
        RECT 54.040 106.940 54.360 107.200 ;
        RECT 55.050 107.185 55.190 107.380 ;
        RECT 54.975 106.955 55.265 107.185 ;
        RECT 57.260 107.140 57.580 107.200 ;
        RECT 58.730 107.185 58.870 107.680 ;
        RECT 66.015 107.480 66.305 107.525 ;
        RECT 65.630 107.340 66.305 107.480 ;
        RECT 65.630 107.200 65.770 107.340 ;
        RECT 66.015 107.295 66.305 107.340 ;
        RECT 57.735 107.140 58.025 107.185 ;
        RECT 57.260 107.000 58.025 107.140 ;
        RECT 57.260 106.940 57.580 107.000 ;
        RECT 57.735 106.955 58.025 107.000 ;
        RECT 58.655 106.955 58.945 107.185 ;
        RECT 60.940 106.940 61.260 107.200 ;
        RECT 65.540 106.940 65.860 107.200 ;
        RECT 66.920 106.940 67.240 107.200 ;
        RECT 67.395 107.140 67.685 107.185 ;
        RECT 67.930 107.140 68.070 107.975 ;
        RECT 70.140 107.960 70.460 108.020 ;
        RECT 144.660 107.960 144.980 108.220 ;
        RECT 85.320 107.820 85.640 107.880 ;
        RECT 110.620 107.820 110.940 107.880 ;
        RECT 85.320 107.680 110.940 107.820 ;
        RECT 85.320 107.620 85.640 107.680 ;
        RECT 110.620 107.620 110.940 107.680 ;
        RECT 71.060 107.480 71.380 107.540 ;
        RECT 71.535 107.480 71.825 107.525 ;
        RECT 117.060 107.480 117.380 107.540 ;
        RECT 117.535 107.480 117.825 107.525 ;
        RECT 125.355 107.480 125.645 107.525 ;
        RECT 71.060 107.340 71.825 107.480 ;
        RECT 71.060 107.280 71.380 107.340 ;
        RECT 71.535 107.295 71.825 107.340 ;
        RECT 81.270 107.340 85.090 107.480 ;
        RECT 67.395 107.000 68.070 107.140 ;
        RECT 70.600 107.140 70.920 107.200 ;
        RECT 74.280 107.140 74.600 107.200 ;
        RECT 70.600 107.000 74.600 107.140 ;
        RECT 67.395 106.955 67.685 107.000 ;
        RECT 70.600 106.940 70.920 107.000 ;
        RECT 74.280 106.940 74.600 107.000 ;
        RECT 80.720 106.940 81.040 107.200 ;
        RECT 81.270 107.185 81.410 107.340 ;
        RECT 84.950 107.200 85.090 107.340 ;
        RECT 117.060 107.340 117.825 107.480 ;
        RECT 117.060 107.280 117.380 107.340 ;
        RECT 117.535 107.295 117.825 107.340 ;
        RECT 123.590 107.340 125.645 107.480 ;
        RECT 81.195 106.955 81.485 107.185 ;
        RECT 82.115 106.955 82.405 107.185 ;
        RECT 82.575 106.955 82.865 107.185 ;
        RECT 84.860 107.140 85.180 107.200 ;
        RECT 85.795 107.140 86.085 107.185 ;
        RECT 84.860 107.000 86.085 107.140 ;
        RECT 55.435 106.800 55.725 106.845 ;
        RECT 46.770 106.660 55.725 106.800 ;
        RECT 37.480 106.600 37.800 106.660 ;
        RECT 55.435 106.615 55.725 106.660 ;
        RECT 56.355 106.615 56.645 106.845 ;
        RECT 66.015 106.800 66.305 106.845 ;
        RECT 68.300 106.800 68.620 106.860 ;
        RECT 66.015 106.660 68.620 106.800 ;
        RECT 66.015 106.615 66.305 106.660 ;
        RECT 31.500 106.460 31.820 106.520 ;
        RECT 31.975 106.460 32.265 106.505 ;
        RECT 31.500 106.320 32.265 106.460 ;
        RECT 31.500 106.260 31.820 106.320 ;
        RECT 31.975 106.275 32.265 106.320 ;
        RECT 35.180 106.260 35.500 106.520 ;
        RECT 40.255 106.460 40.545 106.505 ;
        RECT 40.700 106.460 41.020 106.520 ;
        RECT 40.255 106.320 41.020 106.460 ;
        RECT 40.255 106.275 40.545 106.320 ;
        RECT 40.700 106.260 41.020 106.320 ;
        RECT 43.920 106.260 44.240 106.520 ;
        RECT 45.760 106.460 46.080 106.520 ;
        RECT 51.280 106.460 51.600 106.520 ;
        RECT 45.760 106.320 51.600 106.460 ;
        RECT 45.760 106.260 46.080 106.320 ;
        RECT 51.280 106.260 51.600 106.320 ;
        RECT 51.740 106.260 52.060 106.520 ;
        RECT 52.200 106.460 52.520 106.520 ;
        RECT 56.430 106.460 56.570 106.615 ;
        RECT 68.300 106.600 68.620 106.660 ;
        RECT 52.200 106.320 56.570 106.460 ;
        RECT 52.200 106.260 52.520 106.320 ;
        RECT 60.020 106.260 60.340 106.520 ;
        RECT 73.820 106.460 74.140 106.520 ;
        RECT 74.755 106.460 75.045 106.505 ;
        RECT 73.820 106.320 75.045 106.460 ;
        RECT 73.820 106.260 74.140 106.320 ;
        RECT 74.755 106.275 75.045 106.320 ;
        RECT 79.800 106.260 80.120 106.520 ;
        RECT 82.190 106.460 82.330 106.955 ;
        RECT 82.650 106.800 82.790 106.955 ;
        RECT 84.860 106.940 85.180 107.000 ;
        RECT 85.795 106.955 86.085 107.000 ;
        RECT 86.715 107.140 87.005 107.185 ;
        RECT 88.080 107.140 88.400 107.200 ;
        RECT 86.715 107.000 88.400 107.140 ;
        RECT 86.715 106.955 87.005 107.000 ;
        RECT 88.080 106.940 88.400 107.000 ;
        RECT 94.520 106.940 94.840 107.200 ;
        RECT 96.835 107.140 97.125 107.185 ;
        RECT 97.755 107.140 98.045 107.185 ;
        RECT 98.200 107.140 98.520 107.200 ;
        RECT 96.835 107.000 97.510 107.140 ;
        RECT 96.835 106.955 97.125 107.000 ;
        RECT 87.160 106.800 87.480 106.860 ;
        RECT 82.650 106.660 87.480 106.800 ;
        RECT 87.160 106.600 87.480 106.660 ;
        RECT 97.370 106.520 97.510 107.000 ;
        RECT 97.755 107.000 98.520 107.140 ;
        RECT 97.755 106.955 98.045 107.000 ;
        RECT 98.200 106.940 98.520 107.000 ;
        RECT 100.040 106.940 100.360 107.200 ;
        RECT 112.000 107.140 112.320 107.200 ;
        RECT 113.395 107.140 113.685 107.185 ;
        RECT 112.000 107.000 113.685 107.140 ;
        RECT 112.000 106.940 112.320 107.000 ;
        RECT 113.395 106.955 113.685 107.000 ;
        RECT 114.315 106.955 114.605 107.185 ;
        RECT 114.775 107.140 115.065 107.185 ;
        RECT 115.220 107.140 115.540 107.200 ;
        RECT 114.775 107.000 115.540 107.140 ;
        RECT 114.775 106.955 115.065 107.000 ;
        RECT 112.920 106.800 113.240 106.860 ;
        RECT 114.390 106.800 114.530 106.955 ;
        RECT 115.220 106.940 115.540 107.000 ;
        RECT 115.695 107.140 115.985 107.185 ;
        RECT 116.140 107.140 116.460 107.200 ;
        RECT 115.695 107.000 116.460 107.140 ;
        RECT 115.695 106.955 115.985 107.000 ;
        RECT 115.770 106.800 115.910 106.955 ;
        RECT 116.140 106.940 116.460 107.000 ;
        RECT 118.440 106.940 118.760 107.200 ;
        RECT 123.590 107.185 123.730 107.340 ;
        RECT 125.355 107.295 125.645 107.340 ;
        RECT 126.260 107.480 126.580 107.540 ;
        RECT 128.115 107.480 128.405 107.525 ;
        RECT 126.260 107.340 128.405 107.480 ;
        RECT 126.260 107.280 126.580 107.340 ;
        RECT 128.115 107.295 128.405 107.340 ;
        RECT 131.320 107.280 131.640 107.540 ;
        RECT 142.360 107.480 142.680 107.540 ;
        RECT 142.360 107.340 145.350 107.480 ;
        RECT 142.360 107.280 142.680 107.340 ;
        RECT 123.055 106.955 123.345 107.185 ;
        RECT 123.515 106.955 123.805 107.185 ;
        RECT 123.975 107.140 124.265 107.185 ;
        RECT 124.420 107.140 124.740 107.200 ;
        RECT 123.975 107.000 124.740 107.140 ;
        RECT 123.975 106.955 124.265 107.000 ;
        RECT 112.920 106.660 115.910 106.800 ;
        RECT 112.920 106.600 113.240 106.660 ;
        RECT 121.660 106.600 121.980 106.860 ;
        RECT 123.130 106.800 123.270 106.955 ;
        RECT 124.420 106.940 124.740 107.000 ;
        RECT 124.895 107.140 125.185 107.185 ;
        RECT 127.640 107.140 127.960 107.200 ;
        RECT 124.895 107.000 127.960 107.140 ;
        RECT 124.895 106.955 125.185 107.000 ;
        RECT 127.640 106.940 127.960 107.000 ;
        RECT 129.035 107.140 129.325 107.185 ;
        RECT 129.480 107.140 129.800 107.200 ;
        RECT 129.035 107.000 129.800 107.140 ;
        RECT 129.035 106.955 129.325 107.000 ;
        RECT 129.480 106.940 129.800 107.000 ;
        RECT 130.415 107.140 130.705 107.185 ;
        RECT 130.860 107.140 131.180 107.200 ;
        RECT 130.415 107.000 131.180 107.140 ;
        RECT 130.415 106.955 130.705 107.000 ;
        RECT 130.860 106.940 131.180 107.000 ;
        RECT 143.280 107.140 143.600 107.200 ;
        RECT 145.210 107.185 145.350 107.340 ;
        RECT 144.215 107.140 144.505 107.185 ;
        RECT 143.280 107.000 144.505 107.140 ;
        RECT 143.280 106.940 143.600 107.000 ;
        RECT 144.215 106.955 144.505 107.000 ;
        RECT 145.135 106.955 145.425 107.185 ;
        RECT 123.130 106.660 125.110 106.800 ;
        RECT 124.970 106.520 125.110 106.660 ;
        RECT 84.400 106.460 84.720 106.520 ;
        RECT 85.320 106.460 85.640 106.520 ;
        RECT 82.190 106.320 85.640 106.460 ;
        RECT 84.400 106.260 84.720 106.320 ;
        RECT 85.320 106.260 85.640 106.320 ;
        RECT 86.240 106.260 86.560 106.520 ;
        RECT 93.600 106.260 93.920 106.520 ;
        RECT 95.900 106.260 96.220 106.520 ;
        RECT 97.280 106.260 97.600 106.520 ;
        RECT 100.975 106.460 101.265 106.505 ;
        RECT 103.720 106.460 104.040 106.520 ;
        RECT 100.975 106.320 104.040 106.460 ;
        RECT 100.975 106.275 101.265 106.320 ;
        RECT 103.720 106.260 104.040 106.320 ;
        RECT 113.840 106.260 114.160 106.520 ;
        RECT 114.300 106.460 114.620 106.520 ;
        RECT 115.235 106.460 115.525 106.505 ;
        RECT 114.300 106.320 115.525 106.460 ;
        RECT 114.300 106.260 114.620 106.320 ;
        RECT 115.235 106.275 115.525 106.320 ;
        RECT 119.360 106.260 119.680 106.520 ;
        RECT 124.880 106.260 125.200 106.520 ;
        RECT 125.340 106.460 125.660 106.520 ;
        RECT 129.495 106.460 129.785 106.505 ;
        RECT 125.340 106.320 129.785 106.460 ;
        RECT 125.340 106.260 125.660 106.320 ;
        RECT 129.495 106.275 129.785 106.320 ;
        RECT 22.690 105.640 157.810 106.120 ;
        RECT 29.200 105.240 29.520 105.500 ;
        RECT 33.340 105.440 33.660 105.500 ;
        RECT 38.400 105.440 38.720 105.500 ;
        RECT 33.340 105.300 38.720 105.440 ;
        RECT 33.340 105.240 33.660 105.300 ;
        RECT 38.400 105.240 38.720 105.300 ;
        RECT 44.380 105.240 44.700 105.500 ;
        RECT 51.295 105.440 51.585 105.485 ;
        RECT 53.120 105.440 53.440 105.500 ;
        RECT 51.295 105.300 53.440 105.440 ;
        RECT 51.295 105.255 51.585 105.300 ;
        RECT 53.120 105.240 53.440 105.300 ;
        RECT 57.720 105.240 58.040 105.500 ;
        RECT 60.020 105.240 60.340 105.500 ;
        RECT 64.620 105.240 64.940 105.500 ;
        RECT 66.935 105.440 67.225 105.485 ;
        RECT 70.600 105.440 70.920 105.500 ;
        RECT 66.935 105.300 70.920 105.440 ;
        RECT 66.935 105.255 67.225 105.300 ;
        RECT 70.600 105.240 70.920 105.300 ;
        RECT 73.820 105.240 74.140 105.500 ;
        RECT 87.160 105.240 87.480 105.500 ;
        RECT 89.015 105.440 89.305 105.485 ;
        RECT 92.680 105.440 93.000 105.500 ;
        RECT 89.015 105.300 93.000 105.440 ;
        RECT 89.015 105.255 89.305 105.300 ;
        RECT 92.680 105.240 93.000 105.300 ;
        RECT 99.580 105.240 99.900 105.500 ;
        RECT 100.040 105.440 100.360 105.500 ;
        RECT 100.515 105.440 100.805 105.485 ;
        RECT 109.255 105.440 109.545 105.485 ;
        RECT 100.040 105.300 100.805 105.440 ;
        RECT 100.040 105.240 100.360 105.300 ;
        RECT 100.515 105.255 100.805 105.300 ;
        RECT 101.970 105.300 109.545 105.440 ;
        RECT 35.640 105.100 35.960 105.160 ;
        RECT 26.990 104.960 35.960 105.100 ;
        RECT 26.990 104.805 27.130 104.960 ;
        RECT 35.640 104.900 35.960 104.960 ;
        RECT 37.940 104.900 38.260 105.160 ;
        RECT 48.980 104.900 49.300 105.160 ;
        RECT 57.810 105.100 57.950 105.240 ;
        RECT 55.970 104.960 57.950 105.100 ;
        RECT 25.995 104.575 26.285 104.805 ;
        RECT 26.915 104.575 27.205 104.805 ;
        RECT 27.375 104.575 27.665 104.805 ;
        RECT 27.835 104.760 28.125 104.805 ;
        RECT 29.200 104.760 29.520 104.820 ;
        RECT 31.960 104.805 32.280 104.820 ;
        RECT 27.835 104.620 29.520 104.760 ;
        RECT 27.835 104.575 28.125 104.620 ;
        RECT 26.070 103.740 26.210 104.575 ;
        RECT 26.440 104.420 26.760 104.480 ;
        RECT 27.450 104.420 27.590 104.575 ;
        RECT 29.200 104.560 29.520 104.620 ;
        RECT 31.930 104.575 32.280 104.805 ;
        RECT 31.960 104.560 32.280 104.575 ;
        RECT 50.360 104.560 50.680 104.820 ;
        RECT 52.200 104.560 52.520 104.820 ;
        RECT 54.500 104.760 54.820 104.820 ;
        RECT 55.970 104.805 56.110 104.960 ;
        RECT 54.975 104.760 55.265 104.805 ;
        RECT 54.500 104.620 55.265 104.760 ;
        RECT 54.500 104.560 54.820 104.620 ;
        RECT 54.975 104.575 55.265 104.620 ;
        RECT 55.895 104.575 56.185 104.805 ;
        RECT 57.230 104.760 57.520 104.805 ;
        RECT 60.110 104.760 60.250 105.240 ;
        RECT 64.710 105.100 64.850 105.240 ;
        RECT 65.555 105.100 65.845 105.145 ;
        RECT 64.710 104.960 65.845 105.100 ;
        RECT 65.555 104.915 65.845 104.960 ;
        RECT 72.610 105.100 72.900 105.145 ;
        RECT 73.910 105.100 74.050 105.240 ;
        RECT 72.610 104.960 74.050 105.100 ;
        RECT 74.280 105.100 74.600 105.160 ;
        RECT 93.600 105.145 93.920 105.160 ;
        RECT 74.280 104.960 76.350 105.100 ;
        RECT 72.610 104.915 72.900 104.960 ;
        RECT 74.280 104.900 74.600 104.960 ;
        RECT 57.230 104.620 60.250 104.760 ;
        RECT 64.635 104.760 64.925 104.805 ;
        RECT 67.380 104.760 67.700 104.820 ;
        RECT 64.635 104.620 67.700 104.760 ;
        RECT 57.230 104.575 57.520 104.620 ;
        RECT 64.635 104.575 64.925 104.620 ;
        RECT 26.440 104.280 27.590 104.420 ;
        RECT 26.440 104.220 26.760 104.280 ;
        RECT 30.580 104.220 30.900 104.480 ;
        RECT 31.475 104.420 31.765 104.465 ;
        RECT 32.665 104.420 32.955 104.465 ;
        RECT 35.185 104.420 35.475 104.465 ;
        RECT 31.475 104.280 35.475 104.420 ;
        RECT 31.475 104.235 31.765 104.280 ;
        RECT 32.665 104.235 32.955 104.280 ;
        RECT 35.185 104.235 35.475 104.280 ;
        RECT 49.900 104.420 50.220 104.480 ;
        RECT 52.290 104.420 52.430 104.560 ;
        RECT 49.900 104.280 52.430 104.420 ;
        RECT 56.775 104.420 57.065 104.465 ;
        RECT 57.965 104.420 58.255 104.465 ;
        RECT 60.485 104.420 60.775 104.465 ;
        RECT 56.775 104.280 60.775 104.420 ;
        RECT 49.900 104.220 50.220 104.280 ;
        RECT 56.775 104.235 57.065 104.280 ;
        RECT 57.965 104.235 58.255 104.280 ;
        RECT 60.485 104.235 60.775 104.280 ;
        RECT 31.080 104.080 31.370 104.125 ;
        RECT 33.180 104.080 33.470 104.125 ;
        RECT 34.750 104.080 35.040 104.125 ;
        RECT 31.080 103.940 35.040 104.080 ;
        RECT 31.080 103.895 31.370 103.940 ;
        RECT 33.180 103.895 33.470 103.940 ;
        RECT 34.750 103.895 35.040 103.940 ;
        RECT 56.380 104.080 56.670 104.125 ;
        RECT 58.480 104.080 58.770 104.125 ;
        RECT 60.050 104.080 60.340 104.125 ;
        RECT 56.380 103.940 60.340 104.080 ;
        RECT 56.380 103.895 56.670 103.940 ;
        RECT 58.480 103.895 58.770 103.940 ;
        RECT 60.050 103.895 60.340 103.940 ;
        RECT 62.795 104.080 63.085 104.125 ;
        RECT 64.710 104.080 64.850 104.575 ;
        RECT 67.380 104.560 67.700 104.620 ;
        RECT 73.835 104.760 74.125 104.805 ;
        RECT 74.740 104.760 75.060 104.820 ;
        RECT 73.835 104.620 75.060 104.760 ;
        RECT 73.835 104.575 74.125 104.620 ;
        RECT 74.740 104.560 75.060 104.620 ;
        RECT 75.200 104.560 75.520 104.820 ;
        RECT 76.210 104.805 76.350 104.960 ;
        RECT 84.950 104.960 87.850 105.100 ;
        RECT 84.950 104.820 85.090 104.960 ;
        RECT 76.135 104.575 76.425 104.805 ;
        RECT 80.275 104.760 80.565 104.805 ;
        RECT 84.415 104.760 84.705 104.805 ;
        RECT 80.275 104.620 84.705 104.760 ;
        RECT 80.275 104.575 80.565 104.620 ;
        RECT 84.415 104.575 84.705 104.620 ;
        RECT 69.245 104.420 69.535 104.465 ;
        RECT 71.765 104.420 72.055 104.465 ;
        RECT 72.955 104.420 73.245 104.465 ;
        RECT 69.245 104.280 73.245 104.420 ;
        RECT 84.490 104.420 84.630 104.575 ;
        RECT 84.860 104.560 85.180 104.820 ;
        RECT 85.320 104.760 85.640 104.820 ;
        RECT 85.795 104.760 86.085 104.805 ;
        RECT 85.320 104.620 86.085 104.760 ;
        RECT 85.320 104.560 85.640 104.620 ;
        RECT 85.795 104.575 86.085 104.620 ;
        RECT 86.240 104.560 86.560 104.820 ;
        RECT 86.700 104.560 87.020 104.820 ;
        RECT 87.710 104.805 87.850 104.960 ;
        RECT 90.010 104.960 92.450 105.100 ;
        RECT 90.010 104.805 90.150 104.960 ;
        RECT 87.635 104.575 87.925 104.805 ;
        RECT 89.935 104.575 90.225 104.805 ;
        RECT 90.395 104.760 90.685 104.805 ;
        RECT 90.840 104.760 91.160 104.820 ;
        RECT 90.395 104.620 91.160 104.760 ;
        RECT 90.395 104.575 90.685 104.620 ;
        RECT 90.010 104.420 90.150 104.575 ;
        RECT 90.840 104.560 91.160 104.620 ;
        RECT 91.300 104.560 91.620 104.820 ;
        RECT 91.775 104.575 92.065 104.805 ;
        RECT 92.310 104.760 92.450 104.960 ;
        RECT 93.515 104.915 93.920 105.145 ;
        RECT 99.670 105.100 99.810 105.240 ;
        RECT 101.970 105.100 102.110 105.300 ;
        RECT 109.255 105.255 109.545 105.300 ;
        RECT 113.840 105.240 114.160 105.500 ;
        RECT 116.615 105.255 116.905 105.485 ;
        RECT 118.455 105.440 118.745 105.485 ;
        RECT 119.360 105.440 119.680 105.500 ;
        RECT 118.455 105.300 119.680 105.440 ;
        RECT 118.455 105.255 118.745 105.300 ;
        RECT 99.670 104.960 102.110 105.100 ;
        RECT 102.355 105.100 102.645 105.145 ;
        RECT 102.800 105.100 103.120 105.160 ;
        RECT 113.930 105.100 114.070 105.240 ;
        RECT 102.355 104.960 103.120 105.100 ;
        RECT 102.355 104.915 102.645 104.960 ;
        RECT 93.600 104.900 93.920 104.915 ;
        RECT 102.800 104.900 103.120 104.960 ;
        RECT 104.270 104.960 112.690 105.100 ;
        RECT 113.930 104.960 114.530 105.100 ;
        RECT 104.270 104.760 104.410 104.960 ;
        RECT 92.310 104.620 104.410 104.760 ;
        RECT 84.490 104.280 90.150 104.420 ;
        RECT 69.245 104.235 69.535 104.280 ;
        RECT 71.765 104.235 72.055 104.280 ;
        RECT 72.955 104.235 73.245 104.280 ;
        RECT 62.795 103.940 64.850 104.080 ;
        RECT 69.680 104.080 69.970 104.125 ;
        RECT 71.250 104.080 71.540 104.125 ;
        RECT 73.350 104.080 73.640 104.125 ;
        RECT 69.680 103.940 73.640 104.080 ;
        RECT 62.795 103.895 63.085 103.940 ;
        RECT 69.680 103.895 69.970 103.940 ;
        RECT 71.250 103.895 71.540 103.940 ;
        RECT 73.350 103.895 73.640 103.940 ;
        RECT 30.120 103.740 30.440 103.800 ;
        RECT 32.420 103.740 32.740 103.800 ;
        RECT 26.070 103.600 32.740 103.740 ;
        RECT 30.120 103.540 30.440 103.600 ;
        RECT 32.420 103.540 32.740 103.600 ;
        RECT 35.180 103.740 35.500 103.800 ;
        RECT 37.495 103.740 37.785 103.785 ;
        RECT 48.995 103.740 49.285 103.785 ;
        RECT 35.180 103.600 49.285 103.740 ;
        RECT 35.180 103.540 35.500 103.600 ;
        RECT 37.495 103.555 37.785 103.600 ;
        RECT 48.995 103.555 49.285 103.600 ;
        RECT 52.200 103.540 52.520 103.800 ;
        RECT 63.240 103.740 63.560 103.800 ;
        RECT 63.715 103.740 64.005 103.785 ;
        RECT 63.240 103.600 64.005 103.740 ;
        RECT 63.240 103.540 63.560 103.600 ;
        RECT 63.715 103.555 64.005 103.600 ;
        RECT 77.075 103.740 77.365 103.785 ;
        RECT 77.995 103.740 78.285 103.785 ;
        RECT 77.075 103.600 78.285 103.740 ;
        RECT 77.075 103.555 77.365 103.600 ;
        RECT 77.995 103.555 78.285 103.600 ;
        RECT 83.495 103.740 83.785 103.785 ;
        RECT 85.320 103.740 85.640 103.800 ;
        RECT 83.495 103.600 85.640 103.740 ;
        RECT 91.850 103.740 91.990 104.575 ;
        RECT 108.780 104.560 109.100 104.820 ;
        RECT 112.550 104.805 112.690 104.960 ;
        RECT 112.475 104.575 112.765 104.805 ;
        RECT 112.920 104.560 113.240 104.820 ;
        RECT 114.390 104.805 114.530 104.960 ;
        RECT 113.855 104.760 114.145 104.805 ;
        RECT 113.470 104.620 114.145 104.760 ;
        RECT 113.470 104.480 113.610 104.620 ;
        RECT 113.855 104.575 114.145 104.620 ;
        RECT 114.315 104.575 114.605 104.805 ;
        RECT 116.155 104.760 116.445 104.805 ;
        RECT 116.690 104.760 116.830 105.255 ;
        RECT 119.360 105.240 119.680 105.300 ;
        RECT 126.260 105.240 126.580 105.500 ;
        RECT 125.800 105.100 126.120 105.160 ;
        RECT 116.155 104.620 116.830 104.760 ;
        RECT 123.130 104.960 126.120 105.100 ;
        RECT 116.155 104.575 116.445 104.620 ;
        RECT 92.220 104.220 92.540 104.480 ;
        RECT 93.115 104.420 93.405 104.465 ;
        RECT 94.305 104.420 94.595 104.465 ;
        RECT 96.825 104.420 97.115 104.465 ;
        RECT 93.115 104.280 97.115 104.420 ;
        RECT 93.115 104.235 93.405 104.280 ;
        RECT 94.305 104.235 94.595 104.280 ;
        RECT 96.825 104.235 97.115 104.280 ;
        RECT 97.740 104.220 98.060 104.480 ;
        RECT 98.660 104.220 98.980 104.480 ;
        RECT 99.580 104.420 99.900 104.480 ;
        RECT 102.815 104.420 103.105 104.465 ;
        RECT 99.580 104.280 103.105 104.420 ;
        RECT 99.580 104.220 99.900 104.280 ;
        RECT 102.815 104.235 103.105 104.280 ;
        RECT 103.275 104.235 103.565 104.465 ;
        RECT 109.715 104.235 110.005 104.465 ;
        RECT 113.380 104.420 113.700 104.480 ;
        RECT 115.680 104.420 116.000 104.480 ;
        RECT 113.380 104.280 116.000 104.420 ;
        RECT 92.720 104.080 93.010 104.125 ;
        RECT 94.820 104.080 95.110 104.125 ;
        RECT 96.390 104.080 96.680 104.125 ;
        RECT 97.830 104.080 97.970 104.220 ;
        RECT 92.720 103.940 96.680 104.080 ;
        RECT 92.720 103.895 93.010 103.940 ;
        RECT 94.820 103.895 95.110 103.940 ;
        RECT 96.390 103.895 96.680 103.940 ;
        RECT 96.910 103.940 97.970 104.080 ;
        RECT 98.750 104.080 98.890 104.220 ;
        RECT 103.350 104.080 103.490 104.235 ;
        RECT 98.750 103.940 103.490 104.080 ;
        RECT 108.320 104.080 108.640 104.140 ;
        RECT 109.790 104.080 109.930 104.235 ;
        RECT 113.380 104.220 113.700 104.280 ;
        RECT 115.680 104.220 116.000 104.280 ;
        RECT 116.600 104.420 116.920 104.480 ;
        RECT 118.915 104.420 119.205 104.465 ;
        RECT 116.600 104.280 119.205 104.420 ;
        RECT 116.600 104.220 116.920 104.280 ;
        RECT 118.915 104.235 119.205 104.280 ;
        RECT 119.820 104.220 120.140 104.480 ;
        RECT 108.320 103.940 109.930 104.080 ;
        RECT 111.555 104.080 111.845 104.125 ;
        RECT 123.130 104.080 123.270 104.960 ;
        RECT 125.800 104.900 126.120 104.960 ;
        RECT 123.515 104.575 123.805 104.805 ;
        RECT 126.350 104.760 126.490 105.240 ;
        RECT 124.050 104.620 126.490 104.760 ;
        RECT 130.400 104.760 130.720 104.820 ;
        RECT 131.840 104.760 132.130 104.805 ;
        RECT 130.400 104.620 132.130 104.760 ;
        RECT 111.555 103.940 123.270 104.080 ;
        RECT 123.590 104.080 123.730 104.575 ;
        RECT 124.050 104.465 124.190 104.620 ;
        RECT 130.400 104.560 130.720 104.620 ;
        RECT 131.840 104.575 132.130 104.620 ;
        RECT 133.175 104.760 133.465 104.805 ;
        RECT 138.220 104.760 138.540 104.820 ;
        RECT 133.175 104.620 138.540 104.760 ;
        RECT 133.175 104.575 133.465 104.620 ;
        RECT 138.220 104.560 138.540 104.620 ;
        RECT 143.280 104.560 143.600 104.820 ;
        RECT 123.975 104.235 124.265 104.465 ;
        RECT 125.340 104.220 125.660 104.480 ;
        RECT 128.585 104.420 128.875 104.465 ;
        RECT 131.105 104.420 131.395 104.465 ;
        RECT 132.295 104.420 132.585 104.465 ;
        RECT 128.585 104.280 132.585 104.420 ;
        RECT 128.585 104.235 128.875 104.280 ;
        RECT 131.105 104.235 131.395 104.280 ;
        RECT 132.295 104.235 132.585 104.280 ;
        RECT 129.020 104.080 129.310 104.125 ;
        RECT 130.590 104.080 130.880 104.125 ;
        RECT 132.690 104.080 132.980 104.125 ;
        RECT 123.590 103.940 125.110 104.080 ;
        RECT 92.220 103.740 92.540 103.800 ;
        RECT 96.910 103.740 97.050 103.940 ;
        RECT 108.320 103.880 108.640 103.940 ;
        RECT 111.555 103.895 111.845 103.940 ;
        RECT 124.970 103.800 125.110 103.940 ;
        RECT 129.020 103.940 132.980 104.080 ;
        RECT 129.020 103.895 129.310 103.940 ;
        RECT 130.590 103.895 130.880 103.940 ;
        RECT 132.690 103.895 132.980 103.940 ;
        RECT 91.850 103.600 97.050 103.740 ;
        RECT 97.280 103.740 97.600 103.800 ;
        RECT 99.135 103.740 99.425 103.785 ;
        RECT 97.280 103.600 99.425 103.740 ;
        RECT 83.495 103.555 83.785 103.600 ;
        RECT 85.320 103.540 85.640 103.600 ;
        RECT 92.220 103.540 92.540 103.600 ;
        RECT 97.280 103.540 97.600 103.600 ;
        RECT 99.135 103.555 99.425 103.600 ;
        RECT 106.955 103.740 107.245 103.785 ;
        RECT 107.860 103.740 108.180 103.800 ;
        RECT 106.955 103.600 108.180 103.740 ;
        RECT 106.955 103.555 107.245 103.600 ;
        RECT 107.860 103.540 108.180 103.600 ;
        RECT 115.220 103.540 115.540 103.800 ;
        RECT 124.880 103.540 125.200 103.800 ;
        RECT 144.200 103.540 144.520 103.800 ;
        RECT 22.690 102.920 157.010 103.400 ;
        RECT 31.040 102.720 31.360 102.780 ;
        RECT 33.340 102.720 33.660 102.780 ;
        RECT 31.040 102.580 33.660 102.720 ;
        RECT 31.040 102.520 31.360 102.580 ;
        RECT 33.340 102.520 33.660 102.580 ;
        RECT 37.480 102.720 37.800 102.780 ;
        RECT 38.875 102.720 39.165 102.765 ;
        RECT 44.380 102.720 44.700 102.780 ;
        RECT 48.980 102.720 49.300 102.780 ;
        RECT 49.455 102.720 49.745 102.765 ;
        RECT 37.480 102.580 39.165 102.720 ;
        RECT 37.480 102.520 37.800 102.580 ;
        RECT 38.875 102.535 39.165 102.580 ;
        RECT 42.630 102.580 47.370 102.720 ;
        RECT 26.900 102.380 27.190 102.425 ;
        RECT 28.470 102.380 28.760 102.425 ;
        RECT 30.570 102.380 30.860 102.425 ;
        RECT 26.900 102.240 30.860 102.380 ;
        RECT 26.900 102.195 27.190 102.240 ;
        RECT 28.470 102.195 28.760 102.240 ;
        RECT 30.570 102.195 30.860 102.240 ;
        RECT 34.720 102.380 35.040 102.440 ;
        RECT 35.195 102.380 35.485 102.425 ;
        RECT 34.720 102.240 35.485 102.380 ;
        RECT 34.720 102.180 35.040 102.240 ;
        RECT 35.195 102.195 35.485 102.240 ;
        RECT 38.415 102.380 38.705 102.425 ;
        RECT 41.620 102.380 41.940 102.440 ;
        RECT 38.415 102.240 41.940 102.380 ;
        RECT 38.415 102.195 38.705 102.240 ;
        RECT 41.620 102.180 41.940 102.240 ;
        RECT 42.630 102.085 42.770 102.580 ;
        RECT 44.380 102.520 44.700 102.580 ;
        RECT 43.040 102.380 43.330 102.425 ;
        RECT 45.140 102.380 45.430 102.425 ;
        RECT 46.710 102.380 47.000 102.425 ;
        RECT 43.040 102.240 47.000 102.380 ;
        RECT 47.230 102.380 47.370 102.580 ;
        RECT 48.980 102.580 49.745 102.720 ;
        RECT 48.980 102.520 49.300 102.580 ;
        RECT 49.455 102.535 49.745 102.580 ;
        RECT 54.500 102.720 54.820 102.780 ;
        RECT 56.815 102.720 57.105 102.765 ;
        RECT 54.500 102.580 57.105 102.720 ;
        RECT 54.500 102.520 54.820 102.580 ;
        RECT 56.815 102.535 57.105 102.580 ;
        RECT 57.260 102.720 57.580 102.780 ;
        RECT 60.035 102.720 60.325 102.765 ;
        RECT 57.260 102.580 60.325 102.720 ;
        RECT 57.260 102.520 57.580 102.580 ;
        RECT 60.035 102.535 60.325 102.580 ;
        RECT 60.940 102.520 61.260 102.780 ;
        RECT 70.615 102.720 70.905 102.765 ;
        RECT 74.740 102.720 75.060 102.780 ;
        RECT 70.615 102.580 75.060 102.720 ;
        RECT 70.615 102.535 70.905 102.580 ;
        RECT 50.400 102.380 50.690 102.425 ;
        RECT 52.500 102.380 52.790 102.425 ;
        RECT 54.070 102.380 54.360 102.425 ;
        RECT 47.230 102.240 50.130 102.380 ;
        RECT 43.040 102.195 43.330 102.240 ;
        RECT 45.140 102.195 45.430 102.240 ;
        RECT 46.710 102.195 47.000 102.240 ;
        RECT 49.990 102.085 50.130 102.240 ;
        RECT 50.400 102.240 54.360 102.380 ;
        RECT 50.400 102.195 50.690 102.240 ;
        RECT 52.500 102.195 52.790 102.240 ;
        RECT 54.070 102.195 54.360 102.240 ;
        RECT 64.250 102.240 65.770 102.380 ;
        RECT 64.250 102.100 64.390 102.240 ;
        RECT 26.465 102.040 26.755 102.085 ;
        RECT 28.985 102.040 29.275 102.085 ;
        RECT 30.175 102.040 30.465 102.085 ;
        RECT 42.555 102.040 42.845 102.085 ;
        RECT 26.465 101.900 30.465 102.040 ;
        RECT 26.465 101.855 26.755 101.900 ;
        RECT 28.985 101.855 29.275 101.900 ;
        RECT 30.175 101.855 30.465 101.900 ;
        RECT 39.410 101.900 42.845 102.040 ;
        RECT 39.410 101.760 39.550 101.900 ;
        RECT 42.555 101.855 42.845 101.900 ;
        RECT 43.435 102.040 43.725 102.085 ;
        RECT 44.625 102.040 44.915 102.085 ;
        RECT 47.145 102.040 47.435 102.085 ;
        RECT 43.435 101.900 47.435 102.040 ;
        RECT 43.435 101.855 43.725 101.900 ;
        RECT 44.625 101.855 44.915 101.900 ;
        RECT 47.145 101.855 47.435 101.900 ;
        RECT 49.915 101.855 50.205 102.085 ;
        RECT 50.795 102.040 51.085 102.085 ;
        RECT 51.985 102.040 52.275 102.085 ;
        RECT 54.505 102.040 54.795 102.085 ;
        RECT 50.795 101.900 54.795 102.040 ;
        RECT 50.795 101.855 51.085 101.900 ;
        RECT 51.985 101.855 52.275 101.900 ;
        RECT 54.505 101.855 54.795 101.900 ;
        RECT 64.160 101.840 64.480 102.100 ;
        RECT 65.080 101.840 65.400 102.100 ;
        RECT 65.630 102.040 65.770 102.240 ;
        RECT 66.460 102.180 66.780 102.440 ;
        RECT 70.690 102.380 70.830 102.535 ;
        RECT 74.740 102.520 75.060 102.580 ;
        RECT 75.200 102.520 75.520 102.780 ;
        RECT 76.155 102.720 76.445 102.765 ;
        RECT 77.075 102.720 77.365 102.765 ;
        RECT 76.155 102.580 77.365 102.720 ;
        RECT 76.155 102.535 76.445 102.580 ;
        RECT 77.075 102.535 77.365 102.580 ;
        RECT 94.520 102.520 94.840 102.780 ;
        RECT 108.780 102.720 109.100 102.780 ;
        RECT 109.255 102.720 109.545 102.765 ;
        RECT 116.600 102.720 116.920 102.780 ;
        RECT 101.510 102.580 106.250 102.720 ;
        RECT 68.390 102.240 70.830 102.380 ;
        RECT 68.390 102.040 68.530 102.240 ;
        RECT 65.630 101.900 68.530 102.040 ;
        RECT 30.580 101.700 30.900 101.760 ;
        RECT 31.055 101.700 31.345 101.745 ;
        RECT 30.580 101.560 31.345 101.700 ;
        RECT 30.580 101.500 30.900 101.560 ;
        RECT 31.055 101.515 31.345 101.560 ;
        RECT 31.975 101.700 32.265 101.745 ;
        RECT 32.420 101.700 32.740 101.760 ;
        RECT 31.975 101.560 32.740 101.700 ;
        RECT 31.975 101.515 32.265 101.560 ;
        RECT 29.660 101.405 29.980 101.420 ;
        RECT 29.660 101.175 30.010 101.405 ;
        RECT 31.130 101.360 31.270 101.515 ;
        RECT 32.420 101.500 32.740 101.560 ;
        RECT 32.880 101.500 33.200 101.760 ;
        RECT 33.340 101.500 33.660 101.760 ;
        RECT 33.815 101.700 34.105 101.745 ;
        RECT 36.100 101.700 36.420 101.760 ;
        RECT 33.815 101.560 36.420 101.700 ;
        RECT 33.815 101.515 34.105 101.560 ;
        RECT 36.100 101.500 36.420 101.560 ;
        RECT 36.575 101.700 36.865 101.745 ;
        RECT 37.020 101.700 37.340 101.760 ;
        RECT 36.575 101.560 37.340 101.700 ;
        RECT 36.575 101.515 36.865 101.560 ;
        RECT 37.020 101.500 37.340 101.560 ;
        RECT 39.320 101.500 39.640 101.760 ;
        RECT 43.920 101.745 44.240 101.760 ;
        RECT 42.095 101.515 42.385 101.745 ;
        RECT 43.890 101.700 44.240 101.745 ;
        RECT 43.725 101.560 44.240 101.700 ;
        RECT 43.890 101.515 44.240 101.560 ;
        RECT 58.195 101.700 58.485 101.745 ;
        RECT 59.560 101.700 59.880 101.760 ;
        RECT 58.195 101.560 59.880 101.700 ;
        RECT 58.195 101.515 58.485 101.560 ;
        RECT 31.130 101.220 34.950 101.360 ;
        RECT 29.660 101.160 29.980 101.175 ;
        RECT 34.810 101.080 34.950 101.220 ;
        RECT 37.495 101.175 37.785 101.405 ;
        RECT 42.170 101.360 42.310 101.515 ;
        RECT 43.920 101.500 44.240 101.515 ;
        RECT 59.560 101.500 59.880 101.560 ;
        RECT 63.715 101.515 64.005 101.745 ;
        RECT 64.635 101.700 64.925 101.745 ;
        RECT 67.380 101.700 67.700 101.760 ;
        RECT 64.635 101.560 67.700 101.700 ;
        RECT 64.635 101.515 64.925 101.560 ;
        RECT 49.900 101.360 50.220 101.420 ;
        RECT 42.170 101.220 50.220 101.360 ;
        RECT 24.140 100.820 24.460 101.080 ;
        RECT 31.500 101.020 31.820 101.080 ;
        RECT 32.420 101.020 32.740 101.080 ;
        RECT 31.500 100.880 32.740 101.020 ;
        RECT 31.500 100.820 31.820 100.880 ;
        RECT 32.420 100.820 32.740 100.880 ;
        RECT 34.720 100.820 35.040 101.080 ;
        RECT 37.570 101.020 37.710 101.175 ;
        RECT 49.900 101.160 50.220 101.220 ;
        RECT 51.250 101.360 51.540 101.405 ;
        RECT 51.740 101.360 52.060 101.420 ;
        RECT 51.250 101.220 52.060 101.360 ;
        RECT 51.250 101.175 51.540 101.220 ;
        RECT 51.740 101.160 52.060 101.220 ;
        RECT 60.035 101.360 60.325 101.405 ;
        RECT 63.240 101.360 63.560 101.420 ;
        RECT 60.035 101.220 63.560 101.360 ;
        RECT 63.790 101.360 63.930 101.515 ;
        RECT 67.380 101.500 67.700 101.560 ;
        RECT 67.855 101.700 68.145 101.745 ;
        RECT 68.390 101.700 68.530 101.900 ;
        RECT 69.235 102.040 69.525 102.085 ;
        RECT 70.600 102.040 70.920 102.100 ;
        RECT 69.235 101.900 70.920 102.040 ;
        RECT 75.290 102.040 75.430 102.520 ;
        RECT 83.940 102.380 84.260 102.440 ;
        RECT 85.795 102.380 86.085 102.425 ;
        RECT 101.510 102.380 101.650 102.580 ;
        RECT 83.940 102.240 86.085 102.380 ;
        RECT 83.940 102.180 84.260 102.240 ;
        RECT 85.795 102.195 86.085 102.240 ;
        RECT 96.910 102.240 101.650 102.380 ;
        RECT 101.880 102.380 102.170 102.425 ;
        RECT 103.450 102.380 103.740 102.425 ;
        RECT 105.550 102.380 105.840 102.425 ;
        RECT 101.880 102.240 105.840 102.380 ;
        RECT 106.110 102.380 106.250 102.580 ;
        RECT 108.780 102.580 109.545 102.720 ;
        RECT 108.780 102.520 109.100 102.580 ;
        RECT 109.255 102.535 109.545 102.580 ;
        RECT 114.850 102.580 116.920 102.720 ;
        RECT 108.320 102.380 108.640 102.440 ;
        RECT 114.850 102.380 114.990 102.580 ;
        RECT 116.600 102.520 116.920 102.580 ;
        RECT 118.440 102.720 118.760 102.780 ;
        RECT 121.200 102.720 121.520 102.780 ;
        RECT 121.675 102.720 121.965 102.765 ;
        RECT 118.440 102.580 121.965 102.720 ;
        RECT 118.440 102.520 118.760 102.580 ;
        RECT 121.200 102.520 121.520 102.580 ;
        RECT 121.675 102.535 121.965 102.580 ;
        RECT 124.420 102.520 124.740 102.780 ;
        RECT 125.340 102.520 125.660 102.780 ;
        RECT 106.110 102.240 114.990 102.380 ;
        RECT 115.260 102.380 115.550 102.425 ;
        RECT 117.360 102.380 117.650 102.425 ;
        RECT 118.930 102.380 119.220 102.425 ;
        RECT 115.260 102.240 119.220 102.380 ;
        RECT 75.675 102.040 75.965 102.085 ;
        RECT 75.290 101.900 75.965 102.040 ;
        RECT 69.235 101.855 69.525 101.900 ;
        RECT 70.600 101.840 70.920 101.900 ;
        RECT 75.675 101.855 75.965 101.900 ;
        RECT 79.355 102.040 79.645 102.085 ;
        RECT 80.720 102.040 81.040 102.100 ;
        RECT 96.910 102.085 97.050 102.240 ;
        RECT 101.880 102.195 102.170 102.240 ;
        RECT 103.450 102.195 103.740 102.240 ;
        RECT 105.550 102.195 105.840 102.240 ;
        RECT 108.320 102.180 108.640 102.240 ;
        RECT 115.260 102.195 115.550 102.240 ;
        RECT 117.360 102.195 117.650 102.240 ;
        RECT 118.930 102.195 119.220 102.240 ;
        RECT 123.055 102.380 123.345 102.425 ;
        RECT 124.510 102.380 124.650 102.520 ;
        RECT 123.055 102.240 124.650 102.380 ;
        RECT 123.055 102.195 123.345 102.240 ;
        RECT 79.355 101.900 90.610 102.040 ;
        RECT 79.355 101.855 79.645 101.900 ;
        RECT 80.720 101.840 81.040 101.900 ;
        RECT 67.855 101.560 68.530 101.700 ;
        RECT 67.855 101.515 68.145 101.560 ;
        RECT 75.215 101.515 75.505 101.745 ;
        RECT 81.640 101.700 81.960 101.760 ;
        RECT 82.115 101.700 82.405 101.745 ;
        RECT 81.640 101.560 82.405 101.700 ;
        RECT 68.315 101.360 68.605 101.405 ;
        RECT 71.520 101.360 71.840 101.420 ;
        RECT 75.290 101.360 75.430 101.515 ;
        RECT 81.640 101.500 81.960 101.560 ;
        RECT 82.115 101.515 82.405 101.560 ;
        RECT 63.790 101.220 75.430 101.360 ;
        RECT 82.190 101.360 82.330 101.515 ;
        RECT 83.020 101.500 83.340 101.760 ;
        RECT 85.780 101.500 86.100 101.760 ;
        RECT 90.470 101.745 90.610 101.900 ;
        RECT 96.835 101.855 97.125 102.085 ;
        RECT 97.755 102.040 98.045 102.085 ;
        RECT 98.660 102.040 98.980 102.100 ;
        RECT 97.755 101.900 98.980 102.040 ;
        RECT 97.755 101.855 98.045 101.900 ;
        RECT 98.660 101.840 98.980 101.900 ;
        RECT 101.445 102.040 101.735 102.085 ;
        RECT 103.965 102.040 104.255 102.085 ;
        RECT 105.155 102.040 105.445 102.085 ;
        RECT 114.775 102.040 115.065 102.085 ;
        RECT 101.445 101.900 105.445 102.040 ;
        RECT 101.445 101.855 101.735 101.900 ;
        RECT 103.965 101.855 104.255 101.900 ;
        RECT 105.155 101.855 105.445 101.900 ;
        RECT 106.110 101.900 115.065 102.040 ;
        RECT 86.715 101.515 87.005 101.745 ;
        RECT 90.395 101.515 90.685 101.745 ;
        RECT 84.860 101.360 85.180 101.420 ;
        RECT 86.790 101.360 86.930 101.515 ;
        RECT 82.190 101.220 86.930 101.360 ;
        RECT 90.470 101.360 90.610 101.515 ;
        RECT 90.840 101.500 91.160 101.760 ;
        RECT 91.760 101.500 92.080 101.760 ;
        RECT 92.220 101.500 92.540 101.760 ;
        RECT 95.900 101.700 96.220 101.760 ;
        RECT 96.375 101.700 96.665 101.745 ;
        RECT 95.900 101.560 96.665 101.700 ;
        RECT 95.900 101.500 96.220 101.560 ;
        RECT 96.375 101.515 96.665 101.560 ;
        RECT 103.260 101.700 103.580 101.760 ;
        RECT 105.560 101.700 105.880 101.760 ;
        RECT 106.110 101.745 106.250 101.900 ;
        RECT 114.775 101.855 115.065 101.900 ;
        RECT 115.655 102.040 115.945 102.085 ;
        RECT 116.845 102.040 117.135 102.085 ;
        RECT 119.365 102.040 119.655 102.085 ;
        RECT 115.655 101.900 119.655 102.040 ;
        RECT 125.430 102.040 125.570 102.520 ;
        RECT 128.575 102.380 128.865 102.425 ;
        RECT 130.400 102.380 130.720 102.440 ;
        RECT 137.300 102.380 137.620 102.440 ;
        RECT 142.835 102.380 143.125 102.425 ;
        RECT 128.575 102.240 130.720 102.380 ;
        RECT 128.575 102.195 128.865 102.240 ;
        RECT 130.400 102.180 130.720 102.240 ;
        RECT 134.170 102.240 143.125 102.380 ;
        RECT 134.170 102.085 134.310 102.240 ;
        RECT 137.300 102.180 137.620 102.240 ;
        RECT 142.835 102.195 143.125 102.240 ;
        RECT 145.580 102.380 145.870 102.425 ;
        RECT 147.150 102.380 147.440 102.425 ;
        RECT 149.250 102.380 149.540 102.425 ;
        RECT 145.580 102.240 149.540 102.380 ;
        RECT 145.580 102.195 145.870 102.240 ;
        RECT 147.150 102.195 147.440 102.240 ;
        RECT 149.250 102.195 149.540 102.240 ;
        RECT 126.275 102.040 126.565 102.085 ;
        RECT 125.430 101.900 126.565 102.040 ;
        RECT 115.655 101.855 115.945 101.900 ;
        RECT 116.845 101.855 117.135 101.900 ;
        RECT 119.365 101.855 119.655 101.900 ;
        RECT 126.275 101.855 126.565 101.900 ;
        RECT 134.095 101.855 134.385 102.085 ;
        RECT 140.535 102.040 140.825 102.085 ;
        RECT 141.440 102.040 141.760 102.100 ;
        RECT 140.535 101.900 141.760 102.040 ;
        RECT 140.535 101.855 140.825 101.900 ;
        RECT 141.440 101.840 141.760 101.900 ;
        RECT 145.145 102.040 145.435 102.085 ;
        RECT 147.665 102.040 147.955 102.085 ;
        RECT 148.855 102.040 149.145 102.085 ;
        RECT 145.145 101.900 149.145 102.040 ;
        RECT 145.145 101.855 145.435 101.900 ;
        RECT 147.665 101.855 147.955 101.900 ;
        RECT 148.855 101.855 149.145 101.900 ;
        RECT 149.720 101.840 150.040 102.100 ;
        RECT 106.035 101.700 106.325 101.745 ;
        RECT 103.260 101.560 106.325 101.700 ;
        RECT 103.260 101.500 103.580 101.560 ;
        RECT 105.560 101.500 105.880 101.560 ;
        RECT 106.035 101.515 106.325 101.560 ;
        RECT 107.860 101.500 108.180 101.760 ;
        RECT 110.160 101.500 110.480 101.760 ;
        RECT 110.620 101.500 110.940 101.760 ;
        RECT 115.220 101.700 115.540 101.760 ;
        RECT 116.055 101.700 116.345 101.745 ;
        RECT 115.220 101.560 116.345 101.700 ;
        RECT 115.220 101.500 115.540 101.560 ;
        RECT 116.055 101.515 116.345 101.560 ;
        RECT 123.975 101.515 124.265 101.745 ;
        RECT 125.355 101.700 125.645 101.745 ;
        RECT 125.355 101.560 126.490 101.700 ;
        RECT 125.355 101.515 125.645 101.560 ;
        RECT 103.720 101.360 104.040 101.420 ;
        RECT 104.700 101.360 104.990 101.405 ;
        RECT 124.050 101.360 124.190 101.515 ;
        RECT 126.350 101.420 126.490 101.560 ;
        RECT 126.735 101.515 127.025 101.745 ;
        RECT 127.655 101.700 127.945 101.745 ;
        RECT 130.860 101.700 131.180 101.760 ;
        RECT 127.655 101.560 131.180 101.700 ;
        RECT 127.655 101.515 127.945 101.560 ;
        RECT 90.470 101.220 99.810 101.360 ;
        RECT 60.035 101.175 60.325 101.220 ;
        RECT 63.240 101.160 63.560 101.220 ;
        RECT 68.315 101.175 68.605 101.220 ;
        RECT 71.520 101.160 71.840 101.220 ;
        RECT 84.860 101.160 85.180 101.220 ;
        RECT 52.200 101.020 52.520 101.080 ;
        RECT 37.570 100.880 52.520 101.020 ;
        RECT 52.200 100.820 52.520 100.880 ;
        RECT 66.000 100.820 66.320 101.080 ;
        RECT 67.380 100.820 67.700 101.080 ;
        RECT 69.680 100.820 70.000 101.080 ;
        RECT 70.600 101.065 70.920 101.080 ;
        RECT 70.535 100.835 70.920 101.065 ;
        RECT 70.600 100.820 70.920 100.835 ;
        RECT 82.560 100.820 82.880 101.080 ;
        RECT 89.475 101.020 89.765 101.065 ;
        RECT 93.140 101.020 93.460 101.080 ;
        RECT 89.475 100.880 93.460 101.020 ;
        RECT 89.475 100.835 89.765 100.880 ;
        RECT 93.140 100.820 93.460 100.880 ;
        RECT 96.820 101.020 97.140 101.080 ;
        RECT 99.120 101.020 99.440 101.080 ;
        RECT 96.820 100.880 99.440 101.020 ;
        RECT 99.670 101.020 99.810 101.220 ;
        RECT 103.720 101.220 104.990 101.360 ;
        RECT 103.720 101.160 104.040 101.220 ;
        RECT 104.700 101.175 104.990 101.220 ;
        RECT 105.190 101.220 114.990 101.360 ;
        RECT 124.050 101.220 125.570 101.360 ;
        RECT 105.190 101.020 105.330 101.220 ;
        RECT 114.850 101.080 114.990 101.220 ;
        RECT 99.670 100.880 105.330 101.020 ;
        RECT 96.820 100.820 97.140 100.880 ;
        RECT 99.120 100.820 99.440 100.880 ;
        RECT 106.940 100.820 107.260 101.080 ;
        RECT 114.760 100.820 115.080 101.080 ;
        RECT 124.880 100.820 125.200 101.080 ;
        RECT 125.430 101.020 125.570 101.220 ;
        RECT 126.260 101.160 126.580 101.420 ;
        RECT 126.810 101.360 126.950 101.515 ;
        RECT 130.860 101.500 131.180 101.560 ;
        RECT 133.635 101.700 133.925 101.745 ;
        RECT 135.000 101.700 135.320 101.760 ;
        RECT 133.635 101.560 135.320 101.700 ;
        RECT 133.635 101.515 133.925 101.560 ;
        RECT 135.000 101.500 135.320 101.560 ;
        RECT 140.075 101.515 140.365 101.745 ;
        RECT 144.200 101.700 144.520 101.760 ;
        RECT 148.400 101.700 148.690 101.745 ;
        RECT 144.200 101.560 148.690 101.700 ;
        RECT 129.480 101.360 129.800 101.420 ;
        RECT 126.810 101.220 129.800 101.360 ;
        RECT 126.810 101.020 126.950 101.220 ;
        RECT 129.480 101.160 129.800 101.220 ;
        RECT 125.430 100.880 126.950 101.020 ;
        RECT 135.460 101.020 135.780 101.080 ;
        RECT 140.150 101.020 140.290 101.515 ;
        RECT 144.200 101.500 144.520 101.560 ;
        RECT 148.400 101.515 148.690 101.560 ;
        RECT 135.460 100.880 140.290 101.020 ;
        RECT 135.460 100.820 135.780 100.880 ;
        RECT 141.900 100.820 142.220 101.080 ;
        RECT 22.690 100.200 157.810 100.680 ;
        RECT 25.995 100.000 26.285 100.045 ;
        RECT 26.440 100.000 26.760 100.060 ;
        RECT 33.815 100.000 34.105 100.045 ;
        RECT 25.995 99.860 26.760 100.000 ;
        RECT 25.995 99.815 26.285 99.860 ;
        RECT 26.440 99.800 26.760 99.860 ;
        RECT 29.290 99.860 34.105 100.000 ;
        RECT 29.290 99.380 29.430 99.860 ;
        RECT 33.815 99.815 34.105 99.860 ;
        RECT 35.640 99.800 35.960 100.060 ;
        RECT 36.560 100.000 36.880 100.060 ;
        RECT 37.035 100.000 37.325 100.045 ;
        RECT 36.560 99.860 37.325 100.000 ;
        RECT 36.560 99.800 36.880 99.860 ;
        RECT 37.035 99.815 37.325 99.860 ;
        RECT 46.235 100.000 46.525 100.045 ;
        RECT 49.900 100.000 50.220 100.060 ;
        RECT 46.235 99.860 50.220 100.000 ;
        RECT 46.235 99.815 46.525 99.860 ;
        RECT 49.900 99.800 50.220 99.860 ;
        RECT 59.115 100.000 59.405 100.045 ;
        RECT 59.115 99.860 62.550 100.000 ;
        RECT 59.115 99.815 59.405 99.860 ;
        RECT 32.420 99.660 32.740 99.720 ;
        RECT 37.955 99.660 38.245 99.705 ;
        RECT 62.410 99.660 62.550 99.860 ;
        RECT 64.160 99.800 64.480 100.060 ;
        RECT 65.080 99.800 65.400 100.060 ;
        RECT 66.000 100.000 66.320 100.060 ;
        RECT 66.935 100.000 67.225 100.045 ;
        RECT 66.000 99.860 67.225 100.000 ;
        RECT 66.000 99.800 66.320 99.860 ;
        RECT 66.935 99.815 67.225 99.860 ;
        RECT 83.940 99.800 84.260 100.060 ;
        RECT 84.400 99.800 84.720 100.060 ;
        RECT 90.380 100.000 90.700 100.060 ;
        RECT 86.790 99.860 97.970 100.000 ;
        RECT 64.250 99.660 64.390 99.800 ;
        RECT 65.170 99.660 65.310 99.800 ;
        RECT 31.590 99.520 38.245 99.660 ;
        RECT 24.140 99.320 24.460 99.380 ;
        RECT 28.280 99.320 28.600 99.380 ;
        RECT 28.755 99.320 29.045 99.365 ;
        RECT 24.140 99.180 29.045 99.320 ;
        RECT 24.140 99.120 24.460 99.180 ;
        RECT 28.280 99.120 28.600 99.180 ;
        RECT 28.755 99.135 29.045 99.180 ;
        RECT 28.830 98.300 28.970 99.135 ;
        RECT 29.200 99.120 29.520 99.380 ;
        RECT 29.675 99.320 29.965 99.365 ;
        RECT 30.120 99.320 30.440 99.380 ;
        RECT 29.675 99.180 30.440 99.320 ;
        RECT 29.675 99.135 29.965 99.180 ;
        RECT 30.120 99.120 30.440 99.180 ;
        RECT 30.580 99.120 30.900 99.380 ;
        RECT 31.040 99.120 31.360 99.380 ;
        RECT 31.590 99.365 31.730 99.520 ;
        RECT 32.420 99.460 32.740 99.520 ;
        RECT 37.955 99.475 38.245 99.520 ;
        RECT 60.570 99.520 62.090 99.660 ;
        RECT 31.515 99.135 31.805 99.365 ;
        RECT 33.355 99.135 33.645 99.365 ;
        RECT 34.735 99.135 35.025 99.365 ;
        RECT 35.180 99.320 35.500 99.380 ;
        RECT 37.020 99.320 37.340 99.380 ;
        RECT 40.700 99.365 41.020 99.380 ;
        RECT 38.875 99.320 39.165 99.365 ;
        RECT 40.670 99.320 41.020 99.365 ;
        RECT 35.180 99.180 39.165 99.320 ;
        RECT 40.505 99.180 41.020 99.320 ;
        RECT 31.960 98.980 32.280 99.040 ;
        RECT 32.895 98.980 33.185 99.025 ;
        RECT 31.960 98.840 33.185 98.980 ;
        RECT 33.430 98.980 33.570 99.135 ;
        RECT 34.260 98.980 34.580 99.040 ;
        RECT 34.810 98.980 34.950 99.135 ;
        RECT 35.180 99.120 35.500 99.180 ;
        RECT 37.020 99.120 37.340 99.180 ;
        RECT 38.875 99.135 39.165 99.180 ;
        RECT 40.670 99.135 41.020 99.180 ;
        RECT 40.700 99.120 41.020 99.135 ;
        RECT 57.260 99.120 57.580 99.380 ;
        RECT 59.560 99.365 59.880 99.380 ;
        RECT 59.560 99.320 59.890 99.365 ;
        RECT 60.570 99.320 60.710 99.520 ;
        RECT 59.560 99.180 60.710 99.320 ;
        RECT 59.560 99.135 59.890 99.180 ;
        RECT 60.955 99.135 61.245 99.365 ;
        RECT 59.560 99.120 59.880 99.135 ;
        RECT 33.430 98.840 33.800 98.980 ;
        RECT 31.960 98.780 32.280 98.840 ;
        RECT 32.895 98.795 33.185 98.840 ;
        RECT 33.660 98.300 33.800 98.840 ;
        RECT 34.260 98.840 34.950 98.980 ;
        RECT 34.260 98.780 34.580 98.840 ;
        RECT 39.320 98.780 39.640 99.040 ;
        RECT 40.215 98.980 40.505 99.025 ;
        RECT 41.405 98.980 41.695 99.025 ;
        RECT 43.925 98.980 44.215 99.025 ;
        RECT 40.215 98.840 44.215 98.980 ;
        RECT 40.215 98.795 40.505 98.840 ;
        RECT 41.405 98.795 41.695 98.840 ;
        RECT 43.925 98.795 44.215 98.840 ;
        RECT 34.720 98.640 35.040 98.700 ;
        RECT 39.410 98.640 39.550 98.780 ;
        RECT 34.720 98.500 39.550 98.640 ;
        RECT 39.820 98.640 40.110 98.685 ;
        RECT 41.920 98.640 42.210 98.685 ;
        RECT 43.490 98.640 43.780 98.685 ;
        RECT 39.820 98.500 43.780 98.640 ;
        RECT 57.350 98.640 57.490 99.120 ;
        RECT 58.195 98.980 58.485 99.025 ;
        RECT 61.030 98.980 61.170 99.135 ;
        RECT 58.195 98.840 61.170 98.980 ;
        RECT 58.195 98.795 58.485 98.840 ;
        RECT 61.950 98.685 62.090 99.520 ;
        RECT 62.410 99.520 64.390 99.660 ;
        RECT 64.710 99.520 65.310 99.660 ;
        RECT 67.380 99.660 67.700 99.720 ;
        RECT 67.380 99.520 77.270 99.660 ;
        RECT 62.410 99.365 62.550 99.520 ;
        RECT 62.335 99.135 62.625 99.365 ;
        RECT 63.715 99.320 64.005 99.365 ;
        RECT 64.710 99.320 64.850 99.520 ;
        RECT 67.380 99.460 67.700 99.520 ;
        RECT 63.715 99.180 64.850 99.320 ;
        RECT 65.095 99.320 65.385 99.365 ;
        RECT 66.920 99.320 67.240 99.380 ;
        RECT 69.680 99.320 70.000 99.380 ;
        RECT 65.095 99.180 70.000 99.320 ;
        RECT 63.715 99.135 64.005 99.180 ;
        RECT 65.095 99.135 65.385 99.180 ;
        RECT 66.920 99.120 67.240 99.180 ;
        RECT 69.680 99.120 70.000 99.180 ;
        RECT 70.600 99.120 70.920 99.380 ;
        RECT 75.200 99.120 75.520 99.380 ;
        RECT 77.130 99.365 77.270 99.520 ;
        RECT 77.055 99.135 77.345 99.365 ;
        RECT 84.030 99.320 84.170 99.800 ;
        RECT 84.490 99.660 84.630 99.800 ;
        RECT 84.490 99.520 85.550 99.660 ;
        RECT 85.410 99.365 85.550 99.520 ;
        RECT 86.790 99.380 86.930 99.860 ;
        RECT 90.380 99.800 90.700 99.860 ;
        RECT 90.930 99.520 94.750 99.660 ;
        RECT 90.930 99.380 91.070 99.520 ;
        RECT 84.875 99.320 85.165 99.365 ;
        RECT 84.030 99.180 85.165 99.320 ;
        RECT 84.875 99.135 85.165 99.180 ;
        RECT 85.335 99.135 85.625 99.365 ;
        RECT 85.780 99.320 86.100 99.380 ;
        RECT 86.255 99.320 86.545 99.365 ;
        RECT 85.780 99.180 86.545 99.320 ;
        RECT 85.780 99.120 86.100 99.180 ;
        RECT 86.255 99.135 86.545 99.180 ;
        RECT 86.700 99.120 87.020 99.380 ;
        RECT 88.540 99.320 88.860 99.380 ;
        RECT 89.935 99.320 90.225 99.365 ;
        RECT 88.540 99.180 90.225 99.320 ;
        RECT 88.540 99.120 88.860 99.180 ;
        RECT 89.935 99.135 90.225 99.180 ;
        RECT 90.395 99.320 90.685 99.365 ;
        RECT 90.840 99.320 91.160 99.380 ;
        RECT 90.395 99.180 91.160 99.320 ;
        RECT 90.395 99.135 90.685 99.180 ;
        RECT 90.840 99.120 91.160 99.180 ;
        RECT 91.315 99.135 91.605 99.365 ;
        RECT 91.775 99.320 92.065 99.365 ;
        RECT 92.220 99.320 92.540 99.380 ;
        RECT 93.230 99.365 93.370 99.520 ;
        RECT 94.610 99.380 94.750 99.520 ;
        RECT 91.775 99.180 92.540 99.320 ;
        RECT 91.775 99.135 92.065 99.180 ;
        RECT 64.635 98.980 64.925 99.025 ;
        RECT 67.380 98.980 67.700 99.040 ;
        RECT 64.635 98.840 67.700 98.980 ;
        RECT 64.635 98.795 64.925 98.840 ;
        RECT 67.380 98.780 67.700 98.840 ;
        RECT 61.875 98.640 62.165 98.685 ;
        RECT 62.795 98.640 63.085 98.685 ;
        RECT 70.690 98.640 70.830 99.120 ;
        RECT 75.675 98.980 75.965 99.025 ;
        RECT 80.735 98.980 81.025 99.025 ;
        RECT 75.675 98.840 81.025 98.980 ;
        RECT 75.675 98.795 75.965 98.840 ;
        RECT 80.735 98.795 81.025 98.840 ;
        RECT 82.100 98.980 82.420 99.040 ;
        RECT 84.415 98.980 84.705 99.025 ;
        RECT 88.630 98.980 88.770 99.120 ;
        RECT 82.100 98.840 88.770 98.980 ;
        RECT 91.390 98.980 91.530 99.135 ;
        RECT 92.220 99.120 92.540 99.180 ;
        RECT 93.155 99.135 93.445 99.365 ;
        RECT 94.075 99.135 94.365 99.365 ;
        RECT 94.150 98.980 94.290 99.135 ;
        RECT 94.520 99.120 94.840 99.380 ;
        RECT 95.455 99.320 95.745 99.365 ;
        RECT 97.280 99.320 97.600 99.380 ;
        RECT 95.455 99.180 97.600 99.320 ;
        RECT 95.455 99.135 95.745 99.180 ;
        RECT 97.280 99.120 97.600 99.180 ;
        RECT 96.820 98.980 97.140 99.040 ;
        RECT 91.390 98.840 93.830 98.980 ;
        RECT 94.150 98.840 97.140 98.980 ;
        RECT 82.100 98.780 82.420 98.840 ;
        RECT 84.415 98.795 84.705 98.840 ;
        RECT 57.350 98.500 61.630 98.640 ;
        RECT 34.720 98.440 35.040 98.500 ;
        RECT 39.820 98.455 40.110 98.500 ;
        RECT 41.920 98.455 42.210 98.500 ;
        RECT 43.490 98.455 43.780 98.500 ;
        RECT 28.830 98.160 33.800 98.300 ;
        RECT 60.020 98.100 60.340 98.360 ;
        RECT 61.490 98.300 61.630 98.500 ;
        RECT 61.875 98.500 70.830 98.640 ;
        RECT 61.875 98.455 62.165 98.500 ;
        RECT 62.795 98.455 63.085 98.500 ;
        RECT 93.690 98.360 93.830 98.840 ;
        RECT 96.820 98.780 97.140 98.840 ;
        RECT 65.540 98.300 65.860 98.360 ;
        RECT 66.935 98.300 67.225 98.345 ;
        RECT 61.490 98.160 67.225 98.300 ;
        RECT 65.540 98.100 65.860 98.160 ;
        RECT 66.935 98.115 67.225 98.160 ;
        RECT 67.855 98.300 68.145 98.345 ;
        RECT 68.300 98.300 68.620 98.360 ;
        RECT 67.855 98.160 68.620 98.300 ;
        RECT 67.855 98.115 68.145 98.160 ;
        RECT 68.300 98.100 68.620 98.160 ;
        RECT 87.620 98.100 87.940 98.360 ;
        RECT 89.015 98.300 89.305 98.345 ;
        RECT 91.300 98.300 91.620 98.360 ;
        RECT 89.015 98.160 91.620 98.300 ;
        RECT 89.015 98.115 89.305 98.160 ;
        RECT 91.300 98.100 91.620 98.160 ;
        RECT 93.600 98.300 93.920 98.360 ;
        RECT 94.075 98.300 94.365 98.345 ;
        RECT 93.600 98.160 94.365 98.300 ;
        RECT 93.600 98.100 93.920 98.160 ;
        RECT 94.075 98.115 94.365 98.160 ;
        RECT 95.440 98.100 95.760 98.360 ;
        RECT 97.830 98.300 97.970 99.860 ;
        RECT 99.120 99.800 99.440 100.060 ;
        RECT 102.800 99.800 103.120 100.060 ;
        RECT 110.160 100.000 110.480 100.060 ;
        RECT 112.475 100.000 112.765 100.045 ;
        RECT 110.160 99.860 112.765 100.000 ;
        RECT 110.160 99.800 110.480 99.860 ;
        RECT 112.475 99.815 112.765 99.860 ;
        RECT 114.300 99.800 114.620 100.060 ;
        RECT 116.600 100.000 116.920 100.060 ;
        RECT 115.310 99.860 118.670 100.000 ;
        RECT 99.210 99.660 99.350 99.800 ;
        RECT 106.940 99.705 107.260 99.720 ;
        RECT 99.210 99.520 102.110 99.660 ;
        RECT 98.200 99.320 98.520 99.380 ;
        RECT 101.970 99.365 102.110 99.520 ;
        RECT 106.855 99.475 107.260 99.705 ;
        RECT 114.390 99.660 114.530 99.800 ;
        RECT 106.940 99.460 107.260 99.475 ;
        RECT 113.010 99.520 114.530 99.660 ;
        RECT 100.975 99.320 101.265 99.365 ;
        RECT 98.200 99.180 101.265 99.320 ;
        RECT 98.200 99.120 98.520 99.180 ;
        RECT 100.975 99.135 101.265 99.180 ;
        RECT 101.895 99.135 102.185 99.365 ;
        RECT 110.620 99.320 110.940 99.380 ;
        RECT 113.010 99.365 113.150 99.520 ;
        RECT 104.730 99.180 110.940 99.320 ;
        RECT 101.050 98.980 101.190 99.135 ;
        RECT 104.730 98.980 104.870 99.180 ;
        RECT 110.620 99.120 110.940 99.180 ;
        RECT 112.935 99.135 113.225 99.365 ;
        RECT 113.395 99.320 113.685 99.365 ;
        RECT 113.840 99.320 114.160 99.380 ;
        RECT 113.395 99.180 114.160 99.320 ;
        RECT 113.395 99.135 113.685 99.180 ;
        RECT 113.840 99.120 114.160 99.180 ;
        RECT 114.315 99.135 114.605 99.365 ;
        RECT 101.050 98.840 104.870 98.980 ;
        RECT 105.100 98.980 105.420 99.040 ;
        RECT 105.575 98.980 105.865 99.025 ;
        RECT 105.100 98.840 105.865 98.980 ;
        RECT 105.100 98.780 105.420 98.840 ;
        RECT 105.575 98.795 105.865 98.840 ;
        RECT 106.455 98.980 106.745 99.025 ;
        RECT 107.645 98.980 107.935 99.025 ;
        RECT 110.165 98.980 110.455 99.025 ;
        RECT 114.390 98.980 114.530 99.135 ;
        RECT 114.760 99.120 115.080 99.380 ;
        RECT 115.310 98.980 115.450 99.860 ;
        RECT 116.600 99.800 116.920 99.860 ;
        RECT 115.695 99.660 115.985 99.705 ;
        RECT 117.520 99.660 117.840 99.720 ;
        RECT 115.695 99.520 117.840 99.660 ;
        RECT 115.695 99.475 115.985 99.520 ;
        RECT 117.520 99.460 117.840 99.520 ;
        RECT 118.530 99.660 118.670 99.860 ;
        RECT 135.460 99.800 135.780 100.060 ;
        RECT 137.300 99.800 137.620 100.060 ;
        RECT 141.900 99.800 142.220 100.060 ;
        RECT 143.280 100.000 143.600 100.060 ;
        RECT 143.755 100.000 144.045 100.045 ;
        RECT 143.280 99.860 144.045 100.000 ;
        RECT 143.280 99.800 143.600 99.860 ;
        RECT 143.755 99.815 144.045 99.860 ;
        RECT 135.550 99.660 135.690 99.800 ;
        RECT 118.530 99.520 120.510 99.660 ;
        RECT 118.530 99.365 118.670 99.520 ;
        RECT 120.370 99.365 120.510 99.520 ;
        RECT 134.170 99.520 135.690 99.660 ;
        RECT 106.455 98.840 110.455 98.980 ;
        RECT 106.455 98.795 106.745 98.840 ;
        RECT 107.645 98.795 107.935 98.840 ;
        RECT 110.165 98.795 110.455 98.840 ;
        RECT 113.010 98.840 115.450 98.980 ;
        RECT 115.770 99.180 116.600 99.320 ;
        RECT 113.010 98.700 113.150 98.840 ;
        RECT 106.060 98.640 106.350 98.685 ;
        RECT 108.160 98.640 108.450 98.685 ;
        RECT 109.730 98.640 110.020 98.685 ;
        RECT 106.060 98.500 110.020 98.640 ;
        RECT 106.060 98.455 106.350 98.500 ;
        RECT 108.160 98.455 108.450 98.500 ;
        RECT 109.730 98.455 110.020 98.500 ;
        RECT 112.920 98.440 113.240 98.700 ;
        RECT 115.770 98.300 115.910 99.180 ;
        RECT 116.460 98.980 116.600 99.180 ;
        RECT 117.995 99.135 118.285 99.365 ;
        RECT 118.455 99.135 118.745 99.365 ;
        RECT 119.375 99.135 119.665 99.365 ;
        RECT 119.835 99.135 120.125 99.365 ;
        RECT 120.295 99.135 120.585 99.365 ;
        RECT 118.070 98.980 118.210 99.135 ;
        RECT 116.460 98.840 118.210 98.980 ;
        RECT 116.140 98.640 116.460 98.700 ;
        RECT 119.450 98.640 119.590 99.135 ;
        RECT 119.910 98.980 120.050 99.135 ;
        RECT 121.200 99.120 121.520 99.380 ;
        RECT 133.160 99.120 133.480 99.380 ;
        RECT 134.170 99.365 134.310 99.520 ;
        RECT 134.095 99.135 134.385 99.365 ;
        RECT 134.555 99.135 134.845 99.365 ;
        RECT 135.460 99.320 135.780 99.380 ;
        RECT 137.390 99.365 137.530 99.800 ;
        RECT 136.855 99.320 137.145 99.365 ;
        RECT 135.460 99.180 137.145 99.320 ;
        RECT 120.755 98.980 121.045 99.025 ;
        RECT 119.910 98.840 121.045 98.980 ;
        RECT 120.755 98.795 121.045 98.840 ;
        RECT 123.040 98.980 123.360 99.040 ;
        RECT 131.320 98.980 131.640 99.040 ;
        RECT 123.040 98.840 131.640 98.980 ;
        RECT 123.040 98.780 123.360 98.840 ;
        RECT 131.320 98.780 131.640 98.840 ;
        RECT 116.140 98.500 119.590 98.640 ;
        RECT 133.635 98.640 133.925 98.685 ;
        RECT 134.080 98.640 134.400 98.700 ;
        RECT 133.635 98.500 134.400 98.640 ;
        RECT 116.140 98.440 116.460 98.500 ;
        RECT 133.635 98.455 133.925 98.500 ;
        RECT 134.080 98.440 134.400 98.500 ;
        RECT 134.630 98.360 134.770 99.135 ;
        RECT 135.460 99.120 135.780 99.180 ;
        RECT 136.855 99.135 137.145 99.180 ;
        RECT 137.315 99.135 137.605 99.365 ;
        RECT 137.760 99.120 138.080 99.380 ;
        RECT 138.695 99.135 138.985 99.365 ;
        RECT 141.990 99.320 142.130 99.800 ;
        RECT 142.835 99.320 143.125 99.365 ;
        RECT 141.990 99.180 143.125 99.320 ;
        RECT 142.835 99.135 143.125 99.180 ;
        RECT 137.300 98.640 137.620 98.700 ;
        RECT 138.770 98.640 138.910 99.135 ;
        RECT 141.900 98.780 142.220 99.040 ;
        RECT 137.300 98.500 138.910 98.640 ;
        RECT 137.300 98.440 137.620 98.500 ;
        RECT 97.830 98.160 115.910 98.300 ;
        RECT 117.075 98.300 117.365 98.345 ;
        RECT 125.340 98.300 125.660 98.360 ;
        RECT 117.075 98.160 125.660 98.300 ;
        RECT 117.075 98.115 117.365 98.160 ;
        RECT 125.340 98.100 125.660 98.160 ;
        RECT 129.940 98.300 130.260 98.360 ;
        RECT 132.255 98.300 132.545 98.345 ;
        RECT 129.940 98.160 132.545 98.300 ;
        RECT 129.940 98.100 130.260 98.160 ;
        RECT 132.255 98.115 132.545 98.160 ;
        RECT 134.540 98.100 134.860 98.360 ;
        RECT 135.000 98.300 135.320 98.360 ;
        RECT 135.475 98.300 135.765 98.345 ;
        RECT 135.000 98.160 135.765 98.300 ;
        RECT 135.000 98.100 135.320 98.160 ;
        RECT 135.475 98.115 135.765 98.160 ;
        RECT 22.690 97.480 157.010 97.960 ;
        RECT 26.915 97.280 27.205 97.325 ;
        RECT 23.770 97.140 31.730 97.280 ;
        RECT 23.770 96.260 23.910 97.140 ;
        RECT 26.915 97.095 27.205 97.140 ;
        RECT 25.075 96.940 25.365 96.985 ;
        RECT 25.075 96.800 30.810 96.940 ;
        RECT 25.075 96.755 25.365 96.800 ;
        RECT 24.155 96.600 24.445 96.645 ;
        RECT 27.820 96.600 28.140 96.660 ;
        RECT 24.155 96.460 28.140 96.600 ;
        RECT 24.155 96.415 24.445 96.460 ;
        RECT 27.820 96.400 28.140 96.460 ;
        RECT 28.280 96.400 28.600 96.660 ;
        RECT 29.660 96.600 29.980 96.660 ;
        RECT 30.135 96.600 30.425 96.645 ;
        RECT 29.660 96.460 30.425 96.600 ;
        RECT 29.660 96.400 29.980 96.460 ;
        RECT 30.135 96.415 30.425 96.460 ;
        RECT 25.995 96.260 26.285 96.305 ;
        RECT 23.770 96.120 26.285 96.260 ;
        RECT 25.995 96.075 26.285 96.120 ;
        RECT 26.455 96.075 26.745 96.305 ;
        RECT 28.755 96.260 29.045 96.305 ;
        RECT 29.200 96.260 29.520 96.320 ;
        RECT 28.755 96.120 29.520 96.260 ;
        RECT 30.670 96.260 30.810 96.800 ;
        RECT 31.590 96.600 31.730 97.140 ;
        RECT 32.880 97.080 33.200 97.340 ;
        RECT 60.495 97.280 60.785 97.325 ;
        RECT 64.160 97.280 64.480 97.340 ;
        RECT 60.495 97.140 64.480 97.280 ;
        RECT 60.495 97.095 60.785 97.140 ;
        RECT 64.160 97.080 64.480 97.140 ;
        RECT 71.520 97.280 71.840 97.340 ;
        RECT 72.915 97.280 73.205 97.325 ;
        RECT 71.520 97.140 73.205 97.280 ;
        RECT 71.520 97.080 71.840 97.140 ;
        RECT 72.915 97.095 73.205 97.140 ;
        RECT 75.695 97.280 75.985 97.325 ;
        RECT 76.615 97.280 76.905 97.325 ;
        RECT 75.695 97.140 76.905 97.280 ;
        RECT 75.695 97.095 75.985 97.140 ;
        RECT 76.615 97.095 76.905 97.140 ;
        RECT 110.160 97.280 110.480 97.340 ;
        RECT 128.575 97.280 128.865 97.325 ;
        RECT 129.020 97.280 129.340 97.340 ;
        RECT 130.415 97.280 130.705 97.325 ;
        RECT 110.160 97.140 111.770 97.280 ;
        RECT 110.160 97.080 110.480 97.140 ;
        RECT 31.960 96.940 32.280 97.000 ;
        RECT 34.260 96.940 34.580 97.000 ;
        RECT 31.960 96.800 34.580 96.940 ;
        RECT 31.960 96.740 32.280 96.800 ;
        RECT 34.260 96.740 34.580 96.800 ;
        RECT 36.600 96.940 36.890 96.985 ;
        RECT 38.700 96.940 38.990 96.985 ;
        RECT 40.270 96.940 40.560 96.985 ;
        RECT 36.600 96.800 40.560 96.940 ;
        RECT 36.600 96.755 36.890 96.800 ;
        RECT 38.700 96.755 38.990 96.800 ;
        RECT 40.270 96.755 40.560 96.800 ;
        RECT 46.720 96.940 47.010 96.985 ;
        RECT 48.820 96.940 49.110 96.985 ;
        RECT 50.390 96.940 50.680 96.985 ;
        RECT 46.720 96.800 50.680 96.940 ;
        RECT 46.720 96.755 47.010 96.800 ;
        RECT 48.820 96.755 49.110 96.800 ;
        RECT 50.390 96.755 50.680 96.800 ;
        RECT 54.080 96.940 54.370 96.985 ;
        RECT 56.180 96.940 56.470 96.985 ;
        RECT 57.750 96.940 58.040 96.985 ;
        RECT 54.080 96.800 58.040 96.940 ;
        RECT 54.080 96.755 54.370 96.800 ;
        RECT 56.180 96.755 56.470 96.800 ;
        RECT 57.750 96.755 58.040 96.800 ;
        RECT 66.500 96.940 66.790 96.985 ;
        RECT 68.600 96.940 68.890 96.985 ;
        RECT 70.170 96.940 70.460 96.985 ;
        RECT 66.500 96.800 70.460 96.940 ;
        RECT 66.500 96.755 66.790 96.800 ;
        RECT 68.600 96.755 68.890 96.800 ;
        RECT 70.170 96.755 70.460 96.800 ;
        RECT 84.400 96.740 84.720 97.000 ;
        RECT 90.395 96.940 90.685 96.985 ;
        RECT 91.760 96.940 92.080 97.000 ;
        RECT 90.395 96.800 92.080 96.940 ;
        RECT 90.395 96.755 90.685 96.800 ;
        RECT 91.760 96.740 92.080 96.800 ;
        RECT 101.895 96.940 102.185 96.985 ;
        RECT 104.180 96.940 104.500 97.000 ;
        RECT 101.895 96.800 104.500 96.940 ;
        RECT 101.895 96.755 102.185 96.800 ;
        RECT 104.180 96.740 104.500 96.800 ;
        RECT 107.875 96.940 108.165 96.985 ;
        RECT 110.620 96.940 110.940 97.000 ;
        RECT 107.875 96.800 110.940 96.940 ;
        RECT 107.875 96.755 108.165 96.800 ;
        RECT 110.620 96.740 110.940 96.800 ;
        RECT 32.435 96.600 32.725 96.645 ;
        RECT 31.590 96.460 32.725 96.600 ;
        RECT 32.435 96.415 32.725 96.460 ;
        RECT 36.995 96.600 37.285 96.645 ;
        RECT 38.185 96.600 38.475 96.645 ;
        RECT 40.705 96.600 40.995 96.645 ;
        RECT 36.995 96.460 40.995 96.600 ;
        RECT 36.995 96.415 37.285 96.460 ;
        RECT 38.185 96.415 38.475 96.460 ;
        RECT 40.705 96.415 40.995 96.460 ;
        RECT 47.115 96.600 47.405 96.645 ;
        RECT 48.305 96.600 48.595 96.645 ;
        RECT 50.825 96.600 51.115 96.645 ;
        RECT 47.115 96.460 51.115 96.600 ;
        RECT 47.115 96.415 47.405 96.460 ;
        RECT 48.305 96.415 48.595 96.460 ;
        RECT 50.825 96.415 51.115 96.460 ;
        RECT 54.475 96.600 54.765 96.645 ;
        RECT 55.665 96.600 55.955 96.645 ;
        RECT 58.185 96.600 58.475 96.645 ;
        RECT 54.475 96.460 58.475 96.600 ;
        RECT 54.475 96.415 54.765 96.460 ;
        RECT 55.665 96.415 55.955 96.460 ;
        RECT 58.185 96.415 58.475 96.460 ;
        RECT 66.895 96.600 67.185 96.645 ;
        RECT 68.085 96.600 68.375 96.645 ;
        RECT 70.605 96.600 70.895 96.645 ;
        RECT 66.895 96.460 70.895 96.600 ;
        RECT 66.895 96.415 67.185 96.460 ;
        RECT 68.085 96.415 68.375 96.460 ;
        RECT 70.605 96.415 70.895 96.460 ;
        RECT 75.200 96.400 75.520 96.660 ;
        RECT 82.115 96.600 82.405 96.645 ;
        RECT 82.560 96.600 82.880 96.660 ;
        RECT 82.115 96.460 82.880 96.600 ;
        RECT 82.115 96.415 82.405 96.460 ;
        RECT 82.560 96.400 82.880 96.460 ;
        RECT 83.020 96.600 83.340 96.660 ;
        RECT 84.490 96.600 84.630 96.740 ;
        RECT 93.630 96.645 93.890 96.690 ;
        RECT 83.020 96.460 84.630 96.600 ;
        RECT 90.850 96.600 91.140 96.645 ;
        RECT 93.610 96.600 93.900 96.645 ;
        RECT 90.850 96.460 93.900 96.600 ;
        RECT 83.020 96.400 83.340 96.460 ;
        RECT 90.850 96.415 91.140 96.460 ;
        RECT 93.610 96.415 93.900 96.460 ;
        RECT 93.630 96.370 93.890 96.415 ;
        RECT 31.055 96.260 31.345 96.305 ;
        RECT 30.670 96.120 31.345 96.260 ;
        RECT 28.755 96.075 29.045 96.120 ;
        RECT 26.530 95.580 26.670 96.075 ;
        RECT 29.200 96.060 29.520 96.120 ;
        RECT 31.055 96.075 31.345 96.120 ;
        RECT 31.960 96.060 32.280 96.320 ;
        RECT 34.260 96.260 34.580 96.320 ;
        RECT 36.115 96.260 36.405 96.305 ;
        RECT 46.235 96.260 46.525 96.305 ;
        RECT 34.260 96.120 46.525 96.260 ;
        RECT 34.260 96.060 34.580 96.120 ;
        RECT 36.115 96.075 36.405 96.120 ;
        RECT 46.235 96.075 46.525 96.120 ;
        RECT 50.360 96.260 50.680 96.320 ;
        RECT 53.595 96.260 53.885 96.305 ;
        RECT 66.000 96.260 66.320 96.320 ;
        RECT 50.360 96.120 66.320 96.260 ;
        RECT 50.360 96.060 50.680 96.120 ;
        RECT 53.595 96.075 53.885 96.120 ;
        RECT 66.000 96.060 66.320 96.120 ;
        RECT 74.740 96.060 75.060 96.320 ;
        RECT 81.640 96.260 81.960 96.320 ;
        RECT 84.415 96.260 84.705 96.305 ;
        RECT 85.780 96.260 86.100 96.320 ;
        RECT 81.640 96.120 86.100 96.260 ;
        RECT 81.640 96.060 81.960 96.120 ;
        RECT 84.415 96.075 84.705 96.120 ;
        RECT 85.780 96.060 86.100 96.120 ;
        RECT 86.255 96.075 86.545 96.305 ;
        RECT 33.800 95.720 34.120 95.980 ;
        RECT 34.735 95.920 35.025 95.965 ;
        RECT 35.180 95.920 35.500 95.980 ;
        RECT 34.735 95.780 35.500 95.920 ;
        RECT 34.735 95.735 35.025 95.780 ;
        RECT 35.180 95.720 35.500 95.780 ;
        RECT 35.640 95.920 35.960 95.980 ;
        RECT 37.340 95.920 37.630 95.965 ;
        RECT 35.640 95.780 37.630 95.920 ;
        RECT 35.640 95.720 35.960 95.780 ;
        RECT 37.340 95.735 37.630 95.780 ;
        RECT 47.570 95.920 47.860 95.965 ;
        RECT 51.740 95.920 52.060 95.980 ;
        RECT 47.570 95.780 52.060 95.920 ;
        RECT 47.570 95.735 47.860 95.780 ;
        RECT 51.740 95.720 52.060 95.780 ;
        RECT 54.930 95.920 55.220 95.965 ;
        RECT 60.020 95.920 60.340 95.980 ;
        RECT 67.380 95.965 67.700 95.980 ;
        RECT 54.930 95.780 60.340 95.920 ;
        RECT 54.930 95.735 55.220 95.780 ;
        RECT 60.020 95.720 60.340 95.780 ;
        RECT 67.350 95.735 67.700 95.965 ;
        RECT 67.380 95.720 67.700 95.735 ;
        RECT 83.940 95.720 84.260 95.980 ;
        RECT 86.330 95.920 86.470 96.075 ;
        RECT 92.220 96.060 92.540 96.320 ;
        RECT 94.520 96.060 94.840 96.320 ;
        RECT 97.295 96.075 97.585 96.305 ;
        RECT 88.540 95.920 88.860 95.980 ;
        RECT 97.370 95.920 97.510 96.075 ;
        RECT 100.960 96.060 101.280 96.320 ;
        RECT 106.955 96.260 107.245 96.305 ;
        RECT 107.860 96.260 108.180 96.320 ;
        RECT 111.630 96.305 111.770 97.140 ;
        RECT 128.575 97.140 130.705 97.280 ;
        RECT 128.575 97.095 128.865 97.140 ;
        RECT 129.020 97.080 129.340 97.140 ;
        RECT 130.415 97.095 130.705 97.140 ;
        RECT 134.540 97.080 134.860 97.340 ;
        RECT 139.615 97.280 139.905 97.325 ;
        RECT 136.930 97.140 139.905 97.280 ;
        RECT 129.940 96.940 130.260 97.000 ;
        RECT 136.930 96.940 137.070 97.140 ;
        RECT 139.615 97.095 139.905 97.140 ;
        RECT 140.075 97.280 140.365 97.325 ;
        RECT 140.980 97.280 141.300 97.340 ;
        RECT 140.075 97.140 141.300 97.280 ;
        RECT 140.075 97.095 140.365 97.140 ;
        RECT 125.430 96.800 130.260 96.940 ;
        RECT 117.980 96.600 118.300 96.660 ;
        RECT 123.040 96.600 123.360 96.660 ;
        RECT 125.430 96.600 125.570 96.800 ;
        RECT 129.940 96.740 130.260 96.800 ;
        RECT 134.170 96.800 137.070 96.940 ;
        RECT 134.170 96.660 134.310 96.800 ;
        RECT 137.775 96.755 138.065 96.985 ;
        RECT 139.690 96.940 139.830 97.095 ;
        RECT 140.980 97.080 141.300 97.140 ;
        RECT 141.900 97.280 142.220 97.340 ;
        RECT 141.900 97.140 147.190 97.280 ;
        RECT 141.900 97.080 142.220 97.140 ;
        RECT 141.455 96.940 141.745 96.985 ;
        RECT 139.690 96.800 141.745 96.940 ;
        RECT 141.455 96.755 141.745 96.800 ;
        RECT 129.495 96.600 129.785 96.645 ;
        RECT 130.400 96.600 130.720 96.660 ;
        RECT 117.980 96.460 123.360 96.600 ;
        RECT 117.980 96.400 118.300 96.460 ;
        RECT 123.040 96.400 123.360 96.460 ;
        RECT 124.970 96.460 125.570 96.600 ;
        RECT 129.110 96.460 130.720 96.600 ;
        RECT 106.955 96.120 108.180 96.260 ;
        RECT 106.955 96.075 107.245 96.120 ;
        RECT 107.860 96.060 108.180 96.120 ;
        RECT 111.555 96.075 111.845 96.305 ;
        RECT 112.475 96.260 112.765 96.305 ;
        RECT 112.920 96.260 113.240 96.320 ;
        RECT 112.475 96.120 113.240 96.260 ;
        RECT 112.475 96.075 112.765 96.120 ;
        RECT 112.920 96.060 113.240 96.120 ;
        RECT 115.680 96.060 116.000 96.320 ;
        RECT 122.120 96.060 122.440 96.320 ;
        RECT 124.970 96.305 125.110 96.460 ;
        RECT 124.895 96.075 125.185 96.305 ;
        RECT 125.355 96.260 125.645 96.305 ;
        RECT 128.100 96.260 128.420 96.320 ;
        RECT 129.110 96.305 129.250 96.460 ;
        RECT 129.495 96.415 129.785 96.460 ;
        RECT 130.400 96.400 130.720 96.460 ;
        RECT 134.080 96.400 134.400 96.660 ;
        RECT 136.840 96.600 137.160 96.660 ;
        RECT 136.010 96.460 137.160 96.600 ;
        RECT 137.850 96.600 137.990 96.755 ;
        RECT 145.580 96.740 145.900 97.000 ;
        RECT 140.535 96.600 140.825 96.645 ;
        RECT 137.850 96.460 142.130 96.600 ;
        RECT 125.355 96.120 128.420 96.260 ;
        RECT 125.355 96.075 125.645 96.120 ;
        RECT 128.100 96.060 128.420 96.120 ;
        RECT 129.035 96.075 129.325 96.305 ;
        RECT 129.940 96.260 130.260 96.320 ;
        RECT 130.875 96.260 131.165 96.305 ;
        RECT 129.940 96.120 131.165 96.260 ;
        RECT 129.940 96.060 130.260 96.120 ;
        RECT 130.875 96.075 131.165 96.120 ;
        RECT 134.170 96.120 135.230 96.260 ;
        RECT 115.770 95.920 115.910 96.060 ;
        RECT 86.330 95.780 115.910 95.920 ;
        RECT 122.210 95.920 122.350 96.060 ;
        RECT 134.170 95.920 134.310 96.120 ;
        RECT 122.210 95.780 134.310 95.920 ;
        RECT 88.540 95.720 88.860 95.780 ;
        RECT 134.540 95.720 134.860 95.980 ;
        RECT 135.090 95.920 135.230 96.120 ;
        RECT 135.460 96.060 135.780 96.320 ;
        RECT 136.010 96.305 136.150 96.460 ;
        RECT 136.840 96.400 137.160 96.460 ;
        RECT 140.535 96.415 140.825 96.460 ;
        RECT 135.935 96.075 136.225 96.305 ;
        RECT 137.300 96.060 137.620 96.320 ;
        RECT 137.760 96.260 138.080 96.320 ;
        RECT 138.235 96.260 138.525 96.305 ;
        RECT 137.760 96.120 138.525 96.260 ;
        RECT 137.760 96.060 138.080 96.120 ;
        RECT 138.235 96.075 138.525 96.120 ;
        RECT 138.680 96.260 139.000 96.320 ;
        RECT 139.155 96.260 139.445 96.305 ;
        RECT 138.680 96.120 139.445 96.260 ;
        RECT 138.680 96.060 139.000 96.120 ;
        RECT 139.155 96.075 139.445 96.120 ;
        RECT 140.980 96.060 141.300 96.320 ;
        RECT 141.990 96.305 142.130 96.460 ;
        RECT 143.740 96.400 144.060 96.660 ;
        RECT 147.050 96.645 147.190 97.140 ;
        RECT 146.975 96.415 147.265 96.645 ;
        RECT 141.915 96.075 142.205 96.305 ;
        RECT 143.830 96.260 143.970 96.400 ;
        RECT 142.910 96.120 143.970 96.260 ;
        RECT 142.910 95.980 143.050 96.120 ;
        RECT 147.880 96.060 148.200 96.320 ;
        RECT 142.820 95.920 143.140 95.980 ;
        RECT 135.090 95.780 143.140 95.920 ;
        RECT 142.820 95.720 143.140 95.780 ;
        RECT 143.740 95.720 144.060 95.980 ;
        RECT 148.815 95.920 149.105 95.965 ;
        RECT 151.100 95.920 151.420 95.980 ;
        RECT 148.815 95.780 151.420 95.920 ;
        RECT 148.815 95.735 149.105 95.780 ;
        RECT 151.100 95.720 151.420 95.780 ;
        RECT 31.960 95.580 32.280 95.640 ;
        RECT 26.530 95.440 32.280 95.580 ;
        RECT 31.960 95.380 32.280 95.440 ;
        RECT 40.700 95.580 41.020 95.640 ;
        RECT 43.000 95.580 43.320 95.640 ;
        RECT 40.700 95.440 43.320 95.580 ;
        RECT 40.700 95.380 41.020 95.440 ;
        RECT 43.000 95.380 43.320 95.440 ;
        RECT 53.120 95.380 53.440 95.640 ;
        RECT 78.895 95.580 79.185 95.625 ;
        RECT 86.700 95.580 87.020 95.640 ;
        RECT 78.895 95.440 87.020 95.580 ;
        RECT 78.895 95.395 79.185 95.440 ;
        RECT 86.700 95.380 87.020 95.440 ;
        RECT 88.080 95.580 88.400 95.640 ;
        RECT 94.980 95.580 95.300 95.640 ;
        RECT 110.160 95.580 110.480 95.640 ;
        RECT 88.080 95.440 110.480 95.580 ;
        RECT 88.080 95.380 88.400 95.440 ;
        RECT 94.980 95.380 95.300 95.440 ;
        RECT 110.160 95.380 110.480 95.440 ;
        RECT 112.000 95.380 112.320 95.640 ;
        RECT 115.695 95.580 115.985 95.625 ;
        RECT 117.060 95.580 117.380 95.640 ;
        RECT 115.695 95.440 117.380 95.580 ;
        RECT 115.695 95.395 115.985 95.440 ;
        RECT 117.060 95.380 117.380 95.440 ;
        RECT 124.420 95.380 124.740 95.640 ;
        RECT 126.735 95.580 127.025 95.625 ;
        RECT 128.100 95.580 128.420 95.640 ;
        RECT 126.735 95.440 128.420 95.580 ;
        RECT 126.735 95.395 127.025 95.440 ;
        RECT 128.100 95.380 128.420 95.440 ;
        RECT 129.480 95.380 129.800 95.640 ;
        RECT 146.040 95.380 146.360 95.640 ;
        RECT 22.690 94.760 157.810 95.240 ;
        RECT 30.580 94.560 30.900 94.620 ;
        RECT 36.115 94.560 36.405 94.605 ;
        RECT 30.580 94.420 36.405 94.560 ;
        RECT 30.580 94.360 30.900 94.420 ;
        RECT 36.115 94.375 36.405 94.420 ;
        RECT 38.950 94.420 43.690 94.560 ;
        RECT 32.435 94.220 32.725 94.265 ;
        RECT 34.275 94.220 34.565 94.265 ;
        RECT 32.435 94.080 34.565 94.220 ;
        RECT 32.435 94.035 32.725 94.080 ;
        RECT 34.275 94.035 34.565 94.080 ;
        RECT 35.180 94.020 35.500 94.280 ;
        RECT 36.560 94.220 36.880 94.280 ;
        RECT 37.035 94.220 37.325 94.265 ;
        RECT 36.560 94.080 37.325 94.220 ;
        RECT 36.560 94.020 36.880 94.080 ;
        RECT 37.035 94.035 37.325 94.080 ;
        RECT 37.480 94.220 37.800 94.280 ;
        RECT 38.950 94.265 39.090 94.420 ;
        RECT 37.955 94.220 38.245 94.265 ;
        RECT 37.480 94.080 38.245 94.220 ;
        RECT 37.480 94.020 37.800 94.080 ;
        RECT 37.955 94.035 38.245 94.080 ;
        RECT 38.875 94.035 39.165 94.265 ;
        RECT 39.410 94.080 42.390 94.220 ;
        RECT 33.815 93.880 34.105 93.925 ;
        RECT 35.270 93.880 35.410 94.020 ;
        RECT 33.815 93.740 35.410 93.880 ;
        RECT 35.655 93.880 35.945 93.925 ;
        RECT 36.100 93.880 36.420 93.940 ;
        RECT 35.655 93.740 36.420 93.880 ;
        RECT 33.815 93.695 34.105 93.740 ;
        RECT 35.655 93.695 35.945 93.740 ;
        RECT 36.100 93.680 36.420 93.740 ;
        RECT 32.435 93.540 32.725 93.585 ;
        RECT 34.720 93.540 35.040 93.600 ;
        RECT 32.435 93.400 35.040 93.540 ;
        RECT 32.435 93.355 32.725 93.400 ;
        RECT 34.720 93.340 35.040 93.400 ;
        RECT 34.275 93.200 34.565 93.245 ;
        RECT 35.640 93.200 35.960 93.260 ;
        RECT 34.275 93.060 35.960 93.200 ;
        RECT 34.275 93.015 34.565 93.060 ;
        RECT 35.640 93.000 35.960 93.060 ;
        RECT 33.355 92.860 33.645 92.905 ;
        RECT 36.190 92.860 36.330 93.680 ;
        RECT 37.940 93.540 38.260 93.600 ;
        RECT 39.410 93.540 39.550 94.080 ;
        RECT 39.795 93.695 40.085 93.925 ;
        RECT 37.940 93.400 39.550 93.540 ;
        RECT 37.940 93.340 38.260 93.400 ;
        RECT 39.870 93.200 40.010 93.695 ;
        RECT 40.700 93.680 41.020 93.940 ;
        RECT 42.250 93.925 42.390 94.080 ;
        RECT 42.095 93.760 42.390 93.925 ;
        RECT 43.550 93.880 43.690 94.420 ;
        RECT 43.935 94.375 44.225 94.605 ;
        RECT 44.010 94.220 44.150 94.375 ;
        RECT 51.740 94.360 52.060 94.620 ;
        RECT 67.380 94.360 67.700 94.620 ;
        RECT 68.300 94.360 68.620 94.620 ;
        RECT 82.560 94.360 82.880 94.620 ;
        RECT 90.840 94.360 91.160 94.620 ;
        RECT 94.520 94.560 94.840 94.620 ;
        RECT 91.390 94.420 94.840 94.560 ;
        RECT 44.010 94.080 46.910 94.220 ;
        RECT 44.395 93.880 44.685 93.925 ;
        RECT 42.095 93.695 42.385 93.760 ;
        RECT 43.550 93.740 44.685 93.880 ;
        RECT 44.395 93.695 44.685 93.740 ;
        RECT 45.300 93.680 45.620 93.940 ;
        RECT 46.770 93.925 46.910 94.080 ;
        RECT 46.695 93.695 46.985 93.925 ;
        RECT 52.675 93.880 52.965 93.925 ;
        RECT 53.135 93.880 53.425 93.925 ;
        RECT 52.675 93.740 53.425 93.880 ;
        RECT 52.675 93.695 52.965 93.740 ;
        RECT 53.135 93.695 53.425 93.740 ;
        RECT 54.040 93.680 54.360 93.940 ;
        RECT 68.390 93.925 68.530 94.360 ;
        RECT 82.100 94.220 82.420 94.280 ;
        RECT 81.270 94.080 82.420 94.220 ;
        RECT 82.650 94.220 82.790 94.360 ;
        RECT 82.650 94.080 83.250 94.220 ;
        RECT 68.315 93.695 68.605 93.925 ;
        RECT 79.340 93.680 79.660 93.940 ;
        RECT 81.270 93.925 81.410 94.080 ;
        RECT 82.100 94.020 82.420 94.080 ;
        RECT 79.815 93.695 80.105 93.925 ;
        RECT 81.195 93.695 81.485 93.925 ;
        RECT 41.620 93.340 41.940 93.600 ;
        RECT 47.615 93.540 47.905 93.585 ;
        RECT 54.975 93.540 55.265 93.585 ;
        RECT 64.160 93.540 64.480 93.600 ;
        RECT 47.615 93.400 64.480 93.540 ;
        RECT 47.615 93.355 47.905 93.400 ;
        RECT 54.975 93.355 55.265 93.400 ;
        RECT 64.160 93.340 64.480 93.400 ;
        RECT 77.515 93.355 77.805 93.585 ;
        RECT 79.890 93.540 80.030 93.695 ;
        RECT 81.640 93.680 81.960 93.940 ;
        RECT 82.560 93.680 82.880 93.940 ;
        RECT 83.110 93.925 83.250 94.080 ;
        RECT 90.930 93.925 91.070 94.360 ;
        RECT 91.390 93.925 91.530 94.420 ;
        RECT 94.520 94.360 94.840 94.420 ;
        RECT 112.000 94.560 112.320 94.620 ;
        RECT 112.000 94.420 115.450 94.560 ;
        RECT 112.000 94.360 112.320 94.420 ;
        RECT 92.310 94.080 95.670 94.220 ;
        RECT 92.310 93.925 92.450 94.080 ;
        RECT 95.530 93.940 95.670 94.080 ;
        RECT 104.180 94.020 104.500 94.280 ;
        RECT 105.100 94.220 105.420 94.280 ;
        RECT 105.100 94.080 114.990 94.220 ;
        RECT 105.100 94.020 105.420 94.080 ;
        RECT 83.035 93.695 83.325 93.925 ;
        RECT 90.855 93.695 91.145 93.925 ;
        RECT 91.315 93.695 91.605 93.925 ;
        RECT 92.235 93.695 92.525 93.925 ;
        RECT 92.680 93.680 93.000 93.940 ;
        RECT 94.060 93.680 94.380 93.940 ;
        RECT 95.440 93.680 95.760 93.940 ;
        RECT 95.900 93.880 96.220 93.940 ;
        RECT 97.295 93.880 97.585 93.925 ;
        RECT 95.900 93.740 97.585 93.880 ;
        RECT 104.270 93.880 104.410 94.020 ;
        RECT 107.490 93.925 107.630 94.080 ;
        RECT 106.080 93.880 106.370 93.925 ;
        RECT 104.270 93.740 106.370 93.880 ;
        RECT 95.900 93.680 96.220 93.740 ;
        RECT 97.295 93.695 97.585 93.740 ;
        RECT 106.080 93.695 106.370 93.740 ;
        RECT 107.415 93.695 107.705 93.925 ;
        RECT 110.620 93.880 110.940 93.940 ;
        RECT 113.440 93.880 113.730 93.925 ;
        RECT 110.620 93.740 113.730 93.880 ;
        RECT 110.620 93.680 110.940 93.740 ;
        RECT 113.440 93.695 113.730 93.740 ;
        RECT 80.720 93.540 81.040 93.600 ;
        RECT 84.400 93.540 84.720 93.600 ;
        RECT 79.890 93.400 84.720 93.540 ;
        RECT 42.080 93.200 42.400 93.260 ;
        RECT 77.590 93.200 77.730 93.355 ;
        RECT 80.720 93.340 81.040 93.400 ;
        RECT 84.400 93.340 84.720 93.400 ;
        RECT 94.535 93.355 94.825 93.585 ;
        RECT 92.680 93.200 93.000 93.260 ;
        RECT 39.870 93.060 42.400 93.200 ;
        RECT 42.080 93.000 42.400 93.060 ;
        RECT 44.470 93.060 93.000 93.200 ;
        RECT 94.610 93.200 94.750 93.355 ;
        RECT 96.820 93.340 97.140 93.600 ;
        RECT 114.850 93.585 114.990 94.080 ;
        RECT 115.310 93.940 115.450 94.420 ;
        RECT 115.680 94.360 116.000 94.620 ;
        RECT 124.420 94.360 124.740 94.620 ;
        RECT 129.020 94.560 129.340 94.620 ;
        RECT 129.495 94.560 129.785 94.605 ;
        RECT 129.020 94.420 129.785 94.560 ;
        RECT 129.020 94.360 129.340 94.420 ;
        RECT 129.495 94.375 129.785 94.420 ;
        RECT 130.400 94.560 130.720 94.620 ;
        RECT 130.875 94.560 131.165 94.605 ;
        RECT 130.400 94.420 131.165 94.560 ;
        RECT 130.400 94.360 130.720 94.420 ;
        RECT 130.875 94.375 131.165 94.420 ;
        RECT 133.160 94.560 133.480 94.620 ;
        RECT 133.635 94.560 133.925 94.605 ;
        RECT 138.680 94.560 139.000 94.620 ;
        RECT 133.160 94.420 139.000 94.560 ;
        RECT 133.160 94.360 133.480 94.420 ;
        RECT 133.635 94.375 133.925 94.420 ;
        RECT 115.770 94.220 115.910 94.360 ;
        RECT 124.510 94.220 124.650 94.360 ;
        RECT 132.715 94.220 133.005 94.265 ;
        RECT 134.555 94.220 134.845 94.265 ;
        RECT 115.770 94.080 117.290 94.220 ;
        RECT 124.510 94.080 127.410 94.220 ;
        RECT 115.220 93.680 115.540 93.940 ;
        RECT 115.695 93.880 115.985 93.925 ;
        RECT 116.140 93.880 116.460 93.940 ;
        RECT 115.695 93.740 116.460 93.880 ;
        RECT 115.695 93.695 115.985 93.740 ;
        RECT 116.140 93.680 116.460 93.740 ;
        RECT 116.600 93.680 116.920 93.940 ;
        RECT 117.150 93.925 117.290 94.080 ;
        RECT 127.270 93.925 127.410 94.080 ;
        RECT 128.650 94.080 129.710 94.220 ;
        RECT 117.075 93.695 117.365 93.925 ;
        RECT 119.790 93.880 120.080 93.925 ;
        RECT 126.275 93.880 126.565 93.925 ;
        RECT 119.790 93.740 126.565 93.880 ;
        RECT 119.790 93.695 120.080 93.740 ;
        RECT 126.275 93.695 126.565 93.740 ;
        RECT 127.195 93.695 127.485 93.925 ;
        RECT 128.100 93.680 128.420 93.940 ;
        RECT 128.650 93.925 128.790 94.080 ;
        RECT 129.570 93.940 129.710 94.080 ;
        RECT 130.030 94.080 131.550 94.220 ;
        RECT 128.575 93.695 128.865 93.925 ;
        RECT 129.035 93.695 129.325 93.925 ;
        RECT 102.825 93.540 103.115 93.585 ;
        RECT 105.345 93.540 105.635 93.585 ;
        RECT 106.535 93.540 106.825 93.585 ;
        RECT 102.825 93.400 106.825 93.540 ;
        RECT 102.825 93.355 103.115 93.400 ;
        RECT 105.345 93.355 105.635 93.400 ;
        RECT 106.535 93.355 106.825 93.400 ;
        RECT 110.185 93.540 110.475 93.585 ;
        RECT 112.705 93.540 112.995 93.585 ;
        RECT 113.895 93.540 114.185 93.585 ;
        RECT 110.185 93.400 114.185 93.540 ;
        RECT 110.185 93.355 110.475 93.400 ;
        RECT 112.705 93.355 112.995 93.400 ;
        RECT 113.895 93.355 114.185 93.400 ;
        RECT 114.775 93.540 115.065 93.585 ;
        RECT 118.455 93.540 118.745 93.585 ;
        RECT 114.775 93.400 118.745 93.540 ;
        RECT 114.775 93.355 115.065 93.400 ;
        RECT 117.150 93.260 117.290 93.400 ;
        RECT 118.455 93.355 118.745 93.400 ;
        RECT 119.335 93.540 119.625 93.585 ;
        RECT 120.525 93.540 120.815 93.585 ;
        RECT 123.045 93.540 123.335 93.585 ;
        RECT 119.335 93.400 123.335 93.540 ;
        RECT 119.335 93.355 119.625 93.400 ;
        RECT 120.525 93.355 120.815 93.400 ;
        RECT 123.045 93.355 123.335 93.400 ;
        RECT 129.110 93.540 129.250 93.695 ;
        RECT 129.480 93.680 129.800 93.940 ;
        RECT 130.030 93.925 130.170 94.080 ;
        RECT 131.410 93.925 131.550 94.080 ;
        RECT 132.715 94.080 134.845 94.220 ;
        RECT 135.550 94.220 135.690 94.420 ;
        RECT 138.680 94.360 139.000 94.420 ;
        RECT 139.155 94.560 139.445 94.605 ;
        RECT 140.980 94.560 141.300 94.620 ;
        RECT 139.155 94.420 141.300 94.560 ;
        RECT 139.155 94.375 139.445 94.420 ;
        RECT 140.980 94.360 141.300 94.420 ;
        RECT 149.720 94.360 150.040 94.620 ;
        RECT 151.100 94.560 151.420 94.620 ;
        RECT 151.100 94.420 153.170 94.560 ;
        RECT 151.100 94.360 151.420 94.420 ;
        RECT 135.550 94.080 136.150 94.220 ;
        RECT 132.715 94.035 133.005 94.080 ;
        RECT 134.555 94.035 134.845 94.080 ;
        RECT 129.955 93.695 130.245 93.925 ;
        RECT 130.415 93.695 130.705 93.925 ;
        RECT 131.335 93.880 131.625 93.925 ;
        RECT 132.240 93.880 132.560 93.940 ;
        RECT 131.335 93.740 132.560 93.880 ;
        RECT 131.335 93.695 131.625 93.740 ;
        RECT 130.490 93.540 130.630 93.695 ;
        RECT 132.240 93.680 132.560 93.740 ;
        RECT 133.620 93.680 133.940 93.940 ;
        RECT 134.080 93.880 134.400 93.940 ;
        RECT 136.010 93.925 136.150 94.080 ;
        RECT 137.300 94.020 137.620 94.280 ;
        RECT 135.475 93.880 135.765 93.925 ;
        RECT 134.080 93.740 135.765 93.880 ;
        RECT 134.080 93.680 134.400 93.740 ;
        RECT 135.475 93.695 135.765 93.740 ;
        RECT 135.935 93.695 136.225 93.925 ;
        RECT 137.760 93.880 138.080 93.940 ;
        RECT 138.235 93.880 138.525 93.925 ;
        RECT 137.760 93.740 138.525 93.880 ;
        RECT 137.760 93.680 138.080 93.740 ;
        RECT 138.235 93.695 138.525 93.740 ;
        RECT 129.110 93.400 130.630 93.540 ;
        RECT 133.710 93.540 133.850 93.680 ;
        RECT 134.555 93.540 134.845 93.585 ;
        RECT 133.710 93.400 134.845 93.540 ;
        RECT 94.980 93.200 95.300 93.260 ;
        RECT 100.515 93.200 100.805 93.245 ;
        RECT 94.610 93.060 100.805 93.200 ;
        RECT 33.355 92.720 36.330 92.860 ;
        RECT 41.160 92.860 41.480 92.920 ;
        RECT 44.470 92.860 44.610 93.060 ;
        RECT 92.680 93.000 93.000 93.060 ;
        RECT 94.980 93.000 95.300 93.060 ;
        RECT 100.515 93.015 100.805 93.060 ;
        RECT 103.260 93.200 103.550 93.245 ;
        RECT 104.830 93.200 105.120 93.245 ;
        RECT 106.930 93.200 107.220 93.245 ;
        RECT 103.260 93.060 107.220 93.200 ;
        RECT 103.260 93.015 103.550 93.060 ;
        RECT 104.830 93.015 105.120 93.060 ;
        RECT 106.930 93.015 107.220 93.060 ;
        RECT 110.620 93.200 110.910 93.245 ;
        RECT 112.190 93.200 112.480 93.245 ;
        RECT 114.290 93.200 114.580 93.245 ;
        RECT 110.620 93.060 114.580 93.200 ;
        RECT 110.620 93.015 110.910 93.060 ;
        RECT 112.190 93.015 112.480 93.060 ;
        RECT 114.290 93.015 114.580 93.060 ;
        RECT 117.060 93.000 117.380 93.260 ;
        RECT 118.940 93.200 119.230 93.245 ;
        RECT 121.040 93.200 121.330 93.245 ;
        RECT 122.610 93.200 122.900 93.245 ;
        RECT 118.940 93.060 122.900 93.200 ;
        RECT 118.940 93.015 119.230 93.060 ;
        RECT 121.040 93.015 121.330 93.060 ;
        RECT 122.610 93.015 122.900 93.060 ;
        RECT 125.355 93.200 125.645 93.245 ;
        RECT 129.110 93.200 129.250 93.400 ;
        RECT 134.555 93.355 134.845 93.400 ;
        RECT 125.355 93.060 129.250 93.200 ;
        RECT 125.355 93.015 125.645 93.060 ;
        RECT 41.160 92.720 44.610 92.860 ;
        RECT 33.355 92.675 33.645 92.720 ;
        RECT 41.160 92.660 41.480 92.720 ;
        RECT 44.840 92.660 45.160 92.920 ;
        RECT 45.760 92.660 46.080 92.920 ;
        RECT 78.420 92.660 78.740 92.920 ;
        RECT 80.275 92.860 80.565 92.905 ;
        RECT 81.640 92.860 81.960 92.920 ;
        RECT 80.275 92.720 81.960 92.860 ;
        RECT 80.275 92.675 80.565 92.720 ;
        RECT 81.640 92.660 81.960 92.720 ;
        RECT 89.935 92.860 90.225 92.905 ;
        RECT 90.840 92.860 91.160 92.920 ;
        RECT 89.935 92.720 91.160 92.860 ;
        RECT 89.935 92.675 90.225 92.720 ;
        RECT 90.840 92.660 91.160 92.720 ;
        RECT 95.455 92.860 95.745 92.905 ;
        RECT 95.900 92.860 96.220 92.920 ;
        RECT 95.455 92.720 96.220 92.860 ;
        RECT 95.455 92.675 95.745 92.720 ;
        RECT 95.900 92.660 96.220 92.720 ;
        RECT 98.660 92.660 98.980 92.920 ;
        RECT 104.180 92.860 104.500 92.920 ;
        RECT 107.875 92.860 108.165 92.905 ;
        RECT 104.180 92.720 108.165 92.860 ;
        RECT 104.180 92.660 104.500 92.720 ;
        RECT 107.875 92.675 108.165 92.720 ;
        RECT 117.995 92.860 118.285 92.905 ;
        RECT 122.120 92.860 122.440 92.920 ;
        RECT 117.995 92.720 122.440 92.860 ;
        RECT 117.995 92.675 118.285 92.720 ;
        RECT 122.120 92.660 122.440 92.720 ;
        RECT 132.700 92.660 133.020 92.920 ;
        RECT 138.770 92.860 138.910 94.360 ;
        RECT 140.535 94.220 140.825 94.265 ;
        RECT 143.740 94.220 144.060 94.280 ;
        RECT 140.535 94.080 144.060 94.220 ;
        RECT 149.810 94.220 149.950 94.360 ;
        RECT 149.810 94.080 151.330 94.220 ;
        RECT 140.535 94.035 140.825 94.080 ;
        RECT 143.740 94.020 144.060 94.080 ;
        RECT 140.075 93.695 140.365 93.925 ;
        RECT 140.995 93.880 141.285 93.925 ;
        RECT 142.375 93.880 142.665 93.925 ;
        RECT 145.580 93.880 145.900 93.940 ;
        RECT 147.420 93.880 147.740 93.940 ;
        RECT 151.190 93.925 151.330 94.080 ;
        RECT 153.030 93.925 153.170 94.420 ;
        RECT 140.995 93.740 142.130 93.880 ;
        RECT 140.995 93.695 141.285 93.740 ;
        RECT 140.150 93.540 140.290 93.695 ;
        RECT 141.440 93.540 141.760 93.600 ;
        RECT 140.150 93.400 141.760 93.540 ;
        RECT 141.440 93.340 141.760 93.400 ;
        RECT 141.990 93.200 142.130 93.740 ;
        RECT 142.375 93.740 147.740 93.880 ;
        RECT 142.375 93.695 142.665 93.740 ;
        RECT 145.580 93.680 145.900 93.740 ;
        RECT 147.420 93.680 147.740 93.740 ;
        RECT 149.835 93.880 150.125 93.925 ;
        RECT 149.835 93.740 150.870 93.880 ;
        RECT 149.835 93.695 150.125 93.740 ;
        RECT 143.755 93.540 144.045 93.585 ;
        RECT 145.120 93.540 145.440 93.600 ;
        RECT 143.755 93.400 145.440 93.540 ;
        RECT 143.755 93.355 144.045 93.400 ;
        RECT 145.120 93.340 145.440 93.400 ;
        RECT 146.525 93.540 146.815 93.585 ;
        RECT 149.045 93.540 149.335 93.585 ;
        RECT 150.235 93.540 150.525 93.585 ;
        RECT 146.525 93.400 150.525 93.540 ;
        RECT 150.730 93.540 150.870 93.740 ;
        RECT 151.115 93.695 151.405 93.925 ;
        RECT 152.955 93.695 153.245 93.925 ;
        RECT 150.730 93.400 152.250 93.540 ;
        RECT 146.525 93.355 146.815 93.400 ;
        RECT 149.045 93.355 149.335 93.400 ;
        RECT 150.235 93.355 150.525 93.400 ;
        RECT 152.110 93.245 152.250 93.400 ;
        RECT 146.960 93.200 147.250 93.245 ;
        RECT 148.530 93.200 148.820 93.245 ;
        RECT 150.630 93.200 150.920 93.245 ;
        RECT 141.990 93.060 144.430 93.200 ;
        RECT 141.455 92.860 141.745 92.905 ;
        RECT 138.770 92.720 141.745 92.860 ;
        RECT 141.455 92.675 141.745 92.720 ;
        RECT 143.295 92.860 143.585 92.905 ;
        RECT 143.740 92.860 144.060 92.920 ;
        RECT 144.290 92.905 144.430 93.060 ;
        RECT 146.960 93.060 150.920 93.200 ;
        RECT 146.960 93.015 147.250 93.060 ;
        RECT 148.530 93.015 148.820 93.060 ;
        RECT 150.630 93.015 150.920 93.060 ;
        RECT 152.035 93.015 152.325 93.245 ;
        RECT 143.295 92.720 144.060 92.860 ;
        RECT 143.295 92.675 143.585 92.720 ;
        RECT 143.740 92.660 144.060 92.720 ;
        RECT 144.215 92.860 144.505 92.905 ;
        RECT 146.500 92.860 146.820 92.920 ;
        RECT 144.215 92.720 146.820 92.860 ;
        RECT 144.215 92.675 144.505 92.720 ;
        RECT 146.500 92.660 146.820 92.720 ;
        RECT 22.690 92.040 157.010 92.520 ;
        RECT 31.960 91.640 32.280 91.900 ;
        RECT 36.100 91.840 36.420 91.900 ;
        RECT 41.175 91.840 41.465 91.885 ;
        RECT 41.620 91.840 41.940 91.900 ;
        RECT 36.100 91.700 40.930 91.840 ;
        RECT 36.100 91.640 36.420 91.700 ;
        RECT 37.570 91.545 37.710 91.700 ;
        RECT 40.790 91.560 40.930 91.700 ;
        RECT 41.175 91.700 41.940 91.840 ;
        RECT 41.175 91.655 41.465 91.700 ;
        RECT 41.620 91.640 41.940 91.700 ;
        RECT 42.555 91.840 42.845 91.885 ;
        RECT 45.300 91.840 45.620 91.900 ;
        RECT 42.555 91.700 45.620 91.840 ;
        RECT 42.555 91.655 42.845 91.700 ;
        RECT 37.495 91.315 37.785 91.545 ;
        RECT 37.940 91.300 38.260 91.560 ;
        RECT 40.700 91.300 41.020 91.560 ;
        RECT 26.915 91.160 27.205 91.205 ;
        RECT 27.820 91.160 28.140 91.220 ;
        RECT 41.160 91.160 41.480 91.220 ;
        RECT 26.915 91.020 41.480 91.160 ;
        RECT 26.915 90.975 27.205 91.020 ;
        RECT 27.820 90.960 28.140 91.020 ;
        RECT 41.160 90.960 41.480 91.020 ;
        RECT 41.635 91.160 41.925 91.205 ;
        RECT 42.630 91.160 42.770 91.655 ;
        RECT 45.300 91.640 45.620 91.700 ;
        RECT 45.760 91.640 46.080 91.900 ;
        RECT 53.135 91.840 53.425 91.885 ;
        RECT 54.040 91.840 54.360 91.900 ;
        RECT 53.135 91.700 54.360 91.840 ;
        RECT 53.135 91.655 53.425 91.700 ;
        RECT 54.040 91.640 54.360 91.700 ;
        RECT 78.420 91.840 78.740 91.900 ;
        RECT 78.420 91.700 83.710 91.840 ;
        RECT 78.420 91.640 78.740 91.700 ;
        RECT 43.000 91.300 43.320 91.560 ;
        RECT 41.635 91.020 42.770 91.160 ;
        RECT 41.635 90.975 41.925 91.020 ;
        RECT 29.200 90.620 29.520 90.880 ;
        RECT 30.580 90.620 30.900 90.880 ;
        RECT 31.515 90.820 31.805 90.865 ;
        RECT 36.115 90.820 36.405 90.865 ;
        RECT 31.515 90.680 36.405 90.820 ;
        RECT 31.515 90.635 31.805 90.680 ;
        RECT 36.115 90.635 36.405 90.680 ;
        RECT 37.035 90.635 37.325 90.865 ;
        RECT 28.740 90.480 29.060 90.540 ;
        RECT 31.590 90.480 31.730 90.635 ;
        RECT 28.740 90.340 31.730 90.480 ;
        RECT 28.740 90.280 29.060 90.340 ;
        RECT 32.420 90.280 32.740 90.540 ;
        RECT 35.180 90.480 35.500 90.540 ;
        RECT 37.110 90.480 37.250 90.635 ;
        RECT 38.400 90.620 38.720 90.880 ;
        RECT 40.255 90.635 40.545 90.865 ;
        RECT 40.330 90.480 40.470 90.635 ;
        RECT 40.700 90.620 41.020 90.880 ;
        RECT 42.095 90.820 42.385 90.865 ;
        RECT 42.540 90.820 42.860 90.880 ;
        RECT 43.090 90.865 43.230 91.300 ;
        RECT 42.095 90.680 42.860 90.820 ;
        RECT 42.095 90.635 42.385 90.680 ;
        RECT 42.540 90.620 42.860 90.680 ;
        RECT 43.015 90.635 43.305 90.865 ;
        RECT 45.850 90.820 45.990 91.640 ;
        RECT 77.960 91.500 78.250 91.545 ;
        RECT 79.530 91.500 79.820 91.545 ;
        RECT 81.630 91.500 81.920 91.545 ;
        RECT 77.960 91.360 81.920 91.500 ;
        RECT 77.960 91.315 78.250 91.360 ;
        RECT 79.530 91.315 79.820 91.360 ;
        RECT 81.630 91.315 81.920 91.360 ;
        RECT 54.960 90.960 55.280 91.220 ;
        RECT 64.160 91.160 64.480 91.220 ;
        RECT 77.525 91.160 77.815 91.205 ;
        RECT 80.045 91.160 80.335 91.205 ;
        RECT 81.235 91.160 81.525 91.205 ;
        RECT 83.020 91.160 83.340 91.220 ;
        RECT 64.160 91.020 72.210 91.160 ;
        RECT 64.160 90.960 64.480 91.020 ;
        RECT 46.235 90.820 46.525 90.865 ;
        RECT 45.850 90.680 46.525 90.820 ;
        RECT 46.235 90.635 46.525 90.680 ;
        RECT 54.500 90.620 54.820 90.880 ;
        RECT 63.240 90.620 63.560 90.880 ;
        RECT 70.600 90.620 70.920 90.880 ;
        RECT 71.075 90.635 71.365 90.865 ;
        RECT 57.260 90.480 57.580 90.540 ;
        RECT 35.180 90.340 57.580 90.480 ;
        RECT 35.180 90.280 35.500 90.340 ;
        RECT 57.260 90.280 57.580 90.340 ;
        RECT 69.220 90.280 69.540 90.540 ;
        RECT 28.280 89.940 28.600 90.200 ;
        RECT 40.700 90.140 41.020 90.200 ;
        RECT 44.840 90.140 45.160 90.200 ;
        RECT 40.700 90.000 45.160 90.140 ;
        RECT 40.700 89.940 41.020 90.000 ;
        RECT 44.840 89.940 45.160 90.000 ;
        RECT 46.680 90.140 47.000 90.200 ;
        RECT 47.155 90.140 47.445 90.185 ;
        RECT 46.680 90.000 47.445 90.140 ;
        RECT 46.680 89.940 47.000 90.000 ;
        RECT 47.155 89.955 47.445 90.000 ;
        RECT 62.320 89.940 62.640 90.200 ;
        RECT 68.300 90.140 68.620 90.200 ;
        RECT 71.150 90.140 71.290 90.635 ;
        RECT 71.520 90.620 71.840 90.880 ;
        RECT 72.070 90.480 72.210 91.020 ;
        RECT 77.525 91.020 81.525 91.160 ;
        RECT 77.525 90.975 77.815 91.020 ;
        RECT 80.045 90.975 80.335 91.020 ;
        RECT 81.235 90.975 81.525 91.020 ;
        RECT 81.730 91.020 83.340 91.160 ;
        RECT 72.440 90.820 72.760 90.880 ;
        RECT 81.730 90.820 81.870 91.020 ;
        RECT 83.020 90.960 83.340 91.020 ;
        RECT 72.440 90.680 81.870 90.820 ;
        RECT 72.440 90.620 72.760 90.680 ;
        RECT 82.100 90.620 82.420 90.880 ;
        RECT 83.570 90.865 83.710 91.700 ;
        RECT 84.400 91.640 84.720 91.900 ;
        RECT 88.080 91.640 88.400 91.900 ;
        RECT 92.680 91.640 93.000 91.900 ;
        RECT 98.660 91.640 98.980 91.900 ;
        RECT 100.960 91.840 101.280 91.900 ;
        RECT 101.435 91.840 101.725 91.885 ;
        RECT 100.960 91.700 101.725 91.840 ;
        RECT 100.960 91.640 101.280 91.700 ;
        RECT 101.435 91.655 101.725 91.700 ;
        RECT 107.860 91.640 108.180 91.900 ;
        RECT 110.160 91.840 110.480 91.900 ;
        RECT 137.300 91.840 137.620 91.900 ;
        RECT 138.235 91.840 138.525 91.885 ;
        RECT 110.160 91.700 137.070 91.840 ;
        RECT 110.160 91.640 110.480 91.700 ;
        RECT 88.170 91.160 88.310 91.640 ;
        RECT 84.490 91.020 88.310 91.160 ;
        RECT 83.495 90.635 83.785 90.865 ;
        RECT 80.890 90.480 81.180 90.525 ;
        RECT 82.575 90.480 82.865 90.525 ;
        RECT 72.070 90.340 75.890 90.480 ;
        RECT 68.300 90.000 71.290 90.140 ;
        RECT 68.300 89.940 68.620 90.000 ;
        RECT 75.200 89.940 75.520 90.200 ;
        RECT 75.750 90.140 75.890 90.340 ;
        RECT 80.890 90.340 82.865 90.480 ;
        RECT 80.890 90.295 81.180 90.340 ;
        RECT 82.575 90.295 82.865 90.340 ;
        RECT 84.490 90.140 84.630 91.020 ;
        RECT 84.860 90.820 85.180 90.880 ;
        RECT 92.220 90.820 92.540 90.880 ;
        RECT 84.860 90.680 92.540 90.820 ;
        RECT 92.770 90.820 92.910 91.640 ;
        RECT 98.750 91.160 98.890 91.640 ;
        RECT 117.980 91.500 118.300 91.560 ;
        RECT 106.110 91.360 118.300 91.500 ;
        RECT 98.750 91.020 100.730 91.160 ;
        RECT 100.590 90.865 100.730 91.020 ;
        RECT 106.110 90.865 106.250 91.360 ;
        RECT 117.980 91.300 118.300 91.360 ;
        RECT 131.820 91.500 132.110 91.545 ;
        RECT 133.920 91.500 134.210 91.545 ;
        RECT 135.490 91.500 135.780 91.545 ;
        RECT 131.820 91.360 135.780 91.500 ;
        RECT 136.930 91.500 137.070 91.700 ;
        RECT 137.300 91.700 138.525 91.840 ;
        RECT 137.300 91.640 137.620 91.700 ;
        RECT 138.235 91.655 138.525 91.700 ;
        RECT 146.515 91.840 146.805 91.885 ;
        RECT 147.880 91.840 148.200 91.900 ;
        RECT 146.515 91.700 148.200 91.840 ;
        RECT 146.515 91.655 146.805 91.700 ;
        RECT 147.880 91.640 148.200 91.700 ;
        RECT 141.900 91.500 142.220 91.560 ;
        RECT 136.930 91.360 142.220 91.500 ;
        RECT 131.820 91.315 132.110 91.360 ;
        RECT 133.920 91.315 134.210 91.360 ;
        RECT 135.490 91.315 135.780 91.360 ;
        RECT 141.900 91.300 142.220 91.360 ;
        RECT 115.220 91.160 115.540 91.220 ;
        RECT 118.915 91.160 119.205 91.205 ;
        RECT 115.220 91.020 119.205 91.160 ;
        RECT 115.220 90.960 115.540 91.020 ;
        RECT 118.915 90.975 119.205 91.020 ;
        RECT 132.215 91.160 132.505 91.205 ;
        RECT 133.405 91.160 133.695 91.205 ;
        RECT 135.925 91.160 136.215 91.205 ;
        RECT 132.215 91.020 136.215 91.160 ;
        RECT 132.215 90.975 132.505 91.020 ;
        RECT 133.405 90.975 133.695 91.020 ;
        RECT 135.925 90.975 136.215 91.020 ;
        RECT 141.440 90.960 141.760 91.220 ;
        RECT 145.595 91.160 145.885 91.205 ;
        RECT 146.040 91.160 146.360 91.220 ;
        RECT 145.595 91.020 146.360 91.160 ;
        RECT 145.595 90.975 145.885 91.020 ;
        RECT 146.040 90.960 146.360 91.020 ;
        RECT 146.500 91.160 146.820 91.220 ;
        RECT 146.500 91.020 148.570 91.160 ;
        RECT 146.500 90.960 146.820 91.020 ;
        RECT 99.595 90.820 99.885 90.865 ;
        RECT 92.770 90.680 99.885 90.820 ;
        RECT 84.860 90.620 85.180 90.680 ;
        RECT 92.220 90.620 92.540 90.680 ;
        RECT 99.595 90.635 99.885 90.680 ;
        RECT 100.515 90.635 100.805 90.865 ;
        RECT 106.035 90.820 106.325 90.865 ;
        RECT 104.730 90.680 106.325 90.820 ;
        RECT 99.670 90.480 99.810 90.635 ;
        RECT 104.730 90.480 104.870 90.680 ;
        RECT 106.035 90.635 106.325 90.680 ;
        RECT 106.955 90.635 107.245 90.865 ;
        RECT 114.775 90.820 115.065 90.865 ;
        RECT 115.680 90.820 116.000 90.880 ;
        RECT 114.775 90.680 116.000 90.820 ;
        RECT 114.775 90.635 115.065 90.680 ;
        RECT 99.670 90.340 104.870 90.480 ;
        RECT 105.100 90.480 105.420 90.540 ;
        RECT 107.030 90.480 107.170 90.635 ;
        RECT 115.680 90.620 116.000 90.680 ;
        RECT 116.600 90.620 116.920 90.880 ;
        RECT 117.535 90.635 117.825 90.865 ;
        RECT 105.100 90.340 107.170 90.480 ;
        RECT 116.140 90.480 116.460 90.540 ;
        RECT 117.610 90.480 117.750 90.635 ;
        RECT 128.100 90.620 128.420 90.880 ;
        RECT 131.335 90.820 131.625 90.865 ;
        RECT 138.680 90.820 139.000 90.880 ;
        RECT 131.335 90.680 139.000 90.820 ;
        RECT 131.335 90.635 131.625 90.680 ;
        RECT 138.680 90.620 139.000 90.680 ;
        RECT 132.700 90.525 133.020 90.540 ;
        RECT 132.670 90.480 133.020 90.525 ;
        RECT 116.140 90.340 117.750 90.480 ;
        RECT 132.505 90.340 133.020 90.480 ;
        RECT 141.530 90.480 141.670 90.960 ;
        RECT 145.120 90.820 145.440 90.880 ;
        RECT 146.960 90.820 147.280 90.880 ;
        RECT 148.430 90.865 148.570 91.020 ;
        RECT 145.120 90.680 147.280 90.820 ;
        RECT 145.120 90.620 145.440 90.680 ;
        RECT 146.960 90.620 147.280 90.680 ;
        RECT 147.435 90.635 147.725 90.865 ;
        RECT 148.355 90.635 148.645 90.865 ;
        RECT 147.510 90.480 147.650 90.635 ;
        RECT 141.530 90.340 147.650 90.480 ;
        RECT 105.100 90.280 105.420 90.340 ;
        RECT 116.140 90.280 116.460 90.340 ;
        RECT 132.670 90.295 133.020 90.340 ;
        RECT 132.700 90.280 133.020 90.295 ;
        RECT 75.750 90.000 84.630 90.140 ;
        RECT 118.455 90.140 118.745 90.185 ;
        RECT 121.660 90.140 121.980 90.200 ;
        RECT 118.455 90.000 121.980 90.140 ;
        RECT 118.455 89.955 118.745 90.000 ;
        RECT 121.660 89.940 121.980 90.000 ;
        RECT 147.420 89.940 147.740 90.200 ;
        RECT 22.690 89.320 157.810 89.800 ;
        RECT 29.200 89.120 29.520 89.180 ;
        RECT 31.515 89.120 31.805 89.165 ;
        RECT 29.200 88.980 31.805 89.120 ;
        RECT 29.200 88.920 29.520 88.980 ;
        RECT 31.515 88.935 31.805 88.980 ;
        RECT 34.720 89.120 35.040 89.180 ;
        RECT 54.515 89.120 54.805 89.165 ;
        RECT 54.960 89.120 55.280 89.180 ;
        RECT 34.720 88.980 54.270 89.120 ;
        RECT 34.720 88.920 35.040 88.980 ;
        RECT 34.260 88.780 34.580 88.840 ;
        RECT 42.540 88.780 42.860 88.840 ;
        RECT 46.680 88.825 47.000 88.840 ;
        RECT 46.680 88.780 47.030 88.825 ;
        RECT 24.230 88.640 34.580 88.780 ;
        RECT 24.230 88.485 24.370 88.640 ;
        RECT 34.260 88.580 34.580 88.640 ;
        RECT 36.650 88.640 38.170 88.780 ;
        RECT 25.520 88.485 25.840 88.500 ;
        RECT 24.155 88.255 24.445 88.485 ;
        RECT 25.490 88.255 25.840 88.485 ;
        RECT 25.520 88.240 25.840 88.255 ;
        RECT 32.420 88.440 32.740 88.500 ;
        RECT 33.815 88.440 34.105 88.485 ;
        RECT 32.420 88.300 34.105 88.440 ;
        RECT 32.420 88.240 32.740 88.300 ;
        RECT 33.815 88.255 34.105 88.300 ;
        RECT 35.655 88.255 35.945 88.485 ;
        RECT 36.115 88.440 36.405 88.485 ;
        RECT 36.650 88.440 36.790 88.640 ;
        RECT 38.030 88.500 38.170 88.640 ;
        RECT 39.870 88.640 42.860 88.780 ;
        RECT 46.530 88.640 47.030 88.780 ;
        RECT 54.130 88.780 54.270 88.980 ;
        RECT 54.515 88.980 55.280 89.120 ;
        RECT 54.515 88.935 54.805 88.980 ;
        RECT 54.960 88.920 55.280 88.980 ;
        RECT 57.260 88.920 57.580 89.180 ;
        RECT 70.140 88.920 70.460 89.180 ;
        RECT 71.520 89.120 71.840 89.180 ;
        RECT 71.995 89.120 72.285 89.165 ;
        RECT 71.520 88.980 72.285 89.120 ;
        RECT 71.520 88.920 71.840 88.980 ;
        RECT 71.995 88.935 72.285 88.980 ;
        RECT 79.340 88.920 79.660 89.180 ;
        RECT 80.720 89.120 81.040 89.180 ;
        RECT 82.115 89.120 82.405 89.165 ;
        RECT 80.720 88.980 82.405 89.120 ;
        RECT 80.720 88.920 81.040 88.980 ;
        RECT 82.115 88.935 82.405 88.980 ;
        RECT 83.920 89.120 84.210 89.165 ;
        RECT 83.920 88.980 86.370 89.120 ;
        RECT 83.920 88.935 84.210 88.980 ;
        RECT 70.230 88.780 70.370 88.920 ;
        RECT 72.440 88.780 72.760 88.840 ;
        RECT 54.130 88.640 72.760 88.780 ;
        RECT 36.115 88.300 36.790 88.440 ;
        RECT 37.035 88.440 37.325 88.485 ;
        RECT 37.940 88.440 38.260 88.500 ;
        RECT 39.870 88.485 40.010 88.640 ;
        RECT 42.540 88.580 42.860 88.640 ;
        RECT 46.680 88.595 47.030 88.640 ;
        RECT 46.680 88.580 47.000 88.595 ;
        RECT 72.440 88.580 72.760 88.640 ;
        RECT 75.200 88.780 75.520 88.840 ;
        RECT 75.200 88.640 77.730 88.780 ;
        RECT 75.200 88.580 75.520 88.640 ;
        RECT 38.875 88.440 39.165 88.485 ;
        RECT 37.035 88.300 37.710 88.440 ;
        RECT 36.115 88.255 36.405 88.300 ;
        RECT 37.035 88.255 37.325 88.300 ;
        RECT 25.035 88.100 25.325 88.145 ;
        RECT 26.225 88.100 26.515 88.145 ;
        RECT 28.745 88.100 29.035 88.145 ;
        RECT 25.035 87.960 29.035 88.100 ;
        RECT 35.730 88.100 35.870 88.255 ;
        RECT 37.570 88.145 37.710 88.300 ;
        RECT 37.940 88.300 39.165 88.440 ;
        RECT 37.940 88.240 38.260 88.300 ;
        RECT 38.875 88.255 39.165 88.300 ;
        RECT 39.335 88.255 39.625 88.485 ;
        RECT 39.795 88.255 40.085 88.485 ;
        RECT 40.715 88.440 41.005 88.485 ;
        RECT 43.000 88.440 43.320 88.500 ;
        RECT 40.715 88.300 43.320 88.440 ;
        RECT 40.715 88.255 41.005 88.300 ;
        RECT 35.730 87.960 36.330 88.100 ;
        RECT 25.035 87.915 25.325 87.960 ;
        RECT 26.225 87.915 26.515 87.960 ;
        RECT 28.745 87.915 29.035 87.960 ;
        RECT 24.640 87.760 24.930 87.805 ;
        RECT 26.740 87.760 27.030 87.805 ;
        RECT 28.310 87.760 28.600 87.805 ;
        RECT 24.640 87.620 28.600 87.760 ;
        RECT 24.640 87.575 24.930 87.620 ;
        RECT 26.740 87.575 27.030 87.620 ;
        RECT 28.310 87.575 28.600 87.620 ;
        RECT 30.670 87.620 32.650 87.760 ;
        RECT 30.670 87.480 30.810 87.620 ;
        RECT 30.580 87.220 30.900 87.480 ;
        RECT 31.040 87.220 31.360 87.480 ;
        RECT 32.510 87.465 32.650 87.620 ;
        RECT 32.435 87.235 32.725 87.465 ;
        RECT 36.190 87.420 36.330 87.960 ;
        RECT 37.495 87.915 37.785 88.145 ;
        RECT 38.400 87.900 38.720 88.160 ;
        RECT 39.410 88.100 39.550 88.255 ;
        RECT 43.000 88.240 43.320 88.300 ;
        RECT 48.075 88.440 48.365 88.485 ;
        RECT 50.360 88.440 50.680 88.500 ;
        RECT 48.075 88.300 50.680 88.440 ;
        RECT 48.075 88.255 48.365 88.300 ;
        RECT 50.360 88.240 50.680 88.300 ;
        RECT 50.820 88.240 51.140 88.500 ;
        RECT 51.755 88.440 52.045 88.485 ;
        RECT 53.120 88.440 53.440 88.500 ;
        RECT 51.755 88.300 53.440 88.440 ;
        RECT 51.755 88.255 52.045 88.300 ;
        RECT 53.120 88.240 53.440 88.300 ;
        RECT 54.500 88.440 54.820 88.500 ;
        RECT 54.975 88.440 55.265 88.485 ;
        RECT 54.500 88.300 55.265 88.440 ;
        RECT 54.500 88.240 54.820 88.300 ;
        RECT 54.975 88.255 55.265 88.300 ;
        RECT 56.355 88.255 56.645 88.485 ;
        RECT 58.195 88.440 58.485 88.485 ;
        RECT 62.320 88.440 62.640 88.500 ;
        RECT 58.195 88.300 62.640 88.440 ;
        RECT 58.195 88.255 58.485 88.300 ;
        RECT 43.485 88.100 43.775 88.145 ;
        RECT 46.005 88.100 46.295 88.145 ;
        RECT 47.195 88.100 47.485 88.145 ;
        RECT 39.410 87.960 41.390 88.100 ;
        RECT 37.035 87.760 37.325 87.805 ;
        RECT 38.490 87.760 38.630 87.900 ;
        RECT 37.035 87.620 38.630 87.760 ;
        RECT 37.035 87.575 37.325 87.620 ;
        RECT 39.410 87.420 39.550 87.960 ;
        RECT 41.250 87.820 41.390 87.960 ;
        RECT 43.485 87.960 47.485 88.100 ;
        RECT 43.485 87.915 43.775 87.960 ;
        RECT 46.005 87.915 46.295 87.960 ;
        RECT 47.195 87.915 47.485 87.960 ;
        RECT 51.295 88.100 51.585 88.145 ;
        RECT 52.215 88.100 52.505 88.145 ;
        RECT 55.435 88.100 55.725 88.145 ;
        RECT 51.295 87.960 55.725 88.100 ;
        RECT 51.295 87.915 51.585 87.960 ;
        RECT 52.215 87.915 52.505 87.960 ;
        RECT 55.435 87.915 55.725 87.960 ;
        RECT 41.160 87.560 41.480 87.820 ;
        RECT 43.920 87.760 44.210 87.805 ;
        RECT 45.490 87.760 45.780 87.805 ;
        RECT 47.590 87.760 47.880 87.805 ;
        RECT 53.595 87.760 53.885 87.805 ;
        RECT 56.430 87.760 56.570 88.255 ;
        RECT 62.320 88.240 62.640 88.300 ;
        RECT 62.780 88.440 63.100 88.500 ;
        RECT 65.140 88.440 65.430 88.485 ;
        RECT 62.780 88.300 65.430 88.440 ;
        RECT 62.780 88.240 63.100 88.300 ;
        RECT 65.140 88.255 65.430 88.300 ;
        RECT 66.000 88.440 66.320 88.500 ;
        RECT 66.475 88.440 66.765 88.485 ;
        RECT 69.695 88.440 69.985 88.485 ;
        RECT 66.000 88.300 66.765 88.440 ;
        RECT 66.000 88.240 66.320 88.300 ;
        RECT 66.475 88.255 66.765 88.300 ;
        RECT 68.390 88.300 69.985 88.440 ;
        RECT 68.390 88.160 68.530 88.300 ;
        RECT 69.695 88.255 69.985 88.300 ;
        RECT 70.155 88.440 70.445 88.485 ;
        RECT 70.600 88.440 70.920 88.500 ;
        RECT 70.155 88.300 70.920 88.440 ;
        RECT 70.155 88.255 70.445 88.300 ;
        RECT 70.600 88.240 70.920 88.300 ;
        RECT 71.060 88.240 71.380 88.500 ;
        RECT 77.590 88.485 77.730 88.640 ;
        RECT 76.595 88.255 76.885 88.485 ;
        RECT 77.515 88.440 77.805 88.485 ;
        RECT 78.880 88.440 79.200 88.500 ;
        RECT 79.430 88.485 79.570 88.920 ;
        RECT 84.400 88.580 84.720 88.840 ;
        RECT 77.515 88.300 79.200 88.440 ;
        RECT 77.515 88.255 77.805 88.300 ;
        RECT 61.885 88.100 62.175 88.145 ;
        RECT 64.405 88.100 64.695 88.145 ;
        RECT 65.595 88.100 65.885 88.145 ;
        RECT 61.885 87.960 65.885 88.100 ;
        RECT 61.885 87.915 62.175 87.960 ;
        RECT 64.405 87.915 64.695 87.960 ;
        RECT 65.595 87.915 65.885 87.960 ;
        RECT 68.300 87.900 68.620 88.160 ;
        RECT 43.920 87.620 47.880 87.760 ;
        RECT 43.920 87.575 44.210 87.620 ;
        RECT 45.490 87.575 45.780 87.620 ;
        RECT 47.590 87.575 47.880 87.620 ;
        RECT 53.210 87.620 56.570 87.760 ;
        RECT 59.115 87.760 59.405 87.805 ;
        RECT 62.320 87.760 62.610 87.805 ;
        RECT 63.890 87.760 64.180 87.805 ;
        RECT 65.990 87.760 66.280 87.805 ;
        RECT 59.115 87.620 62.090 87.760 ;
        RECT 53.210 87.480 53.350 87.620 ;
        RECT 53.595 87.575 53.885 87.620 ;
        RECT 59.115 87.575 59.405 87.620 ;
        RECT 36.190 87.280 39.550 87.420 ;
        RECT 53.120 87.220 53.440 87.480 ;
        RECT 59.560 87.220 59.880 87.480 ;
        RECT 61.950 87.420 62.090 87.620 ;
        RECT 62.320 87.620 66.280 87.760 ;
        RECT 62.320 87.575 62.610 87.620 ;
        RECT 63.890 87.575 64.180 87.620 ;
        RECT 65.990 87.575 66.280 87.620 ;
        RECT 62.780 87.420 63.100 87.480 ;
        RECT 61.950 87.280 63.100 87.420 ;
        RECT 71.150 87.420 71.290 88.240 ;
        RECT 76.120 88.100 76.440 88.160 ;
        RECT 76.670 88.100 76.810 88.255 ;
        RECT 78.880 88.240 79.200 88.300 ;
        RECT 79.355 88.255 79.645 88.485 ;
        RECT 79.815 88.255 80.105 88.485 ;
        RECT 82.560 88.440 82.880 88.500 ;
        RECT 83.035 88.440 83.325 88.485 ;
        RECT 82.560 88.300 83.325 88.440 ;
        RECT 76.120 87.960 76.810 88.100 ;
        RECT 77.055 88.100 77.345 88.145 ;
        RECT 77.975 88.100 78.265 88.145 ;
        RECT 79.890 88.100 80.030 88.255 ;
        RECT 82.560 88.240 82.880 88.300 ;
        RECT 83.035 88.255 83.325 88.300 ;
        RECT 83.480 88.240 83.800 88.500 ;
        RECT 86.230 88.485 86.370 88.980 ;
        RECT 92.220 88.920 92.540 89.180 ;
        RECT 95.455 89.120 95.745 89.165 ;
        RECT 96.820 89.120 97.140 89.180 ;
        RECT 95.455 88.980 97.140 89.120 ;
        RECT 95.455 88.935 95.745 88.980 ;
        RECT 96.820 88.920 97.140 88.980 ;
        RECT 133.620 88.920 133.940 89.180 ;
        RECT 94.150 88.640 95.210 88.780 ;
        RECT 84.875 88.430 85.165 88.485 ;
        RECT 84.030 88.290 85.165 88.430 ;
        RECT 84.030 88.100 84.170 88.290 ;
        RECT 84.875 88.255 85.165 88.290 ;
        RECT 86.155 88.255 86.445 88.485 ;
        RECT 93.155 88.440 93.445 88.485 ;
        RECT 94.150 88.440 94.290 88.640 ;
        RECT 92.770 88.300 94.290 88.440 ;
        RECT 77.055 87.960 80.030 88.100 ;
        RECT 82.190 87.960 84.170 88.100 ;
        RECT 85.755 88.100 86.045 88.145 ;
        RECT 86.945 88.100 87.235 88.145 ;
        RECT 89.465 88.100 89.755 88.145 ;
        RECT 92.770 88.100 92.910 88.300 ;
        RECT 93.155 88.255 93.445 88.300 ;
        RECT 94.535 88.255 94.825 88.485 ;
        RECT 95.070 88.440 95.210 88.640 ;
        RECT 104.180 88.580 104.500 88.840 ;
        RECT 119.360 88.780 119.680 88.840 ;
        RECT 122.120 88.780 122.440 88.840 ;
        RECT 133.710 88.780 133.850 88.920 ;
        RECT 119.360 88.640 123.730 88.780 ;
        RECT 119.360 88.580 119.680 88.640 ;
        RECT 122.120 88.580 122.440 88.640 ;
        RECT 96.820 88.440 97.140 88.500 ;
        RECT 95.070 88.300 97.140 88.440 ;
        RECT 94.610 88.100 94.750 88.255 ;
        RECT 96.820 88.240 97.140 88.300 ;
        RECT 102.800 88.240 103.120 88.500 ;
        RECT 103.735 88.440 104.025 88.485 ;
        RECT 104.270 88.440 104.410 88.580 ;
        RECT 103.735 88.300 104.410 88.440 ;
        RECT 110.160 88.440 110.480 88.500 ;
        RECT 114.315 88.440 114.605 88.485 ;
        RECT 110.160 88.300 114.605 88.440 ;
        RECT 103.735 88.255 104.025 88.300 ;
        RECT 110.160 88.240 110.480 88.300 ;
        RECT 114.315 88.255 114.605 88.300 ;
        RECT 115.220 88.240 115.540 88.500 ;
        RECT 116.155 88.440 116.445 88.485 ;
        RECT 116.615 88.440 116.905 88.485 ;
        RECT 116.155 88.300 116.905 88.440 ;
        RECT 116.155 88.255 116.445 88.300 ;
        RECT 116.615 88.255 116.905 88.300 ;
        RECT 117.520 88.440 117.840 88.500 ;
        RECT 118.900 88.440 119.220 88.500 ;
        RECT 123.590 88.485 123.730 88.640 ;
        RECT 126.810 88.640 128.790 88.780 ;
        RECT 133.710 88.640 139.830 88.780 ;
        RECT 126.810 88.485 126.950 88.640 ;
        RECT 123.055 88.440 123.345 88.485 ;
        RECT 117.520 88.300 123.345 88.440 ;
        RECT 117.520 88.240 117.840 88.300 ;
        RECT 118.900 88.240 119.220 88.300 ;
        RECT 123.055 88.255 123.345 88.300 ;
        RECT 123.515 88.255 123.805 88.485 ;
        RECT 124.435 88.255 124.725 88.485 ;
        RECT 125.355 88.440 125.645 88.485 ;
        RECT 126.275 88.440 126.565 88.485 ;
        RECT 125.355 88.300 126.565 88.440 ;
        RECT 125.355 88.255 125.645 88.300 ;
        RECT 126.275 88.255 126.565 88.300 ;
        RECT 126.735 88.255 127.025 88.485 ;
        RECT 127.195 88.255 127.485 88.485 ;
        RECT 85.755 87.960 89.755 88.100 ;
        RECT 76.120 87.900 76.440 87.960 ;
        RECT 77.055 87.915 77.345 87.960 ;
        RECT 77.975 87.915 78.265 87.960 ;
        RECT 82.190 87.820 82.330 87.960 ;
        RECT 85.755 87.915 86.045 87.960 ;
        RECT 86.945 87.915 87.235 87.960 ;
        RECT 89.465 87.915 89.755 87.960 ;
        RECT 91.390 87.960 92.910 88.100 ;
        RECT 93.230 87.960 94.750 88.100 ;
        RECT 71.520 87.760 71.840 87.820 ;
        RECT 82.100 87.760 82.420 87.820 ;
        RECT 71.520 87.620 82.420 87.760 ;
        RECT 71.520 87.560 71.840 87.620 ;
        RECT 82.100 87.560 82.420 87.620 ;
        RECT 83.480 87.560 83.800 87.820 ;
        RECT 85.360 87.760 85.650 87.805 ;
        RECT 87.460 87.760 87.750 87.805 ;
        RECT 89.030 87.760 89.320 87.805 ;
        RECT 85.360 87.620 89.320 87.760 ;
        RECT 85.360 87.575 85.650 87.620 ;
        RECT 87.460 87.575 87.750 87.620 ;
        RECT 89.030 87.575 89.320 87.620 ;
        RECT 78.420 87.420 78.740 87.480 ;
        RECT 71.150 87.280 78.740 87.420 ;
        RECT 62.780 87.220 63.100 87.280 ;
        RECT 78.420 87.220 78.740 87.280 ;
        RECT 78.895 87.420 79.185 87.465 ;
        RECT 80.260 87.420 80.580 87.480 ;
        RECT 78.895 87.280 80.580 87.420 ;
        RECT 83.570 87.420 83.710 87.560 ;
        RECT 91.390 87.420 91.530 87.960 ;
        RECT 93.230 87.480 93.370 87.960 ;
        RECT 95.440 87.900 95.760 88.160 ;
        RECT 109.700 87.900 110.020 88.160 ;
        RECT 124.510 88.100 124.650 88.255 ;
        RECT 125.800 88.100 126.120 88.160 ;
        RECT 127.270 88.100 127.410 88.255 ;
        RECT 128.100 88.240 128.420 88.500 ;
        RECT 128.650 88.440 128.790 88.640 ;
        RECT 139.690 88.485 139.830 88.640 ;
        RECT 147.510 88.640 149.490 88.780 ;
        RECT 129.495 88.440 129.785 88.485 ;
        RECT 128.650 88.300 129.785 88.440 ;
        RECT 129.495 88.255 129.785 88.300 ;
        RECT 139.615 88.255 139.905 88.485 ;
        RECT 140.535 88.255 140.825 88.485 ;
        RECT 141.455 88.440 141.745 88.485 ;
        RECT 141.915 88.440 142.205 88.485 ;
        RECT 141.455 88.300 142.205 88.440 ;
        RECT 141.455 88.255 141.745 88.300 ;
        RECT 141.915 88.255 142.205 88.300 ;
        RECT 145.120 88.440 145.440 88.500 ;
        RECT 147.510 88.485 147.650 88.640 ;
        RECT 147.435 88.440 147.725 88.485 ;
        RECT 148.355 88.440 148.645 88.485 ;
        RECT 148.815 88.440 149.105 88.485 ;
        RECT 145.120 88.300 147.725 88.440 ;
        RECT 127.640 88.100 127.960 88.160 ;
        RECT 124.510 87.960 125.570 88.100 ;
        RECT 125.430 87.820 125.570 87.960 ;
        RECT 125.800 87.960 127.960 88.100 ;
        RECT 125.800 87.900 126.120 87.960 ;
        RECT 127.640 87.900 127.960 87.960 ;
        RECT 128.580 88.100 128.870 88.145 ;
        RECT 130.920 88.100 131.210 88.145 ;
        RECT 128.580 87.960 131.210 88.100 ;
        RECT 140.610 88.100 140.750 88.255 ;
        RECT 145.120 88.240 145.440 88.300 ;
        RECT 147.435 88.255 147.725 88.300 ;
        RECT 147.970 88.300 149.105 88.440 ;
        RECT 149.350 88.440 149.490 88.640 ;
        RECT 149.735 88.440 150.025 88.485 ;
        RECT 149.350 88.300 150.025 88.440 ;
        RECT 144.660 88.100 144.980 88.160 ;
        RECT 140.610 87.960 144.980 88.100 ;
        RECT 128.580 87.915 128.870 87.960 ;
        RECT 130.920 87.915 131.210 87.960 ;
        RECT 144.660 87.900 144.980 87.960 ;
        RECT 93.615 87.575 93.905 87.805 ;
        RECT 94.075 87.760 94.365 87.805 ;
        RECT 95.900 87.760 96.220 87.820 ;
        RECT 94.075 87.620 96.220 87.760 ;
        RECT 94.075 87.575 94.365 87.620 ;
        RECT 83.570 87.280 91.530 87.420 ;
        RECT 78.895 87.235 79.185 87.280 ;
        RECT 80.260 87.220 80.580 87.280 ;
        RECT 91.760 87.220 92.080 87.480 ;
        RECT 93.140 87.220 93.460 87.480 ;
        RECT 93.690 87.420 93.830 87.575 ;
        RECT 95.900 87.560 96.220 87.620 ;
        RECT 111.540 87.560 111.860 87.820 ;
        RECT 125.340 87.560 125.660 87.820 ;
        RECT 129.040 87.760 129.330 87.805 ;
        RECT 130.415 87.760 130.705 87.805 ;
        RECT 129.040 87.620 130.705 87.760 ;
        RECT 129.040 87.575 129.330 87.620 ;
        RECT 130.415 87.575 130.705 87.620 ;
        RECT 133.175 87.760 133.465 87.805 ;
        RECT 135.460 87.760 135.780 87.820 ;
        RECT 133.175 87.620 135.780 87.760 ;
        RECT 133.175 87.575 133.465 87.620 ;
        RECT 135.460 87.560 135.780 87.620 ;
        RECT 147.970 87.480 148.110 88.300 ;
        RECT 148.355 88.255 148.645 88.300 ;
        RECT 148.815 88.255 149.105 88.300 ;
        RECT 149.735 88.255 150.025 88.300 ;
        RECT 96.360 87.420 96.680 87.480 ;
        RECT 93.690 87.280 96.680 87.420 ;
        RECT 96.360 87.220 96.680 87.280 ;
        RECT 103.260 87.220 103.580 87.480 ;
        RECT 112.000 87.220 112.320 87.480 ;
        RECT 117.520 87.220 117.840 87.480 ;
        RECT 119.820 87.220 120.140 87.480 ;
        RECT 142.360 87.420 142.680 87.480 ;
        RECT 142.835 87.420 143.125 87.465 ;
        RECT 142.360 87.280 143.125 87.420 ;
        RECT 142.360 87.220 142.680 87.280 ;
        RECT 142.835 87.235 143.125 87.280 ;
        RECT 147.880 87.220 148.200 87.480 ;
        RECT 148.340 87.220 148.660 87.480 ;
        RECT 148.800 87.420 149.120 87.480 ;
        RECT 149.275 87.420 149.565 87.465 ;
        RECT 148.800 87.280 149.565 87.420 ;
        RECT 148.800 87.220 149.120 87.280 ;
        RECT 149.275 87.235 149.565 87.280 ;
        RECT 22.690 86.600 157.010 87.080 ;
        RECT 25.520 86.400 25.840 86.460 ;
        RECT 26.915 86.400 27.205 86.445 ;
        RECT 25.520 86.260 27.205 86.400 ;
        RECT 25.520 86.200 25.840 86.260 ;
        RECT 26.915 86.215 27.205 86.260 ;
        RECT 28.755 86.400 29.045 86.445 ;
        RECT 29.200 86.400 29.520 86.460 ;
        RECT 28.755 86.260 29.520 86.400 ;
        RECT 28.755 86.215 29.045 86.260 ;
        RECT 29.200 86.200 29.520 86.260 ;
        RECT 30.580 86.200 30.900 86.460 ;
        RECT 31.040 86.200 31.360 86.460 ;
        RECT 31.515 86.400 31.805 86.445 ;
        RECT 32.420 86.400 32.740 86.460 ;
        RECT 31.515 86.260 32.740 86.400 ;
        RECT 31.515 86.215 31.805 86.260 ;
        RECT 32.420 86.200 32.740 86.260 ;
        RECT 37.940 86.200 38.260 86.460 ;
        RECT 41.160 86.200 41.480 86.460 ;
        RECT 50.820 86.200 51.140 86.460 ;
        RECT 53.120 86.200 53.440 86.460 ;
        RECT 54.500 86.400 54.820 86.460 ;
        RECT 55.895 86.400 56.185 86.445 ;
        RECT 54.500 86.260 56.185 86.400 ;
        RECT 54.500 86.200 54.820 86.260 ;
        RECT 55.895 86.215 56.185 86.260 ;
        RECT 63.240 86.400 63.560 86.460 ;
        RECT 64.175 86.400 64.465 86.445 ;
        RECT 63.240 86.260 64.465 86.400 ;
        RECT 63.240 86.200 63.560 86.260 ;
        RECT 64.175 86.215 64.465 86.260 ;
        RECT 66.000 86.400 66.320 86.460 ;
        RECT 71.520 86.400 71.840 86.460 ;
        RECT 66.000 86.260 71.840 86.400 ;
        RECT 66.000 86.200 66.320 86.260 ;
        RECT 71.520 86.200 71.840 86.260 ;
        RECT 78.420 86.200 78.740 86.460 ;
        RECT 80.260 86.400 80.580 86.460 ;
        RECT 81.655 86.400 81.945 86.445 ;
        RECT 80.260 86.260 81.945 86.400 ;
        RECT 80.260 86.200 80.580 86.260 ;
        RECT 81.655 86.215 81.945 86.260 ;
        RECT 84.400 86.400 84.720 86.460 ;
        RECT 88.095 86.400 88.385 86.445 ;
        RECT 84.400 86.260 88.385 86.400 ;
        RECT 84.400 86.200 84.720 86.260 ;
        RECT 88.095 86.215 88.385 86.260 ;
        RECT 90.380 86.400 90.700 86.460 ;
        RECT 90.855 86.400 91.145 86.445 ;
        RECT 90.380 86.260 91.145 86.400 ;
        RECT 90.380 86.200 90.700 86.260 ;
        RECT 90.855 86.215 91.145 86.260 ;
        RECT 91.760 86.200 92.080 86.460 ;
        RECT 93.140 86.200 93.460 86.460 ;
        RECT 94.980 86.200 95.300 86.460 ;
        RECT 96.820 86.400 97.140 86.460 ;
        RECT 100.055 86.400 100.345 86.445 ;
        RECT 96.820 86.260 100.345 86.400 ;
        RECT 96.820 86.200 97.140 86.260 ;
        RECT 100.055 86.215 100.345 86.260 ;
        RECT 105.100 86.200 105.420 86.460 ;
        RECT 112.000 86.200 112.320 86.460 ;
        RECT 115.220 86.200 115.540 86.460 ;
        RECT 119.820 86.400 120.140 86.460 ;
        RECT 124.880 86.400 125.200 86.460 ;
        RECT 126.735 86.400 127.025 86.445 ;
        RECT 119.820 86.260 121.890 86.400 ;
        RECT 119.820 86.200 120.140 86.260 ;
        RECT 28.740 85.720 29.060 85.780 ;
        RECT 29.215 85.720 29.505 85.765 ;
        RECT 28.740 85.580 29.505 85.720 ;
        RECT 28.740 85.520 29.060 85.580 ;
        RECT 29.215 85.535 29.505 85.580 ;
        RECT 27.835 85.380 28.125 85.425 ;
        RECT 28.280 85.380 28.600 85.440 ;
        RECT 31.130 85.425 31.270 86.200 ;
        RECT 27.835 85.240 28.600 85.380 ;
        RECT 27.835 85.195 28.125 85.240 ;
        RECT 28.280 85.180 28.600 85.240 ;
        RECT 29.675 85.195 29.965 85.425 ;
        RECT 30.595 85.380 30.885 85.425 ;
        RECT 31.055 85.380 31.345 85.425 ;
        RECT 30.595 85.240 31.345 85.380 ;
        RECT 30.595 85.195 30.885 85.240 ;
        RECT 31.055 85.195 31.345 85.240 ;
        RECT 31.975 85.195 32.265 85.425 ;
        RECT 29.750 85.040 29.890 85.195 ;
        RECT 32.050 85.040 32.190 85.195 ;
        RECT 33.340 85.180 33.660 85.440 ;
        RECT 37.480 85.180 37.800 85.440 ;
        RECT 38.030 85.425 38.170 86.200 ;
        RECT 38.415 85.720 38.705 85.765 ;
        RECT 41.250 85.720 41.390 86.200 ;
        RECT 38.415 85.580 41.390 85.720 ;
        RECT 50.910 85.720 51.050 86.200 ;
        RECT 60.480 86.060 60.800 86.120 ;
        RECT 57.350 85.920 60.800 86.060 ;
        RECT 50.910 85.580 53.810 85.720 ;
        RECT 38.415 85.535 38.705 85.580 ;
        RECT 53.670 85.440 53.810 85.580 ;
        RECT 37.955 85.195 38.245 85.425 ;
        RECT 43.920 85.180 44.240 85.440 ;
        RECT 48.980 85.180 49.300 85.440 ;
        RECT 52.660 85.180 52.980 85.440 ;
        RECT 53.580 85.180 53.900 85.440 ;
        RECT 56.815 85.380 57.105 85.425 ;
        RECT 57.350 85.380 57.490 85.920 ;
        RECT 60.480 85.860 60.800 85.920 ;
        RECT 61.400 86.060 61.720 86.120 ;
        RECT 91.850 86.060 91.990 86.200 ;
        RECT 61.400 85.920 82.330 86.060 ;
        RECT 61.400 85.860 61.720 85.920 ;
        RECT 57.735 85.720 58.025 85.765 ;
        RECT 58.640 85.720 58.960 85.780 ;
        RECT 57.735 85.580 58.960 85.720 ;
        RECT 57.735 85.535 58.025 85.580 ;
        RECT 58.640 85.520 58.960 85.580 ;
        RECT 60.955 85.720 61.245 85.765 ;
        RECT 62.335 85.720 62.625 85.765 ;
        RECT 60.955 85.580 62.625 85.720 ;
        RECT 60.955 85.535 61.245 85.580 ;
        RECT 62.335 85.535 62.625 85.580 ;
        RECT 76.210 85.580 80.950 85.720 ;
        RECT 76.210 85.440 76.350 85.580 ;
        RECT 56.815 85.240 57.490 85.380 ;
        RECT 58.195 85.380 58.485 85.425 ;
        RECT 62.795 85.380 63.085 85.425 ;
        RECT 58.195 85.240 63.085 85.380 ;
        RECT 56.815 85.195 57.105 85.240 ;
        RECT 58.195 85.195 58.485 85.240 ;
        RECT 29.750 84.900 32.190 85.040 ;
        RECT 31.130 84.760 31.270 84.900 ;
        RECT 31.040 84.500 31.360 84.760 ;
        RECT 37.570 84.700 37.710 85.180 ;
        RECT 61.030 84.760 61.170 85.240 ;
        RECT 62.795 85.195 63.085 85.240 ;
        RECT 76.120 85.180 76.440 85.440 ;
        RECT 77.500 85.180 77.820 85.440 ;
        RECT 77.975 85.195 78.265 85.425 ;
        RECT 78.050 85.040 78.190 85.195 ;
        RECT 78.880 85.180 79.200 85.440 ;
        RECT 79.340 85.180 79.660 85.440 ;
        RECT 80.810 85.425 80.950 85.580 ;
        RECT 80.735 85.195 81.025 85.425 ;
        RECT 81.655 85.195 81.945 85.425 ;
        RECT 77.590 84.900 78.190 85.040 ;
        RECT 78.970 85.040 79.110 85.180 ;
        RECT 81.730 85.040 81.870 85.195 ;
        RECT 78.970 84.900 81.870 85.040 ;
        RECT 77.590 84.760 77.730 84.900 ;
        RECT 39.795 84.700 40.085 84.745 ;
        RECT 37.570 84.560 40.085 84.700 ;
        RECT 39.795 84.515 40.085 84.560 ;
        RECT 60.940 84.500 61.260 84.760 ;
        RECT 71.075 84.700 71.365 84.745 ;
        RECT 71.520 84.700 71.840 84.760 ;
        RECT 71.075 84.560 71.840 84.700 ;
        RECT 71.075 84.515 71.365 84.560 ;
        RECT 71.520 84.500 71.840 84.560 ;
        RECT 77.500 84.500 77.820 84.760 ;
        RECT 77.960 84.700 78.280 84.760 ;
        RECT 80.275 84.700 80.565 84.745 ;
        RECT 77.960 84.560 80.565 84.700 ;
        RECT 82.190 84.700 82.330 85.920 ;
        RECT 90.470 85.920 91.990 86.060 ;
        RECT 82.560 85.520 82.880 85.780 ;
        RECT 83.020 85.720 83.340 85.780 ;
        RECT 87.635 85.720 87.925 85.765 ;
        RECT 83.020 85.580 87.925 85.720 ;
        RECT 83.020 85.520 83.340 85.580 ;
        RECT 87.635 85.535 87.925 85.580 ;
        RECT 82.650 85.380 82.790 85.520 ;
        RECT 88.540 85.380 88.860 85.440 ;
        RECT 90.470 85.425 90.610 85.920 ;
        RECT 95.070 85.720 95.210 86.200 ;
        RECT 95.900 86.060 96.220 86.120 ;
        RECT 103.260 86.060 103.580 86.120 ;
        RECT 106.495 86.060 106.785 86.105 ;
        RECT 95.900 85.920 97.510 86.060 ;
        RECT 95.900 85.860 96.220 85.920 ;
        RECT 91.850 85.580 95.670 85.720 ;
        RECT 91.850 85.425 91.990 85.580 ;
        RECT 82.650 85.240 88.860 85.380 ;
        RECT 88.540 85.180 88.860 85.240 ;
        RECT 89.015 85.195 89.305 85.425 ;
        RECT 90.395 85.195 90.685 85.425 ;
        RECT 91.315 85.195 91.605 85.425 ;
        RECT 91.775 85.195 92.065 85.425 ;
        RECT 83.480 85.040 83.800 85.100 ;
        RECT 89.090 85.040 89.230 85.195 ;
        RECT 83.480 84.900 89.230 85.040 ;
        RECT 91.390 85.040 91.530 85.195 ;
        RECT 94.980 85.180 95.300 85.440 ;
        RECT 95.530 85.425 95.670 85.580 ;
        RECT 97.370 85.425 97.510 85.920 ;
        RECT 101.050 85.920 106.785 86.060 ;
        RECT 101.050 85.425 101.190 85.920 ;
        RECT 103.260 85.860 103.580 85.920 ;
        RECT 106.495 85.875 106.785 85.920 ;
        RECT 104.195 85.720 104.485 85.765 ;
        RECT 106.035 85.720 106.325 85.765 ;
        RECT 104.195 85.580 106.325 85.720 ;
        RECT 104.195 85.535 104.485 85.580 ;
        RECT 106.035 85.535 106.325 85.580 ;
        RECT 111.095 85.720 111.385 85.765 ;
        RECT 112.090 85.720 112.230 86.200 ;
        RECT 112.475 86.060 112.765 86.105 ;
        RECT 115.310 86.060 115.450 86.200 ;
        RECT 112.475 85.920 115.450 86.060 ;
        RECT 117.060 86.060 117.350 86.105 ;
        RECT 118.630 86.060 118.920 86.105 ;
        RECT 120.730 86.060 121.020 86.105 ;
        RECT 117.060 85.920 121.020 86.060 ;
        RECT 112.475 85.875 112.765 85.920 ;
        RECT 117.060 85.875 117.350 85.920 ;
        RECT 118.630 85.875 118.920 85.920 ;
        RECT 120.730 85.875 121.020 85.920 ;
        RECT 121.750 85.765 121.890 86.260 ;
        RECT 124.880 86.260 127.025 86.400 ;
        RECT 124.880 86.200 125.200 86.260 ;
        RECT 126.735 86.215 127.025 86.260 ;
        RECT 132.240 86.200 132.560 86.460 ;
        RECT 137.760 86.200 138.080 86.460 ;
        RECT 144.660 86.400 144.980 86.460 ;
        RECT 144.660 86.260 145.810 86.400 ;
        RECT 144.660 86.200 144.980 86.260 ;
        RECT 122.600 86.060 122.890 86.105 ;
        RECT 123.975 86.060 124.265 86.105 ;
        RECT 122.600 85.920 124.265 86.060 ;
        RECT 122.600 85.875 122.890 85.920 ;
        RECT 123.975 85.875 124.265 85.920 ;
        RECT 128.120 86.060 128.410 86.105 ;
        RECT 129.495 86.060 129.785 86.105 ;
        RECT 128.120 85.920 129.785 86.060 ;
        RECT 128.120 85.875 128.410 85.920 ;
        RECT 129.495 85.875 129.785 85.920 ;
        RECT 133.640 86.060 133.930 86.105 ;
        RECT 135.015 86.060 135.305 86.105 ;
        RECT 133.640 85.920 135.305 86.060 ;
        RECT 133.640 85.875 133.930 85.920 ;
        RECT 135.015 85.875 135.305 85.920 ;
        RECT 141.480 86.060 141.770 86.105 ;
        RECT 143.580 86.060 143.870 86.105 ;
        RECT 145.150 86.060 145.440 86.105 ;
        RECT 141.480 85.920 145.440 86.060 ;
        RECT 145.670 86.060 145.810 86.260 ;
        RECT 147.880 86.200 148.200 86.460 ;
        RECT 149.735 86.400 150.025 86.445 ;
        RECT 148.430 86.260 150.025 86.400 ;
        RECT 148.430 86.060 148.570 86.260 ;
        RECT 149.735 86.215 150.025 86.260 ;
        RECT 145.670 85.920 148.570 86.060 ;
        RECT 148.800 86.060 149.120 86.120 ;
        RECT 152.955 86.060 153.245 86.105 ;
        RECT 148.800 85.920 153.245 86.060 ;
        RECT 141.480 85.875 141.770 85.920 ;
        RECT 143.580 85.875 143.870 85.920 ;
        RECT 145.150 85.875 145.440 85.920 ;
        RECT 148.800 85.860 149.120 85.920 ;
        RECT 152.955 85.875 153.245 85.920 ;
        RECT 111.095 85.580 112.230 85.720 ;
        RECT 116.625 85.720 116.915 85.765 ;
        RECT 119.145 85.720 119.435 85.765 ;
        RECT 120.335 85.720 120.625 85.765 ;
        RECT 116.625 85.580 120.625 85.720 ;
        RECT 111.095 85.535 111.385 85.580 ;
        RECT 116.625 85.535 116.915 85.580 ;
        RECT 119.145 85.535 119.435 85.580 ;
        RECT 120.335 85.535 120.625 85.580 ;
        RECT 121.675 85.535 121.965 85.765 ;
        RECT 122.140 85.720 122.430 85.765 ;
        RECT 124.480 85.720 124.770 85.765 ;
        RECT 122.140 85.580 124.770 85.720 ;
        RECT 122.140 85.535 122.430 85.580 ;
        RECT 124.480 85.535 124.770 85.580 ;
        RECT 127.660 85.720 127.950 85.765 ;
        RECT 130.000 85.720 130.290 85.765 ;
        RECT 127.660 85.580 130.290 85.720 ;
        RECT 127.660 85.535 127.950 85.580 ;
        RECT 130.000 85.535 130.290 85.580 ;
        RECT 133.180 85.720 133.470 85.765 ;
        RECT 135.520 85.720 135.810 85.765 ;
        RECT 133.180 85.580 135.810 85.720 ;
        RECT 133.180 85.535 133.470 85.580 ;
        RECT 135.520 85.535 135.810 85.580 ;
        RECT 138.680 85.720 139.000 85.780 ;
        RECT 140.995 85.720 141.285 85.765 ;
        RECT 138.680 85.580 141.285 85.720 ;
        RECT 138.680 85.520 139.000 85.580 ;
        RECT 140.995 85.535 141.285 85.580 ;
        RECT 141.875 85.720 142.165 85.765 ;
        RECT 143.065 85.720 143.355 85.765 ;
        RECT 145.585 85.720 145.875 85.765 ;
        RECT 141.875 85.580 145.875 85.720 ;
        RECT 141.875 85.535 142.165 85.580 ;
        RECT 143.065 85.535 143.355 85.580 ;
        RECT 145.585 85.535 145.875 85.580 ;
        RECT 151.575 85.720 151.865 85.765 ;
        RECT 152.495 85.720 152.785 85.765 ;
        RECT 151.575 85.580 152.785 85.720 ;
        RECT 151.575 85.535 151.865 85.580 ;
        RECT 152.495 85.535 152.785 85.580 ;
        RECT 95.455 85.195 95.745 85.425 ;
        RECT 95.915 85.195 96.205 85.425 ;
        RECT 96.835 85.380 97.125 85.425 ;
        RECT 97.295 85.380 97.585 85.425 ;
        RECT 96.835 85.240 97.585 85.380 ;
        RECT 96.835 85.195 97.125 85.240 ;
        RECT 97.295 85.195 97.585 85.240 ;
        RECT 100.975 85.195 101.265 85.425 ;
        RECT 101.895 85.195 102.185 85.425 ;
        RECT 102.355 85.380 102.645 85.425 ;
        RECT 103.735 85.380 104.025 85.425 ;
        RECT 107.860 85.380 108.180 85.440 ;
        RECT 102.355 85.240 108.180 85.380 ;
        RECT 102.355 85.195 102.645 85.240 ;
        RECT 103.735 85.195 104.025 85.240 ;
        RECT 93.155 85.040 93.445 85.085 ;
        RECT 93.615 85.040 93.905 85.085 ;
        RECT 91.390 84.900 92.910 85.040 ;
        RECT 83.480 84.840 83.800 84.900 ;
        RECT 91.300 84.700 91.620 84.760 ;
        RECT 82.190 84.560 91.620 84.700 ;
        RECT 77.960 84.500 78.280 84.560 ;
        RECT 80.275 84.515 80.565 84.560 ;
        RECT 91.300 84.500 91.620 84.560 ;
        RECT 92.220 84.500 92.540 84.760 ;
        RECT 92.770 84.700 92.910 84.900 ;
        RECT 93.155 84.900 93.905 85.040 ;
        RECT 93.155 84.855 93.445 84.900 ;
        RECT 93.615 84.855 93.905 84.900 ;
        RECT 95.990 85.040 96.130 85.195 ;
        RECT 98.215 85.040 98.505 85.085 ;
        RECT 95.990 84.900 98.505 85.040 ;
        RECT 101.970 85.040 102.110 85.195 ;
        RECT 107.860 85.180 108.180 85.240 ;
        RECT 110.160 85.380 110.480 85.440 ;
        RECT 110.635 85.380 110.925 85.425 ;
        RECT 110.160 85.240 110.925 85.380 ;
        RECT 110.160 85.180 110.480 85.240 ;
        RECT 110.635 85.195 110.925 85.240 ;
        RECT 117.060 85.380 117.380 85.440 ;
        RECT 121.215 85.380 121.505 85.425 ;
        RECT 123.055 85.380 123.345 85.425 ;
        RECT 117.060 85.240 121.505 85.380 ;
        RECT 117.060 85.180 117.380 85.240 ;
        RECT 121.215 85.195 121.505 85.240 ;
        RECT 122.210 85.240 123.345 85.380 ;
        RECT 108.320 85.040 108.640 85.100 ;
        RECT 101.970 84.900 108.640 85.040 ;
        RECT 95.990 84.760 96.130 84.900 ;
        RECT 98.215 84.855 98.505 84.900 ;
        RECT 108.320 84.840 108.640 84.900 ;
        RECT 117.520 85.040 117.840 85.100 ;
        RECT 119.880 85.040 120.170 85.085 ;
        RECT 117.520 84.900 120.170 85.040 ;
        RECT 117.520 84.840 117.840 84.900 ;
        RECT 119.880 84.855 120.170 84.900 ;
        RECT 122.210 84.760 122.350 85.240 ;
        RECT 123.055 85.195 123.345 85.240 ;
        RECT 127.180 85.180 127.500 85.440 ;
        RECT 128.575 85.195 128.865 85.425 ;
        RECT 128.650 84.760 128.790 85.195 ;
        RECT 132.700 85.180 133.020 85.440 ;
        RECT 134.080 85.180 134.400 85.440 ;
        RECT 137.300 85.380 137.620 85.440 ;
        RECT 142.360 85.425 142.680 85.440 ;
        RECT 139.155 85.380 139.445 85.425 ;
        RECT 142.330 85.380 142.680 85.425 ;
        RECT 137.300 85.240 139.445 85.380 ;
        RECT 142.165 85.240 142.680 85.380 ;
        RECT 137.300 85.180 137.620 85.240 ;
        RECT 139.155 85.195 139.445 85.240 ;
        RECT 142.330 85.195 142.680 85.240 ;
        RECT 142.360 85.180 142.680 85.195 ;
        RECT 150.640 85.380 150.960 85.440 ;
        RECT 151.115 85.380 151.405 85.425 ;
        RECT 150.640 85.240 151.405 85.380 ;
        RECT 150.640 85.180 150.960 85.240 ;
        RECT 151.115 85.195 151.405 85.240 ;
        RECT 148.340 85.040 148.660 85.100 ;
        RECT 154.795 85.040 155.085 85.085 ;
        RECT 148.340 84.900 155.085 85.040 ;
        RECT 148.340 84.840 148.660 84.900 ;
        RECT 154.795 84.855 155.085 84.900 ;
        RECT 95.900 84.700 96.220 84.760 ;
        RECT 92.770 84.560 96.220 84.700 ;
        RECT 95.900 84.500 96.220 84.560 ;
        RECT 99.120 84.500 99.440 84.760 ;
        RECT 114.300 84.500 114.620 84.760 ;
        RECT 122.120 84.500 122.440 84.760 ;
        RECT 128.560 84.500 128.880 84.760 ;
        RECT 22.690 83.880 157.810 84.360 ;
        RECT 33.340 83.480 33.660 83.740 ;
        RECT 37.940 83.680 38.260 83.740 ;
        RECT 38.415 83.680 38.705 83.725 ;
        RECT 37.940 83.540 38.705 83.680 ;
        RECT 37.940 83.480 38.260 83.540 ;
        RECT 38.415 83.495 38.705 83.540 ;
        RECT 42.540 83.480 42.860 83.740 ;
        RECT 43.920 83.480 44.240 83.740 ;
        RECT 48.980 83.480 49.300 83.740 ;
        RECT 53.580 83.680 53.900 83.740 ;
        RECT 54.055 83.680 54.345 83.725 ;
        RECT 53.580 83.540 54.345 83.680 ;
        RECT 53.580 83.480 53.900 83.540 ;
        RECT 54.055 83.495 54.345 83.540 ;
        RECT 58.640 83.680 58.960 83.740 ;
        RECT 59.115 83.680 59.405 83.725 ;
        RECT 58.640 83.540 59.405 83.680 ;
        RECT 58.640 83.480 58.960 83.540 ;
        RECT 59.115 83.495 59.405 83.540 ;
        RECT 60.480 83.480 60.800 83.740 ;
        RECT 65.555 83.680 65.845 83.725 ;
        RECT 68.300 83.680 68.620 83.740 ;
        RECT 90.840 83.680 91.160 83.740 ;
        RECT 94.995 83.680 95.285 83.725 ;
        RECT 65.555 83.540 68.620 83.680 ;
        RECT 65.555 83.495 65.845 83.540 ;
        RECT 68.300 83.480 68.620 83.540 ;
        RECT 68.850 83.540 91.160 83.680 ;
        RECT 31.500 82.800 31.820 83.060 ;
        RECT 33.430 83.045 33.570 83.480 ;
        RECT 44.010 83.340 44.150 83.480 ;
        RECT 44.010 83.200 47.830 83.340 ;
        RECT 33.355 82.815 33.645 83.045 ;
        RECT 34.720 82.800 35.040 83.060 ;
        RECT 46.220 82.800 46.540 83.060 ;
        RECT 47.690 83.045 47.830 83.200 ;
        RECT 49.070 83.045 49.210 83.480 ;
        RECT 67.380 83.340 67.700 83.400 ;
        RECT 68.850 83.340 68.990 83.540 ;
        RECT 90.840 83.480 91.160 83.540 ;
        RECT 94.150 83.540 95.285 83.680 ;
        RECT 58.730 83.200 60.250 83.340 ;
        RECT 47.615 82.815 47.905 83.045 ;
        RECT 48.995 82.815 49.285 83.045 ;
        RECT 50.360 82.800 50.680 83.060 ;
        RECT 58.180 83.000 58.500 83.060 ;
        RECT 58.730 83.045 58.870 83.200 ;
        RECT 58.655 83.000 58.945 83.045 ;
        RECT 58.180 82.860 58.945 83.000 ;
        RECT 58.180 82.800 58.500 82.860 ;
        RECT 58.655 82.815 58.945 82.860 ;
        RECT 59.560 82.800 59.880 83.060 ;
        RECT 60.110 83.045 60.250 83.200 ;
        RECT 67.380 83.200 68.990 83.340 ;
        RECT 71.230 83.340 71.520 83.385 ;
        RECT 77.960 83.340 78.280 83.400 ;
        RECT 87.620 83.340 87.940 83.400 ;
        RECT 71.230 83.200 78.280 83.340 ;
        RECT 67.380 83.140 67.700 83.200 ;
        RECT 71.230 83.155 71.520 83.200 ;
        RECT 77.960 83.140 78.280 83.200 ;
        RECT 82.650 83.200 87.940 83.340 ;
        RECT 82.650 83.060 82.790 83.200 ;
        RECT 87.620 83.140 87.940 83.200 ;
        RECT 88.540 83.340 88.860 83.400 ;
        RECT 94.150 83.340 94.290 83.540 ;
        RECT 94.995 83.495 95.285 83.540 ;
        RECT 95.440 83.480 95.760 83.740 ;
        RECT 99.120 83.480 99.440 83.740 ;
        RECT 107.860 83.480 108.180 83.740 ;
        RECT 108.320 83.480 108.640 83.740 ;
        RECT 111.540 83.680 111.860 83.740 ;
        RECT 112.015 83.680 112.305 83.725 ;
        RECT 109.330 83.540 112.305 83.680 ;
        RECT 95.530 83.340 95.670 83.480 ;
        RECT 88.540 83.200 94.290 83.340 ;
        RECT 88.540 83.140 88.860 83.200 ;
        RECT 60.035 82.815 60.325 83.045 ;
        RECT 60.955 82.815 61.245 83.045 ;
        RECT 32.880 82.460 33.200 82.720 ;
        RECT 33.820 82.660 34.110 82.705 ;
        RECT 36.160 82.660 36.450 82.705 ;
        RECT 33.820 82.520 36.450 82.660 ;
        RECT 33.820 82.475 34.110 82.520 ;
        RECT 36.160 82.475 36.450 82.520 ;
        RECT 44.810 82.660 45.100 82.705 ;
        RECT 47.150 82.660 47.440 82.705 ;
        RECT 44.810 82.520 47.440 82.660 ;
        RECT 44.810 82.475 45.100 82.520 ;
        RECT 47.150 82.475 47.440 82.520 ;
        RECT 49.460 82.660 49.750 82.705 ;
        RECT 51.800 82.660 52.090 82.705 ;
        RECT 49.460 82.520 52.090 82.660 ;
        RECT 59.650 82.660 59.790 82.800 ;
        RECT 61.030 82.660 61.170 82.815 ;
        RECT 61.400 82.800 61.720 83.060 ;
        RECT 68.300 83.000 68.620 83.060 ;
        RECT 68.300 82.860 75.430 83.000 ;
        RECT 68.300 82.800 68.620 82.860 ;
        RECT 59.650 82.520 61.170 82.660 ;
        RECT 49.460 82.475 49.750 82.520 ;
        RECT 51.800 82.475 52.090 82.520 ;
        RECT 34.280 82.320 34.570 82.365 ;
        RECT 35.655 82.320 35.945 82.365 ;
        RECT 34.280 82.180 35.945 82.320 ;
        RECT 34.280 82.135 34.570 82.180 ;
        RECT 35.655 82.135 35.945 82.180 ;
        RECT 45.315 82.320 45.605 82.365 ;
        RECT 46.690 82.320 46.980 82.365 ;
        RECT 45.315 82.180 46.980 82.320 ;
        RECT 45.315 82.135 45.605 82.180 ;
        RECT 46.690 82.135 46.980 82.180 ;
        RECT 49.920 82.320 50.210 82.365 ;
        RECT 51.295 82.320 51.585 82.365 ;
        RECT 61.490 82.320 61.630 82.800 ;
        RECT 67.865 82.660 68.155 82.705 ;
        RECT 70.385 82.660 70.675 82.705 ;
        RECT 71.575 82.660 71.865 82.705 ;
        RECT 67.865 82.520 71.865 82.660 ;
        RECT 67.865 82.475 68.155 82.520 ;
        RECT 70.385 82.475 70.675 82.520 ;
        RECT 71.575 82.475 71.865 82.520 ;
        RECT 72.440 82.460 72.760 82.720 ;
        RECT 75.290 82.705 75.430 82.860 ;
        RECT 75.675 82.815 75.965 83.045 ;
        RECT 78.880 83.000 79.200 83.060 ;
        RECT 79.800 83.000 80.120 83.060 ;
        RECT 81.180 83.000 81.500 83.060 ;
        RECT 78.880 82.860 81.500 83.000 ;
        RECT 75.215 82.475 75.505 82.705 ;
        RECT 49.920 82.180 51.585 82.320 ;
        RECT 49.920 82.135 50.210 82.180 ;
        RECT 51.295 82.135 51.585 82.180 ;
        RECT 51.830 82.180 61.630 82.320 ;
        RECT 68.300 82.320 68.590 82.365 ;
        RECT 69.870 82.320 70.160 82.365 ;
        RECT 71.970 82.320 72.260 82.365 ;
        RECT 68.300 82.180 72.260 82.320 ;
        RECT 25.980 81.980 26.300 82.040 ;
        RECT 26.455 81.980 26.745 82.025 ;
        RECT 25.980 81.840 26.745 81.980 ;
        RECT 25.980 81.780 26.300 81.840 ;
        RECT 26.455 81.795 26.745 81.840 ;
        RECT 30.580 81.780 30.900 82.040 ;
        RECT 32.435 81.980 32.725 82.025 ;
        RECT 36.100 81.980 36.420 82.040 ;
        RECT 51.830 81.980 51.970 82.180 ;
        RECT 68.300 82.135 68.590 82.180 ;
        RECT 69.870 82.135 70.160 82.180 ;
        RECT 71.970 82.135 72.260 82.180 ;
        RECT 32.435 81.840 51.970 81.980 ;
        RECT 32.435 81.795 32.725 81.840 ;
        RECT 36.100 81.780 36.420 81.840 ;
        RECT 54.500 81.780 54.820 82.040 ;
        RECT 68.760 81.980 69.080 82.040 ;
        RECT 70.600 81.980 70.920 82.040 ;
        RECT 75.750 81.980 75.890 82.815 ;
        RECT 78.880 82.800 79.200 82.860 ;
        RECT 79.800 82.800 80.120 82.860 ;
        RECT 81.180 82.800 81.500 82.860 ;
        RECT 81.640 82.800 81.960 83.060 ;
        RECT 82.560 82.800 82.880 83.060 ;
        RECT 84.400 83.000 84.720 83.060 ;
        RECT 86.255 83.000 86.545 83.045 ;
        RECT 84.400 82.860 86.545 83.000 ;
        RECT 84.400 82.800 84.720 82.860 ;
        RECT 86.255 82.815 86.545 82.860 ;
        RECT 84.860 82.460 85.180 82.720 ;
        RECT 85.340 82.660 85.630 82.705 ;
        RECT 87.680 82.660 87.970 82.705 ;
        RECT 85.340 82.520 87.970 82.660 ;
        RECT 94.150 82.660 94.290 83.200 ;
        RECT 94.610 83.200 95.670 83.340 ;
        RECT 94.610 83.045 94.750 83.200 ;
        RECT 94.535 82.815 94.825 83.045 ;
        RECT 95.455 83.000 95.745 83.045 ;
        RECT 99.210 83.000 99.350 83.480 ;
        RECT 103.275 83.340 103.565 83.385 ;
        RECT 108.410 83.340 108.550 83.480 ;
        RECT 103.275 83.200 108.550 83.340 ;
        RECT 103.275 83.155 103.565 83.200 ;
        RECT 95.455 82.860 99.350 83.000 ;
        RECT 95.455 82.815 95.745 82.860 ;
        RECT 102.800 82.800 103.120 83.060 ;
        RECT 103.735 83.000 104.025 83.045 ;
        RECT 104.180 83.000 104.500 83.060 ;
        RECT 103.735 82.860 104.500 83.000 ;
        RECT 103.735 82.815 104.025 82.860 ;
        RECT 104.180 82.800 104.500 82.860 ;
        RECT 108.795 83.000 109.085 83.045 ;
        RECT 109.330 83.000 109.470 83.540 ;
        RECT 111.540 83.480 111.860 83.540 ;
        RECT 112.015 83.495 112.305 83.540 ;
        RECT 114.300 83.480 114.620 83.740 ;
        RECT 127.180 83.480 127.500 83.740 ;
        RECT 132.700 83.480 133.020 83.740 ;
        RECT 134.080 83.480 134.400 83.740 ;
        RECT 136.855 83.495 137.145 83.725 ;
        RECT 141.440 83.680 141.760 83.740 ;
        RECT 142.375 83.680 142.665 83.725 ;
        RECT 141.440 83.540 142.665 83.680 ;
        RECT 111.630 83.200 113.150 83.340 ;
        RECT 108.795 82.860 109.470 83.000 ;
        RECT 108.795 82.815 109.085 82.860 ;
        RECT 109.700 82.800 110.020 83.060 ;
        RECT 110.160 82.800 110.480 83.060 ;
        RECT 110.620 82.800 110.940 83.060 ;
        RECT 111.630 83.045 111.770 83.200 ;
        RECT 113.010 83.045 113.150 83.200 ;
        RECT 111.555 82.815 111.845 83.045 ;
        RECT 112.015 82.815 112.305 83.045 ;
        RECT 112.935 83.000 113.225 83.045 ;
        RECT 114.390 83.000 114.530 83.480 ;
        RECT 112.935 82.860 114.530 83.000 ;
        RECT 124.895 83.000 125.185 83.045 ;
        RECT 127.270 83.000 127.410 83.480 ;
        RECT 132.790 83.045 132.930 83.480 ;
        RECT 124.895 82.860 127.410 83.000 ;
        RECT 112.935 82.815 113.225 82.860 ;
        RECT 124.895 82.815 125.185 82.860 ;
        RECT 132.715 82.815 133.005 83.045 ;
        RECT 96.360 82.660 96.680 82.720 ;
        RECT 94.150 82.520 96.680 82.660 ;
        RECT 109.790 82.660 109.930 82.800 ;
        RECT 111.095 82.660 111.385 82.705 ;
        RECT 109.790 82.520 111.385 82.660 ;
        RECT 85.340 82.475 85.630 82.520 ;
        RECT 87.680 82.475 87.970 82.520 ;
        RECT 96.360 82.460 96.680 82.520 ;
        RECT 111.095 82.475 111.385 82.520 ;
        RECT 85.800 82.320 86.090 82.365 ;
        RECT 87.175 82.320 87.465 82.365 ;
        RECT 85.800 82.180 87.465 82.320 ;
        RECT 85.800 82.135 86.090 82.180 ;
        RECT 87.175 82.135 87.465 82.180 ;
        RECT 89.935 82.320 90.225 82.365 ;
        RECT 92.220 82.320 92.540 82.380 ;
        RECT 94.980 82.320 95.300 82.380 ;
        RECT 89.935 82.180 95.300 82.320 ;
        RECT 89.935 82.135 90.225 82.180 ;
        RECT 92.220 82.120 92.540 82.180 ;
        RECT 94.980 82.120 95.300 82.180 ;
        RECT 110.620 82.320 110.940 82.380 ;
        RECT 112.090 82.320 112.230 82.815 ;
        RECT 135.000 82.800 135.320 83.060 ;
        RECT 135.920 82.800 136.240 83.060 ;
        RECT 136.930 83.000 137.070 83.495 ;
        RECT 141.440 83.480 141.760 83.540 ;
        RECT 142.375 83.495 142.665 83.540 ;
        RECT 146.960 83.480 147.280 83.740 ;
        RECT 138.695 83.000 138.985 83.045 ;
        RECT 136.930 82.860 138.985 83.000 ;
        RECT 138.695 82.815 138.985 82.860 ;
        RECT 147.895 83.000 148.185 83.045 ;
        RECT 148.800 83.000 149.120 83.060 ;
        RECT 147.895 82.860 149.120 83.000 ;
        RECT 147.895 82.815 148.185 82.860 ;
        RECT 148.800 82.800 149.120 82.860 ;
        RECT 137.300 82.460 137.620 82.720 ;
        RECT 137.780 82.660 138.070 82.705 ;
        RECT 140.120 82.660 140.410 82.705 ;
        RECT 137.780 82.520 140.410 82.660 ;
        RECT 137.780 82.475 138.070 82.520 ;
        RECT 140.120 82.475 140.410 82.520 ;
        RECT 148.340 82.460 148.660 82.720 ;
        RECT 149.275 82.660 149.565 82.705 ;
        RECT 150.640 82.660 150.960 82.720 ;
        RECT 149.275 82.520 150.960 82.660 ;
        RECT 149.275 82.475 149.565 82.520 ;
        RECT 150.640 82.460 150.960 82.520 ;
        RECT 110.620 82.180 112.230 82.320 ;
        RECT 138.240 82.320 138.530 82.365 ;
        RECT 139.615 82.320 139.905 82.365 ;
        RECT 138.240 82.180 139.905 82.320 ;
        RECT 110.620 82.120 110.940 82.180 ;
        RECT 138.240 82.135 138.530 82.180 ;
        RECT 139.615 82.135 139.905 82.180 ;
        RECT 141.440 82.320 141.760 82.380 ;
        RECT 142.835 82.320 143.125 82.365 ;
        RECT 141.440 82.180 143.125 82.320 ;
        RECT 148.430 82.320 148.570 82.460 ;
        RECT 148.815 82.320 149.105 82.365 ;
        RECT 148.430 82.180 149.105 82.320 ;
        RECT 141.440 82.120 141.760 82.180 ;
        RECT 142.835 82.135 143.125 82.180 ;
        RECT 148.815 82.135 149.105 82.180 ;
        RECT 68.760 81.840 75.890 81.980 ;
        RECT 68.760 81.780 69.080 81.840 ;
        RECT 70.600 81.780 70.920 81.840 ;
        RECT 77.500 81.780 77.820 82.040 ;
        RECT 78.895 81.980 79.185 82.025 ;
        RECT 80.260 81.980 80.580 82.040 ;
        RECT 78.895 81.840 80.580 81.980 ;
        RECT 78.895 81.795 79.185 81.840 ;
        RECT 80.260 81.780 80.580 81.840 ;
        RECT 83.480 81.780 83.800 82.040 ;
        RECT 90.840 81.780 91.160 82.040 ;
        RECT 97.740 81.980 98.060 82.040 ;
        RECT 98.215 81.980 98.505 82.025 ;
        RECT 97.740 81.840 98.505 81.980 ;
        RECT 97.740 81.780 98.060 81.840 ;
        RECT 98.215 81.795 98.505 81.840 ;
        RECT 123.500 81.980 123.820 82.040 ;
        RECT 127.640 81.980 127.960 82.040 ;
        RECT 123.500 81.840 127.960 81.980 ;
        RECT 123.500 81.780 123.820 81.840 ;
        RECT 127.640 81.780 127.960 81.840 ;
        RECT 22.690 81.160 157.010 81.640 ;
        RECT 31.040 80.760 31.360 81.020 ;
        RECT 33.355 80.960 33.645 81.005 ;
        RECT 34.720 80.960 35.040 81.020 ;
        RECT 33.355 80.820 35.040 80.960 ;
        RECT 33.355 80.775 33.645 80.820 ;
        RECT 34.720 80.760 35.040 80.820 ;
        RECT 45.315 80.960 45.605 81.005 ;
        RECT 46.220 80.960 46.540 81.020 ;
        RECT 45.315 80.820 46.540 80.960 ;
        RECT 45.315 80.775 45.605 80.820 ;
        RECT 46.220 80.760 46.540 80.820 ;
        RECT 49.455 80.960 49.745 81.005 ;
        RECT 50.360 80.960 50.680 81.020 ;
        RECT 54.500 80.960 54.820 81.020 ;
        RECT 49.455 80.820 50.680 80.960 ;
        RECT 49.455 80.775 49.745 80.820 ;
        RECT 50.360 80.760 50.680 80.820 ;
        RECT 53.210 80.820 54.820 80.960 ;
        RECT 26.920 80.620 27.210 80.665 ;
        RECT 28.295 80.620 28.585 80.665 ;
        RECT 26.920 80.480 28.585 80.620 ;
        RECT 26.920 80.435 27.210 80.480 ;
        RECT 28.295 80.435 28.585 80.480 ;
        RECT 53.210 80.325 53.350 80.820 ;
        RECT 54.500 80.760 54.820 80.820 ;
        RECT 58.180 80.760 58.500 81.020 ;
        RECT 71.075 80.960 71.365 81.005 ;
        RECT 79.340 80.960 79.660 81.020 ;
        RECT 71.075 80.820 79.660 80.960 ;
        RECT 71.075 80.775 71.365 80.820 ;
        RECT 79.340 80.760 79.660 80.820 ;
        RECT 79.800 80.960 80.120 81.020 ;
        RECT 83.495 80.960 83.785 81.005 ;
        RECT 84.400 80.960 84.720 81.020 ;
        RECT 79.800 80.820 82.100 80.960 ;
        RECT 79.800 80.760 80.120 80.820 ;
        RECT 54.060 80.620 54.350 80.665 ;
        RECT 55.435 80.620 55.725 80.665 ;
        RECT 54.060 80.480 55.725 80.620 ;
        RECT 54.060 80.435 54.350 80.480 ;
        RECT 55.435 80.435 55.725 80.480 ;
        RECT 76.120 80.420 76.440 80.680 ;
        RECT 78.895 80.620 79.185 80.665 ;
        RECT 80.270 80.620 80.560 80.665 ;
        RECT 78.895 80.480 80.560 80.620 ;
        RECT 81.960 80.620 82.100 80.820 ;
        RECT 83.495 80.820 84.720 80.960 ;
        RECT 83.495 80.775 83.785 80.820 ;
        RECT 84.400 80.760 84.720 80.820 ;
        RECT 84.860 80.760 85.180 81.020 ;
        RECT 91.390 80.820 95.670 80.960 ;
        RECT 91.390 80.620 91.530 80.820 ;
        RECT 81.960 80.480 91.530 80.620 ;
        RECT 91.780 80.620 92.070 80.665 ;
        RECT 93.155 80.620 93.445 80.665 ;
        RECT 91.780 80.480 93.445 80.620 ;
        RECT 95.530 80.620 95.670 80.820 ;
        RECT 95.900 80.760 96.220 81.020 ;
        RECT 98.290 80.820 102.570 80.960 ;
        RECT 98.290 80.620 98.430 80.820 ;
        RECT 95.530 80.480 98.430 80.620 ;
        RECT 98.680 80.620 98.970 80.665 ;
        RECT 100.055 80.620 100.345 80.665 ;
        RECT 98.680 80.480 100.345 80.620 ;
        RECT 102.430 80.620 102.570 80.820 ;
        RECT 102.800 80.760 103.120 81.020 ;
        RECT 119.820 80.960 120.140 81.020 ;
        RECT 123.500 80.960 123.820 81.020 ;
        RECT 118.070 80.820 123.820 80.960 ;
        RECT 113.380 80.620 113.700 80.680 ;
        RECT 102.430 80.480 113.700 80.620 ;
        RECT 78.895 80.435 79.185 80.480 ;
        RECT 80.270 80.435 80.560 80.480 ;
        RECT 91.780 80.435 92.070 80.480 ;
        RECT 93.155 80.435 93.445 80.480 ;
        RECT 98.680 80.435 98.970 80.480 ;
        RECT 100.055 80.435 100.345 80.480 ;
        RECT 113.380 80.420 113.700 80.480 ;
        RECT 26.460 80.280 26.750 80.325 ;
        RECT 28.800 80.280 29.090 80.325 ;
        RECT 26.460 80.140 29.090 80.280 ;
        RECT 26.460 80.095 26.750 80.140 ;
        RECT 28.800 80.095 29.090 80.140 ;
        RECT 53.135 80.095 53.425 80.325 ;
        RECT 53.600 80.280 53.890 80.325 ;
        RECT 55.940 80.280 56.230 80.325 ;
        RECT 53.600 80.140 56.230 80.280 ;
        RECT 53.600 80.095 53.890 80.140 ;
        RECT 55.940 80.095 56.230 80.140 ;
        RECT 63.715 80.280 64.005 80.325 ;
        RECT 64.160 80.280 64.480 80.340 ;
        RECT 63.715 80.140 64.480 80.280 ;
        RECT 63.715 80.095 64.005 80.140 ;
        RECT 64.160 80.080 64.480 80.140 ;
        RECT 78.390 80.280 78.680 80.325 ;
        RECT 80.730 80.280 81.020 80.325 ;
        RECT 78.390 80.140 81.020 80.280 ;
        RECT 78.390 80.095 78.680 80.140 ;
        RECT 80.730 80.095 81.020 80.140 ;
        RECT 90.840 80.080 91.160 80.340 ;
        RECT 91.320 80.280 91.610 80.325 ;
        RECT 93.660 80.280 93.950 80.325 ;
        RECT 91.320 80.140 93.950 80.280 ;
        RECT 91.320 80.095 91.610 80.140 ;
        RECT 93.660 80.095 93.950 80.140 ;
        RECT 98.220 80.280 98.510 80.325 ;
        RECT 100.560 80.280 100.850 80.325 ;
        RECT 98.220 80.140 100.850 80.280 ;
        RECT 98.220 80.095 98.510 80.140 ;
        RECT 100.560 80.095 100.850 80.140 ;
        RECT 25.520 79.740 25.840 80.000 ;
        RECT 25.980 79.740 26.300 80.000 ;
        RECT 27.375 79.755 27.665 79.985 ;
        RECT 30.580 79.940 30.900 80.000 ;
        RECT 33.355 79.940 33.645 79.985 ;
        RECT 30.580 79.800 33.645 79.940 ;
        RECT 27.450 79.600 27.590 79.755 ;
        RECT 30.580 79.740 30.900 79.800 ;
        RECT 33.355 79.755 33.645 79.800 ;
        RECT 34.275 79.940 34.565 79.985 ;
        RECT 36.560 79.940 36.880 80.000 ;
        RECT 34.275 79.800 36.880 79.940 ;
        RECT 34.275 79.755 34.565 79.800 ;
        RECT 36.560 79.740 36.880 79.800 ;
        RECT 44.395 79.940 44.685 79.985 ;
        RECT 45.300 79.940 45.620 80.000 ;
        RECT 44.395 79.800 45.620 79.940 ;
        RECT 44.395 79.755 44.685 79.800 ;
        RECT 45.300 79.740 45.620 79.800 ;
        RECT 48.520 79.740 48.840 80.000 ;
        RECT 51.740 79.740 52.060 80.000 ;
        RECT 54.515 79.755 54.805 79.985 ;
        RECT 62.335 79.755 62.625 79.985 ;
        RECT 54.590 79.600 54.730 79.755 ;
        RECT 27.450 79.460 33.800 79.600 ;
        RECT 33.660 79.260 33.800 79.460 ;
        RECT 52.750 79.460 54.730 79.600 ;
        RECT 37.020 79.260 37.340 79.320 ;
        RECT 52.750 79.305 52.890 79.460 ;
        RECT 62.410 79.320 62.550 79.755 ;
        RECT 62.780 79.740 63.100 80.000 ;
        RECT 70.155 79.755 70.445 79.985 ;
        RECT 71.060 79.940 71.380 80.000 ;
        RECT 72.455 79.940 72.745 79.985 ;
        RECT 71.060 79.800 72.745 79.940 ;
        RECT 33.660 79.120 37.340 79.260 ;
        RECT 37.020 79.060 37.340 79.120 ;
        RECT 52.675 79.075 52.965 79.305 ;
        RECT 62.320 79.060 62.640 79.320 ;
        RECT 63.700 79.060 64.020 79.320 ;
        RECT 67.840 79.260 68.160 79.320 ;
        RECT 70.230 79.260 70.370 79.755 ;
        RECT 71.060 79.740 71.380 79.800 ;
        RECT 72.455 79.755 72.745 79.800 ;
        RECT 73.820 79.740 74.140 80.000 ;
        RECT 79.815 79.755 80.105 79.985 ;
        RECT 80.260 79.940 80.580 80.000 ;
        RECT 81.195 79.940 81.485 79.985 ;
        RECT 80.260 79.800 81.485 79.940 ;
        RECT 71.995 79.600 72.285 79.645 ;
        RECT 77.500 79.600 77.820 79.660 ;
        RECT 71.995 79.460 77.820 79.600 ;
        RECT 79.890 79.600 80.030 79.755 ;
        RECT 80.260 79.740 80.580 79.800 ;
        RECT 81.195 79.755 81.485 79.800 ;
        RECT 82.575 79.755 82.865 79.985 ;
        RECT 80.720 79.600 81.040 79.660 ;
        RECT 82.650 79.600 82.790 79.755 ;
        RECT 83.480 79.740 83.800 80.000 ;
        RECT 85.320 79.740 85.640 80.000 ;
        RECT 92.220 79.740 92.540 80.000 ;
        RECT 96.360 79.740 96.680 80.000 ;
        RECT 97.740 79.740 98.060 80.000 ;
        RECT 118.070 79.985 118.210 80.820 ;
        RECT 119.820 80.760 120.140 80.820 ;
        RECT 123.500 80.760 123.820 80.820 ;
        RECT 124.895 80.960 125.185 81.005 ;
        RECT 128.560 80.960 128.880 81.020 ;
        RECT 133.635 80.960 133.925 81.005 ;
        RECT 124.895 80.820 133.925 80.960 ;
        RECT 124.895 80.775 125.185 80.820 ;
        RECT 128.560 80.760 128.880 80.820 ;
        RECT 133.635 80.775 133.925 80.820 ;
        RECT 135.475 80.960 135.765 81.005 ;
        RECT 135.920 80.960 136.240 81.020 ;
        RECT 135.475 80.820 136.240 80.960 ;
        RECT 135.475 80.775 135.765 80.820 ;
        RECT 135.920 80.760 136.240 80.820 ;
        RECT 138.680 80.960 139.000 81.020 ;
        RECT 142.360 80.960 142.680 81.020 ;
        RECT 149.275 80.960 149.565 81.005 ;
        RECT 151.560 80.960 151.880 81.020 ;
        RECT 138.680 80.820 151.880 80.960 ;
        RECT 138.680 80.760 139.000 80.820 ;
        RECT 142.360 80.760 142.680 80.820 ;
        RECT 149.275 80.775 149.565 80.820 ;
        RECT 151.560 80.760 151.880 80.820 ;
        RECT 152.035 80.775 152.325 81.005 ;
        RECT 118.990 80.480 126.030 80.620 ;
        RECT 118.990 80.000 119.130 80.480 ;
        RECT 125.890 80.340 126.030 80.480 ;
        RECT 127.640 80.420 127.960 80.680 ;
        RECT 148.800 80.620 149.120 80.680 ;
        RECT 152.110 80.620 152.250 80.775 ;
        RECT 148.800 80.480 152.250 80.620 ;
        RECT 148.800 80.420 149.120 80.480 ;
        RECT 121.290 80.140 124.190 80.280 ;
        RECT 99.135 79.755 99.425 79.985 ;
        RECT 117.995 79.755 118.285 79.985 ;
        RECT 85.410 79.600 85.550 79.740 ;
        RECT 99.210 79.600 99.350 79.755 ;
        RECT 118.900 79.740 119.220 80.000 ;
        RECT 121.290 79.645 121.430 80.140 ;
        RECT 121.660 79.940 121.980 80.000 ;
        RECT 122.595 79.940 122.885 79.985 ;
        RECT 121.660 79.800 122.885 79.940 ;
        RECT 121.660 79.740 121.980 79.800 ;
        RECT 122.595 79.755 122.885 79.800 ;
        RECT 123.500 79.740 123.820 80.000 ;
        RECT 124.050 79.985 124.190 80.140 ;
        RECT 125.800 80.080 126.120 80.340 ;
        RECT 128.115 80.280 128.405 80.325 ;
        RECT 152.495 80.280 152.785 80.325 ;
        RECT 128.115 80.140 130.170 80.280 ;
        RECT 128.115 80.095 128.405 80.140 ;
        RECT 123.975 79.755 124.265 79.985 ;
        RECT 124.895 79.940 125.185 79.985 ;
        RECT 127.180 79.940 127.500 80.000 ;
        RECT 128.575 79.940 128.865 79.985 ;
        RECT 124.510 79.800 128.865 79.940 ;
        RECT 124.510 79.660 124.650 79.800 ;
        RECT 124.895 79.755 125.185 79.800 ;
        RECT 127.180 79.740 127.500 79.800 ;
        RECT 128.575 79.755 128.865 79.800 ;
        RECT 129.495 79.940 129.785 79.985 ;
        RECT 130.030 79.940 130.170 80.140 ;
        RECT 147.970 80.140 152.785 80.280 ;
        RECT 147.970 80.000 148.110 80.140 ;
        RECT 152.495 80.095 152.785 80.140 ;
        RECT 130.875 79.940 131.165 79.985 ;
        RECT 129.495 79.800 131.165 79.940 ;
        RECT 129.495 79.755 129.785 79.800 ;
        RECT 130.875 79.755 131.165 79.800 ;
        RECT 133.620 79.740 133.940 80.000 ;
        RECT 134.540 79.740 134.860 80.000 ;
        RECT 138.680 79.940 139.000 80.000 ;
        RECT 140.535 79.940 140.825 79.985 ;
        RECT 138.680 79.800 140.825 79.940 ;
        RECT 138.680 79.740 139.000 79.800 ;
        RECT 140.535 79.755 140.825 79.800 ;
        RECT 142.820 79.740 143.140 80.000 ;
        RECT 147.880 79.740 148.200 80.000 ;
        RECT 150.180 79.940 150.500 80.000 ;
        RECT 152.035 79.940 152.325 79.985 ;
        RECT 150.180 79.800 152.325 79.940 ;
        RECT 150.180 79.740 150.500 79.800 ;
        RECT 152.035 79.755 152.325 79.800 ;
        RECT 79.890 79.460 80.490 79.600 ;
        RECT 71.995 79.415 72.285 79.460 ;
        RECT 77.500 79.400 77.820 79.460 ;
        RECT 80.350 79.320 80.490 79.460 ;
        RECT 80.720 79.460 85.550 79.600 ;
        RECT 97.370 79.460 99.350 79.600 ;
        RECT 119.835 79.600 120.125 79.645 ;
        RECT 121.215 79.600 121.505 79.645 ;
        RECT 119.835 79.460 121.505 79.600 ;
        RECT 80.720 79.400 81.040 79.460 ;
        RECT 76.580 79.260 76.900 79.320 ;
        RECT 79.340 79.260 79.660 79.320 ;
        RECT 67.840 79.120 79.660 79.260 ;
        RECT 67.840 79.060 68.160 79.120 ;
        RECT 76.580 79.060 76.900 79.120 ;
        RECT 79.340 79.060 79.660 79.120 ;
        RECT 80.260 79.060 80.580 79.320 ;
        RECT 97.370 79.305 97.510 79.460 ;
        RECT 119.835 79.415 120.125 79.460 ;
        RECT 121.215 79.415 121.505 79.460 ;
        RECT 122.135 79.415 122.425 79.645 ;
        RECT 123.055 79.600 123.345 79.645 ;
        RECT 124.420 79.600 124.740 79.660 ;
        RECT 123.055 79.460 124.740 79.600 ;
        RECT 123.055 79.415 123.345 79.460 ;
        RECT 97.295 79.075 97.585 79.305 ;
        RECT 120.280 79.060 120.600 79.320 ;
        RECT 120.740 79.260 121.060 79.320 ;
        RECT 122.210 79.260 122.350 79.415 ;
        RECT 124.420 79.400 124.740 79.460 ;
        RECT 125.340 79.400 125.660 79.660 ;
        RECT 123.500 79.260 123.820 79.320 ;
        RECT 125.430 79.260 125.570 79.400 ;
        RECT 120.740 79.120 125.570 79.260 ;
        RECT 120.740 79.060 121.060 79.120 ;
        RECT 123.500 79.060 123.820 79.120 ;
        RECT 130.400 79.060 130.720 79.320 ;
        RECT 130.860 79.260 131.180 79.320 ;
        RECT 131.335 79.260 131.625 79.305 ;
        RECT 130.860 79.120 131.625 79.260 ;
        RECT 130.860 79.060 131.180 79.120 ;
        RECT 131.335 79.075 131.625 79.120 ;
        RECT 153.860 79.060 154.180 79.320 ;
        RECT 22.690 78.440 157.810 78.920 ;
        RECT 25.520 78.040 25.840 78.300 ;
        RECT 29.660 78.240 29.980 78.300 ;
        RECT 31.055 78.240 31.345 78.285 ;
        RECT 29.660 78.100 31.345 78.240 ;
        RECT 29.660 78.040 29.980 78.100 ;
        RECT 31.055 78.055 31.345 78.100 ;
        RECT 48.520 78.240 48.840 78.300 ;
        RECT 48.995 78.240 49.285 78.285 ;
        RECT 48.520 78.100 49.285 78.240 ;
        RECT 48.520 78.040 48.840 78.100 ;
        RECT 48.995 78.055 49.285 78.100 ;
        RECT 60.940 78.040 61.260 78.300 ;
        RECT 63.700 78.240 64.020 78.300 ;
        RECT 65.635 78.240 65.925 78.285 ;
        RECT 63.700 78.100 65.925 78.240 ;
        RECT 63.700 78.040 64.020 78.100 ;
        RECT 65.635 78.055 65.925 78.100 ;
        RECT 68.760 78.040 69.080 78.300 ;
        RECT 73.820 78.040 74.140 78.300 ;
        RECT 81.180 78.240 81.500 78.300 ;
        RECT 91.775 78.240 92.065 78.285 ;
        RECT 92.220 78.240 92.540 78.300 ;
        RECT 81.180 78.100 83.710 78.240 ;
        RECT 81.180 78.040 81.500 78.100 ;
        RECT 25.610 77.560 25.750 78.040 ;
        RECT 32.880 77.900 33.200 77.960 ;
        RECT 35.655 77.900 35.945 77.945 ;
        RECT 40.700 77.900 41.020 77.960 ;
        RECT 61.400 77.900 61.720 77.960 ;
        RECT 62.780 77.900 63.100 77.960 ;
        RECT 32.880 77.760 34.950 77.900 ;
        RECT 32.880 77.700 33.200 77.760 ;
        RECT 25.995 77.560 26.285 77.605 ;
        RECT 25.610 77.420 26.285 77.560 ;
        RECT 25.995 77.375 26.285 77.420 ;
        RECT 27.375 77.560 27.665 77.605 ;
        RECT 30.580 77.560 30.900 77.620 ;
        RECT 34.810 77.605 34.950 77.760 ;
        RECT 35.655 77.760 36.790 77.900 ;
        RECT 35.655 77.715 35.945 77.760 ;
        RECT 36.650 77.620 36.790 77.760 ;
        RECT 37.110 77.760 45.070 77.900 ;
        RECT 27.375 77.420 30.900 77.560 ;
        RECT 27.375 77.375 27.665 77.420 ;
        RECT 30.580 77.360 30.900 77.420 ;
        RECT 34.735 77.560 35.025 77.605 ;
        RECT 35.180 77.560 35.500 77.620 ;
        RECT 34.735 77.420 35.500 77.560 ;
        RECT 34.735 77.375 35.025 77.420 ;
        RECT 35.180 77.360 35.500 77.420 ;
        RECT 36.115 77.375 36.405 77.605 ;
        RECT 26.460 77.220 26.750 77.265 ;
        RECT 28.800 77.220 29.090 77.265 ;
        RECT 26.460 77.080 29.090 77.220 ;
        RECT 26.460 77.035 26.750 77.080 ;
        RECT 28.800 77.035 29.090 77.080 ;
        RECT 32.880 77.220 33.200 77.280 ;
        RECT 33.815 77.220 34.105 77.265 ;
        RECT 36.190 77.220 36.330 77.375 ;
        RECT 36.560 77.360 36.880 77.620 ;
        RECT 37.110 77.605 37.250 77.760 ;
        RECT 40.700 77.700 41.020 77.760 ;
        RECT 37.035 77.375 37.325 77.605 ;
        RECT 32.880 77.080 36.330 77.220 ;
        RECT 37.110 77.220 37.250 77.375 ;
        RECT 37.480 77.360 37.800 77.620 ;
        RECT 38.415 77.560 38.705 77.605 ;
        RECT 41.620 77.560 41.940 77.620 ;
        RECT 43.920 77.560 44.240 77.620 ;
        RECT 44.395 77.560 44.685 77.605 ;
        RECT 38.415 77.420 41.940 77.560 ;
        RECT 38.415 77.375 38.705 77.420 ;
        RECT 41.620 77.360 41.940 77.420 ;
        RECT 43.090 77.420 44.685 77.560 ;
        RECT 37.955 77.220 38.245 77.265 ;
        RECT 37.110 77.080 38.245 77.220 ;
        RECT 32.880 77.020 33.200 77.080 ;
        RECT 33.815 77.035 34.105 77.080 ;
        RECT 37.955 77.035 38.245 77.080 ;
        RECT 40.715 77.220 41.005 77.265 ;
        RECT 41.160 77.220 41.480 77.280 ;
        RECT 43.090 77.265 43.230 77.420 ;
        RECT 43.920 77.360 44.240 77.420 ;
        RECT 44.395 77.375 44.685 77.420 ;
        RECT 40.715 77.080 41.480 77.220 ;
        RECT 40.715 77.035 41.005 77.080 ;
        RECT 41.160 77.020 41.480 77.080 ;
        RECT 43.015 77.035 43.305 77.265 ;
        RECT 43.475 77.220 43.765 77.265 ;
        RECT 44.930 77.220 45.070 77.760 ;
        RECT 59.650 77.760 61.720 77.900 ;
        RECT 45.315 77.560 45.605 77.605 ;
        RECT 45.775 77.560 46.065 77.605 ;
        RECT 45.315 77.420 46.065 77.560 ;
        RECT 45.315 77.375 45.605 77.420 ;
        RECT 45.775 77.375 46.065 77.420 ;
        RECT 47.600 77.560 47.920 77.620 ;
        RECT 59.650 77.605 59.790 77.760 ;
        RECT 61.400 77.700 61.720 77.760 ;
        RECT 61.950 77.760 63.100 77.900 ;
        RECT 61.950 77.605 62.090 77.760 ;
        RECT 62.780 77.700 63.100 77.760 ;
        RECT 64.635 77.900 64.925 77.945 ;
        RECT 65.080 77.900 65.400 77.960 ;
        RECT 67.840 77.900 68.160 77.960 ;
        RECT 64.635 77.760 68.160 77.900 ;
        RECT 64.635 77.715 64.925 77.760 ;
        RECT 65.080 77.700 65.400 77.760 ;
        RECT 67.840 77.700 68.160 77.760 ;
        RECT 73.360 77.700 73.680 77.960 ;
        RECT 50.835 77.560 51.125 77.605 ;
        RECT 47.600 77.420 51.125 77.560 ;
        RECT 47.600 77.360 47.920 77.420 ;
        RECT 50.835 77.375 51.125 77.420 ;
        RECT 57.275 77.375 57.565 77.605 ;
        RECT 58.195 77.560 58.485 77.605 ;
        RECT 59.575 77.560 59.865 77.605 ;
        RECT 58.195 77.420 59.865 77.560 ;
        RECT 58.195 77.375 58.485 77.420 ;
        RECT 59.575 77.375 59.865 77.420 ;
        RECT 60.495 77.560 60.785 77.605 ;
        RECT 61.875 77.560 62.165 77.605 ;
        RECT 63.255 77.560 63.545 77.605 ;
        RECT 60.495 77.420 62.165 77.560 ;
        RECT 60.495 77.375 60.785 77.420 ;
        RECT 61.875 77.375 62.165 77.420 ;
        RECT 62.410 77.420 63.545 77.560 ;
        RECT 43.475 77.080 45.070 77.220 ;
        RECT 49.900 77.220 50.220 77.280 ;
        RECT 50.375 77.220 50.665 77.265 ;
        RECT 49.900 77.080 50.665 77.220 ;
        RECT 57.350 77.220 57.490 77.375 ;
        RECT 58.655 77.220 58.945 77.265 ;
        RECT 60.020 77.220 60.340 77.280 ;
        RECT 57.350 77.080 60.340 77.220 ;
        RECT 43.475 77.035 43.765 77.080 ;
        RECT 49.900 77.020 50.220 77.080 ;
        RECT 50.375 77.035 50.665 77.080 ;
        RECT 58.655 77.035 58.945 77.080 ;
        RECT 60.020 77.020 60.340 77.080 ;
        RECT 62.410 76.940 62.550 77.420 ;
        RECT 63.255 77.375 63.545 77.420 ;
        RECT 64.160 77.360 64.480 77.620 ;
        RECT 66.935 77.560 67.225 77.605 ;
        RECT 66.550 77.420 67.225 77.560 ;
        RECT 26.920 76.880 27.210 76.925 ;
        RECT 28.295 76.880 28.585 76.925 ;
        RECT 26.920 76.740 28.585 76.880 ;
        RECT 26.920 76.695 27.210 76.740 ;
        RECT 28.295 76.695 28.585 76.740 ;
        RECT 37.020 76.880 37.340 76.940 ;
        RECT 37.020 76.740 40.470 76.880 ;
        RECT 37.020 76.680 37.340 76.740 ;
        RECT 40.330 76.540 40.470 76.740 ;
        RECT 42.080 76.680 42.400 76.940 ;
        RECT 58.195 76.880 58.485 76.925 ;
        RECT 62.320 76.880 62.640 76.940 ;
        RECT 66.550 76.925 66.690 77.420 ;
        RECT 66.935 77.375 67.225 77.420 ;
        RECT 72.455 77.560 72.745 77.605 ;
        RECT 73.450 77.560 73.590 77.700 ;
        RECT 73.910 77.605 74.050 78.040 ;
        RECT 75.675 77.900 75.965 77.945 ;
        RECT 77.515 77.900 77.805 77.945 ;
        RECT 80.260 77.900 80.580 77.960 ;
        RECT 83.570 77.945 83.710 78.100 ;
        RECT 91.775 78.100 92.540 78.240 ;
        RECT 91.775 78.055 92.065 78.100 ;
        RECT 92.220 78.040 92.540 78.100 ;
        RECT 95.455 78.240 95.745 78.285 ;
        RECT 96.360 78.240 96.680 78.300 ;
        RECT 95.455 78.100 96.680 78.240 ;
        RECT 95.455 78.055 95.745 78.100 ;
        RECT 96.360 78.040 96.680 78.100 ;
        RECT 110.160 78.240 110.480 78.300 ;
        RECT 127.180 78.285 127.500 78.300 ;
        RECT 110.635 78.240 110.925 78.285 ;
        RECT 110.160 78.100 110.925 78.240 ;
        RECT 110.160 78.040 110.480 78.100 ;
        RECT 110.635 78.055 110.925 78.100 ;
        RECT 127.180 78.055 127.565 78.285 ;
        RECT 127.180 78.040 127.500 78.055 ;
        RECT 130.400 78.040 130.720 78.300 ;
        RECT 137.315 78.055 137.605 78.285 ;
        RECT 139.615 78.055 139.905 78.285 ;
        RECT 75.675 77.760 80.030 77.900 ;
        RECT 75.675 77.715 75.965 77.760 ;
        RECT 77.515 77.715 77.805 77.760 ;
        RECT 72.455 77.420 73.590 77.560 ;
        RECT 72.455 77.375 72.745 77.420 ;
        RECT 73.835 77.375 74.125 77.605 ;
        RECT 76.120 77.560 76.440 77.620 ;
        RECT 76.595 77.560 76.885 77.605 ;
        RECT 76.120 77.420 76.885 77.560 ;
        RECT 76.120 77.360 76.440 77.420 ;
        RECT 76.595 77.375 76.885 77.420 ;
        RECT 78.435 77.560 78.725 77.605 ;
        RECT 78.880 77.560 79.200 77.620 ;
        RECT 79.890 77.605 80.030 77.760 ;
        RECT 80.260 77.760 83.250 77.900 ;
        RECT 80.260 77.700 80.580 77.760 ;
        RECT 78.435 77.420 79.200 77.560 ;
        RECT 78.435 77.375 78.725 77.420 ;
        RECT 78.880 77.360 79.200 77.420 ;
        RECT 79.355 77.375 79.645 77.605 ;
        RECT 79.815 77.375 80.105 77.605 ;
        RECT 80.735 77.375 81.025 77.605 ;
        RECT 81.195 77.375 81.485 77.605 ;
        RECT 82.115 77.560 82.405 77.605 ;
        RECT 82.560 77.560 82.880 77.620 ;
        RECT 82.115 77.420 82.880 77.560 ;
        RECT 83.110 77.560 83.250 77.760 ;
        RECT 83.495 77.715 83.785 77.945 ;
        RECT 120.280 77.900 120.600 77.960 ;
        RECT 84.895 77.760 87.850 77.900 ;
        RECT 84.895 77.560 85.035 77.760 ;
        RECT 87.160 77.560 87.480 77.620 ;
        RECT 83.110 77.420 85.035 77.560 ;
        RECT 85.870 77.420 87.480 77.560 ;
        RECT 82.115 77.375 82.405 77.420 ;
        RECT 71.030 77.220 71.320 77.265 ;
        RECT 73.370 77.220 73.660 77.265 ;
        RECT 71.030 77.080 73.660 77.220 ;
        RECT 79.430 77.220 79.570 77.375 ;
        RECT 80.260 77.220 80.580 77.280 ;
        RECT 79.430 77.080 80.580 77.220 ;
        RECT 71.030 77.035 71.320 77.080 ;
        RECT 73.370 77.035 73.660 77.080 ;
        RECT 80.260 77.020 80.580 77.080 ;
        RECT 42.630 76.740 50.130 76.880 ;
        RECT 42.630 76.540 42.770 76.740 ;
        RECT 40.330 76.400 42.770 76.540 ;
        RECT 46.695 76.540 46.985 76.585 ;
        RECT 47.140 76.540 47.460 76.600 ;
        RECT 49.990 76.585 50.130 76.740 ;
        RECT 58.195 76.740 62.640 76.880 ;
        RECT 58.195 76.695 58.485 76.740 ;
        RECT 62.320 76.680 62.640 76.740 ;
        RECT 66.475 76.695 66.765 76.925 ;
        RECT 71.535 76.880 71.825 76.925 ;
        RECT 72.910 76.880 73.200 76.925 ;
        RECT 71.535 76.740 73.200 76.880 ;
        RECT 80.810 76.880 80.950 77.375 ;
        RECT 81.270 77.220 81.410 77.375 ;
        RECT 82.560 77.360 82.880 77.420 ;
        RECT 83.940 77.220 84.260 77.280 ;
        RECT 85.870 77.265 86.010 77.420 ;
        RECT 87.160 77.360 87.480 77.420 ;
        RECT 81.270 77.080 84.260 77.220 ;
        RECT 83.940 77.020 84.260 77.080 ;
        RECT 85.795 77.035 86.085 77.265 ;
        RECT 86.255 77.035 86.545 77.265 ;
        RECT 87.710 77.220 87.850 77.760 ;
        RECT 119.450 77.760 120.600 77.900 ;
        RECT 88.095 77.560 88.385 77.605 ;
        RECT 88.555 77.560 88.845 77.605 ;
        RECT 88.095 77.420 88.845 77.560 ;
        RECT 88.095 77.375 88.385 77.420 ;
        RECT 88.555 77.375 88.845 77.420 ;
        RECT 90.840 77.360 91.160 77.620 ;
        RECT 93.600 77.360 93.920 77.620 ;
        RECT 94.520 77.360 94.840 77.620 ;
        RECT 102.800 77.360 103.120 77.620 ;
        RECT 107.415 77.560 107.705 77.605 ;
        RECT 107.860 77.560 108.180 77.620 ;
        RECT 107.415 77.420 108.180 77.560 ;
        RECT 107.415 77.375 107.705 77.420 ;
        RECT 107.860 77.360 108.180 77.420 ;
        RECT 108.320 77.360 108.640 77.620 ;
        RECT 116.600 77.605 116.920 77.620 ;
        RECT 109.715 77.560 110.005 77.605 ;
        RECT 109.330 77.420 110.005 77.560 ;
        RECT 109.330 77.280 109.470 77.420 ;
        RECT 109.715 77.375 110.005 77.420 ;
        RECT 116.600 77.375 116.950 77.605 ;
        RECT 118.440 77.560 118.760 77.620 ;
        RECT 119.450 77.605 119.590 77.760 ;
        RECT 120.280 77.700 120.600 77.760 ;
        RECT 125.800 77.900 126.120 77.960 ;
        RECT 126.275 77.900 126.565 77.945 ;
        RECT 130.490 77.900 130.630 78.040 ;
        RECT 125.800 77.760 126.565 77.900 ;
        RECT 125.800 77.700 126.120 77.760 ;
        RECT 126.275 77.715 126.565 77.760 ;
        RECT 130.030 77.760 130.630 77.900 ;
        RECT 135.015 77.900 135.305 77.945 ;
        RECT 135.015 77.760 137.070 77.900 ;
        RECT 130.030 77.605 130.170 77.760 ;
        RECT 135.015 77.715 135.305 77.760 ;
        RECT 136.930 77.620 137.070 77.760 ;
        RECT 119.375 77.560 119.665 77.605 ;
        RECT 118.440 77.420 119.665 77.560 ;
        RECT 116.600 77.360 116.920 77.375 ;
        RECT 118.440 77.360 118.760 77.420 ;
        RECT 119.375 77.375 119.665 77.420 ;
        RECT 129.915 77.375 130.205 77.605 ;
        RECT 131.335 77.375 131.625 77.605 ;
        RECT 136.395 77.375 136.685 77.605 ;
        RECT 99.595 77.220 99.885 77.265 ;
        RECT 101.435 77.220 101.725 77.265 ;
        RECT 87.710 77.080 93.830 77.220 ;
        RECT 81.195 76.880 81.485 76.925 ;
        RECT 80.810 76.740 81.485 76.880 ;
        RECT 71.535 76.695 71.825 76.740 ;
        RECT 72.910 76.695 73.200 76.740 ;
        RECT 81.195 76.695 81.485 76.740 ;
        RECT 46.695 76.400 47.460 76.540 ;
        RECT 46.695 76.355 46.985 76.400 ;
        RECT 47.140 76.340 47.460 76.400 ;
        RECT 49.915 76.355 50.205 76.585 ;
        RECT 54.960 76.540 55.280 76.600 ;
        RECT 55.435 76.540 55.725 76.585 ;
        RECT 54.960 76.400 55.725 76.540 ;
        RECT 54.960 76.340 55.280 76.400 ;
        RECT 55.435 76.355 55.725 76.400 ;
        RECT 65.540 76.340 65.860 76.600 ;
        RECT 67.855 76.540 68.145 76.585 ;
        RECT 68.300 76.540 68.620 76.600 ;
        RECT 67.855 76.400 68.620 76.540 ;
        RECT 67.855 76.355 68.145 76.400 ;
        RECT 68.300 76.340 68.620 76.400 ;
        RECT 74.740 76.340 75.060 76.600 ;
        RECT 81.270 76.540 81.410 76.695 ;
        RECT 85.320 76.680 85.640 76.940 ;
        RECT 83.940 76.540 84.260 76.600 ;
        RECT 85.780 76.540 86.100 76.600 ;
        RECT 86.330 76.540 86.470 77.035 ;
        RECT 81.270 76.400 86.470 76.540 ;
        RECT 89.475 76.540 89.765 76.585 ;
        RECT 91.300 76.540 91.620 76.600 ;
        RECT 93.690 76.585 93.830 77.080 ;
        RECT 99.595 77.080 101.725 77.220 ;
        RECT 99.595 77.035 99.885 77.080 ;
        RECT 101.435 77.035 101.725 77.080 ;
        RECT 101.900 77.220 102.190 77.265 ;
        RECT 104.240 77.220 104.530 77.265 ;
        RECT 101.900 77.080 104.530 77.220 ;
        RECT 101.900 77.035 102.190 77.080 ;
        RECT 104.240 77.035 104.530 77.080 ;
        RECT 109.240 77.020 109.560 77.280 ;
        RECT 113.405 77.220 113.695 77.265 ;
        RECT 115.925 77.220 116.215 77.265 ;
        RECT 117.115 77.220 117.405 77.265 ;
        RECT 113.405 77.080 117.405 77.220 ;
        RECT 113.405 77.035 113.695 77.080 ;
        RECT 115.925 77.035 116.215 77.080 ;
        RECT 117.115 77.035 117.405 77.080 ;
        RECT 117.995 77.035 118.285 77.265 ;
        RECT 131.410 77.220 131.550 77.375 ;
        RECT 128.190 77.080 131.550 77.220 ;
        RECT 132.700 77.220 133.020 77.280 ;
        RECT 135.475 77.220 135.765 77.265 ;
        RECT 132.700 77.080 135.765 77.220 ;
        RECT 102.360 76.880 102.650 76.925 ;
        RECT 103.735 76.880 104.025 76.925 ;
        RECT 102.360 76.740 104.025 76.880 ;
        RECT 102.360 76.695 102.650 76.740 ;
        RECT 103.735 76.695 104.025 76.740 ;
        RECT 106.495 76.880 106.785 76.925 ;
        RECT 110.620 76.880 110.940 76.940 ;
        RECT 106.495 76.740 110.940 76.880 ;
        RECT 106.495 76.695 106.785 76.740 ;
        RECT 110.620 76.680 110.940 76.740 ;
        RECT 113.840 76.880 114.130 76.925 ;
        RECT 115.410 76.880 115.700 76.925 ;
        RECT 117.510 76.880 117.800 76.925 ;
        RECT 113.840 76.740 117.800 76.880 ;
        RECT 113.840 76.695 114.130 76.740 ;
        RECT 115.410 76.695 115.700 76.740 ;
        RECT 117.510 76.695 117.800 76.740 ;
        RECT 89.475 76.400 91.620 76.540 ;
        RECT 83.940 76.340 84.260 76.400 ;
        RECT 85.780 76.340 86.100 76.400 ;
        RECT 89.475 76.355 89.765 76.400 ;
        RECT 91.300 76.340 91.620 76.400 ;
        RECT 93.615 76.355 93.905 76.585 ;
        RECT 111.080 76.340 111.400 76.600 ;
        RECT 117.060 76.540 117.380 76.600 ;
        RECT 118.070 76.540 118.210 77.035 ;
        RECT 119.835 76.880 120.125 76.925 ;
        RECT 122.120 76.880 122.440 76.940 ;
        RECT 128.190 76.925 128.330 77.080 ;
        RECT 132.700 77.020 133.020 77.080 ;
        RECT 135.475 77.035 135.765 77.080 ;
        RECT 119.835 76.740 127.870 76.880 ;
        RECT 119.835 76.695 120.125 76.740 ;
        RECT 122.120 76.680 122.440 76.740 ;
        RECT 117.060 76.400 118.210 76.540 ;
        RECT 126.720 76.540 127.040 76.600 ;
        RECT 127.195 76.540 127.485 76.585 ;
        RECT 126.720 76.400 127.485 76.540 ;
        RECT 127.730 76.540 127.870 76.740 ;
        RECT 128.115 76.695 128.405 76.925 ;
        RECT 136.470 76.880 136.610 77.375 ;
        RECT 136.840 77.360 137.160 77.620 ;
        RECT 137.390 77.560 137.530 78.055 ;
        RECT 138.695 77.560 138.985 77.605 ;
        RECT 137.390 77.420 138.985 77.560 ;
        RECT 139.690 77.560 139.830 78.055 ;
        RECT 145.120 78.040 145.440 78.300 ;
        RECT 148.800 78.240 149.120 78.300 ;
        RECT 145.670 78.100 149.120 78.240 ;
        RECT 145.670 77.605 145.810 78.100 ;
        RECT 148.800 78.040 149.120 78.100 ;
        RECT 150.640 78.040 150.960 78.300 ;
        RECT 153.035 78.240 153.325 78.285 ;
        RECT 151.190 78.100 153.325 78.240 ;
        RECT 146.975 77.900 147.265 77.945 ;
        RECT 151.190 77.900 151.330 78.100 ;
        RECT 153.035 78.055 153.325 78.100 ;
        RECT 153.875 78.055 154.165 78.285 ;
        RECT 146.975 77.760 151.330 77.900 ;
        RECT 146.975 77.715 147.265 77.760 ;
        RECT 152.020 77.700 152.340 77.960 ;
        RECT 141.455 77.560 141.745 77.605 ;
        RECT 139.690 77.420 141.745 77.560 ;
        RECT 138.695 77.375 138.985 77.420 ;
        RECT 141.455 77.375 141.745 77.420 ;
        RECT 145.595 77.375 145.885 77.605 ;
        RECT 147.435 77.560 147.725 77.605 ;
        RECT 147.880 77.560 148.200 77.620 ;
        RECT 147.050 77.420 148.200 77.560 ;
        RECT 147.050 77.265 147.190 77.420 ;
        RECT 147.435 77.375 147.725 77.420 ;
        RECT 147.880 77.360 148.200 77.420 ;
        RECT 148.355 77.560 148.645 77.605 ;
        RECT 148.800 77.560 149.120 77.620 ;
        RECT 148.355 77.420 149.120 77.560 ;
        RECT 148.355 77.375 148.645 77.420 ;
        RECT 148.800 77.360 149.120 77.420 ;
        RECT 149.735 77.560 150.025 77.605 ;
        RECT 150.180 77.560 150.500 77.620 ;
        RECT 149.735 77.420 150.500 77.560 ;
        RECT 153.950 77.560 154.090 78.055 ;
        RECT 155.255 77.560 155.545 77.605 ;
        RECT 153.950 77.420 155.545 77.560 ;
        RECT 149.735 77.375 150.025 77.420 ;
        RECT 140.075 77.035 140.365 77.265 ;
        RECT 140.540 77.220 140.830 77.265 ;
        RECT 142.880 77.220 143.170 77.265 ;
        RECT 140.540 77.080 143.170 77.220 ;
        RECT 140.540 77.035 140.830 77.080 ;
        RECT 142.880 77.035 143.170 77.080 ;
        RECT 146.975 77.035 147.265 77.265 ;
        RECT 130.260 76.740 136.610 76.880 ;
        RECT 130.260 76.540 130.400 76.740 ;
        RECT 127.730 76.400 130.400 76.540 ;
        RECT 130.875 76.540 131.165 76.585 ;
        RECT 131.320 76.540 131.640 76.600 ;
        RECT 130.875 76.400 131.640 76.540 ;
        RECT 117.060 76.340 117.380 76.400 ;
        RECT 126.720 76.340 127.040 76.400 ;
        RECT 127.195 76.355 127.485 76.400 ;
        RECT 130.875 76.355 131.165 76.400 ;
        RECT 131.320 76.340 131.640 76.400 ;
        RECT 132.240 76.340 132.560 76.600 ;
        RECT 135.460 76.340 135.780 76.600 ;
        RECT 140.150 76.540 140.290 77.035 ;
        RECT 141.000 76.880 141.290 76.925 ;
        RECT 142.375 76.880 142.665 76.925 ;
        RECT 141.000 76.740 142.665 76.880 ;
        RECT 141.000 76.695 141.290 76.740 ;
        RECT 142.375 76.695 142.665 76.740 ;
        RECT 146.055 76.880 146.345 76.925 ;
        RECT 147.420 76.880 147.740 76.940 ;
        RECT 149.810 76.880 149.950 77.375 ;
        RECT 150.180 77.360 150.500 77.420 ;
        RECT 155.255 77.375 155.545 77.420 ;
        RECT 153.860 77.020 154.180 77.280 ;
        RECT 146.055 76.740 149.950 76.880 ;
        RECT 146.055 76.695 146.345 76.740 ;
        RECT 147.420 76.680 147.740 76.740 ;
        RECT 141.440 76.540 141.760 76.600 ;
        RECT 140.150 76.400 141.760 76.540 ;
        RECT 141.440 76.340 141.760 76.400 ;
        RECT 152.955 76.540 153.245 76.585 ;
        RECT 153.950 76.540 154.090 77.020 ;
        RECT 152.955 76.400 154.090 76.540 ;
        RECT 152.955 76.355 153.245 76.400 ;
        RECT 154.320 76.340 154.640 76.600 ;
        RECT 22.690 75.720 157.010 76.200 ;
        RECT 41.160 75.520 41.480 75.580 ;
        RECT 37.570 75.380 41.480 75.520 ;
        RECT 35.180 75.180 35.500 75.240 ;
        RECT 37.020 75.180 37.340 75.240 ;
        RECT 37.570 75.225 37.710 75.380 ;
        RECT 41.160 75.320 41.480 75.380 ;
        RECT 42.080 75.320 42.400 75.580 ;
        RECT 43.015 75.520 43.305 75.565 ;
        RECT 44.380 75.520 44.700 75.580 ;
        RECT 43.015 75.380 44.700 75.520 ;
        RECT 43.015 75.335 43.305 75.380 ;
        RECT 44.380 75.320 44.700 75.380 ;
        RECT 51.295 75.335 51.585 75.565 ;
        RECT 51.740 75.520 52.060 75.580 ;
        RECT 52.675 75.520 52.965 75.565 ;
        RECT 51.740 75.380 52.965 75.520 ;
        RECT 37.495 75.180 37.785 75.225 ;
        RECT 42.170 75.180 42.310 75.320 ;
        RECT 44.840 75.180 45.160 75.240 ;
        RECT 35.180 75.040 37.785 75.180 ;
        RECT 35.180 74.980 35.500 75.040 ;
        RECT 37.020 74.980 37.340 75.040 ;
        RECT 37.495 74.995 37.785 75.040 ;
        RECT 38.030 75.040 45.160 75.180 ;
        RECT 51.370 75.180 51.510 75.335 ;
        RECT 51.740 75.320 52.060 75.380 ;
        RECT 52.675 75.335 52.965 75.380 ;
        RECT 60.020 75.320 60.340 75.580 ;
        RECT 62.320 75.520 62.640 75.580 ;
        RECT 62.795 75.520 63.085 75.565 ;
        RECT 62.320 75.380 63.085 75.520 ;
        RECT 62.320 75.320 62.640 75.380 ;
        RECT 62.795 75.335 63.085 75.380 ;
        RECT 64.635 75.520 64.925 75.565 ;
        RECT 65.540 75.520 65.860 75.580 ;
        RECT 64.635 75.380 65.860 75.520 ;
        RECT 64.635 75.335 64.925 75.380 ;
        RECT 65.540 75.320 65.860 75.380 ;
        RECT 85.320 75.320 85.640 75.580 ;
        RECT 107.415 75.520 107.705 75.565 ;
        RECT 108.320 75.520 108.640 75.580 ;
        RECT 110.175 75.520 110.465 75.565 ;
        RECT 107.415 75.380 110.465 75.520 ;
        RECT 107.415 75.335 107.705 75.380 ;
        RECT 108.320 75.320 108.640 75.380 ;
        RECT 110.175 75.335 110.465 75.380 ;
        RECT 112.015 75.520 112.305 75.565 ;
        RECT 114.315 75.520 114.605 75.565 ;
        RECT 112.015 75.380 114.605 75.520 ;
        RECT 112.015 75.335 112.305 75.380 ;
        RECT 114.315 75.335 114.605 75.380 ;
        RECT 116.600 75.320 116.920 75.580 ;
        RECT 132.700 75.520 133.020 75.580 ;
        RECT 126.350 75.380 133.020 75.520 ;
        RECT 52.200 75.180 52.520 75.240 ;
        RECT 51.370 75.040 52.520 75.180 ;
        RECT 36.115 74.840 36.405 74.885 ;
        RECT 36.560 74.840 36.880 74.900 ;
        RECT 38.030 74.840 38.170 75.040 ;
        RECT 44.840 74.980 45.160 75.040 ;
        RECT 52.200 74.980 52.520 75.040 ;
        RECT 55.900 75.180 56.190 75.225 ;
        RECT 57.275 75.180 57.565 75.225 ;
        RECT 55.900 75.040 57.565 75.180 ;
        RECT 55.900 74.995 56.190 75.040 ;
        RECT 57.275 74.995 57.565 75.040 ;
        RECT 68.300 75.180 68.590 75.225 ;
        RECT 69.870 75.180 70.160 75.225 ;
        RECT 71.970 75.180 72.260 75.225 ;
        RECT 68.300 75.040 72.260 75.180 ;
        RECT 68.300 74.995 68.590 75.040 ;
        RECT 69.870 74.995 70.160 75.040 ;
        RECT 71.970 74.995 72.260 75.040 ;
        RECT 73.375 75.180 73.665 75.225 ;
        RECT 74.280 75.180 74.600 75.240 ;
        RECT 94.980 75.180 95.300 75.240 ;
        RECT 73.375 75.040 95.300 75.180 ;
        RECT 73.375 74.995 73.665 75.040 ;
        RECT 74.280 74.980 74.600 75.040 ;
        RECT 94.980 74.980 95.300 75.040 ;
        RECT 101.440 75.180 101.730 75.225 ;
        RECT 102.815 75.180 103.105 75.225 ;
        RECT 101.440 75.040 103.105 75.180 ;
        RECT 101.440 74.995 101.730 75.040 ;
        RECT 102.815 74.995 103.105 75.040 ;
        RECT 111.080 74.980 111.400 75.240 ;
        RECT 122.135 75.180 122.425 75.225 ;
        RECT 125.800 75.180 126.120 75.240 ;
        RECT 122.135 75.040 126.120 75.180 ;
        RECT 122.135 74.995 122.425 75.040 ;
        RECT 36.115 74.700 38.170 74.840 ;
        RECT 38.415 74.840 38.705 74.885 ;
        RECT 50.835 74.840 51.125 74.885 ;
        RECT 38.415 74.700 51.125 74.840 ;
        RECT 36.115 74.655 36.405 74.700 ;
        RECT 36.560 74.640 36.880 74.700 ;
        RECT 38.415 74.655 38.705 74.700 ;
        RECT 30.135 74.500 30.425 74.545 ;
        RECT 31.040 74.500 31.360 74.560 ;
        RECT 31.975 74.500 32.265 74.545 ;
        RECT 30.135 74.360 32.265 74.500 ;
        RECT 30.135 74.315 30.425 74.360 ;
        RECT 31.040 74.300 31.360 74.360 ;
        RECT 31.975 74.315 32.265 74.360 ;
        RECT 32.880 74.300 33.200 74.560 ;
        RECT 37.480 74.500 37.800 74.560 ;
        RECT 39.870 74.545 40.010 74.700 ;
        RECT 38.875 74.500 39.165 74.545 ;
        RECT 37.480 74.360 39.165 74.500 ;
        RECT 37.480 74.300 37.800 74.360 ;
        RECT 38.875 74.315 39.165 74.360 ;
        RECT 39.795 74.315 40.085 74.545 ;
        RECT 40.700 74.500 41.020 74.560 ;
        RECT 40.700 74.360 41.850 74.500 ;
        RECT 40.700 74.300 41.020 74.360 ;
        RECT 41.710 74.220 41.850 74.360 ;
        RECT 43.920 74.300 44.240 74.560 ;
        RECT 44.380 74.500 44.700 74.560 ;
        RECT 46.770 74.545 46.910 74.700 ;
        RECT 50.835 74.655 51.125 74.700 ;
        RECT 55.440 74.840 55.730 74.885 ;
        RECT 57.780 74.840 58.070 74.885 ;
        RECT 55.440 74.700 58.070 74.840 ;
        RECT 55.440 74.655 55.730 74.700 ;
        RECT 57.780 74.655 58.070 74.700 ;
        RECT 67.865 74.840 68.155 74.885 ;
        RECT 70.385 74.840 70.675 74.885 ;
        RECT 71.575 74.840 71.865 74.885 ;
        RECT 74.740 74.840 75.060 74.900 ;
        RECT 67.865 74.700 71.865 74.840 ;
        RECT 67.865 74.655 68.155 74.700 ;
        RECT 70.385 74.655 70.675 74.700 ;
        RECT 71.575 74.655 71.865 74.700 ;
        RECT 72.990 74.700 75.060 74.840 ;
        RECT 72.990 74.560 73.130 74.700 ;
        RECT 74.740 74.640 75.060 74.700 ;
        RECT 100.980 74.840 101.270 74.885 ;
        RECT 103.320 74.840 103.610 74.885 ;
        RECT 107.875 74.840 108.165 74.885 ;
        RECT 111.170 74.840 111.310 74.980 ;
        RECT 122.210 74.840 122.350 74.995 ;
        RECT 125.800 74.980 126.120 75.040 ;
        RECT 100.980 74.700 103.610 74.840 ;
        RECT 100.980 74.655 101.270 74.700 ;
        RECT 103.320 74.655 103.610 74.700 ;
        RECT 106.570 74.700 108.165 74.840 ;
        RECT 45.315 74.500 45.605 74.545 ;
        RECT 44.380 74.360 45.605 74.500 ;
        RECT 44.380 74.300 44.700 74.360 ;
        RECT 45.315 74.315 45.605 74.360 ;
        RECT 46.695 74.315 46.985 74.545 ;
        RECT 47.140 74.500 47.460 74.560 ;
        RECT 48.075 74.500 48.365 74.545 ;
        RECT 48.980 74.500 49.300 74.560 ;
        RECT 51.755 74.500 52.045 74.545 ;
        RECT 47.140 74.360 49.300 74.500 ;
        RECT 47.140 74.300 47.460 74.360 ;
        RECT 48.075 74.315 48.365 74.360 ;
        RECT 48.980 74.300 49.300 74.360 ;
        RECT 49.530 74.360 52.045 74.500 ;
        RECT 31.500 74.160 31.820 74.220 ;
        RECT 33.800 74.160 34.120 74.220 ;
        RECT 40.240 74.160 40.560 74.220 ;
        RECT 31.500 74.020 40.560 74.160 ;
        RECT 31.500 73.960 31.820 74.020 ;
        RECT 33.800 73.960 34.120 74.020 ;
        RECT 40.240 73.960 40.560 74.020 ;
        RECT 41.160 73.960 41.480 74.220 ;
        RECT 41.620 74.160 41.940 74.220 ;
        RECT 42.175 74.160 42.465 74.205 ;
        RECT 49.530 74.160 49.670 74.360 ;
        RECT 51.755 74.315 52.045 74.360 ;
        RECT 53.580 74.300 53.900 74.560 ;
        RECT 54.960 74.300 55.280 74.560 ;
        RECT 56.355 74.315 56.645 74.545 ;
        RECT 41.620 74.020 42.465 74.160 ;
        RECT 41.620 73.960 41.940 74.020 ;
        RECT 42.175 73.975 42.465 74.020 ;
        RECT 42.630 74.020 49.670 74.160 ;
        RECT 50.375 74.160 50.665 74.205 ;
        RECT 50.820 74.160 51.140 74.220 ;
        RECT 56.430 74.160 56.570 74.315 ;
        RECT 62.780 74.300 63.100 74.560 ;
        RECT 63.715 74.500 64.005 74.545 ;
        RECT 64.160 74.500 64.480 74.560 ;
        RECT 65.540 74.500 65.860 74.560 ;
        RECT 63.715 74.360 65.860 74.500 ;
        RECT 63.715 74.315 64.005 74.360 ;
        RECT 64.160 74.300 64.480 74.360 ;
        RECT 65.540 74.300 65.860 74.360 ;
        RECT 68.300 74.500 68.620 74.560 ;
        RECT 71.120 74.500 71.410 74.545 ;
        RECT 68.300 74.360 71.410 74.500 ;
        RECT 68.300 74.300 68.620 74.360 ;
        RECT 71.120 74.315 71.410 74.360 ;
        RECT 72.455 74.315 72.745 74.545 ;
        RECT 50.375 74.020 51.140 74.160 ;
        RECT 30.580 73.820 30.900 73.880 ;
        RECT 42.630 73.820 42.770 74.020 ;
        RECT 50.375 73.975 50.665 74.020 ;
        RECT 50.820 73.960 51.140 74.020 ;
        RECT 54.590 74.020 56.570 74.160 ;
        RECT 69.680 74.160 70.000 74.220 ;
        RECT 71.520 74.160 71.840 74.220 ;
        RECT 72.530 74.160 72.670 74.315 ;
        RECT 72.900 74.300 73.220 74.560 ;
        RECT 78.435 74.500 78.725 74.545 ;
        RECT 78.880 74.500 79.200 74.560 ;
        RECT 78.435 74.360 79.200 74.500 ;
        RECT 78.435 74.315 78.725 74.360 ;
        RECT 78.880 74.300 79.200 74.360 ;
        RECT 79.355 74.500 79.645 74.545 ;
        RECT 80.260 74.500 80.580 74.560 ;
        RECT 86.700 74.500 87.020 74.560 ;
        RECT 79.355 74.360 80.580 74.500 ;
        RECT 79.355 74.315 79.645 74.360 ;
        RECT 80.260 74.300 80.580 74.360 ;
        RECT 84.490 74.360 87.020 74.500 ;
        RECT 69.680 74.020 72.670 74.160 ;
        RECT 78.970 74.160 79.110 74.300 ;
        RECT 84.490 74.205 84.630 74.360 ;
        RECT 86.700 74.300 87.020 74.360 ;
        RECT 87.160 74.500 87.480 74.560 ;
        RECT 87.635 74.500 87.925 74.545 ;
        RECT 87.160 74.360 87.925 74.500 ;
        RECT 87.160 74.300 87.480 74.360 ;
        RECT 87.635 74.315 87.925 74.360 ;
        RECT 89.475 74.315 89.765 74.545 ;
        RECT 85.780 74.205 86.100 74.220 ;
        RECT 84.415 74.160 84.705 74.205 ;
        RECT 78.970 74.020 84.705 74.160 ;
        RECT 30.580 73.680 42.770 73.820 ;
        RECT 30.580 73.620 30.900 73.680 ;
        RECT 44.380 73.620 44.700 73.880 ;
        RECT 46.220 73.620 46.540 73.880 ;
        RECT 47.140 73.620 47.460 73.880 ;
        RECT 48.995 73.820 49.285 73.865 ;
        RECT 49.900 73.820 50.220 73.880 ;
        RECT 53.120 73.820 53.440 73.880 ;
        RECT 54.590 73.865 54.730 74.020 ;
        RECT 69.680 73.960 70.000 74.020 ;
        RECT 71.520 73.960 71.840 74.020 ;
        RECT 84.415 73.975 84.705 74.020 ;
        RECT 85.495 73.975 86.100 74.205 ;
        RECT 89.550 74.160 89.690 74.315 ;
        RECT 96.360 74.300 96.680 74.560 ;
        RECT 97.740 74.300 98.060 74.560 ;
        RECT 100.055 74.500 100.345 74.545 ;
        RECT 100.515 74.500 100.805 74.545 ;
        RECT 100.055 74.360 100.805 74.500 ;
        RECT 100.055 74.315 100.345 74.360 ;
        RECT 100.515 74.315 100.805 74.360 ;
        RECT 101.895 74.315 102.185 74.545 ;
        RECT 101.970 74.160 102.110 74.315 ;
        RECT 102.800 74.300 103.120 74.560 ;
        RECT 106.570 74.545 106.710 74.700 ;
        RECT 107.875 74.655 108.165 74.700 ;
        RECT 108.870 74.700 111.310 74.840 ;
        RECT 118.530 74.700 122.350 74.840 ;
        RECT 122.595 74.840 122.885 74.885 ;
        RECT 126.350 74.840 126.490 75.380 ;
        RECT 132.700 75.320 133.020 75.380 ;
        RECT 134.540 75.320 134.860 75.580 ;
        RECT 135.920 75.320 136.240 75.580 ;
        RECT 146.975 75.520 147.265 75.565 ;
        RECT 147.420 75.520 147.740 75.580 ;
        RECT 146.975 75.380 147.740 75.520 ;
        RECT 146.975 75.335 147.265 75.380 ;
        RECT 147.420 75.320 147.740 75.380 ;
        RECT 151.560 75.520 151.880 75.580 ;
        RECT 151.560 75.380 155.470 75.520 ;
        RECT 151.560 75.320 151.880 75.380 ;
        RECT 126.720 75.180 127.040 75.240 ;
        RECT 131.320 75.180 131.640 75.240 ;
        RECT 133.160 75.180 133.480 75.240 ;
        RECT 126.720 75.040 127.410 75.180 ;
        RECT 126.720 74.980 127.040 75.040 ;
        RECT 122.595 74.700 126.490 74.840 ;
        RECT 108.870 74.545 109.010 74.700 ;
        RECT 106.495 74.500 106.785 74.545 ;
        RECT 105.650 74.360 106.785 74.500 ;
        RECT 85.780 73.960 86.100 73.975 ;
        RECT 86.330 74.020 89.690 74.160 ;
        RECT 97.370 74.020 102.110 74.160 ;
        RECT 48.995 73.680 53.440 73.820 ;
        RECT 48.995 73.635 49.285 73.680 ;
        RECT 49.900 73.620 50.220 73.680 ;
        RECT 53.120 73.620 53.440 73.680 ;
        RECT 54.515 73.635 54.805 73.865 ;
        RECT 61.400 73.820 61.720 73.880 ;
        RECT 65.555 73.820 65.845 73.865 ;
        RECT 61.400 73.680 65.845 73.820 ;
        RECT 61.400 73.620 61.720 73.680 ;
        RECT 65.555 73.635 65.845 73.680 ;
        RECT 75.200 73.820 75.520 73.880 ;
        RECT 78.895 73.820 79.185 73.865 ;
        RECT 84.860 73.820 85.180 73.880 ;
        RECT 86.330 73.865 86.470 74.020 ;
        RECT 75.200 73.680 85.180 73.820 ;
        RECT 75.200 73.620 75.520 73.680 ;
        RECT 78.895 73.635 79.185 73.680 ;
        RECT 84.860 73.620 85.180 73.680 ;
        RECT 86.255 73.635 86.545 73.865 ;
        RECT 88.080 73.620 88.400 73.880 ;
        RECT 90.395 73.820 90.685 73.865 ;
        RECT 96.820 73.820 97.140 73.880 ;
        RECT 97.370 73.865 97.510 74.020 ;
        RECT 90.395 73.680 97.140 73.820 ;
        RECT 90.395 73.635 90.685 73.680 ;
        RECT 96.820 73.620 97.140 73.680 ;
        RECT 97.295 73.635 97.585 73.865 ;
        RECT 98.675 73.820 98.965 73.865 ;
        RECT 102.890 73.820 103.030 74.300 ;
        RECT 105.650 73.865 105.790 74.360 ;
        RECT 106.495 74.315 106.785 74.360 ;
        RECT 107.415 74.500 107.705 74.545 ;
        RECT 108.795 74.500 109.085 74.545 ;
        RECT 107.415 74.360 109.085 74.500 ;
        RECT 107.415 74.315 107.705 74.360 ;
        RECT 108.795 74.315 109.085 74.360 ;
        RECT 109.240 74.500 109.560 74.560 ;
        RECT 118.530 74.545 118.670 74.700 ;
        RECT 122.595 74.655 122.885 74.700 ;
        RECT 110.175 74.500 110.465 74.545 ;
        RECT 109.240 74.360 110.465 74.500 ;
        RECT 109.240 74.300 109.560 74.360 ;
        RECT 110.175 74.315 110.465 74.360 ;
        RECT 110.635 74.315 110.925 74.545 ;
        RECT 115.695 74.500 115.985 74.545 ;
        RECT 115.310 74.360 115.985 74.500 ;
        RECT 107.860 74.160 108.180 74.220 ;
        RECT 110.710 74.160 110.850 74.315 ;
        RECT 107.860 74.020 110.850 74.160 ;
        RECT 107.860 73.960 108.180 74.020 ;
        RECT 113.380 73.960 113.700 74.220 ;
        RECT 98.675 73.680 103.030 73.820 ;
        RECT 98.675 73.635 98.965 73.680 ;
        RECT 105.575 73.635 105.865 73.865 ;
        RECT 109.240 73.820 109.560 73.880 ;
        RECT 109.715 73.820 110.005 73.865 ;
        RECT 109.240 73.680 110.005 73.820 ;
        RECT 109.240 73.620 109.560 73.680 ;
        RECT 109.715 73.635 110.005 73.680 ;
        RECT 110.160 73.820 110.480 73.880 ;
        RECT 115.310 73.865 115.450 74.360 ;
        RECT 115.695 74.315 115.985 74.360 ;
        RECT 118.455 74.315 118.745 74.545 ;
        RECT 119.375 74.500 119.665 74.545 ;
        RECT 119.820 74.500 120.140 74.560 ;
        RECT 120.295 74.500 120.585 74.545 ;
        RECT 119.375 74.360 120.585 74.500 ;
        RECT 119.375 74.315 119.665 74.360 ;
        RECT 119.820 74.300 120.140 74.360 ;
        RECT 120.295 74.315 120.585 74.360 ;
        RECT 121.200 74.500 121.520 74.560 ;
        RECT 124.050 74.545 124.190 74.700 ;
        RECT 123.055 74.500 123.345 74.545 ;
        RECT 121.200 74.360 123.345 74.500 ;
        RECT 121.200 74.300 121.520 74.360 ;
        RECT 123.055 74.315 123.345 74.360 ;
        RECT 123.975 74.315 124.265 74.545 ;
        RECT 124.420 74.300 124.740 74.560 ;
        RECT 125.800 74.500 126.120 74.560 ;
        RECT 127.270 74.545 127.410 75.040 ;
        RECT 130.490 75.040 133.480 75.180 ;
        RECT 128.115 74.840 128.405 74.885 ;
        RECT 128.115 74.700 130.170 74.840 ;
        RECT 128.115 74.655 128.405 74.700 ;
        RECT 126.425 74.500 126.715 74.545 ;
        RECT 125.800 74.360 126.715 74.500 ;
        RECT 125.800 74.300 126.120 74.360 ;
        RECT 126.425 74.315 126.715 74.360 ;
        RECT 127.195 74.315 127.485 74.545 ;
        RECT 127.655 74.315 127.945 74.545 ;
        RECT 128.575 74.315 128.865 74.545 ;
        RECT 127.730 74.160 127.870 74.315 ;
        RECT 125.890 74.020 127.870 74.160 ;
        RECT 125.890 73.880 126.030 74.020 ;
        RECT 114.395 73.820 114.685 73.865 ;
        RECT 110.160 73.680 114.685 73.820 ;
        RECT 110.160 73.620 110.480 73.680 ;
        RECT 114.395 73.635 114.685 73.680 ;
        RECT 115.235 73.635 115.525 73.865 ;
        RECT 118.900 73.620 119.220 73.880 ;
        RECT 125.355 73.820 125.645 73.865 ;
        RECT 125.800 73.820 126.120 73.880 ;
        RECT 125.355 73.680 126.120 73.820 ;
        RECT 125.355 73.635 125.645 73.680 ;
        RECT 125.800 73.620 126.120 73.680 ;
        RECT 127.180 73.820 127.500 73.880 ;
        RECT 128.650 73.820 128.790 74.315 ;
        RECT 129.020 74.300 129.340 74.560 ;
        RECT 130.030 74.220 130.170 74.700 ;
        RECT 130.490 74.545 130.630 75.040 ;
        RECT 131.320 74.980 131.640 75.040 ;
        RECT 133.160 74.980 133.480 75.040 ;
        RECT 140.540 75.180 140.830 75.225 ;
        RECT 141.915 75.180 142.205 75.225 ;
        RECT 140.540 75.040 142.205 75.180 ;
        RECT 140.540 74.995 140.830 75.040 ;
        RECT 141.915 74.995 142.205 75.040 ;
        RECT 151.100 75.180 151.390 75.225 ;
        RECT 152.670 75.180 152.960 75.225 ;
        RECT 154.770 75.180 155.060 75.225 ;
        RECT 151.100 75.040 155.060 75.180 ;
        RECT 151.100 74.995 151.390 75.040 ;
        RECT 152.670 74.995 152.960 75.040 ;
        RECT 154.770 74.995 155.060 75.040 ;
        RECT 135.475 74.840 135.765 74.885 ;
        RECT 131.870 74.700 135.765 74.840 ;
        RECT 130.415 74.315 130.705 74.545 ;
        RECT 131.870 74.500 132.010 74.700 ;
        RECT 135.475 74.655 135.765 74.700 ;
        RECT 138.680 74.840 139.000 74.900 ;
        RECT 139.615 74.840 139.905 74.885 ;
        RECT 138.680 74.700 139.905 74.840 ;
        RECT 138.680 74.640 139.000 74.700 ;
        RECT 139.615 74.655 139.905 74.700 ;
        RECT 140.080 74.840 140.370 74.885 ;
        RECT 142.420 74.840 142.710 74.885 ;
        RECT 140.080 74.700 142.710 74.840 ;
        RECT 140.080 74.655 140.370 74.700 ;
        RECT 142.420 74.655 142.710 74.700 ;
        RECT 150.665 74.840 150.955 74.885 ;
        RECT 153.185 74.840 153.475 74.885 ;
        RECT 154.375 74.840 154.665 74.885 ;
        RECT 150.665 74.700 154.665 74.840 ;
        RECT 150.665 74.655 150.955 74.700 ;
        RECT 153.185 74.655 153.475 74.700 ;
        RECT 154.375 74.655 154.665 74.700 ;
        RECT 130.950 74.360 132.010 74.500 ;
        RECT 132.255 74.500 132.545 74.545 ;
        RECT 132.700 74.500 133.020 74.560 ;
        RECT 132.255 74.360 133.020 74.500 ;
        RECT 129.940 74.160 130.260 74.220 ;
        RECT 130.950 74.160 131.090 74.360 ;
        RECT 132.255 74.315 132.545 74.360 ;
        RECT 132.700 74.300 133.020 74.360 ;
        RECT 133.160 74.500 133.480 74.560 ;
        RECT 133.635 74.500 133.925 74.545 ;
        RECT 133.160 74.360 133.925 74.500 ;
        RECT 133.160 74.300 133.480 74.360 ;
        RECT 133.635 74.315 133.925 74.360 ;
        RECT 136.380 74.300 136.700 74.560 ;
        RECT 140.980 74.300 141.300 74.560 ;
        RECT 155.330 74.545 155.470 75.380 ;
        RECT 145.135 74.500 145.425 74.545 ;
        RECT 144.750 74.360 145.425 74.500 ;
        RECT 129.940 74.020 131.090 74.160 ;
        RECT 131.335 74.160 131.625 74.205 ;
        RECT 135.015 74.160 135.305 74.205 ;
        RECT 131.335 74.020 135.305 74.160 ;
        RECT 129.940 73.960 130.260 74.020 ;
        RECT 131.335 73.975 131.625 74.020 ;
        RECT 135.015 73.975 135.305 74.020 ;
        RECT 144.750 73.880 144.890 74.360 ;
        RECT 145.135 74.315 145.425 74.360 ;
        RECT 146.055 74.500 146.345 74.545 ;
        RECT 146.055 74.360 148.570 74.500 ;
        RECT 146.055 74.315 146.345 74.360 ;
        RECT 148.430 73.880 148.570 74.360 ;
        RECT 153.920 74.315 154.210 74.545 ;
        RECT 155.255 74.315 155.545 74.545 ;
        RECT 153.950 74.160 154.090 74.315 ;
        RECT 154.320 74.160 154.640 74.220 ;
        RECT 153.950 74.020 154.640 74.160 ;
        RECT 154.320 73.960 154.640 74.020 ;
        RECT 127.180 73.680 128.790 73.820 ;
        RECT 129.020 73.820 129.340 73.880 ;
        RECT 129.495 73.820 129.785 73.865 ;
        RECT 129.020 73.680 129.785 73.820 ;
        RECT 127.180 73.620 127.500 73.680 ;
        RECT 129.020 73.620 129.340 73.680 ;
        RECT 129.495 73.635 129.785 73.680 ;
        RECT 132.700 73.620 133.020 73.880 ;
        RECT 137.300 73.620 137.620 73.880 ;
        RECT 144.660 73.620 144.980 73.880 ;
        RECT 148.340 73.620 148.660 73.880 ;
        RECT 22.690 73.000 157.810 73.480 ;
        RECT 34.720 72.800 35.040 72.860 ;
        RECT 33.660 72.660 35.040 72.800 ;
        RECT 30.120 71.440 30.440 71.500 ;
        RECT 33.660 71.440 33.800 72.660 ;
        RECT 34.720 72.600 35.040 72.660 ;
        RECT 35.180 72.800 35.500 72.860 ;
        RECT 35.180 72.660 44.610 72.800 ;
        RECT 35.180 72.600 35.500 72.660 ;
        RECT 38.415 72.460 38.705 72.505 ;
        RECT 44.470 72.460 44.610 72.660 ;
        RECT 45.300 72.600 45.620 72.860 ;
        RECT 52.675 72.800 52.965 72.845 ;
        RECT 53.580 72.800 53.900 72.860 ;
        RECT 52.675 72.660 53.900 72.800 ;
        RECT 52.675 72.615 52.965 72.660 ;
        RECT 53.580 72.600 53.900 72.660 ;
        RECT 68.760 72.800 69.080 72.860 ;
        RECT 73.375 72.800 73.665 72.845 ;
        RECT 73.820 72.800 74.140 72.860 ;
        RECT 80.260 72.800 80.580 72.860 ;
        RECT 68.760 72.660 74.140 72.800 ;
        RECT 68.760 72.600 69.080 72.660 ;
        RECT 73.375 72.615 73.665 72.660 ;
        RECT 73.820 72.600 74.140 72.660 ;
        RECT 78.510 72.660 80.580 72.800 ;
        RECT 78.510 72.505 78.650 72.660 ;
        RECT 80.260 72.600 80.580 72.660 ;
        RECT 83.940 72.600 84.260 72.860 ;
        RECT 84.860 72.800 85.180 72.860 ;
        RECT 88.095 72.800 88.385 72.845 ;
        RECT 88.540 72.800 88.860 72.860 ;
        RECT 84.860 72.660 88.860 72.800 ;
        RECT 84.860 72.600 85.180 72.660 ;
        RECT 88.095 72.615 88.385 72.660 ;
        RECT 88.540 72.600 88.860 72.660 ;
        RECT 94.520 72.800 94.840 72.860 ;
        RECT 96.360 72.800 96.680 72.860 ;
        RECT 97.295 72.800 97.585 72.845 ;
        RECT 94.520 72.660 96.130 72.800 ;
        RECT 94.520 72.600 94.840 72.660 ;
        RECT 46.235 72.460 46.525 72.505 ;
        RECT 78.435 72.460 78.725 72.505 ;
        RECT 34.810 72.320 36.790 72.460 ;
        RECT 34.810 72.165 34.950 72.320 ;
        RECT 36.650 72.180 36.790 72.320 ;
        RECT 38.415 72.320 42.770 72.460 ;
        RECT 38.415 72.275 38.705 72.320 ;
        RECT 42.630 72.180 42.770 72.320 ;
        RECT 44.470 72.320 46.525 72.460 ;
        RECT 34.735 71.935 35.025 72.165 ;
        RECT 35.655 71.935 35.945 72.165 ;
        RECT 35.730 71.780 35.870 71.935 ;
        RECT 36.560 71.920 36.880 72.180 ;
        RECT 37.020 72.120 37.340 72.180 ;
        RECT 40.255 72.120 40.545 72.165 ;
        RECT 37.020 71.980 37.535 72.120 ;
        RECT 39.870 71.980 40.545 72.120 ;
        RECT 37.020 71.920 37.340 71.980 ;
        RECT 37.110 71.780 37.250 71.920 ;
        RECT 35.730 71.640 37.250 71.780 ;
        RECT 30.120 71.300 33.800 71.440 ;
        RECT 36.100 71.440 36.420 71.500 ;
        RECT 39.870 71.440 40.010 71.980 ;
        RECT 40.255 71.935 40.545 71.980 ;
        RECT 40.700 72.120 41.020 72.180 ;
        RECT 41.175 72.120 41.465 72.165 ;
        RECT 40.700 71.980 41.465 72.120 ;
        RECT 40.700 71.920 41.020 71.980 ;
        RECT 41.175 71.935 41.465 71.980 ;
        RECT 41.250 71.780 41.390 71.935 ;
        RECT 41.620 71.920 41.940 72.180 ;
        RECT 42.540 71.920 42.860 72.180 ;
        RECT 43.460 71.920 43.780 72.180 ;
        RECT 44.470 72.165 44.610 72.320 ;
        RECT 46.235 72.275 46.525 72.320 ;
        RECT 46.770 72.320 54.270 72.460 ;
        RECT 44.395 71.935 44.685 72.165 ;
        RECT 45.775 72.120 46.065 72.165 ;
        RECT 46.770 72.120 46.910 72.320 ;
        RECT 54.130 72.180 54.270 72.320 ;
        RECT 63.330 72.320 66.690 72.460 ;
        RECT 45.775 71.980 46.910 72.120 ;
        RECT 45.775 71.935 46.065 71.980 ;
        RECT 47.155 71.935 47.445 72.165 ;
        RECT 48.075 72.120 48.365 72.165 ;
        RECT 50.375 72.120 50.665 72.165 ;
        RECT 48.075 71.980 50.665 72.120 ;
        RECT 48.075 71.935 48.365 71.980 ;
        RECT 50.375 71.935 50.665 71.980 ;
        RECT 51.755 71.935 52.045 72.165 ;
        RECT 42.080 71.780 42.400 71.840 ;
        RECT 45.850 71.780 45.990 71.935 ;
        RECT 41.250 71.640 45.990 71.780 ;
        RECT 47.230 71.780 47.370 71.935 ;
        RECT 48.980 71.780 49.300 71.840 ;
        RECT 50.835 71.780 51.125 71.825 ;
        RECT 47.230 71.640 49.300 71.780 ;
        RECT 42.080 71.580 42.400 71.640 ;
        RECT 48.980 71.580 49.300 71.640 ;
        RECT 49.530 71.640 51.125 71.780 ;
        RECT 36.100 71.300 40.010 71.440 ;
        RECT 42.555 71.440 42.845 71.485 ;
        RECT 49.530 71.440 49.670 71.640 ;
        RECT 50.835 71.595 51.125 71.640 ;
        RECT 51.280 71.780 51.600 71.840 ;
        RECT 51.830 71.780 51.970 71.935 ;
        RECT 53.120 71.920 53.440 72.180 ;
        RECT 54.040 71.920 54.360 72.180 ;
        RECT 55.435 72.120 55.725 72.165 ;
        RECT 55.050 71.980 55.725 72.120 ;
        RECT 53.595 71.780 53.885 71.825 ;
        RECT 51.280 71.640 53.885 71.780 ;
        RECT 51.280 71.580 51.600 71.640 ;
        RECT 53.595 71.595 53.885 71.640 ;
        RECT 55.050 71.485 55.190 71.980 ;
        RECT 55.435 71.935 55.725 71.980 ;
        RECT 62.780 72.120 63.100 72.180 ;
        RECT 63.330 72.165 63.470 72.320 ;
        RECT 66.550 72.165 66.690 72.320 ;
        RECT 78.050 72.320 78.725 72.460 ;
        RECT 84.030 72.460 84.170 72.600 ;
        RECT 84.030 72.320 85.550 72.460 ;
        RECT 63.255 72.120 63.545 72.165 ;
        RECT 62.780 71.980 63.545 72.120 ;
        RECT 62.780 71.920 63.100 71.980 ;
        RECT 63.255 71.935 63.545 71.980 ;
        RECT 64.175 72.120 64.465 72.165 ;
        RECT 65.555 72.120 65.845 72.165 ;
        RECT 64.175 71.980 65.845 72.120 ;
        RECT 64.175 71.935 64.465 71.980 ;
        RECT 65.555 71.935 65.845 71.980 ;
        RECT 66.475 71.935 66.765 72.165 ;
        RECT 71.060 72.120 71.380 72.180 ;
        RECT 72.900 72.120 73.220 72.180 ;
        RECT 78.050 72.165 78.190 72.320 ;
        RECT 78.435 72.275 78.725 72.320 ;
        RECT 71.060 71.980 73.220 72.120 ;
        RECT 60.940 71.780 61.260 71.840 ;
        RECT 64.250 71.780 64.390 71.935 ;
        RECT 71.060 71.920 71.380 71.980 ;
        RECT 72.900 71.920 73.220 71.980 ;
        RECT 73.835 71.935 74.125 72.165 ;
        RECT 77.510 71.935 77.800 72.165 ;
        RECT 77.975 71.935 78.265 72.165 ;
        RECT 82.115 71.935 82.405 72.165 ;
        RECT 82.560 72.120 82.880 72.180 ;
        RECT 85.410 72.165 85.550 72.320 ;
        RECT 86.240 72.260 86.560 72.520 ;
        RECT 87.620 72.275 87.940 72.520 ;
        RECT 89.935 72.460 90.225 72.505 ;
        RECT 94.995 72.460 95.285 72.505 ;
        RECT 89.935 72.320 95.285 72.460 ;
        RECT 95.990 72.460 96.130 72.660 ;
        RECT 96.360 72.660 97.585 72.800 ;
        RECT 96.360 72.600 96.680 72.660 ;
        RECT 97.295 72.615 97.585 72.660 ;
        RECT 108.320 72.600 108.640 72.860 ;
        RECT 110.160 72.600 110.480 72.860 ;
        RECT 116.600 72.800 116.920 72.860 ;
        RECT 118.440 72.800 118.760 72.860 ;
        RECT 116.600 72.660 118.760 72.800 ;
        RECT 116.600 72.600 116.920 72.660 ;
        RECT 118.440 72.600 118.760 72.660 ;
        RECT 118.900 72.600 119.220 72.860 ;
        RECT 129.020 72.600 129.340 72.860 ;
        RECT 129.480 72.800 129.800 72.860 ;
        RECT 132.700 72.800 133.020 72.860 ;
        RECT 129.480 72.660 133.020 72.800 ;
        RECT 129.480 72.600 129.800 72.660 ;
        RECT 132.700 72.600 133.020 72.660 ;
        RECT 134.540 72.600 134.860 72.860 ;
        RECT 136.380 72.600 136.700 72.860 ;
        RECT 137.300 72.600 137.620 72.860 ;
        RECT 139.155 72.800 139.445 72.845 ;
        RECT 140.980 72.800 141.300 72.860 ;
        RECT 139.155 72.660 141.300 72.800 ;
        RECT 139.155 72.615 139.445 72.660 ;
        RECT 140.980 72.600 141.300 72.660 ;
        RECT 144.660 72.600 144.980 72.860 ;
        RECT 148.340 72.600 148.660 72.860 ;
        RECT 95.990 72.320 100.730 72.460 ;
        RECT 89.935 72.275 90.225 72.320 ;
        RECT 94.995 72.275 95.285 72.320 ;
        RECT 87.620 72.260 88.005 72.275 ;
        RECT 84.415 72.120 84.705 72.165 ;
        RECT 82.560 71.980 84.705 72.120 ;
        RECT 60.940 71.640 64.390 71.780 ;
        RECT 73.910 71.780 74.050 71.935 ;
        RECT 76.580 71.780 76.900 71.840 ;
        RECT 73.910 71.640 76.900 71.780 ;
        RECT 77.590 71.780 77.730 71.935 ;
        RECT 80.735 71.780 81.025 71.825 ;
        RECT 82.190 71.780 82.330 71.935 ;
        RECT 82.560 71.920 82.880 71.980 ;
        RECT 84.415 71.935 84.705 71.980 ;
        RECT 85.335 71.935 85.625 72.165 ;
        RECT 85.780 71.920 86.100 72.180 ;
        RECT 86.700 71.920 87.020 72.180 ;
        RECT 87.715 72.045 88.005 72.260 ;
        RECT 89.015 72.120 89.305 72.165 ;
        RECT 91.760 72.120 92.080 72.180 ;
        RECT 92.235 72.120 92.525 72.165 ;
        RECT 89.015 71.980 91.070 72.120 ;
        RECT 89.015 71.935 89.305 71.980 ;
        RECT 83.035 71.780 83.325 71.825 ;
        RECT 83.940 71.780 84.260 71.840 ;
        RECT 77.590 71.640 79.110 71.780 ;
        RECT 60.940 71.580 61.260 71.640 ;
        RECT 76.580 71.580 76.900 71.640 ;
        RECT 78.970 71.500 79.110 71.640 ;
        RECT 80.735 71.640 82.790 71.780 ;
        RECT 80.735 71.595 81.025 71.640 ;
        RECT 42.555 71.300 49.670 71.440 ;
        RECT 30.120 71.240 30.440 71.300 ;
        RECT 36.100 71.240 36.420 71.300 ;
        RECT 42.555 71.255 42.845 71.300 ;
        RECT 40.715 71.100 41.005 71.145 ;
        RECT 42.080 71.100 42.400 71.160 ;
        RECT 44.470 71.145 44.610 71.300 ;
        RECT 54.975 71.255 55.265 71.485 ;
        RECT 78.880 71.440 79.200 71.500 ;
        RECT 79.815 71.440 80.105 71.485 ;
        RECT 82.650 71.440 82.790 71.640 ;
        RECT 83.035 71.640 84.260 71.780 ;
        RECT 83.035 71.595 83.325 71.640 ;
        RECT 83.940 71.580 84.260 71.640 ;
        RECT 84.875 71.780 85.165 71.825 ;
        RECT 89.460 71.780 89.780 71.840 ;
        RECT 84.875 71.640 89.780 71.780 ;
        RECT 90.930 71.780 91.070 71.980 ;
        RECT 91.760 71.980 92.525 72.120 ;
        RECT 91.760 71.920 92.080 71.980 ;
        RECT 92.235 71.935 92.525 71.980 ;
        RECT 92.680 71.920 93.000 72.180 ;
        RECT 93.615 72.120 93.905 72.165 ;
        RECT 94.060 72.120 94.380 72.180 ;
        RECT 93.615 71.980 94.380 72.120 ;
        RECT 93.615 71.935 93.905 71.980 ;
        RECT 91.300 71.780 91.620 71.840 ;
        RECT 93.690 71.780 93.830 71.935 ;
        RECT 94.060 71.920 94.380 71.980 ;
        RECT 96.375 71.935 96.665 72.165 ;
        RECT 96.820 72.120 97.140 72.180 ;
        RECT 97.755 72.120 98.045 72.165 ;
        RECT 98.200 72.120 98.520 72.180 ;
        RECT 96.820 71.980 98.520 72.120 ;
        RECT 90.930 71.640 93.830 71.780 ;
        RECT 94.520 71.780 94.840 71.840 ;
        RECT 95.455 71.780 95.745 71.825 ;
        RECT 94.520 71.640 95.745 71.780 ;
        RECT 96.450 71.780 96.590 71.935 ;
        RECT 96.820 71.920 97.140 71.980 ;
        RECT 97.755 71.935 98.045 71.980 ;
        RECT 98.200 71.920 98.520 71.980 ;
        RECT 98.660 71.920 98.980 72.180 ;
        RECT 100.590 72.165 100.730 72.320 ;
        RECT 100.515 71.935 100.805 72.165 ;
        RECT 108.410 72.120 108.550 72.600 ;
        RECT 118.990 72.460 119.130 72.600 ;
        RECT 129.110 72.460 129.250 72.600 ;
        RECT 118.990 72.320 131.090 72.460 ;
        RECT 108.795 72.120 109.085 72.165 ;
        RECT 108.410 71.980 109.085 72.120 ;
        RECT 108.795 71.935 109.085 71.980 ;
        RECT 109.240 71.920 109.560 72.180 ;
        RECT 117.535 71.935 117.825 72.165 ;
        RECT 118.455 72.120 118.745 72.165 ;
        RECT 118.990 72.120 119.130 72.320 ;
        RECT 118.455 71.980 119.130 72.120 ;
        RECT 118.455 71.935 118.745 71.980 ;
        RECT 99.595 71.780 99.885 71.825 ;
        RECT 100.975 71.780 101.265 71.825 ;
        RECT 96.450 71.640 101.265 71.780 ;
        RECT 84.875 71.595 85.165 71.640 ;
        RECT 89.460 71.580 89.780 71.640 ;
        RECT 91.300 71.580 91.620 71.640 ;
        RECT 94.520 71.580 94.840 71.640 ;
        RECT 95.455 71.595 95.745 71.640 ;
        RECT 99.595 71.595 99.885 71.640 ;
        RECT 100.975 71.595 101.265 71.640 ;
        RECT 107.860 71.780 108.180 71.840 ;
        RECT 110.175 71.780 110.465 71.825 ;
        RECT 107.860 71.640 110.465 71.780 ;
        RECT 117.610 71.780 117.750 71.935 ;
        RECT 120.740 71.920 121.060 72.180 ;
        RECT 126.260 72.120 126.580 72.180 ;
        RECT 126.735 72.120 127.025 72.165 ;
        RECT 126.260 71.980 127.025 72.120 ;
        RECT 126.260 71.920 126.580 71.980 ;
        RECT 126.735 71.935 127.025 71.980 ;
        RECT 127.180 72.120 127.500 72.180 ;
        RECT 127.655 72.120 127.945 72.165 ;
        RECT 127.180 71.980 127.945 72.120 ;
        RECT 127.180 71.920 127.500 71.980 ;
        RECT 127.655 71.935 127.945 71.980 ;
        RECT 128.115 71.935 128.405 72.165 ;
        RECT 129.035 72.120 129.325 72.165 ;
        RECT 128.650 71.980 129.325 72.120 ;
        RECT 120.830 71.780 120.970 71.920 ;
        RECT 117.610 71.640 120.970 71.780 ;
        RECT 125.340 71.780 125.660 71.840 ;
        RECT 128.190 71.780 128.330 71.935 ;
        RECT 128.650 71.840 128.790 71.980 ;
        RECT 129.035 71.935 129.325 71.980 ;
        RECT 130.400 71.920 130.720 72.180 ;
        RECT 130.950 72.165 131.090 72.320 ;
        RECT 130.875 71.935 131.165 72.165 ;
        RECT 132.240 72.120 132.560 72.180 ;
        RECT 133.175 72.120 133.465 72.165 ;
        RECT 133.620 72.120 133.940 72.180 ;
        RECT 132.240 71.980 133.940 72.120 ;
        RECT 132.240 71.920 132.560 71.980 ;
        RECT 133.175 71.935 133.465 71.980 ;
        RECT 133.620 71.920 133.940 71.980 ;
        RECT 134.095 71.935 134.385 72.165 ;
        RECT 134.630 72.120 134.770 72.600 ;
        RECT 135.015 72.460 135.305 72.505 ;
        RECT 136.470 72.460 136.610 72.600 ;
        RECT 135.015 72.320 136.610 72.460 ;
        RECT 135.015 72.275 135.305 72.320 ;
        RECT 136.470 72.165 136.610 72.320 ;
        RECT 135.475 72.120 135.765 72.165 ;
        RECT 134.630 71.980 135.765 72.120 ;
        RECT 135.475 71.935 135.765 71.980 ;
        RECT 136.395 71.935 136.685 72.165 ;
        RECT 137.390 72.120 137.530 72.600 ;
        RECT 138.235 72.120 138.525 72.165 ;
        RECT 137.390 71.980 138.525 72.120 ;
        RECT 138.235 71.935 138.525 71.980 ;
        RECT 139.615 71.935 139.905 72.165 ;
        RECT 144.750 72.120 144.890 72.600 ;
        RECT 146.975 72.120 147.265 72.165 ;
        RECT 144.750 71.980 147.265 72.120 ;
        RECT 146.975 71.935 147.265 71.980 ;
        RECT 147.895 72.120 148.185 72.165 ;
        RECT 148.430 72.120 148.570 72.600 ;
        RECT 147.895 71.980 148.570 72.120 ;
        RECT 147.895 71.935 148.185 71.980 ;
        RECT 125.340 71.640 128.330 71.780 ;
        RECT 107.860 71.580 108.180 71.640 ;
        RECT 110.175 71.595 110.465 71.640 ;
        RECT 125.340 71.580 125.660 71.640 ;
        RECT 128.560 71.580 128.880 71.840 ;
        RECT 91.760 71.440 92.080 71.500 ;
        RECT 117.520 71.440 117.840 71.500 ;
        RECT 134.170 71.440 134.310 71.935 ;
        RECT 135.000 71.580 135.320 71.840 ;
        RECT 139.690 71.780 139.830 71.935 ;
        RECT 147.435 71.780 147.725 71.825 ;
        RECT 148.800 71.780 149.120 71.840 ;
        RECT 137.390 71.640 139.830 71.780 ;
        RECT 140.150 71.640 147.190 71.780 ;
        RECT 55.510 71.300 77.730 71.440 ;
        RECT 40.715 70.960 42.400 71.100 ;
        RECT 40.715 70.915 41.005 70.960 ;
        RECT 42.080 70.900 42.400 70.960 ;
        RECT 44.395 70.915 44.685 71.145 ;
        RECT 51.740 70.900 52.060 71.160 ;
        RECT 52.200 71.100 52.520 71.160 ;
        RECT 53.135 71.100 53.425 71.145 ;
        RECT 52.200 70.960 53.425 71.100 ;
        RECT 52.200 70.900 52.520 70.960 ;
        RECT 53.135 70.915 53.425 70.960 ;
        RECT 54.500 71.100 54.820 71.160 ;
        RECT 55.510 71.100 55.650 71.300 ;
        RECT 54.500 70.960 55.650 71.100 ;
        RECT 56.355 71.100 56.645 71.145 ;
        RECT 56.800 71.100 57.120 71.160 ;
        RECT 56.355 70.960 57.120 71.100 ;
        RECT 54.500 70.900 54.820 70.960 ;
        RECT 56.355 70.915 56.645 70.960 ;
        RECT 56.800 70.900 57.120 70.960 ;
        RECT 57.260 70.900 57.580 71.160 ;
        RECT 64.160 71.100 64.480 71.160 ;
        RECT 65.095 71.100 65.385 71.145 ;
        RECT 64.160 70.960 65.385 71.100 ;
        RECT 64.160 70.900 64.480 70.960 ;
        RECT 65.095 70.915 65.385 70.960 ;
        RECT 65.540 71.100 65.860 71.160 ;
        RECT 66.015 71.100 66.305 71.145 ;
        RECT 65.540 70.960 66.305 71.100 ;
        RECT 65.540 70.900 65.860 70.960 ;
        RECT 66.015 70.915 66.305 70.960 ;
        RECT 77.040 70.900 77.360 71.160 ;
        RECT 77.590 71.100 77.730 71.300 ;
        RECT 78.880 71.300 80.105 71.440 ;
        RECT 78.880 71.240 79.200 71.300 ;
        RECT 79.815 71.255 80.105 71.300 ;
        RECT 80.350 71.300 82.100 71.440 ;
        RECT 82.650 71.300 92.080 71.440 ;
        RECT 80.350 71.100 80.490 71.300 ;
        RECT 77.590 70.960 80.490 71.100 ;
        RECT 81.180 70.900 81.500 71.160 ;
        RECT 81.960 71.100 82.100 71.300 ;
        RECT 91.760 71.240 92.080 71.300 ;
        RECT 95.530 71.300 105.330 71.440 ;
        RECT 95.530 71.160 95.670 71.300 ;
        RECT 105.190 71.160 105.330 71.300 ;
        RECT 117.520 71.300 134.310 71.440 ;
        RECT 117.520 71.240 117.840 71.300 ;
        RECT 92.220 71.100 92.540 71.160 ;
        RECT 81.960 70.960 92.540 71.100 ;
        RECT 92.220 70.900 92.540 70.960 ;
        RECT 95.440 70.900 95.760 71.160 ;
        RECT 97.280 71.100 97.600 71.160 ;
        RECT 100.515 71.100 100.805 71.145 ;
        RECT 97.280 70.960 100.805 71.100 ;
        RECT 97.280 70.900 97.600 70.960 ;
        RECT 100.515 70.915 100.805 70.960 ;
        RECT 102.340 70.900 102.660 71.160 ;
        RECT 105.100 70.900 105.420 71.160 ;
        RECT 108.320 71.100 108.640 71.160 ;
        RECT 117.060 71.100 117.380 71.160 ;
        RECT 108.320 70.960 117.380 71.100 ;
        RECT 108.320 70.900 108.640 70.960 ;
        RECT 117.060 70.900 117.380 70.960 ;
        RECT 117.995 71.100 118.285 71.145 ;
        RECT 118.440 71.100 118.760 71.160 ;
        RECT 117.995 70.960 118.760 71.100 ;
        RECT 117.995 70.915 118.285 70.960 ;
        RECT 118.440 70.900 118.760 70.960 ;
        RECT 127.180 70.900 127.500 71.160 ;
        RECT 128.575 71.100 128.865 71.145 ;
        RECT 129.020 71.100 129.340 71.160 ;
        RECT 128.575 70.960 129.340 71.100 ;
        RECT 128.575 70.915 128.865 70.960 ;
        RECT 129.020 70.900 129.340 70.960 ;
        RECT 129.940 71.100 130.260 71.160 ;
        RECT 130.415 71.100 130.705 71.145 ;
        RECT 129.940 70.960 130.705 71.100 ;
        RECT 129.940 70.900 130.260 70.960 ;
        RECT 130.415 70.915 130.705 70.960 ;
        RECT 132.255 71.100 132.545 71.145 ;
        RECT 135.090 71.100 135.230 71.580 ;
        RECT 137.390 71.485 137.530 71.640 ;
        RECT 137.315 71.255 137.605 71.485 ;
        RECT 140.150 71.440 140.290 71.640 ;
        RECT 138.770 71.300 140.290 71.440 ;
        RECT 140.535 71.440 140.825 71.485 ;
        RECT 141.440 71.440 141.760 71.500 ;
        RECT 140.535 71.300 141.760 71.440 ;
        RECT 147.050 71.440 147.190 71.640 ;
        RECT 147.435 71.640 149.120 71.780 ;
        RECT 147.435 71.595 147.725 71.640 ;
        RECT 148.800 71.580 149.120 71.640 ;
        RECT 148.340 71.440 148.660 71.500 ;
        RECT 152.020 71.440 152.340 71.500 ;
        RECT 147.050 71.300 152.340 71.440 ;
        RECT 138.770 71.160 138.910 71.300 ;
        RECT 140.535 71.255 140.825 71.300 ;
        RECT 141.440 71.240 141.760 71.300 ;
        RECT 148.340 71.240 148.660 71.300 ;
        RECT 152.020 71.240 152.340 71.300 ;
        RECT 132.255 70.960 135.230 71.100 ;
        RECT 132.255 70.915 132.545 70.960 ;
        RECT 135.460 70.900 135.780 71.160 ;
        RECT 138.680 70.900 139.000 71.160 ;
        RECT 140.995 71.100 141.285 71.145 ;
        RECT 142.820 71.100 143.140 71.160 ;
        RECT 140.995 70.960 143.140 71.100 ;
        RECT 140.995 70.915 141.285 70.960 ;
        RECT 142.820 70.900 143.140 70.960 ;
        RECT 22.690 70.280 157.010 70.760 ;
        RECT 31.040 69.880 31.360 70.140 ;
        RECT 49.915 70.080 50.205 70.125 ;
        RECT 51.280 70.080 51.600 70.140 ;
        RECT 54.960 70.080 55.280 70.140 ;
        RECT 57.260 70.080 57.580 70.140 ;
        RECT 49.915 69.940 51.600 70.080 ;
        RECT 49.915 69.895 50.205 69.940 ;
        RECT 51.280 69.880 51.600 69.940 ;
        RECT 54.130 69.940 55.280 70.080 ;
        RECT 31.130 69.400 31.270 69.880 ;
        RECT 46.220 69.740 46.540 69.800 ;
        RECT 54.130 69.740 54.270 69.940 ;
        RECT 54.960 69.880 55.280 69.940 ;
        RECT 55.970 69.940 57.580 70.080 ;
        RECT 29.290 69.260 31.270 69.400 ;
        RECT 29.290 69.105 29.430 69.260 ;
        RECT 28.295 68.875 28.585 69.105 ;
        RECT 29.215 68.875 29.505 69.105 ;
        RECT 29.675 69.060 29.965 69.105 ;
        RECT 30.120 69.060 30.440 69.120 ;
        RECT 31.130 69.105 31.270 69.260 ;
        RECT 32.050 69.600 36.330 69.740 ;
        RECT 32.050 69.120 32.190 69.600 ;
        RECT 33.800 69.200 34.120 69.460 ;
        RECT 35.180 69.400 35.500 69.460 ;
        RECT 34.350 69.260 35.500 69.400 ;
        RECT 29.675 68.920 30.440 69.060 ;
        RECT 29.675 68.875 29.965 68.920 ;
        RECT 28.370 68.720 28.510 68.875 ;
        RECT 29.750 68.720 29.890 68.875 ;
        RECT 30.120 68.860 30.440 68.920 ;
        RECT 30.595 68.875 30.885 69.105 ;
        RECT 31.055 68.875 31.345 69.105 ;
        RECT 28.370 68.580 29.890 68.720 ;
        RECT 26.440 68.380 26.760 68.440 ;
        RECT 28.755 68.380 29.045 68.425 ;
        RECT 26.440 68.240 29.045 68.380 ;
        RECT 26.440 68.180 26.760 68.240 ;
        RECT 28.755 68.195 29.045 68.240 ;
        RECT 30.120 68.180 30.440 68.440 ;
        RECT 30.670 68.380 30.810 68.875 ;
        RECT 31.960 68.860 32.280 69.120 ;
        RECT 33.355 69.060 33.645 69.105 ;
        RECT 33.890 69.060 34.030 69.200 ;
        RECT 34.350 69.105 34.490 69.260 ;
        RECT 35.180 69.200 35.500 69.260 ;
        RECT 36.190 69.120 36.330 69.600 ;
        RECT 46.220 69.600 54.270 69.740 ;
        RECT 46.220 69.540 46.540 69.600 ;
        RECT 54.500 69.540 54.820 69.800 ;
        RECT 38.860 69.400 39.180 69.460 ;
        RECT 54.590 69.400 54.730 69.540 ;
        RECT 55.970 69.445 56.110 69.940 ;
        RECT 57.260 69.880 57.580 69.940 ;
        RECT 60.940 69.880 61.260 70.140 ;
        RECT 62.780 69.880 63.100 70.140 ;
        RECT 71.060 69.880 71.380 70.140 ;
        RECT 79.340 70.080 79.660 70.140 ;
        RECT 72.990 69.940 74.050 70.080 ;
        RECT 56.820 69.740 57.110 69.785 ;
        RECT 58.195 69.740 58.485 69.785 ;
        RECT 56.820 69.600 58.485 69.740 ;
        RECT 56.820 69.555 57.110 69.600 ;
        RECT 58.195 69.555 58.485 69.600 ;
        RECT 65.540 69.740 65.830 69.785 ;
        RECT 67.110 69.740 67.400 69.785 ;
        RECT 69.210 69.740 69.500 69.785 ;
        RECT 65.540 69.600 69.500 69.740 ;
        RECT 71.150 69.740 71.290 69.880 ;
        RECT 71.150 69.600 72.210 69.740 ;
        RECT 65.540 69.555 65.830 69.600 ;
        RECT 67.110 69.555 67.400 69.600 ;
        RECT 69.210 69.555 69.500 69.600 ;
        RECT 38.860 69.260 51.050 69.400 ;
        RECT 38.860 69.200 39.180 69.260 ;
        RECT 33.355 68.920 34.030 69.060 ;
        RECT 33.355 68.875 33.645 68.920 ;
        RECT 34.275 68.875 34.565 69.105 ;
        RECT 36.100 69.060 36.420 69.120 ;
        RECT 50.910 69.105 51.050 69.260 ;
        RECT 51.325 69.260 54.730 69.400 ;
        RECT 37.035 69.060 37.325 69.105 ;
        RECT 36.100 68.920 37.325 69.060 ;
        RECT 36.100 68.860 36.420 68.920 ;
        RECT 37.035 68.875 37.325 68.920 ;
        RECT 37.570 68.920 49.210 69.060 ;
        RECT 31.515 68.720 31.805 68.765 ;
        RECT 32.420 68.720 32.740 68.780 ;
        RECT 37.570 68.720 37.710 68.920 ;
        RECT 31.515 68.580 37.710 68.720 ;
        RECT 37.955 68.720 38.245 68.765 ;
        RECT 41.620 68.720 41.940 68.780 ;
        RECT 37.955 68.580 41.940 68.720 ;
        RECT 31.515 68.535 31.805 68.580 ;
        RECT 32.420 68.520 32.740 68.580 ;
        RECT 37.955 68.535 38.245 68.580 ;
        RECT 41.620 68.520 41.940 68.580 ;
        RECT 46.220 68.720 46.540 68.780 ;
        RECT 49.070 68.765 49.210 68.920 ;
        RECT 50.835 68.875 51.125 69.105 ;
        RECT 48.075 68.720 48.365 68.765 ;
        RECT 46.220 68.580 48.365 68.720 ;
        RECT 46.220 68.520 46.540 68.580 ;
        RECT 48.075 68.535 48.365 68.580 ;
        RECT 48.995 68.535 49.285 68.765 ;
        RECT 51.325 68.720 51.465 69.260 ;
        RECT 51.755 69.060 52.045 69.105 ;
        RECT 52.215 69.060 52.505 69.105 ;
        RECT 51.755 68.920 52.505 69.060 ;
        RECT 51.755 68.875 52.045 68.920 ;
        RECT 52.215 68.875 52.505 68.920 ;
        RECT 49.530 68.580 51.465 68.720 ;
        RECT 52.290 68.720 52.430 68.875 ;
        RECT 53.120 68.860 53.440 69.120 ;
        RECT 53.670 69.105 53.810 69.260 ;
        RECT 55.895 69.215 56.185 69.445 ;
        RECT 56.360 69.400 56.650 69.445 ;
        RECT 58.700 69.400 58.990 69.445 ;
        RECT 56.360 69.260 58.990 69.400 ;
        RECT 56.360 69.215 56.650 69.260 ;
        RECT 58.700 69.215 58.990 69.260 ;
        RECT 65.105 69.400 65.395 69.445 ;
        RECT 67.625 69.400 67.915 69.445 ;
        RECT 68.815 69.400 69.105 69.445 ;
        RECT 65.105 69.260 69.105 69.400 ;
        RECT 65.105 69.215 65.395 69.260 ;
        RECT 67.625 69.215 67.915 69.260 ;
        RECT 68.815 69.215 69.105 69.260 ;
        RECT 69.680 69.200 70.000 69.460 ;
        RECT 53.595 68.875 53.885 69.105 ;
        RECT 54.515 68.875 54.805 69.105 ;
        RECT 56.800 69.060 57.120 69.120 ;
        RECT 72.070 69.105 72.210 69.600 ;
        RECT 57.275 69.060 57.565 69.105 ;
        RECT 56.800 68.920 57.565 69.060 ;
        RECT 54.055 68.720 54.345 68.765 ;
        RECT 52.290 68.580 54.345 68.720 ;
        RECT 54.590 68.720 54.730 68.875 ;
        RECT 56.800 68.860 57.120 68.920 ;
        RECT 57.275 68.875 57.565 68.920 ;
        RECT 71.075 68.875 71.365 69.105 ;
        RECT 71.995 68.875 72.285 69.105 ;
        RECT 72.455 69.060 72.745 69.105 ;
        RECT 72.990 69.060 73.130 69.940 ;
        RECT 73.360 69.540 73.680 69.800 ;
        RECT 73.910 69.740 74.050 69.940 ;
        RECT 79.340 69.940 85.035 70.080 ;
        RECT 79.340 69.880 79.660 69.940 ;
        RECT 84.400 69.740 84.720 69.800 ;
        RECT 73.910 69.600 84.720 69.740 ;
        RECT 84.895 69.740 85.035 69.940 ;
        RECT 89.000 69.880 89.320 70.140 ;
        RECT 90.840 69.880 91.160 70.140 ;
        RECT 91.315 70.080 91.605 70.125 ;
        RECT 95.440 70.080 95.760 70.140 ;
        RECT 91.315 69.940 95.760 70.080 ;
        RECT 91.315 69.895 91.605 69.940 ;
        RECT 95.440 69.880 95.760 69.940 ;
        RECT 97.280 69.880 97.600 70.140 ;
        RECT 97.740 70.080 98.060 70.140 ;
        RECT 98.215 70.080 98.505 70.125 ;
        RECT 102.340 70.080 102.660 70.140 ;
        RECT 97.740 69.940 98.505 70.080 ;
        RECT 97.740 69.880 98.060 69.940 ;
        RECT 98.215 69.895 98.505 69.940 ;
        RECT 99.670 69.940 102.660 70.080 ;
        RECT 90.380 69.740 90.700 69.800 ;
        RECT 84.895 69.600 90.700 69.740 ;
        RECT 84.400 69.540 84.720 69.600 ;
        RECT 90.380 69.540 90.700 69.600 ;
        RECT 91.760 69.740 92.080 69.800 ;
        RECT 91.760 69.600 96.590 69.740 ;
        RECT 91.760 69.540 92.080 69.600 ;
        RECT 75.675 69.400 75.965 69.445 ;
        RECT 86.240 69.400 86.560 69.460 ;
        RECT 96.450 69.445 96.590 69.600 ;
        RECT 73.450 69.260 75.965 69.400 ;
        RECT 73.450 69.105 73.590 69.260 ;
        RECT 72.455 68.920 73.130 69.060 ;
        RECT 72.455 68.875 72.745 68.920 ;
        RECT 73.375 68.875 73.665 69.105 ;
        RECT 55.880 68.720 56.200 68.780 ;
        RECT 54.590 68.580 56.200 68.720 ;
        RECT 33.340 68.380 33.660 68.440 ;
        RECT 33.815 68.380 34.105 68.425 ;
        RECT 30.670 68.240 34.105 68.380 ;
        RECT 33.340 68.180 33.660 68.240 ;
        RECT 33.815 68.195 34.105 68.240 ;
        RECT 41.160 68.380 41.480 68.440 ;
        RECT 49.530 68.380 49.670 68.580 ;
        RECT 54.055 68.535 54.345 68.580 ;
        RECT 55.880 68.520 56.200 68.580 ;
        RECT 68.300 68.765 68.620 68.780 ;
        RECT 68.300 68.535 68.650 68.765 ;
        RECT 71.150 68.720 71.290 68.875 ;
        RECT 72.530 68.720 72.670 68.875 ;
        RECT 73.820 68.860 74.140 69.120 ;
        RECT 74.370 69.070 74.510 69.260 ;
        RECT 75.675 69.215 75.965 69.260 ;
        RECT 78.510 69.260 85.090 69.400 ;
        RECT 74.755 69.070 75.045 69.105 ;
        RECT 74.370 68.930 75.045 69.070 ;
        RECT 74.755 68.875 75.045 68.930 ;
        RECT 75.200 68.860 75.520 69.120 ;
        RECT 76.120 69.060 76.440 69.120 ;
        RECT 78.510 69.105 78.650 69.260 ;
        RECT 78.435 69.060 78.725 69.105 ;
        RECT 76.120 68.920 78.725 69.060 ;
        RECT 76.120 68.860 76.440 68.920 ;
        RECT 78.435 68.875 78.725 68.920 ;
        RECT 81.640 69.060 81.960 69.120 ;
        RECT 83.570 69.105 83.710 69.260 ;
        RECT 82.575 69.060 82.865 69.105 ;
        RECT 81.640 68.920 82.865 69.060 ;
        RECT 81.640 68.860 81.960 68.920 ;
        RECT 82.575 68.875 82.865 68.920 ;
        RECT 83.495 68.875 83.785 69.105 ;
        RECT 83.955 69.060 84.245 69.105 ;
        RECT 84.400 69.060 84.720 69.120 ;
        RECT 84.950 69.105 85.090 69.260 ;
        RECT 86.240 69.260 92.450 69.400 ;
        RECT 86.240 69.200 86.560 69.260 ;
        RECT 83.955 68.920 84.720 69.060 ;
        RECT 83.955 68.875 84.245 68.920 ;
        RECT 84.400 68.860 84.720 68.920 ;
        RECT 84.875 69.060 85.165 69.105 ;
        RECT 87.620 69.060 87.940 69.120 ;
        RECT 84.875 68.920 87.940 69.060 ;
        RECT 84.875 68.875 85.165 68.920 ;
        RECT 87.620 68.860 87.940 68.920 ;
        RECT 88.540 68.860 88.860 69.120 ;
        RECT 89.000 68.860 89.320 69.120 ;
        RECT 89.475 68.875 89.765 69.105 ;
        RECT 71.150 68.580 72.670 68.720 ;
        RECT 76.580 68.720 76.900 68.780 ;
        RECT 77.515 68.720 77.805 68.765 ;
        RECT 81.730 68.720 81.870 68.860 ;
        RECT 76.580 68.580 81.870 68.720 ;
        RECT 88.630 68.720 88.770 68.860 ;
        RECT 89.550 68.720 89.690 68.875 ;
        RECT 91.300 68.860 91.620 69.120 ;
        RECT 92.310 69.105 92.450 69.260 ;
        RECT 96.375 69.215 96.665 69.445 ;
        RECT 92.235 69.060 92.525 69.105 ;
        RECT 92.695 69.060 92.985 69.105 ;
        RECT 92.235 68.920 92.985 69.060 ;
        RECT 92.235 68.875 92.525 68.920 ;
        RECT 92.695 68.875 92.985 68.920 ;
        RECT 93.615 68.875 93.905 69.105 ;
        RECT 94.980 69.060 95.300 69.120 ;
        RECT 99.670 69.105 99.810 69.940 ;
        RECT 102.340 69.880 102.660 69.940 ;
        RECT 107.860 70.080 108.180 70.140 ;
        RECT 109.255 70.080 109.545 70.125 ;
        RECT 111.095 70.080 111.385 70.125 ;
        RECT 107.860 69.940 111.385 70.080 ;
        RECT 107.860 69.880 108.180 69.940 ;
        RECT 109.255 69.895 109.545 69.940 ;
        RECT 111.095 69.895 111.385 69.940 ;
        RECT 113.380 70.080 113.700 70.140 ;
        RECT 138.680 70.080 139.000 70.140 ;
        RECT 142.820 70.080 143.140 70.140 ;
        RECT 113.380 69.940 139.000 70.080 ;
        RECT 113.380 69.880 113.700 69.940 ;
        RECT 138.680 69.880 139.000 69.940 ;
        RECT 139.690 69.940 143.140 70.080 ;
        RECT 101.900 69.740 102.190 69.785 ;
        RECT 103.275 69.740 103.565 69.785 ;
        RECT 101.900 69.600 103.565 69.740 ;
        RECT 101.900 69.555 102.190 69.600 ;
        RECT 103.275 69.555 103.565 69.600 ;
        RECT 106.035 69.555 106.325 69.785 ;
        RECT 101.440 69.400 101.730 69.445 ;
        RECT 103.780 69.400 104.070 69.445 ;
        RECT 101.440 69.260 104.070 69.400 ;
        RECT 101.440 69.215 101.730 69.260 ;
        RECT 103.780 69.215 104.070 69.260 ;
        RECT 97.295 69.060 97.585 69.105 ;
        RECT 94.980 68.920 97.585 69.060 ;
        RECT 88.630 68.580 89.690 68.720 ;
        RECT 90.840 68.720 91.160 68.780 ;
        RECT 93.690 68.720 93.830 68.875 ;
        RECT 94.980 68.860 95.300 68.920 ;
        RECT 97.295 68.875 97.585 68.920 ;
        RECT 99.595 68.875 99.885 69.105 ;
        RECT 100.960 68.860 101.280 69.120 ;
        RECT 102.355 68.875 102.645 69.105 ;
        RECT 106.110 69.060 106.250 69.555 ;
        RECT 116.140 69.540 116.460 69.800 ;
        RECT 116.600 69.740 116.920 69.800 ;
        RECT 119.360 69.740 119.680 69.800 ;
        RECT 125.340 69.740 125.660 69.800 ;
        RECT 116.600 69.600 117.290 69.740 ;
        RECT 116.600 69.540 116.920 69.600 ;
        RECT 110.620 69.060 110.940 69.120 ;
        RECT 106.110 68.920 110.940 69.060 ;
        RECT 90.840 68.580 93.830 68.720 ;
        RECT 95.915 68.720 96.205 68.765 ;
        RECT 99.120 68.720 99.440 68.780 ;
        RECT 102.430 68.720 102.570 68.875 ;
        RECT 110.620 68.860 110.940 68.920 ;
        RECT 111.540 68.860 111.860 69.120 ;
        RECT 116.230 69.105 116.370 69.540 ;
        RECT 117.150 69.445 117.290 69.600 ;
        RECT 119.360 69.600 125.660 69.740 ;
        RECT 119.360 69.540 119.680 69.600 ;
        RECT 125.340 69.540 125.660 69.600 ;
        RECT 127.180 69.740 127.500 69.800 ;
        RECT 132.700 69.740 133.020 69.800 ;
        RECT 133.620 69.740 133.940 69.800 ;
        RECT 127.180 69.600 132.470 69.740 ;
        RECT 127.180 69.540 127.500 69.600 ;
        RECT 117.075 69.215 117.365 69.445 ;
        RECT 119.450 69.400 119.590 69.540 ;
        RECT 118.070 69.260 119.590 69.400 ;
        RECT 122.135 69.400 122.425 69.445 ;
        RECT 124.880 69.400 125.200 69.460 ;
        RECT 122.135 69.260 125.200 69.400 ;
        RECT 118.070 69.105 118.210 69.260 ;
        RECT 122.135 69.215 122.425 69.260 ;
        RECT 124.880 69.200 125.200 69.260 ;
        RECT 115.235 68.875 115.525 69.105 ;
        RECT 116.155 69.060 116.445 69.105 ;
        RECT 116.615 69.060 116.905 69.105 ;
        RECT 116.155 68.920 116.905 69.060 ;
        RECT 116.155 68.875 116.445 68.920 ;
        RECT 116.615 68.875 116.905 68.920 ;
        RECT 117.535 69.070 117.825 69.105 ;
        RECT 117.995 69.070 118.285 69.105 ;
        RECT 117.535 68.930 118.285 69.070 ;
        RECT 117.535 68.875 117.825 68.930 ;
        RECT 117.995 68.875 118.285 68.930 ;
        RECT 118.440 69.060 118.760 69.120 ;
        RECT 121.660 69.105 121.980 69.120 ;
        RECT 125.430 69.105 125.570 69.540 ;
        RECT 130.400 69.200 130.720 69.460 ;
        RECT 118.915 69.060 119.205 69.105 ;
        RECT 119.375 69.060 119.665 69.105 ;
        RECT 118.440 68.920 119.665 69.060 ;
        RECT 95.915 68.580 99.440 68.720 ;
        RECT 68.300 68.520 68.620 68.535 ;
        RECT 76.580 68.520 76.900 68.580 ;
        RECT 77.515 68.535 77.805 68.580 ;
        RECT 90.840 68.520 91.160 68.580 ;
        RECT 95.915 68.535 96.205 68.580 ;
        RECT 41.160 68.240 49.670 68.380 ;
        RECT 41.160 68.180 41.480 68.240 ;
        RECT 51.280 68.180 51.600 68.440 ;
        RECT 51.740 68.380 52.060 68.440 ;
        RECT 52.675 68.380 52.965 68.425 ;
        RECT 61.400 68.380 61.720 68.440 ;
        RECT 51.740 68.240 61.720 68.380 ;
        RECT 51.740 68.180 52.060 68.240 ;
        RECT 52.675 68.195 52.965 68.240 ;
        RECT 61.400 68.180 61.720 68.240 ;
        RECT 70.140 68.380 70.460 68.440 ;
        RECT 71.535 68.380 71.825 68.425 ;
        RECT 70.140 68.240 71.825 68.380 ;
        RECT 70.140 68.180 70.460 68.240 ;
        RECT 71.535 68.195 71.825 68.240 ;
        RECT 74.295 68.380 74.585 68.425 ;
        RECT 74.740 68.380 75.060 68.440 ;
        RECT 74.295 68.240 75.060 68.380 ;
        RECT 74.295 68.195 74.585 68.240 ;
        RECT 74.740 68.180 75.060 68.240 ;
        RECT 83.480 68.180 83.800 68.440 ;
        RECT 84.400 68.180 84.720 68.440 ;
        RECT 93.155 68.380 93.445 68.425 ;
        RECT 95.990 68.380 96.130 68.535 ;
        RECT 99.120 68.520 99.440 68.580 ;
        RECT 100.590 68.580 102.570 68.720 ;
        RECT 110.175 68.720 110.465 68.765 ;
        RECT 113.380 68.720 113.700 68.780 ;
        RECT 110.175 68.580 113.700 68.720 ;
        RECT 115.310 68.720 115.450 68.875 ;
        RECT 118.440 68.860 118.760 68.920 ;
        RECT 118.915 68.875 119.205 68.920 ;
        RECT 119.375 68.875 119.665 68.920 ;
        RECT 120.295 69.060 120.585 69.105 ;
        RECT 121.660 69.060 121.995 69.105 ;
        RECT 120.295 68.920 122.175 69.060 ;
        RECT 120.295 68.875 120.585 68.920 ;
        RECT 121.660 68.875 121.995 68.920 ;
        RECT 122.595 68.875 122.885 69.105 ;
        RECT 125.355 68.875 125.645 69.105 ;
        RECT 129.955 69.060 130.245 69.105 ;
        RECT 129.955 68.920 130.355 69.060 ;
        RECT 129.955 68.875 130.245 68.920 ;
        RECT 120.370 68.720 120.510 68.875 ;
        RECT 121.660 68.860 121.980 68.875 ;
        RECT 115.310 68.580 120.510 68.720 ;
        RECT 120.740 68.720 121.060 68.780 ;
        RECT 122.670 68.720 122.810 68.875 ;
        RECT 124.435 68.720 124.725 68.765 ;
        RECT 128.560 68.720 128.880 68.780 ;
        RECT 120.740 68.580 128.880 68.720 ;
        RECT 100.590 68.425 100.730 68.580 ;
        RECT 110.175 68.535 110.465 68.580 ;
        RECT 113.380 68.520 113.700 68.580 ;
        RECT 120.740 68.520 121.060 68.580 ;
        RECT 124.435 68.535 124.725 68.580 ;
        RECT 128.560 68.520 128.880 68.580 ;
        RECT 130.030 68.720 130.170 68.875 ;
        RECT 130.860 68.860 131.180 69.120 ;
        RECT 132.330 69.105 132.470 69.600 ;
        RECT 132.700 69.600 133.390 69.740 ;
        RECT 132.700 69.540 133.020 69.600 ;
        RECT 133.250 69.400 133.390 69.600 ;
        RECT 133.620 69.600 138.450 69.740 ;
        RECT 133.620 69.540 133.940 69.600 ;
        RECT 133.250 69.260 133.850 69.400 ;
        RECT 133.710 69.105 133.850 69.260 ;
        RECT 131.335 68.875 131.625 69.105 ;
        RECT 132.255 69.060 132.545 69.105 ;
        RECT 132.715 69.060 133.005 69.105 ;
        RECT 132.255 68.920 133.005 69.060 ;
        RECT 132.255 68.875 132.545 68.920 ;
        RECT 132.715 68.875 133.005 68.920 ;
        RECT 133.635 68.875 133.925 69.105 ;
        RECT 131.410 68.720 131.550 68.875 ;
        RECT 136.840 68.860 137.160 69.120 ;
        RECT 130.030 68.580 131.550 68.720 ;
        RECT 131.795 68.720 132.085 68.765 ;
        RECT 137.760 68.720 138.080 68.780 ;
        RECT 131.795 68.580 138.080 68.720 ;
        RECT 138.310 68.720 138.450 69.600 ;
        RECT 139.690 69.445 139.830 69.940 ;
        RECT 142.820 69.880 143.140 69.940 ;
        RECT 147.435 70.080 147.725 70.125 ;
        RECT 147.880 70.080 148.200 70.140 ;
        RECT 151.575 70.080 151.865 70.125 ;
        RECT 147.435 69.940 151.865 70.080 ;
        RECT 147.435 69.895 147.725 69.940 ;
        RECT 147.880 69.880 148.200 69.940 ;
        RECT 151.575 69.895 151.865 69.940 ;
        RECT 140.540 69.740 140.830 69.785 ;
        RECT 141.915 69.740 142.205 69.785 ;
        RECT 140.540 69.600 142.205 69.740 ;
        RECT 140.540 69.555 140.830 69.600 ;
        RECT 141.915 69.555 142.205 69.600 ;
        RECT 144.675 69.555 144.965 69.785 ;
        RECT 139.615 69.215 139.905 69.445 ;
        RECT 140.080 69.400 140.370 69.445 ;
        RECT 142.420 69.400 142.710 69.445 ;
        RECT 140.080 69.260 142.710 69.400 ;
        RECT 144.750 69.400 144.890 69.555 ;
        RECT 144.750 69.260 152.250 69.400 ;
        RECT 140.080 69.215 140.370 69.260 ;
        RECT 142.420 69.215 142.710 69.260 ;
        RECT 140.995 69.060 141.285 69.105 ;
        RECT 141.440 69.060 141.760 69.120 ;
        RECT 140.995 68.920 141.760 69.060 ;
        RECT 140.995 68.875 141.285 68.920 ;
        RECT 141.440 68.860 141.760 68.920 ;
        RECT 145.580 68.860 145.900 69.120 ;
        RECT 149.810 69.105 149.950 69.260 ;
        RECT 152.110 69.105 152.250 69.260 ;
        RECT 146.055 69.060 146.345 69.105 ;
        RECT 146.055 68.920 146.730 69.060 ;
        RECT 146.055 68.875 146.345 68.920 ;
        RECT 145.670 68.720 145.810 68.860 ;
        RECT 138.310 68.580 145.810 68.720 ;
        RECT 93.155 68.240 96.130 68.380 ;
        RECT 93.155 68.195 93.445 68.240 ;
        RECT 100.515 68.195 100.805 68.425 ;
        RECT 108.320 68.180 108.640 68.440 ;
        RECT 109.175 68.380 109.465 68.425 ;
        RECT 110.620 68.380 110.940 68.440 ;
        RECT 109.175 68.240 110.940 68.380 ;
        RECT 109.175 68.195 109.465 68.240 ;
        RECT 110.620 68.180 110.940 68.240 ;
        RECT 115.680 68.180 116.000 68.440 ;
        RECT 118.440 68.180 118.760 68.440 ;
        RECT 119.820 68.180 120.140 68.440 ;
        RECT 123.500 68.380 123.820 68.440 ;
        RECT 130.030 68.380 130.170 68.580 ;
        RECT 131.795 68.535 132.085 68.580 ;
        RECT 137.760 68.520 138.080 68.580 ;
        RECT 123.500 68.240 130.170 68.380 ;
        RECT 133.175 68.380 133.465 68.425 ;
        RECT 135.920 68.380 136.240 68.440 ;
        RECT 144.200 68.380 144.520 68.440 ;
        RECT 133.175 68.240 144.520 68.380 ;
        RECT 123.500 68.180 123.820 68.240 ;
        RECT 133.175 68.195 133.465 68.240 ;
        RECT 135.920 68.180 136.240 68.240 ;
        RECT 144.200 68.180 144.520 68.240 ;
        RECT 145.120 68.180 145.440 68.440 ;
        RECT 146.590 68.425 146.730 68.920 ;
        RECT 149.735 68.875 150.025 69.105 ;
        RECT 151.115 68.875 151.405 69.105 ;
        RECT 152.035 68.875 152.325 69.105 ;
        RECT 148.340 68.520 148.660 68.780 ;
        RECT 150.180 68.720 150.500 68.780 ;
        RECT 150.655 68.720 150.945 68.765 ;
        RECT 151.190 68.720 151.330 68.875 ;
        RECT 150.180 68.580 151.330 68.720 ;
        RECT 150.180 68.520 150.500 68.580 ;
        RECT 150.655 68.535 150.945 68.580 ;
        RECT 146.515 68.195 146.805 68.425 ;
        RECT 147.355 68.380 147.645 68.425 ;
        RECT 148.815 68.380 149.105 68.425 ;
        RECT 147.355 68.240 149.105 68.380 ;
        RECT 147.355 68.195 147.645 68.240 ;
        RECT 148.815 68.195 149.105 68.240 ;
        RECT 22.690 67.560 157.810 68.040 ;
        RECT 43.460 67.360 43.780 67.420 ;
        RECT 45.315 67.360 45.605 67.405 ;
        RECT 43.460 67.220 45.605 67.360 ;
        RECT 43.460 67.160 43.780 67.220 ;
        RECT 45.315 67.175 45.605 67.220 ;
        RECT 50.835 67.360 51.125 67.405 ;
        RECT 52.200 67.360 52.520 67.420 ;
        RECT 50.835 67.220 52.520 67.360 ;
        RECT 50.835 67.175 51.125 67.220 ;
        RECT 52.200 67.160 52.520 67.220 ;
        RECT 53.120 67.360 53.440 67.420 ;
        RECT 64.160 67.405 64.480 67.420 ;
        RECT 53.595 67.360 53.885 67.405 ;
        RECT 53.120 67.220 53.885 67.360 ;
        RECT 53.120 67.160 53.440 67.220 ;
        RECT 53.595 67.175 53.885 67.220 ;
        RECT 64.160 67.175 64.595 67.405 ;
        RECT 65.095 67.175 65.385 67.405 ;
        RECT 66.475 67.360 66.765 67.405 ;
        RECT 68.300 67.360 68.620 67.420 ;
        RECT 66.475 67.220 68.620 67.360 ;
        RECT 66.475 67.175 66.765 67.220 ;
        RECT 64.160 67.160 64.480 67.175 ;
        RECT 49.915 67.020 50.205 67.065 ;
        RECT 37.110 66.880 42.770 67.020 ;
        RECT 31.960 66.680 32.280 66.740 ;
        RECT 32.435 66.680 32.725 66.725 ;
        RECT 31.960 66.540 32.725 66.680 ;
        RECT 31.960 66.480 32.280 66.540 ;
        RECT 32.435 66.495 32.725 66.540 ;
        RECT 33.340 66.480 33.660 66.740 ;
        RECT 37.110 66.725 37.250 66.880 ;
        RECT 42.630 66.740 42.770 66.880 ;
        RECT 47.230 66.880 49.670 67.020 ;
        RECT 37.035 66.495 37.325 66.725 ;
        RECT 37.955 66.495 38.245 66.725 ;
        RECT 38.030 66.340 38.170 66.495 ;
        RECT 41.620 66.480 41.940 66.740 ;
        RECT 42.540 66.680 42.860 66.740 ;
        RECT 43.015 66.680 43.305 66.725 ;
        RECT 42.540 66.540 43.305 66.680 ;
        RECT 42.540 66.480 42.860 66.540 ;
        RECT 43.015 66.495 43.305 66.540 ;
        RECT 43.935 66.680 44.225 66.725 ;
        RECT 44.380 66.680 44.700 66.740 ;
        RECT 43.935 66.540 44.700 66.680 ;
        RECT 43.935 66.495 44.225 66.540 ;
        RECT 44.380 66.480 44.700 66.540 ;
        RECT 44.855 66.495 45.145 66.725 ;
        RECT 45.300 66.680 45.620 66.740 ;
        RECT 45.775 66.680 46.065 66.725 ;
        RECT 46.695 66.680 46.985 66.725 ;
        RECT 47.230 66.680 47.370 66.880 ;
        RECT 45.300 66.540 47.370 66.680 ;
        RECT 47.615 66.680 47.905 66.725 ;
        RECT 48.060 66.680 48.380 66.740 ;
        RECT 47.615 66.540 48.380 66.680 ;
        RECT 38.860 66.340 39.180 66.400 ;
        RECT 44.930 66.340 45.070 66.495 ;
        RECT 45.300 66.480 45.620 66.540 ;
        RECT 45.775 66.495 46.065 66.540 ;
        RECT 46.695 66.495 46.985 66.540 ;
        RECT 47.615 66.495 47.905 66.540 ;
        RECT 48.060 66.480 48.380 66.540 ;
        RECT 48.995 66.495 49.285 66.725 ;
        RECT 49.530 66.680 49.670 66.880 ;
        RECT 49.915 66.880 52.890 67.020 ;
        RECT 49.915 66.835 50.205 66.880 ;
        RECT 51.295 66.710 51.585 66.725 ;
        RECT 50.910 66.680 51.585 66.710 ;
        RECT 49.530 66.570 51.585 66.680 ;
        RECT 49.530 66.540 51.050 66.570 ;
        RECT 51.295 66.495 51.585 66.570 ;
        RECT 49.070 66.340 49.210 66.495 ;
        RECT 52.200 66.480 52.520 66.740 ;
        RECT 38.030 66.200 45.070 66.340 ;
        RECT 48.610 66.200 49.210 66.340 ;
        RECT 38.860 66.140 39.180 66.200 ;
        RECT 33.340 66.000 33.660 66.060 ;
        RECT 48.610 66.000 48.750 66.200 ;
        RECT 33.340 65.860 48.750 66.000 ;
        RECT 52.215 66.000 52.505 66.045 ;
        RECT 52.750 66.000 52.890 66.880 ;
        RECT 63.255 66.835 63.545 67.065 ;
        RECT 53.595 66.495 53.885 66.725 ;
        RECT 54.515 66.680 54.805 66.725 ;
        RECT 58.180 66.680 58.500 66.740 ;
        RECT 54.515 66.540 58.500 66.680 ;
        RECT 54.515 66.495 54.805 66.540 ;
        RECT 53.670 66.340 53.810 66.495 ;
        RECT 58.180 66.480 58.500 66.540 ;
        RECT 54.040 66.340 54.360 66.400 ;
        RECT 63.330 66.340 63.470 66.835 ;
        RECT 65.170 66.680 65.310 67.175 ;
        RECT 68.300 67.160 68.620 67.220 ;
        RECT 73.820 67.360 74.140 67.420 ;
        RECT 76.580 67.360 76.900 67.420 ;
        RECT 73.820 67.220 76.900 67.360 ;
        RECT 73.820 67.160 74.140 67.220 ;
        RECT 76.580 67.160 76.900 67.220 ;
        RECT 83.480 67.360 83.800 67.420 ;
        RECT 84.400 67.360 84.720 67.420 ;
        RECT 83.480 67.220 84.720 67.360 ;
        RECT 83.480 67.160 83.800 67.220 ;
        RECT 84.400 67.160 84.720 67.220 ;
        RECT 88.540 67.160 88.860 67.420 ;
        RECT 96.375 67.360 96.665 67.405 ;
        RECT 97.280 67.360 97.600 67.420 ;
        RECT 96.375 67.220 97.600 67.360 ;
        RECT 96.375 67.175 96.665 67.220 ;
        RECT 97.280 67.160 97.600 67.220 ;
        RECT 111.095 67.360 111.385 67.405 ;
        RECT 111.095 67.220 111.770 67.360 ;
        RECT 111.095 67.175 111.385 67.220 ;
        RECT 111.630 67.080 111.770 67.220 ;
        RECT 130.875 67.175 131.165 67.405 ;
        RECT 132.255 67.360 132.545 67.405 ;
        RECT 134.080 67.360 134.400 67.420 ;
        RECT 132.255 67.220 134.400 67.360 ;
        RECT 132.255 67.175 132.545 67.220 ;
        RECT 93.155 67.020 93.445 67.065 ;
        RECT 95.455 67.020 95.745 67.065 ;
        RECT 96.820 67.020 97.140 67.080 ;
        RECT 107.860 67.020 108.180 67.080 ;
        RECT 83.570 66.880 87.390 67.020 ;
        RECT 83.570 66.740 83.710 66.880 ;
        RECT 65.555 66.680 65.845 66.725 ;
        RECT 65.170 66.540 65.845 66.680 ;
        RECT 65.555 66.495 65.845 66.540 ;
        RECT 77.040 66.680 77.360 66.740 ;
        RECT 78.435 66.680 78.725 66.725 ;
        RECT 77.040 66.540 78.725 66.680 ;
        RECT 77.040 66.480 77.360 66.540 ;
        RECT 78.435 66.495 78.725 66.540 ;
        RECT 65.080 66.340 65.400 66.400 ;
        RECT 53.670 66.200 56.110 66.340 ;
        RECT 63.330 66.200 65.400 66.340 ;
        RECT 54.040 66.140 54.360 66.200 ;
        RECT 55.970 66.000 56.110 66.200 ;
        RECT 65.080 66.140 65.400 66.200 ;
        RECT 67.380 66.140 67.700 66.400 ;
        RECT 78.510 66.340 78.650 66.495 ;
        RECT 79.340 66.480 79.660 66.740 ;
        RECT 80.720 66.480 81.040 66.740 ;
        RECT 82.560 66.480 82.880 66.740 ;
        RECT 83.480 66.480 83.800 66.740 ;
        RECT 83.955 66.495 84.245 66.725 ;
        RECT 84.400 66.680 84.720 66.740 ;
        RECT 84.875 66.680 85.165 66.725 ;
        RECT 84.400 66.540 85.165 66.680 ;
        RECT 82.650 66.340 82.790 66.480 ;
        RECT 84.030 66.340 84.170 66.495 ;
        RECT 84.400 66.480 84.720 66.540 ;
        RECT 84.875 66.495 85.165 66.540 ;
        RECT 78.510 66.200 84.170 66.340 ;
        RECT 67.470 66.000 67.610 66.140 ;
        RECT 52.215 65.860 55.650 66.000 ;
        RECT 55.970 65.860 67.610 66.000 ;
        RECT 70.600 66.000 70.920 66.060 ;
        RECT 74.740 66.000 75.060 66.060 ;
        RECT 70.600 65.860 75.060 66.000 ;
        RECT 33.340 65.800 33.660 65.860 ;
        RECT 52.215 65.815 52.505 65.860 ;
        RECT 55.510 65.720 55.650 65.860 ;
        RECT 70.600 65.800 70.920 65.860 ;
        RECT 74.740 65.800 75.060 65.860 ;
        RECT 83.020 66.000 83.340 66.060 ;
        RECT 83.955 66.000 84.245 66.045 ;
        RECT 83.020 65.860 84.245 66.000 ;
        RECT 84.950 66.000 85.090 66.495 ;
        RECT 87.250 66.340 87.390 66.880 ;
        RECT 88.170 66.880 92.450 67.020 ;
        RECT 88.170 66.740 88.310 66.880 ;
        RECT 88.080 66.480 88.400 66.740 ;
        RECT 89.015 66.680 89.305 66.725 ;
        RECT 90.840 66.680 91.160 66.740 ;
        RECT 89.015 66.540 91.160 66.680 ;
        RECT 89.015 66.495 89.305 66.540 ;
        RECT 90.840 66.480 91.160 66.540 ;
        RECT 91.300 66.480 91.620 66.740 ;
        RECT 92.310 66.725 92.450 66.880 ;
        RECT 93.155 66.880 97.140 67.020 ;
        RECT 93.155 66.835 93.445 66.880 ;
        RECT 95.455 66.835 95.745 66.880 ;
        RECT 96.820 66.820 97.140 66.880 ;
        RECT 104.270 66.880 108.180 67.020 ;
        RECT 92.235 66.680 92.525 66.725 ;
        RECT 92.695 66.680 92.985 66.725 ;
        RECT 93.615 66.680 93.905 66.725 ;
        RECT 92.235 66.540 92.985 66.680 ;
        RECT 92.235 66.495 92.525 66.540 ;
        RECT 92.695 66.495 92.985 66.540 ;
        RECT 93.230 66.540 93.905 66.680 ;
        RECT 91.390 66.340 91.530 66.480 ;
        RECT 87.250 66.200 91.530 66.340 ;
        RECT 93.230 66.060 93.370 66.540 ;
        RECT 93.615 66.495 93.905 66.540 ;
        RECT 94.535 66.680 94.825 66.725 ;
        RECT 94.980 66.680 95.300 66.740 ;
        RECT 94.535 66.540 95.300 66.680 ;
        RECT 94.535 66.495 94.825 66.540 ;
        RECT 94.980 66.480 95.300 66.540 ;
        RECT 100.960 66.480 101.280 66.740 ;
        RECT 104.270 66.725 104.410 66.880 ;
        RECT 107.860 66.820 108.180 66.880 ;
        RECT 111.540 66.820 111.860 67.080 ;
        RECT 112.475 66.835 112.765 67.065 ;
        RECT 124.420 67.020 124.740 67.080 ;
        RECT 130.950 67.020 131.090 67.175 ;
        RECT 134.080 67.160 134.400 67.220 ;
        RECT 135.460 67.360 135.780 67.420 ;
        RECT 135.935 67.360 136.225 67.405 ;
        RECT 135.460 67.220 136.225 67.360 ;
        RECT 135.460 67.160 135.780 67.220 ;
        RECT 135.935 67.175 136.225 67.220 ;
        RECT 149.275 67.360 149.565 67.405 ;
        RECT 150.180 67.360 150.500 67.420 ;
        RECT 149.275 67.220 150.500 67.360 ;
        RECT 149.275 67.175 149.565 67.220 ;
        RECT 150.180 67.160 150.500 67.220 ;
        RECT 135.015 67.020 135.305 67.065 ;
        RECT 143.710 67.020 144.000 67.065 ;
        RECT 145.120 67.020 145.440 67.080 ;
        RECT 122.670 66.880 124.740 67.020 ;
        RECT 104.195 66.495 104.485 66.725 ;
        RECT 104.640 66.680 104.960 66.740 ;
        RECT 105.475 66.680 105.765 66.725 ;
        RECT 104.640 66.540 105.765 66.680 ;
        RECT 104.640 66.480 104.960 66.540 ;
        RECT 105.475 66.495 105.765 66.540 ;
        RECT 111.080 66.680 111.400 66.740 ;
        RECT 112.550 66.680 112.690 66.835 ;
        RECT 111.080 66.540 112.690 66.680 ;
        RECT 111.080 66.480 111.400 66.540 ;
        RECT 121.200 66.480 121.520 66.740 ;
        RECT 122.670 66.725 122.810 66.880 ;
        RECT 124.420 66.820 124.740 66.880 ;
        RECT 124.970 66.880 126.950 67.020 ;
        RECT 130.950 66.880 137.990 67.020 ;
        RECT 124.970 66.740 125.110 66.880 ;
        RECT 122.595 66.495 122.885 66.725 ;
        RECT 123.515 66.680 123.805 66.725 ;
        RECT 123.975 66.680 124.265 66.725 ;
        RECT 123.515 66.540 124.265 66.680 ;
        RECT 123.515 66.495 123.805 66.540 ;
        RECT 123.975 66.495 124.265 66.540 ;
        RECT 105.075 66.340 105.365 66.385 ;
        RECT 106.265 66.340 106.555 66.385 ;
        RECT 108.785 66.340 109.075 66.385 ;
        RECT 105.075 66.200 109.075 66.340 ;
        RECT 105.075 66.155 105.365 66.200 ;
        RECT 106.265 66.155 106.555 66.200 ;
        RECT 108.785 66.155 109.075 66.200 ;
        RECT 110.620 66.340 110.940 66.400 ;
        RECT 113.395 66.340 113.685 66.385 ;
        RECT 124.050 66.340 124.190 66.495 ;
        RECT 124.880 66.480 125.200 66.740 ;
        RECT 125.800 66.680 126.120 66.740 ;
        RECT 126.275 66.680 126.565 66.725 ;
        RECT 125.800 66.540 126.565 66.680 ;
        RECT 125.800 66.480 126.120 66.540 ;
        RECT 126.275 66.495 126.565 66.540 ;
        RECT 125.890 66.340 126.030 66.480 ;
        RECT 110.620 66.200 113.685 66.340 ;
        RECT 110.620 66.140 110.940 66.200 ;
        RECT 113.395 66.155 113.685 66.200 ;
        RECT 118.530 66.200 123.270 66.340 ;
        RECT 124.050 66.200 126.030 66.340 ;
        RECT 126.810 66.340 126.950 66.880 ;
        RECT 135.015 66.835 135.305 66.880 ;
        RECT 127.195 66.680 127.485 66.725 ;
        RECT 129.020 66.680 129.340 66.740 ;
        RECT 130.415 66.680 130.705 66.725 ;
        RECT 127.195 66.540 130.705 66.680 ;
        RECT 127.195 66.495 127.485 66.540 ;
        RECT 129.020 66.480 129.340 66.540 ;
        RECT 130.415 66.495 130.705 66.540 ;
        RECT 130.860 66.680 131.180 66.740 ;
        RECT 131.335 66.680 131.625 66.725 ;
        RECT 131.795 66.680 132.085 66.725 ;
        RECT 130.860 66.540 132.085 66.680 ;
        RECT 130.860 66.480 131.180 66.540 ;
        RECT 131.335 66.495 131.625 66.540 ;
        RECT 131.795 66.495 132.085 66.540 ;
        RECT 132.700 66.480 133.020 66.740 ;
        RECT 137.850 66.725 137.990 66.880 ;
        RECT 143.710 66.880 145.440 67.020 ;
        RECT 143.710 66.835 144.000 66.880 ;
        RECT 145.120 66.820 145.440 66.880 ;
        RECT 134.095 66.495 134.385 66.725 ;
        RECT 137.775 66.495 138.065 66.725 ;
        RECT 132.790 66.340 132.930 66.480 ;
        RECT 126.810 66.200 132.930 66.340 ;
        RECT 118.530 66.060 118.670 66.200 ;
        RECT 93.140 66.000 93.460 66.060 ;
        RECT 84.950 65.860 93.460 66.000 ;
        RECT 83.020 65.800 83.340 65.860 ;
        RECT 83.955 65.815 84.245 65.860 ;
        RECT 93.140 65.800 93.460 65.860 ;
        RECT 104.680 66.000 104.970 66.045 ;
        RECT 106.780 66.000 107.070 66.045 ;
        RECT 108.350 66.000 108.640 66.045 ;
        RECT 104.680 65.860 108.640 66.000 ;
        RECT 104.680 65.815 104.970 65.860 ;
        RECT 106.780 65.815 107.070 65.860 ;
        RECT 108.350 65.815 108.640 65.860 ;
        RECT 118.440 65.800 118.760 66.060 ;
        RECT 121.660 66.000 121.980 66.060 ;
        RECT 122.595 66.000 122.885 66.045 ;
        RECT 121.660 65.860 122.885 66.000 ;
        RECT 123.130 66.000 123.270 66.200 ;
        RECT 134.170 66.000 134.310 66.495 ;
        RECT 141.900 66.480 142.220 66.740 ;
        RECT 142.360 66.480 142.680 66.740 ;
        RECT 136.380 66.140 136.700 66.400 ;
        RECT 136.860 66.340 137.150 66.385 ;
        RECT 139.200 66.340 139.490 66.385 ;
        RECT 136.860 66.200 139.490 66.340 ;
        RECT 136.860 66.155 137.150 66.200 ;
        RECT 139.200 66.155 139.490 66.200 ;
        RECT 143.255 66.340 143.545 66.385 ;
        RECT 144.445 66.340 144.735 66.385 ;
        RECT 146.965 66.340 147.255 66.385 ;
        RECT 143.255 66.200 147.255 66.340 ;
        RECT 143.255 66.155 143.545 66.200 ;
        RECT 144.445 66.155 144.735 66.200 ;
        RECT 146.965 66.155 147.255 66.200 ;
        RECT 123.130 65.860 134.310 66.000 ;
        RECT 137.320 66.000 137.610 66.045 ;
        RECT 138.740 66.000 139.030 66.045 ;
        RECT 137.320 65.860 139.030 66.000 ;
        RECT 121.660 65.800 121.980 65.860 ;
        RECT 122.595 65.815 122.885 65.860 ;
        RECT 137.320 65.815 137.610 65.860 ;
        RECT 138.740 65.815 139.030 65.860 ;
        RECT 142.860 66.000 143.150 66.045 ;
        RECT 144.960 66.000 145.250 66.045 ;
        RECT 146.530 66.000 146.820 66.045 ;
        RECT 142.860 65.860 146.820 66.000 ;
        RECT 142.860 65.815 143.150 65.860 ;
        RECT 144.960 65.815 145.250 65.860 ;
        RECT 146.530 65.815 146.820 65.860 ;
        RECT 37.940 65.460 38.260 65.720 ;
        RECT 40.255 65.660 40.545 65.705 ;
        RECT 40.700 65.660 41.020 65.720 ;
        RECT 40.255 65.520 41.020 65.660 ;
        RECT 40.255 65.475 40.545 65.520 ;
        RECT 40.700 65.460 41.020 65.520 ;
        RECT 42.555 65.660 42.845 65.705 ;
        RECT 43.000 65.660 43.320 65.720 ;
        RECT 42.555 65.520 43.320 65.660 ;
        RECT 42.555 65.475 42.845 65.520 ;
        RECT 43.000 65.460 43.320 65.520 ;
        RECT 43.920 65.460 44.240 65.720 ;
        RECT 47.600 65.660 47.920 65.720 ;
        RECT 50.360 65.660 50.680 65.720 ;
        RECT 47.600 65.520 50.680 65.660 ;
        RECT 47.600 65.460 47.920 65.520 ;
        RECT 50.360 65.460 50.680 65.520 ;
        RECT 54.960 65.460 55.280 65.720 ;
        RECT 55.420 65.460 55.740 65.720 ;
        RECT 64.175 65.660 64.465 65.705 ;
        RECT 65.540 65.660 65.860 65.720 ;
        RECT 64.175 65.520 65.860 65.660 ;
        RECT 64.175 65.475 64.465 65.520 ;
        RECT 65.540 65.460 65.860 65.520 ;
        RECT 71.520 65.460 71.840 65.720 ;
        RECT 79.340 65.460 79.660 65.720 ;
        RECT 79.800 65.460 80.120 65.720 ;
        RECT 83.480 65.460 83.800 65.720 ;
        RECT 91.315 65.660 91.605 65.705 ;
        RECT 93.600 65.660 93.920 65.720 ;
        RECT 94.520 65.660 94.840 65.720 ;
        RECT 91.315 65.520 94.840 65.660 ;
        RECT 91.315 65.475 91.605 65.520 ;
        RECT 93.600 65.460 93.920 65.520 ;
        RECT 94.520 65.460 94.840 65.520 ;
        RECT 122.120 65.460 122.440 65.720 ;
        RECT 124.880 65.460 125.200 65.720 ;
        RECT 126.275 65.660 126.565 65.705 ;
        RECT 127.640 65.660 127.960 65.720 ;
        RECT 126.275 65.520 127.960 65.660 ;
        RECT 126.275 65.475 126.565 65.520 ;
        RECT 127.640 65.460 127.960 65.520 ;
        RECT 22.690 64.840 157.010 65.320 ;
        RECT 40.240 64.440 40.560 64.700 ;
        RECT 43.920 64.440 44.240 64.700 ;
        RECT 44.380 64.640 44.700 64.700 ;
        RECT 48.060 64.640 48.380 64.700 ;
        RECT 53.120 64.640 53.440 64.700 ;
        RECT 54.960 64.640 55.280 64.700 ;
        RECT 44.380 64.500 53.440 64.640 ;
        RECT 44.380 64.440 44.700 64.500 ;
        RECT 48.060 64.440 48.380 64.500 ;
        RECT 53.120 64.440 53.440 64.500 ;
        RECT 53.670 64.500 55.280 64.640 ;
        RECT 30.140 64.300 30.430 64.345 ;
        RECT 31.560 64.300 31.850 64.345 ;
        RECT 30.140 64.160 31.850 64.300 ;
        RECT 30.140 64.115 30.430 64.160 ;
        RECT 31.560 64.115 31.850 64.160 ;
        RECT 40.330 64.005 40.470 64.440 ;
        RECT 41.180 64.300 41.470 64.345 ;
        RECT 42.600 64.300 42.890 64.345 ;
        RECT 41.180 64.160 42.890 64.300 ;
        RECT 41.180 64.115 41.470 64.160 ;
        RECT 42.600 64.115 42.890 64.160 ;
        RECT 29.680 63.960 29.970 64.005 ;
        RECT 32.020 63.960 32.310 64.005 ;
        RECT 29.680 63.820 32.310 63.960 ;
        RECT 29.680 63.775 29.970 63.820 ;
        RECT 32.020 63.775 32.310 63.820 ;
        RECT 40.255 63.775 40.545 64.005 ;
        RECT 40.720 63.960 41.010 64.005 ;
        RECT 43.060 63.960 43.350 64.005 ;
        RECT 40.720 63.820 43.350 63.960 ;
        RECT 40.720 63.775 41.010 63.820 ;
        RECT 43.060 63.775 43.350 63.820 ;
        RECT 24.600 63.420 24.920 63.680 ;
        RECT 25.520 63.620 25.840 63.680 ;
        RECT 26.455 63.620 26.745 63.665 ;
        RECT 25.520 63.480 26.745 63.620 ;
        RECT 25.520 63.420 25.840 63.480 ;
        RECT 26.455 63.435 26.745 63.480 ;
        RECT 28.755 63.620 29.045 63.665 ;
        RECT 29.215 63.620 29.505 63.665 ;
        RECT 28.755 63.480 29.505 63.620 ;
        RECT 28.755 63.435 29.045 63.480 ;
        RECT 29.215 63.435 29.505 63.480 ;
        RECT 30.595 63.620 30.885 63.665 ;
        RECT 33.340 63.620 33.660 63.680 ;
        RECT 30.595 63.480 33.660 63.620 ;
        RECT 30.595 63.435 30.885 63.480 ;
        RECT 33.340 63.420 33.660 63.480 ;
        RECT 34.720 63.420 35.040 63.680 ;
        RECT 36.115 63.620 36.405 63.665 ;
        RECT 36.560 63.620 36.880 63.680 ;
        RECT 36.115 63.480 36.880 63.620 ;
        RECT 36.115 63.435 36.405 63.480 ;
        RECT 36.560 63.420 36.880 63.480 ;
        RECT 37.480 63.620 37.800 63.680 ;
        RECT 38.415 63.620 38.705 63.665 ;
        RECT 37.480 63.480 38.705 63.620 ;
        RECT 37.480 63.420 37.800 63.480 ;
        RECT 38.415 63.435 38.705 63.480 ;
        RECT 39.795 63.435 40.085 63.665 ;
        RECT 41.635 63.620 41.925 63.665 ;
        RECT 44.010 63.620 44.150 64.440 ;
        RECT 48.540 64.300 48.830 64.345 ;
        RECT 49.960 64.300 50.250 64.345 ;
        RECT 48.540 64.160 50.250 64.300 ;
        RECT 48.540 64.115 48.830 64.160 ;
        RECT 49.960 64.115 50.250 64.160 ;
        RECT 53.670 64.005 53.810 64.500 ;
        RECT 54.960 64.440 55.280 64.500 ;
        RECT 71.520 64.440 71.840 64.700 ;
        RECT 75.200 64.640 75.520 64.700 ;
        RECT 94.980 64.640 95.300 64.700 ;
        RECT 75.200 64.500 95.300 64.640 ;
        RECT 75.200 64.440 75.520 64.500 ;
        RECT 94.980 64.440 95.300 64.500 ;
        RECT 104.640 64.640 104.960 64.700 ;
        RECT 107.415 64.640 107.705 64.685 ;
        RECT 126.735 64.640 127.025 64.685 ;
        RECT 104.640 64.500 107.705 64.640 ;
        RECT 104.640 64.440 104.960 64.500 ;
        RECT 107.415 64.455 107.705 64.500 ;
        RECT 120.830 64.500 127.025 64.640 ;
        RECT 54.520 64.300 54.810 64.345 ;
        RECT 55.940 64.300 56.230 64.345 ;
        RECT 54.520 64.160 56.230 64.300 ;
        RECT 54.520 64.115 54.810 64.160 ;
        RECT 55.940 64.115 56.230 64.160 ;
        RECT 69.650 64.300 69.940 64.345 ;
        RECT 71.070 64.300 71.360 64.345 ;
        RECT 69.650 64.160 71.360 64.300 ;
        RECT 71.610 64.300 71.750 64.440 ;
        RECT 73.380 64.300 73.670 64.345 ;
        RECT 74.800 64.300 75.090 64.345 ;
        RECT 71.610 64.160 72.210 64.300 ;
        RECT 69.650 64.115 69.940 64.160 ;
        RECT 71.070 64.115 71.360 64.160 ;
        RECT 72.070 64.005 72.210 64.160 ;
        RECT 73.380 64.160 75.090 64.300 ;
        RECT 73.380 64.115 73.670 64.160 ;
        RECT 74.800 64.115 75.090 64.160 ;
        RECT 79.360 64.300 79.650 64.345 ;
        RECT 80.780 64.300 81.070 64.345 ;
        RECT 79.360 64.160 81.070 64.300 ;
        RECT 79.360 64.115 79.650 64.160 ;
        RECT 80.780 64.115 81.070 64.160 ;
        RECT 96.840 64.300 97.130 64.345 ;
        RECT 98.260 64.300 98.550 64.345 ;
        RECT 96.840 64.160 98.550 64.300 ;
        RECT 96.840 64.115 97.130 64.160 ;
        RECT 98.260 64.115 98.550 64.160 ;
        RECT 115.700 64.300 115.990 64.345 ;
        RECT 117.120 64.300 117.410 64.345 ;
        RECT 115.700 64.160 117.410 64.300 ;
        RECT 115.700 64.115 115.990 64.160 ;
        RECT 117.120 64.115 117.410 64.160 ;
        RECT 120.830 64.005 120.970 64.500 ;
        RECT 126.735 64.455 127.025 64.500 ;
        RECT 121.680 64.300 121.970 64.345 ;
        RECT 123.100 64.300 123.390 64.345 ;
        RECT 121.680 64.160 123.390 64.300 ;
        RECT 121.680 64.115 121.970 64.160 ;
        RECT 123.100 64.115 123.390 64.160 ;
        RECT 132.720 64.300 133.010 64.345 ;
        RECT 134.140 64.300 134.430 64.345 ;
        RECT 132.720 64.160 134.430 64.300 ;
        RECT 132.720 64.115 133.010 64.160 ;
        RECT 134.140 64.115 134.430 64.160 ;
        RECT 143.760 64.300 144.050 64.345 ;
        RECT 145.180 64.300 145.470 64.345 ;
        RECT 143.760 64.160 145.470 64.300 ;
        RECT 143.760 64.115 144.050 64.160 ;
        RECT 145.180 64.115 145.470 64.160 ;
        RECT 48.080 63.960 48.370 64.005 ;
        RECT 50.420 63.960 50.710 64.005 ;
        RECT 48.080 63.820 50.710 63.960 ;
        RECT 48.080 63.775 48.370 63.820 ;
        RECT 50.420 63.775 50.710 63.820 ;
        RECT 53.595 63.775 53.885 64.005 ;
        RECT 54.060 63.960 54.350 64.005 ;
        RECT 56.400 63.960 56.690 64.005 ;
        RECT 54.060 63.820 56.690 63.960 ;
        RECT 54.060 63.775 54.350 63.820 ;
        RECT 56.400 63.775 56.690 63.820 ;
        RECT 69.190 63.960 69.480 64.005 ;
        RECT 71.530 63.960 71.820 64.005 ;
        RECT 69.190 63.820 71.820 63.960 ;
        RECT 69.190 63.775 69.480 63.820 ;
        RECT 71.530 63.775 71.820 63.820 ;
        RECT 71.995 63.775 72.285 64.005 ;
        RECT 72.920 63.960 73.210 64.005 ;
        RECT 75.260 63.960 75.550 64.005 ;
        RECT 72.920 63.820 75.550 63.960 ;
        RECT 72.920 63.775 73.210 63.820 ;
        RECT 75.260 63.775 75.550 63.820 ;
        RECT 78.900 63.960 79.190 64.005 ;
        RECT 81.240 63.960 81.530 64.005 ;
        RECT 78.900 63.820 81.530 63.960 ;
        RECT 78.900 63.775 79.190 63.820 ;
        RECT 81.240 63.775 81.530 63.820 ;
        RECT 96.380 63.960 96.670 64.005 ;
        RECT 98.720 63.960 99.010 64.005 ;
        RECT 96.380 63.820 99.010 63.960 ;
        RECT 96.380 63.775 96.670 63.820 ;
        RECT 98.720 63.775 99.010 63.820 ;
        RECT 115.240 63.960 115.530 64.005 ;
        RECT 117.580 63.960 117.870 64.005 ;
        RECT 115.240 63.820 117.870 63.960 ;
        RECT 115.240 63.775 115.530 63.820 ;
        RECT 117.580 63.775 117.870 63.820 ;
        RECT 120.755 63.775 121.045 64.005 ;
        RECT 121.220 63.960 121.510 64.005 ;
        RECT 123.560 63.960 123.850 64.005 ;
        RECT 121.220 63.820 123.850 63.960 ;
        RECT 121.220 63.775 121.510 63.820 ;
        RECT 123.560 63.775 123.850 63.820 ;
        RECT 132.260 63.960 132.550 64.005 ;
        RECT 134.600 63.960 134.890 64.005 ;
        RECT 132.260 63.820 134.890 63.960 ;
        RECT 132.260 63.775 132.550 63.820 ;
        RECT 134.600 63.775 134.890 63.820 ;
        RECT 143.300 63.960 143.590 64.005 ;
        RECT 145.640 63.960 145.930 64.005 ;
        RECT 143.300 63.820 145.930 63.960 ;
        RECT 143.300 63.775 143.590 63.820 ;
        RECT 145.640 63.775 145.930 63.820 ;
        RECT 41.635 63.480 44.150 63.620 ;
        RECT 41.635 63.435 41.925 63.480 ;
        RECT 39.870 63.280 40.010 63.435 ;
        RECT 45.760 63.420 46.080 63.680 ;
        RECT 46.220 63.420 46.540 63.680 ;
        RECT 47.615 63.620 47.905 63.665 ;
        RECT 48.520 63.620 48.840 63.680 ;
        RECT 47.615 63.480 48.840 63.620 ;
        RECT 47.615 63.435 47.905 63.480 ;
        RECT 48.520 63.420 48.840 63.480 ;
        RECT 48.980 63.420 49.300 63.680 ;
        RECT 53.120 63.420 53.440 63.680 ;
        RECT 54.975 63.620 55.265 63.665 ;
        RECT 55.420 63.620 55.740 63.680 ;
        RECT 54.975 63.480 55.740 63.620 ;
        RECT 54.975 63.435 55.265 63.480 ;
        RECT 55.420 63.420 55.740 63.480 ;
        RECT 59.100 63.420 59.420 63.680 ;
        RECT 59.560 63.420 59.880 63.680 ;
        RECT 66.000 63.420 66.320 63.680 ;
        RECT 66.475 63.435 66.765 63.665 ;
        RECT 40.240 63.280 40.560 63.340 ;
        RECT 39.870 63.140 40.560 63.280 ;
        RECT 40.240 63.080 40.560 63.140 ;
        RECT 37.480 62.740 37.800 63.000 ;
        RECT 66.550 62.940 66.690 63.435 ;
        RECT 70.600 63.420 70.920 63.680 ;
        RECT 72.455 63.435 72.745 63.665 ;
        RECT 71.520 63.280 71.840 63.340 ;
        RECT 72.530 63.280 72.670 63.435 ;
        RECT 73.820 63.420 74.140 63.680 ;
        RECT 77.960 63.420 78.280 63.680 ;
        RECT 78.420 63.420 78.740 63.680 ;
        RECT 79.800 63.420 80.120 63.680 ;
        RECT 83.940 63.420 84.260 63.680 ;
        RECT 84.400 63.420 84.720 63.680 ;
        RECT 85.780 63.420 86.100 63.680 ;
        RECT 90.840 63.420 91.160 63.680 ;
        RECT 93.140 63.420 93.460 63.680 ;
        RECT 95.455 63.620 95.745 63.665 ;
        RECT 95.915 63.620 96.205 63.665 ;
        RECT 95.455 63.480 96.205 63.620 ;
        RECT 95.455 63.435 95.745 63.480 ;
        RECT 95.915 63.435 96.205 63.480 ;
        RECT 96.820 63.620 97.140 63.680 ;
        RECT 97.295 63.620 97.585 63.665 ;
        RECT 96.820 63.480 97.585 63.620 ;
        RECT 96.820 63.420 97.140 63.480 ;
        RECT 97.295 63.435 97.585 63.480 ;
        RECT 101.420 63.420 101.740 63.680 ;
        RECT 101.880 63.420 102.200 63.680 ;
        RECT 104.195 63.620 104.485 63.665 ;
        RECT 106.480 63.620 106.800 63.680 ;
        RECT 104.195 63.480 106.800 63.620 ;
        RECT 104.195 63.435 104.485 63.480 ;
        RECT 106.480 63.420 106.800 63.480 ;
        RECT 108.320 63.420 108.640 63.680 ;
        RECT 114.315 63.620 114.605 63.665 ;
        RECT 114.775 63.620 115.065 63.665 ;
        RECT 114.315 63.480 115.065 63.620 ;
        RECT 114.315 63.435 114.605 63.480 ;
        RECT 114.775 63.435 115.065 63.480 ;
        RECT 116.155 63.620 116.445 63.665 ;
        RECT 118.900 63.620 119.220 63.680 ;
        RECT 116.155 63.480 119.220 63.620 ;
        RECT 116.155 63.435 116.445 63.480 ;
        RECT 118.900 63.420 119.220 63.480 ;
        RECT 120.280 63.420 120.600 63.680 ;
        RECT 122.120 63.420 122.440 63.680 ;
        RECT 126.260 63.420 126.580 63.680 ;
        RECT 127.180 63.620 127.500 63.680 ;
        RECT 128.115 63.620 128.405 63.665 ;
        RECT 127.180 63.480 128.405 63.620 ;
        RECT 127.180 63.420 127.500 63.480 ;
        RECT 128.115 63.435 128.405 63.480 ;
        RECT 129.480 63.420 129.800 63.680 ;
        RECT 131.795 63.620 132.085 63.665 ;
        RECT 132.700 63.620 133.020 63.680 ;
        RECT 131.795 63.480 133.020 63.620 ;
        RECT 131.795 63.435 132.085 63.480 ;
        RECT 132.700 63.420 133.020 63.480 ;
        RECT 133.160 63.420 133.480 63.680 ;
        RECT 136.380 63.620 136.700 63.680 ;
        RECT 137.315 63.620 137.605 63.665 ;
        RECT 136.380 63.480 137.605 63.620 ;
        RECT 136.380 63.420 136.700 63.480 ;
        RECT 137.315 63.435 137.605 63.480 ;
        RECT 138.680 63.620 139.000 63.680 ;
        RECT 139.155 63.620 139.445 63.665 ;
        RECT 138.680 63.480 139.445 63.620 ;
        RECT 138.680 63.420 139.000 63.480 ;
        RECT 139.155 63.435 139.445 63.480 ;
        RECT 142.835 63.435 143.125 63.665 ;
        RECT 71.520 63.140 72.670 63.280 ;
        RECT 142.910 63.280 143.050 63.435 ;
        RECT 144.200 63.420 144.520 63.680 ;
        RECT 148.355 63.620 148.645 63.665 ;
        RECT 150.180 63.620 150.500 63.680 ;
        RECT 148.355 63.480 150.500 63.620 ;
        RECT 148.355 63.435 148.645 63.480 ;
        RECT 150.180 63.420 150.500 63.480 ;
        RECT 146.500 63.280 146.820 63.340 ;
        RECT 142.910 63.140 146.820 63.280 ;
        RECT 71.520 63.080 71.840 63.140 ;
        RECT 146.500 63.080 146.820 63.140 ;
        RECT 75.660 62.940 75.980 63.000 ;
        RECT 66.550 62.800 75.980 62.940 ;
        RECT 75.660 62.740 75.980 62.800 ;
        RECT 22.690 62.120 157.810 62.600 ;
        RECT 26.440 61.720 26.760 61.980 ;
        RECT 30.120 61.720 30.440 61.980 ;
        RECT 37.480 61.720 37.800 61.980 ;
        RECT 51.280 61.920 51.600 61.980 ;
        RECT 56.800 61.920 57.120 61.980 ;
        RECT 51.280 61.780 57.120 61.920 ;
        RECT 51.280 61.720 51.600 61.780 ;
        RECT 56.800 61.720 57.120 61.780 ;
        RECT 59.560 61.720 59.880 61.980 ;
        RECT 79.340 61.720 79.660 61.980 ;
        RECT 118.440 61.720 118.760 61.980 ;
        RECT 124.880 61.720 125.200 61.980 ;
        RECT 134.080 61.720 134.400 61.980 ;
        RECT 24.615 61.240 24.905 61.285 ;
        RECT 25.520 61.240 25.840 61.300 ;
        RECT 24.615 61.100 25.840 61.240 ;
        RECT 24.615 61.055 24.905 61.100 ;
        RECT 25.520 61.040 25.840 61.100 ;
        RECT 25.995 61.240 26.285 61.285 ;
        RECT 26.530 61.240 26.670 61.720 ;
        RECT 30.210 61.580 30.350 61.720 ;
        RECT 30.210 61.440 32.190 61.580 ;
        RECT 25.995 61.100 26.670 61.240 ;
        RECT 30.135 61.240 30.425 61.285 ;
        RECT 31.500 61.240 31.820 61.300 ;
        RECT 32.050 61.285 32.190 61.440 ;
        RECT 30.135 61.100 31.820 61.240 ;
        RECT 25.995 61.055 26.285 61.100 ;
        RECT 30.135 61.055 30.425 61.100 ;
        RECT 31.500 61.040 31.820 61.100 ;
        RECT 31.975 61.055 32.265 61.285 ;
        RECT 36.100 61.040 36.420 61.300 ;
        RECT 37.570 61.240 37.710 61.720 ;
        RECT 50.820 61.580 51.140 61.640 ;
        RECT 59.650 61.580 59.790 61.720 ;
        RECT 64.620 61.580 64.940 61.640 ;
        RECT 42.630 61.440 46.450 61.580 ;
        RECT 37.955 61.240 38.245 61.285 ;
        RECT 37.570 61.100 38.245 61.240 ;
        RECT 37.955 61.055 38.245 61.100 ;
        RECT 42.080 61.040 42.400 61.300 ;
        RECT 42.630 61.285 42.770 61.440 ;
        RECT 46.310 61.300 46.450 61.440 ;
        RECT 48.150 61.440 51.140 61.580 ;
        RECT 42.555 61.055 42.845 61.285 ;
        RECT 43.460 61.240 43.780 61.300 ;
        RECT 43.935 61.240 44.225 61.285 ;
        RECT 43.460 61.100 44.225 61.240 ;
        RECT 43.460 61.040 43.780 61.100 ;
        RECT 43.935 61.055 44.225 61.100 ;
        RECT 46.220 61.040 46.540 61.300 ;
        RECT 48.150 61.285 48.290 61.440 ;
        RECT 50.820 61.380 51.140 61.440 ;
        RECT 55.050 61.440 59.790 61.580 ;
        RECT 61.030 61.440 64.940 61.580 ;
        RECT 48.075 61.055 48.365 61.285 ;
        RECT 48.520 61.240 48.840 61.300 ;
        RECT 48.995 61.240 49.285 61.285 ;
        RECT 55.050 61.240 55.190 61.440 ;
        RECT 48.520 61.100 49.285 61.240 ;
        RECT 48.520 61.040 48.840 61.100 ;
        RECT 48.995 61.055 49.285 61.100 ;
        RECT 54.130 61.100 55.190 61.240 ;
        RECT 25.080 60.900 25.370 60.945 ;
        RECT 27.420 60.900 27.710 60.945 ;
        RECT 25.080 60.760 27.710 60.900 ;
        RECT 25.080 60.715 25.370 60.760 ;
        RECT 27.420 60.715 27.710 60.760 ;
        RECT 30.580 60.700 30.900 60.960 ;
        RECT 31.060 60.900 31.350 60.945 ;
        RECT 33.400 60.900 33.690 60.945 ;
        RECT 31.060 60.760 33.690 60.900 ;
        RECT 31.060 60.715 31.350 60.760 ;
        RECT 33.400 60.715 33.690 60.760 ;
        RECT 36.560 60.700 36.880 60.960 ;
        RECT 54.130 60.945 54.270 61.100 ;
        RECT 55.420 61.040 55.740 61.300 ;
        RECT 59.575 61.240 59.865 61.285 ;
        RECT 61.030 61.240 61.170 61.440 ;
        RECT 64.620 61.380 64.940 61.440 ;
        RECT 59.575 61.100 61.170 61.240 ;
        RECT 59.575 61.055 59.865 61.100 ;
        RECT 61.400 61.040 61.720 61.300 ;
        RECT 65.555 61.240 65.845 61.285 ;
        RECT 66.460 61.240 66.780 61.300 ;
        RECT 65.555 61.100 66.780 61.240 ;
        RECT 65.555 61.055 65.845 61.100 ;
        RECT 66.460 61.040 66.780 61.100 ;
        RECT 69.220 61.040 69.540 61.300 ;
        RECT 73.360 61.040 73.680 61.300 ;
        RECT 76.595 61.240 76.885 61.285 ;
        RECT 79.430 61.240 79.570 61.720 ;
        RECT 105.100 61.580 105.420 61.640 ;
        RECT 81.960 61.440 84.630 61.580 ;
        RECT 76.595 61.100 79.570 61.240 ;
        RECT 76.595 61.055 76.885 61.100 ;
        RECT 80.720 61.040 81.040 61.300 ;
        RECT 81.960 61.240 82.100 61.440 ;
        RECT 84.490 61.300 84.630 61.440 ;
        RECT 105.100 61.440 108.090 61.580 ;
        RECT 105.100 61.380 105.420 61.440 ;
        RECT 81.270 61.100 82.100 61.240 ;
        RECT 82.575 61.240 82.865 61.285 ;
        RECT 83.020 61.240 83.340 61.300 ;
        RECT 82.575 61.100 83.340 61.240 ;
        RECT 37.040 60.900 37.330 60.945 ;
        RECT 39.380 60.900 39.670 60.945 ;
        RECT 37.040 60.760 39.670 60.900 ;
        RECT 37.040 60.715 37.330 60.760 ;
        RECT 39.380 60.715 39.670 60.760 ;
        RECT 43.020 60.900 43.310 60.945 ;
        RECT 45.360 60.900 45.650 60.945 ;
        RECT 43.020 60.760 45.650 60.900 ;
        RECT 43.020 60.715 43.310 60.760 ;
        RECT 45.360 60.715 45.650 60.760 ;
        RECT 54.055 60.715 54.345 60.945 ;
        RECT 54.520 60.900 54.810 60.945 ;
        RECT 56.860 60.900 57.150 60.945 ;
        RECT 54.520 60.760 57.150 60.900 ;
        RECT 54.520 60.715 54.810 60.760 ;
        RECT 56.860 60.715 57.150 60.760 ;
        RECT 60.020 60.700 60.340 60.960 ;
        RECT 60.500 60.900 60.790 60.945 ;
        RECT 62.840 60.900 63.130 60.945 ;
        RECT 60.500 60.760 63.130 60.900 ;
        RECT 60.500 60.715 60.790 60.760 ;
        RECT 62.840 60.715 63.130 60.760 ;
        RECT 67.395 60.900 67.685 60.945 ;
        RECT 67.855 60.900 68.145 60.945 ;
        RECT 67.395 60.760 68.145 60.900 ;
        RECT 67.395 60.715 67.685 60.760 ;
        RECT 67.855 60.715 68.145 60.760 ;
        RECT 68.320 60.900 68.610 60.945 ;
        RECT 70.660 60.900 70.950 60.945 ;
        RECT 68.320 60.760 70.950 60.900 ;
        RECT 68.320 60.715 68.610 60.760 ;
        RECT 70.660 60.715 70.950 60.760 ;
        RECT 75.200 60.700 75.520 60.960 ;
        RECT 81.270 60.945 81.410 61.100 ;
        RECT 82.575 61.055 82.865 61.100 ;
        RECT 83.020 61.040 83.340 61.100 ;
        RECT 84.400 61.040 84.720 61.300 ;
        RECT 86.715 61.240 87.005 61.285 ;
        RECT 88.080 61.240 88.400 61.300 ;
        RECT 86.715 61.100 88.400 61.240 ;
        RECT 86.715 61.055 87.005 61.100 ;
        RECT 88.080 61.040 88.400 61.100 ;
        RECT 88.540 61.040 88.860 61.300 ;
        RECT 92.680 61.040 93.000 61.300 ;
        RECT 93.140 61.040 93.460 61.300 ;
        RECT 94.520 61.040 94.840 61.300 ;
        RECT 98.660 61.040 98.980 61.300 ;
        RECT 99.120 61.240 99.440 61.300 ;
        RECT 101.895 61.240 102.185 61.285 ;
        RECT 99.120 61.100 102.185 61.240 ;
        RECT 99.120 61.040 99.440 61.100 ;
        RECT 101.895 61.055 102.185 61.100 ;
        RECT 103.720 61.240 104.040 61.300 ;
        RECT 106.035 61.240 106.325 61.285 ;
        RECT 103.720 61.100 106.325 61.240 ;
        RECT 103.720 61.040 104.040 61.100 ;
        RECT 106.035 61.055 106.325 61.100 ;
        RECT 106.480 61.040 106.800 61.300 ;
        RECT 107.950 61.285 108.090 61.440 ;
        RECT 107.875 61.055 108.165 61.285 ;
        RECT 108.780 61.240 109.100 61.300 ;
        RECT 112.015 61.240 112.305 61.285 ;
        RECT 108.780 61.100 112.305 61.240 ;
        RECT 108.780 61.040 109.100 61.100 ;
        RECT 112.015 61.055 112.305 61.100 ;
        RECT 112.460 61.040 112.780 61.300 ;
        RECT 116.600 61.040 116.920 61.300 ;
        RECT 118.530 61.240 118.670 61.720 ;
        RECT 119.360 61.580 119.680 61.640 ;
        RECT 124.970 61.580 125.110 61.720 ;
        RECT 130.400 61.580 130.720 61.640 ;
        RECT 134.170 61.580 134.310 61.720 ;
        RECT 119.360 61.440 124.190 61.580 ;
        RECT 124.970 61.440 127.870 61.580 ;
        RECT 119.360 61.380 119.680 61.440 ;
        RECT 124.050 61.285 124.190 61.440 ;
        RECT 119.835 61.240 120.125 61.285 ;
        RECT 118.530 61.100 120.125 61.240 ;
        RECT 119.835 61.055 120.125 61.100 ;
        RECT 123.975 61.055 124.265 61.285 ;
        RECT 126.275 61.240 126.565 61.285 ;
        RECT 127.180 61.240 127.500 61.300 ;
        RECT 127.730 61.285 127.870 61.440 ;
        RECT 130.400 61.440 133.850 61.580 ;
        RECT 134.170 61.440 139.830 61.580 ;
        RECT 130.400 61.380 130.720 61.440 ;
        RECT 126.275 61.100 127.500 61.240 ;
        RECT 126.275 61.055 126.565 61.100 ;
        RECT 127.180 61.040 127.500 61.100 ;
        RECT 127.655 61.055 127.945 61.285 ;
        RECT 129.940 61.240 130.260 61.300 ;
        RECT 133.710 61.285 133.850 61.440 ;
        RECT 131.795 61.240 132.085 61.285 ;
        RECT 129.940 61.100 132.085 61.240 ;
        RECT 129.940 61.040 130.260 61.100 ;
        RECT 131.795 61.055 132.085 61.100 ;
        RECT 133.635 61.055 133.925 61.285 ;
        RECT 134.080 61.240 134.400 61.300 ;
        RECT 139.690 61.285 139.830 61.440 ;
        RECT 137.775 61.240 138.065 61.285 ;
        RECT 134.080 61.100 138.065 61.240 ;
        RECT 134.080 61.040 134.400 61.100 ;
        RECT 137.775 61.055 138.065 61.100 ;
        RECT 139.615 61.055 139.905 61.285 ;
        RECT 141.440 61.240 141.760 61.300 ;
        RECT 143.755 61.240 144.045 61.285 ;
        RECT 141.440 61.100 144.045 61.240 ;
        RECT 141.440 61.040 141.760 61.100 ;
        RECT 143.755 61.055 144.045 61.100 ;
        RECT 145.580 61.040 145.900 61.300 ;
        RECT 147.420 61.240 147.740 61.300 ;
        RECT 149.735 61.240 150.025 61.285 ;
        RECT 147.420 61.100 150.025 61.240 ;
        RECT 147.420 61.040 147.740 61.100 ;
        RECT 149.735 61.055 150.025 61.100 ;
        RECT 75.680 60.900 75.970 60.945 ;
        RECT 78.020 60.900 78.310 60.945 ;
        RECT 75.680 60.760 78.310 60.900 ;
        RECT 75.680 60.715 75.970 60.760 ;
        RECT 78.020 60.715 78.310 60.760 ;
        RECT 81.195 60.715 81.485 60.945 ;
        RECT 81.660 60.900 81.950 60.945 ;
        RECT 84.000 60.900 84.290 60.945 ;
        RECT 81.660 60.760 84.290 60.900 ;
        RECT 81.660 60.715 81.950 60.760 ;
        RECT 84.000 60.715 84.290 60.760 ;
        RECT 87.160 60.700 87.480 60.960 ;
        RECT 87.640 60.900 87.930 60.945 ;
        RECT 89.980 60.900 90.270 60.945 ;
        RECT 87.640 60.760 90.270 60.900 ;
        RECT 87.640 60.715 87.930 60.760 ;
        RECT 89.980 60.715 90.270 60.760 ;
        RECT 93.620 60.900 93.910 60.945 ;
        RECT 95.960 60.900 96.250 60.945 ;
        RECT 93.620 60.760 96.250 60.900 ;
        RECT 93.620 60.715 93.910 60.760 ;
        RECT 95.960 60.715 96.250 60.760 ;
        RECT 100.500 60.700 100.820 60.960 ;
        RECT 100.980 60.900 101.270 60.945 ;
        RECT 103.320 60.900 103.610 60.945 ;
        RECT 100.980 60.760 103.610 60.900 ;
        RECT 100.980 60.715 101.270 60.760 ;
        RECT 103.320 60.715 103.610 60.760 ;
        RECT 106.960 60.900 107.250 60.945 ;
        RECT 109.300 60.900 109.590 60.945 ;
        RECT 106.960 60.760 109.590 60.900 ;
        RECT 106.960 60.715 107.250 60.760 ;
        RECT 109.300 60.715 109.590 60.760 ;
        RECT 115.190 60.900 115.480 60.945 ;
        RECT 117.530 60.900 117.820 60.945 ;
        RECT 115.190 60.760 117.820 60.900 ;
        RECT 115.190 60.715 115.480 60.760 ;
        RECT 117.530 60.715 117.820 60.760 ;
        RECT 117.995 60.715 118.285 60.945 ;
        RECT 25.540 60.560 25.830 60.605 ;
        RECT 26.960 60.560 27.250 60.605 ;
        RECT 25.540 60.420 27.250 60.560 ;
        RECT 25.540 60.375 25.830 60.420 ;
        RECT 26.960 60.375 27.250 60.420 ;
        RECT 31.520 60.560 31.810 60.605 ;
        RECT 32.940 60.560 33.230 60.605 ;
        RECT 31.520 60.420 33.230 60.560 ;
        RECT 31.520 60.375 31.810 60.420 ;
        RECT 32.940 60.375 33.230 60.420 ;
        RECT 37.500 60.560 37.790 60.605 ;
        RECT 38.920 60.560 39.210 60.605 ;
        RECT 37.500 60.420 39.210 60.560 ;
        RECT 37.500 60.375 37.790 60.420 ;
        RECT 38.920 60.375 39.210 60.420 ;
        RECT 43.480 60.560 43.770 60.605 ;
        RECT 44.900 60.560 45.190 60.605 ;
        RECT 43.480 60.420 45.190 60.560 ;
        RECT 43.480 60.375 43.770 60.420 ;
        RECT 44.900 60.375 45.190 60.420 ;
        RECT 54.980 60.560 55.270 60.605 ;
        RECT 56.400 60.560 56.690 60.605 ;
        RECT 54.980 60.420 56.690 60.560 ;
        RECT 54.980 60.375 55.270 60.420 ;
        RECT 56.400 60.375 56.690 60.420 ;
        RECT 60.960 60.560 61.250 60.605 ;
        RECT 62.380 60.560 62.670 60.605 ;
        RECT 60.960 60.420 62.670 60.560 ;
        RECT 60.960 60.375 61.250 60.420 ;
        RECT 62.380 60.375 62.670 60.420 ;
        RECT 68.780 60.560 69.070 60.605 ;
        RECT 70.200 60.560 70.490 60.605 ;
        RECT 68.780 60.420 70.490 60.560 ;
        RECT 68.780 60.375 69.070 60.420 ;
        RECT 70.200 60.375 70.490 60.420 ;
        RECT 76.140 60.560 76.430 60.605 ;
        RECT 77.560 60.560 77.850 60.605 ;
        RECT 76.140 60.420 77.850 60.560 ;
        RECT 76.140 60.375 76.430 60.420 ;
        RECT 77.560 60.375 77.850 60.420 ;
        RECT 82.120 60.560 82.410 60.605 ;
        RECT 83.540 60.560 83.830 60.605 ;
        RECT 82.120 60.420 83.830 60.560 ;
        RECT 82.120 60.375 82.410 60.420 ;
        RECT 83.540 60.375 83.830 60.420 ;
        RECT 88.100 60.560 88.390 60.605 ;
        RECT 89.520 60.560 89.810 60.605 ;
        RECT 88.100 60.420 89.810 60.560 ;
        RECT 88.100 60.375 88.390 60.420 ;
        RECT 89.520 60.375 89.810 60.420 ;
        RECT 94.080 60.560 94.370 60.605 ;
        RECT 95.500 60.560 95.790 60.605 ;
        RECT 94.080 60.420 95.790 60.560 ;
        RECT 94.080 60.375 94.370 60.420 ;
        RECT 95.500 60.375 95.790 60.420 ;
        RECT 101.440 60.560 101.730 60.605 ;
        RECT 102.860 60.560 103.150 60.605 ;
        RECT 101.440 60.420 103.150 60.560 ;
        RECT 101.440 60.375 101.730 60.420 ;
        RECT 102.860 60.375 103.150 60.420 ;
        RECT 107.420 60.560 107.710 60.605 ;
        RECT 108.840 60.560 109.130 60.605 ;
        RECT 107.420 60.420 109.130 60.560 ;
        RECT 107.420 60.375 107.710 60.420 ;
        RECT 108.840 60.375 109.130 60.420 ;
        RECT 115.650 60.560 115.940 60.605 ;
        RECT 117.070 60.560 117.360 60.605 ;
        RECT 115.650 60.420 117.360 60.560 ;
        RECT 115.650 60.375 115.940 60.420 ;
        RECT 117.070 60.375 117.360 60.420 ;
        RECT 51.280 60.020 51.600 60.280 ;
        RECT 53.580 60.020 53.900 60.280 ;
        RECT 109.240 60.220 109.560 60.280 ;
        RECT 118.070 60.220 118.210 60.715 ;
        RECT 118.440 60.700 118.760 60.960 ;
        RECT 118.920 60.900 119.210 60.945 ;
        RECT 121.260 60.900 121.550 60.945 ;
        RECT 118.920 60.760 121.550 60.900 ;
        RECT 118.920 60.715 119.210 60.760 ;
        RECT 121.260 60.715 121.550 60.760 ;
        RECT 126.740 60.900 127.030 60.945 ;
        RECT 129.080 60.900 129.370 60.945 ;
        RECT 126.740 60.760 129.370 60.900 ;
        RECT 126.740 60.715 127.030 60.760 ;
        RECT 129.080 60.715 129.370 60.760 ;
        RECT 132.240 60.700 132.560 60.960 ;
        RECT 132.720 60.900 133.010 60.945 ;
        RECT 135.060 60.900 135.350 60.945 ;
        RECT 132.720 60.760 135.350 60.900 ;
        RECT 132.720 60.715 133.010 60.760 ;
        RECT 135.060 60.715 135.350 60.760 ;
        RECT 138.220 60.700 138.540 60.960 ;
        RECT 138.700 60.900 138.990 60.945 ;
        RECT 141.040 60.900 141.330 60.945 ;
        RECT 138.700 60.760 141.330 60.900 ;
        RECT 138.700 60.715 138.990 60.760 ;
        RECT 141.040 60.715 141.330 60.760 ;
        RECT 144.200 60.700 144.520 60.960 ;
        RECT 144.680 60.900 144.970 60.945 ;
        RECT 147.020 60.900 147.310 60.945 ;
        RECT 144.680 60.760 147.310 60.900 ;
        RECT 144.680 60.715 144.970 60.760 ;
        RECT 147.020 60.715 147.310 60.760 ;
        RECT 119.380 60.560 119.670 60.605 ;
        RECT 120.800 60.560 121.090 60.605 ;
        RECT 119.380 60.420 121.090 60.560 ;
        RECT 119.380 60.375 119.670 60.420 ;
        RECT 120.800 60.375 121.090 60.420 ;
        RECT 127.200 60.560 127.490 60.605 ;
        RECT 128.620 60.560 128.910 60.605 ;
        RECT 127.200 60.420 128.910 60.560 ;
        RECT 127.200 60.375 127.490 60.420 ;
        RECT 128.620 60.375 128.910 60.420 ;
        RECT 133.180 60.560 133.470 60.605 ;
        RECT 134.600 60.560 134.890 60.605 ;
        RECT 133.180 60.420 134.890 60.560 ;
        RECT 133.180 60.375 133.470 60.420 ;
        RECT 134.600 60.375 134.890 60.420 ;
        RECT 139.160 60.560 139.450 60.605 ;
        RECT 140.580 60.560 140.870 60.605 ;
        RECT 139.160 60.420 140.870 60.560 ;
        RECT 139.160 60.375 139.450 60.420 ;
        RECT 140.580 60.375 140.870 60.420 ;
        RECT 145.140 60.560 145.430 60.605 ;
        RECT 146.560 60.560 146.850 60.605 ;
        RECT 145.140 60.420 146.850 60.560 ;
        RECT 145.140 60.375 145.430 60.420 ;
        RECT 146.560 60.375 146.850 60.420 ;
        RECT 109.240 60.080 118.210 60.220 ;
        RECT 109.240 60.020 109.560 60.080 ;
        RECT 125.340 60.020 125.660 60.280 ;
        RECT 22.690 59.400 157.010 59.880 ;
        RECT 30.580 59.200 30.900 59.260 ;
        RECT 31.055 59.200 31.345 59.245 ;
        RECT 30.580 59.060 31.345 59.200 ;
        RECT 30.580 59.000 30.900 59.060 ;
        RECT 31.055 59.015 31.345 59.060 ;
        RECT 40.700 59.000 41.020 59.260 ;
        RECT 51.280 59.200 51.600 59.260 ;
        RECT 49.530 59.060 51.600 59.200 ;
        RECT 25.540 58.860 25.830 58.905 ;
        RECT 26.960 58.860 27.250 58.905 ;
        RECT 25.540 58.720 27.250 58.860 ;
        RECT 25.540 58.675 25.830 58.720 ;
        RECT 26.960 58.675 27.250 58.720 ;
        RECT 37.040 58.860 37.330 58.905 ;
        RECT 38.460 58.860 38.750 58.905 ;
        RECT 37.040 58.720 38.750 58.860 ;
        RECT 37.040 58.675 37.330 58.720 ;
        RECT 38.460 58.675 38.750 58.720 ;
        RECT 24.600 58.320 24.920 58.580 ;
        RECT 25.080 58.520 25.370 58.565 ;
        RECT 27.420 58.520 27.710 58.565 ;
        RECT 25.080 58.380 27.710 58.520 ;
        RECT 25.080 58.335 25.370 58.380 ;
        RECT 27.420 58.335 27.710 58.380 ;
        RECT 36.580 58.520 36.870 58.565 ;
        RECT 38.920 58.520 39.210 58.565 ;
        RECT 36.580 58.380 39.210 58.520 ;
        RECT 40.790 58.520 40.930 59.000 ;
        RECT 43.020 58.860 43.310 58.905 ;
        RECT 44.440 58.860 44.730 58.905 ;
        RECT 43.020 58.720 44.730 58.860 ;
        RECT 43.020 58.675 43.310 58.720 ;
        RECT 44.440 58.675 44.730 58.720 ;
        RECT 49.530 58.565 49.670 59.060 ;
        RECT 51.280 59.000 51.600 59.060 ;
        RECT 53.580 59.000 53.900 59.260 ;
        RECT 60.020 59.200 60.340 59.260 ;
        RECT 61.875 59.200 62.165 59.245 ;
        RECT 60.020 59.060 62.165 59.200 ;
        RECT 60.020 59.000 60.340 59.060 ;
        RECT 61.875 59.015 62.165 59.060 ;
        RECT 71.520 59.200 71.840 59.260 ;
        RECT 72.915 59.200 73.205 59.245 ;
        RECT 71.520 59.060 73.205 59.200 ;
        RECT 71.520 59.000 71.840 59.060 ;
        RECT 72.915 59.015 73.205 59.060 ;
        RECT 75.200 59.200 75.520 59.260 ;
        RECT 76.135 59.200 76.425 59.245 ;
        RECT 75.200 59.060 76.425 59.200 ;
        RECT 75.200 59.000 75.520 59.060 ;
        RECT 76.135 59.015 76.425 59.060 ;
        RECT 78.420 59.000 78.740 59.260 ;
        RECT 85.780 59.200 86.100 59.260 ;
        RECT 81.270 59.060 86.100 59.200 ;
        RECT 50.380 58.860 50.670 58.905 ;
        RECT 51.800 58.860 52.090 58.905 ;
        RECT 50.380 58.720 52.090 58.860 ;
        RECT 50.380 58.675 50.670 58.720 ;
        RECT 51.800 58.675 52.090 58.720 ;
        RECT 42.095 58.520 42.385 58.565 ;
        RECT 40.790 58.380 42.385 58.520 ;
        RECT 36.580 58.335 36.870 58.380 ;
        RECT 38.920 58.335 39.210 58.380 ;
        RECT 42.095 58.335 42.385 58.380 ;
        RECT 42.560 58.520 42.850 58.565 ;
        RECT 44.900 58.520 45.190 58.565 ;
        RECT 42.560 58.380 45.190 58.520 ;
        RECT 42.560 58.335 42.850 58.380 ;
        RECT 44.900 58.335 45.190 58.380 ;
        RECT 49.455 58.335 49.745 58.565 ;
        RECT 49.920 58.520 50.210 58.565 ;
        RECT 52.260 58.520 52.550 58.565 ;
        RECT 49.920 58.380 52.550 58.520 ;
        RECT 53.670 58.520 53.810 59.000 ;
        RECT 56.360 58.860 56.650 58.905 ;
        RECT 57.780 58.860 58.070 58.905 ;
        RECT 56.360 58.720 58.070 58.860 ;
        RECT 56.360 58.675 56.650 58.720 ;
        RECT 57.780 58.675 58.070 58.720 ;
        RECT 66.940 58.860 67.230 58.905 ;
        RECT 68.360 58.860 68.650 58.905 ;
        RECT 66.940 58.720 68.650 58.860 ;
        RECT 66.940 58.675 67.230 58.720 ;
        RECT 68.360 58.675 68.650 58.720 ;
        RECT 55.435 58.520 55.725 58.565 ;
        RECT 53.670 58.380 55.725 58.520 ;
        RECT 49.920 58.335 50.210 58.380 ;
        RECT 52.260 58.335 52.550 58.380 ;
        RECT 55.435 58.335 55.725 58.380 ;
        RECT 55.900 58.520 56.190 58.565 ;
        RECT 58.240 58.520 58.530 58.565 ;
        RECT 55.900 58.380 58.530 58.520 ;
        RECT 55.900 58.335 56.190 58.380 ;
        RECT 58.240 58.335 58.530 58.380 ;
        RECT 66.000 58.320 66.320 58.580 ;
        RECT 81.270 58.565 81.410 59.060 ;
        RECT 85.780 59.000 86.100 59.060 ;
        RECT 87.160 59.200 87.480 59.260 ;
        RECT 87.635 59.200 87.925 59.245 ;
        RECT 87.160 59.060 87.925 59.200 ;
        RECT 87.160 59.000 87.480 59.060 ;
        RECT 87.635 59.015 87.925 59.060 ;
        RECT 90.840 59.000 91.160 59.260 ;
        RECT 98.675 59.200 98.965 59.245 ;
        RECT 100.500 59.200 100.820 59.260 ;
        RECT 98.675 59.060 100.820 59.200 ;
        RECT 98.675 59.015 98.965 59.060 ;
        RECT 100.500 59.000 100.820 59.060 ;
        RECT 109.240 59.000 109.560 59.260 ;
        RECT 112.475 59.200 112.765 59.245 ;
        RECT 118.440 59.200 118.760 59.260 ;
        RECT 112.475 59.060 118.760 59.200 ;
        RECT 112.475 59.015 112.765 59.060 ;
        RECT 118.440 59.000 118.760 59.060 ;
        RECT 125.340 59.000 125.660 59.260 ;
        RECT 129.480 59.200 129.800 59.260 ;
        RECT 126.350 59.060 129.800 59.200 ;
        RECT 82.120 58.860 82.410 58.905 ;
        RECT 83.540 58.860 83.830 58.905 ;
        RECT 90.930 58.860 91.070 59.000 ;
        RECT 82.120 58.720 83.830 58.860 ;
        RECT 82.120 58.675 82.410 58.720 ;
        RECT 83.540 58.675 83.830 58.720 ;
        RECT 90.470 58.720 91.070 58.860 ;
        RECT 91.320 58.860 91.610 58.905 ;
        RECT 92.740 58.860 93.030 58.905 ;
        RECT 91.320 58.720 93.030 58.860 ;
        RECT 90.470 58.565 90.610 58.720 ;
        RECT 91.320 58.675 91.610 58.720 ;
        RECT 92.740 58.675 93.030 58.720 ;
        RECT 101.900 58.860 102.190 58.905 ;
        RECT 103.320 58.860 103.610 58.905 ;
        RECT 101.900 58.720 103.610 58.860 ;
        RECT 101.900 58.675 102.190 58.720 ;
        RECT 103.320 58.675 103.610 58.720 ;
        RECT 114.320 58.860 114.610 58.905 ;
        RECT 115.740 58.860 116.030 58.905 ;
        RECT 114.320 58.720 116.030 58.860 ;
        RECT 114.320 58.675 114.610 58.720 ;
        RECT 115.740 58.675 116.030 58.720 ;
        RECT 122.550 58.860 122.840 58.905 ;
        RECT 123.970 58.860 124.260 58.905 ;
        RECT 122.550 58.720 124.260 58.860 ;
        RECT 122.550 58.675 122.840 58.720 ;
        RECT 123.970 58.675 124.260 58.720 ;
        RECT 66.480 58.520 66.770 58.565 ;
        RECT 68.820 58.520 69.110 58.565 ;
        RECT 66.480 58.380 69.110 58.520 ;
        RECT 66.480 58.335 66.770 58.380 ;
        RECT 68.820 58.335 69.110 58.380 ;
        RECT 81.195 58.335 81.485 58.565 ;
        RECT 81.660 58.520 81.950 58.565 ;
        RECT 84.000 58.520 84.290 58.565 ;
        RECT 81.660 58.380 84.290 58.520 ;
        RECT 81.660 58.335 81.950 58.380 ;
        RECT 84.000 58.335 84.290 58.380 ;
        RECT 90.395 58.335 90.685 58.565 ;
        RECT 90.860 58.520 91.150 58.565 ;
        RECT 93.200 58.520 93.490 58.565 ;
        RECT 90.860 58.380 93.490 58.520 ;
        RECT 90.860 58.335 91.150 58.380 ;
        RECT 93.200 58.335 93.490 58.380 ;
        RECT 101.440 58.520 101.730 58.565 ;
        RECT 103.780 58.520 104.070 58.565 ;
        RECT 101.440 58.380 104.070 58.520 ;
        RECT 101.440 58.335 101.730 58.380 ;
        RECT 103.780 58.335 104.070 58.380 ;
        RECT 111.095 58.520 111.385 58.565 ;
        RECT 113.395 58.520 113.685 58.565 ;
        RECT 111.095 58.380 113.685 58.520 ;
        RECT 111.095 58.335 111.385 58.380 ;
        RECT 113.395 58.335 113.685 58.380 ;
        RECT 113.860 58.520 114.150 58.565 ;
        RECT 116.200 58.520 116.490 58.565 ;
        RECT 113.860 58.380 116.490 58.520 ;
        RECT 113.860 58.335 114.150 58.380 ;
        RECT 116.200 58.335 116.490 58.380 ;
        RECT 122.090 58.520 122.380 58.565 ;
        RECT 124.430 58.520 124.720 58.565 ;
        RECT 122.090 58.380 124.720 58.520 ;
        RECT 122.090 58.335 122.380 58.380 ;
        RECT 124.430 58.335 124.720 58.380 ;
        RECT 124.895 58.520 125.185 58.565 ;
        RECT 125.430 58.520 125.570 59.000 ;
        RECT 126.350 58.565 126.490 59.060 ;
        RECT 129.480 59.000 129.800 59.060 ;
        RECT 132.240 59.000 132.560 59.260 ;
        RECT 132.700 59.200 133.020 59.260 ;
        RECT 133.635 59.200 133.925 59.245 ;
        RECT 132.700 59.060 133.925 59.200 ;
        RECT 132.700 59.000 133.020 59.060 ;
        RECT 133.635 59.015 133.925 59.060 ;
        RECT 135.935 59.200 136.225 59.245 ;
        RECT 138.220 59.200 138.540 59.260 ;
        RECT 135.935 59.060 138.540 59.200 ;
        RECT 135.935 59.015 136.225 59.060 ;
        RECT 138.220 59.000 138.540 59.060 ;
        RECT 144.200 59.200 144.520 59.260 ;
        RECT 145.135 59.200 145.425 59.245 ;
        RECT 144.200 59.060 145.425 59.200 ;
        RECT 144.200 59.000 144.520 59.060 ;
        RECT 145.135 59.015 145.425 59.060 ;
        RECT 146.500 59.000 146.820 59.260 ;
        RECT 127.200 58.860 127.490 58.905 ;
        RECT 128.620 58.860 128.910 58.905 ;
        RECT 127.200 58.720 128.910 58.860 ;
        RECT 127.200 58.675 127.490 58.720 ;
        RECT 128.620 58.675 128.910 58.720 ;
        RECT 140.080 58.860 140.370 58.905 ;
        RECT 141.500 58.860 141.790 58.905 ;
        RECT 140.080 58.720 141.790 58.860 ;
        RECT 140.080 58.675 140.370 58.720 ;
        RECT 141.500 58.675 141.790 58.720 ;
        RECT 124.895 58.380 125.570 58.520 ;
        RECT 124.895 58.335 125.185 58.380 ;
        RECT 126.275 58.335 126.565 58.565 ;
        RECT 126.740 58.520 127.030 58.565 ;
        RECT 129.080 58.520 129.370 58.565 ;
        RECT 126.740 58.380 129.370 58.520 ;
        RECT 126.740 58.335 127.030 58.380 ;
        RECT 129.080 58.335 129.370 58.380 ;
        RECT 138.680 58.520 139.000 58.580 ;
        RECT 139.155 58.520 139.445 58.565 ;
        RECT 138.680 58.380 139.445 58.520 ;
        RECT 138.680 58.320 139.000 58.380 ;
        RECT 139.155 58.335 139.445 58.380 ;
        RECT 139.620 58.520 139.910 58.565 ;
        RECT 141.960 58.520 142.250 58.565 ;
        RECT 139.620 58.380 142.250 58.520 ;
        RECT 139.620 58.335 139.910 58.380 ;
        RECT 141.960 58.335 142.250 58.380 ;
        RECT 25.995 57.995 26.285 58.225 ;
        RECT 28.740 58.180 29.060 58.240 ;
        RECT 30.135 58.180 30.425 58.225 ;
        RECT 28.740 58.040 30.425 58.180 ;
        RECT 26.070 57.840 26.210 57.995 ;
        RECT 28.740 57.980 29.060 58.040 ;
        RECT 30.135 57.995 30.425 58.040 ;
        RECT 32.420 57.980 32.740 58.240 ;
        RECT 35.195 58.180 35.485 58.225 ;
        RECT 36.115 58.180 36.405 58.225 ;
        RECT 35.195 58.040 36.405 58.180 ;
        RECT 35.195 57.995 35.485 58.040 ;
        RECT 36.115 57.995 36.405 58.040 ;
        RECT 37.495 58.180 37.785 58.225 ;
        RECT 37.940 58.180 38.260 58.240 ;
        RECT 37.495 58.040 38.260 58.180 ;
        RECT 37.495 57.995 37.785 58.040 ;
        RECT 37.940 57.980 38.260 58.040 ;
        RECT 40.240 58.180 40.560 58.240 ;
        RECT 41.635 58.180 41.925 58.225 ;
        RECT 40.240 58.040 41.925 58.180 ;
        RECT 40.240 57.980 40.560 58.040 ;
        RECT 41.635 57.995 41.925 58.040 ;
        RECT 43.000 58.180 43.320 58.240 ;
        RECT 43.475 58.180 43.765 58.225 ;
        RECT 43.000 58.040 43.765 58.180 ;
        RECT 43.000 57.980 43.320 58.040 ;
        RECT 43.475 57.995 43.765 58.040 ;
        RECT 47.600 57.980 47.920 58.240 ;
        RECT 50.360 58.180 50.680 58.240 ;
        RECT 50.835 58.180 51.125 58.225 ;
        RECT 50.360 58.040 51.125 58.180 ;
        RECT 50.360 57.980 50.680 58.040 ;
        RECT 50.835 57.995 51.125 58.040 ;
        RECT 54.960 57.980 55.280 58.240 ;
        RECT 56.800 57.980 57.120 58.240 ;
        RECT 60.955 58.180 61.245 58.225 ;
        RECT 61.400 58.180 61.720 58.240 ;
        RECT 60.955 58.040 61.720 58.180 ;
        RECT 60.955 57.995 61.245 58.040 ;
        RECT 61.400 57.980 61.720 58.040 ;
        RECT 67.395 58.180 67.685 58.225 ;
        RECT 68.300 58.180 68.620 58.240 ;
        RECT 67.395 58.040 68.620 58.180 ;
        RECT 67.395 57.995 67.685 58.040 ;
        RECT 68.300 57.980 68.620 58.040 ;
        RECT 70.140 58.180 70.460 58.240 ;
        RECT 71.535 58.180 71.825 58.225 ;
        RECT 70.140 58.040 71.825 58.180 ;
        RECT 70.140 57.980 70.460 58.040 ;
        RECT 71.535 57.995 71.825 58.040 ;
        RECT 82.575 58.180 82.865 58.225 ;
        RECT 83.480 58.180 83.800 58.240 ;
        RECT 82.575 58.040 83.800 58.180 ;
        RECT 82.575 57.995 82.865 58.040 ;
        RECT 83.480 57.980 83.800 58.040 ;
        RECT 86.700 57.980 87.020 58.240 ;
        RECT 91.775 58.180 92.065 58.225 ;
        RECT 94.060 58.180 94.380 58.240 ;
        RECT 91.775 58.040 94.380 58.180 ;
        RECT 91.775 57.995 92.065 58.040 ;
        RECT 94.060 57.980 94.380 58.040 ;
        RECT 94.980 58.180 95.300 58.240 ;
        RECT 95.915 58.180 96.205 58.225 ;
        RECT 94.980 58.040 96.205 58.180 ;
        RECT 94.980 57.980 95.300 58.040 ;
        RECT 95.915 57.995 96.205 58.040 ;
        RECT 100.975 58.180 101.265 58.225 ;
        RECT 101.880 58.180 102.200 58.240 ;
        RECT 100.975 58.040 102.200 58.180 ;
        RECT 100.975 57.995 101.265 58.040 ;
        RECT 101.880 57.980 102.200 58.040 ;
        RECT 102.355 57.995 102.645 58.225 ;
        RECT 32.510 57.840 32.650 57.980 ;
        RECT 26.070 57.700 32.650 57.840 ;
        RECT 99.580 57.840 99.900 57.900 ;
        RECT 102.430 57.840 102.570 57.995 ;
        RECT 106.480 57.980 106.800 58.240 ;
        RECT 114.760 57.980 115.080 58.240 ;
        RECT 116.600 58.180 116.920 58.240 ;
        RECT 118.915 58.180 119.205 58.225 ;
        RECT 116.600 58.040 119.205 58.180 ;
        RECT 116.600 57.980 116.920 58.040 ;
        RECT 118.915 57.995 119.205 58.040 ;
        RECT 119.375 58.180 119.665 58.225 ;
        RECT 121.200 58.180 121.520 58.240 ;
        RECT 119.375 58.040 121.520 58.180 ;
        RECT 119.375 57.995 119.665 58.040 ;
        RECT 121.200 57.980 121.520 58.040 ;
        RECT 121.660 58.180 121.980 58.240 ;
        RECT 123.515 58.180 123.805 58.225 ;
        RECT 121.660 58.040 123.805 58.180 ;
        RECT 121.660 57.980 121.980 58.040 ;
        RECT 123.515 57.995 123.805 58.040 ;
        RECT 127.640 57.980 127.960 58.240 ;
        RECT 131.780 57.980 132.100 58.240 ;
        RECT 137.760 58.180 138.080 58.240 ;
        RECT 140.535 58.180 140.825 58.225 ;
        RECT 137.760 58.040 140.825 58.180 ;
        RECT 137.760 57.980 138.080 58.040 ;
        RECT 140.535 57.995 140.825 58.040 ;
        RECT 144.660 57.980 144.980 58.240 ;
        RECT 99.580 57.700 102.570 57.840 ;
        RECT 99.580 57.640 99.900 57.700 ;
        RECT 22.690 56.680 157.810 57.160 ;
        RECT 114.980 52.000 115.830 52.015 ;
        RECT 120.065 52.000 120.875 52.055 ;
        RECT 122.030 52.000 122.780 52.005 ;
        RECT 124.675 52.000 125.485 52.025 ;
        RECT 132.755 52.000 133.505 52.005 ;
        RECT 136.755 52.000 137.505 52.055 ;
        RECT 138.620 52.000 139.430 52.025 ;
        RECT 142.555 52.000 143.305 52.055 ;
        RECT 75.100 50.600 75.950 50.615 ;
        RECT 80.185 50.600 80.995 50.655 ;
        RECT 82.150 50.600 82.900 50.605 ;
        RECT 84.795 50.600 85.605 50.625 ;
        RECT 92.875 50.600 93.625 50.605 ;
        RECT 96.875 50.600 97.625 50.655 ;
        RECT 98.740 50.600 99.550 50.625 ;
        RECT 102.675 50.600 103.425 50.655 ;
        RECT 33.880 49.760 34.730 49.775 ;
        RECT 38.965 49.760 39.775 49.815 ;
        RECT 40.930 49.760 41.680 49.765 ;
        RECT 43.575 49.760 44.385 49.785 ;
        RECT 51.655 49.760 52.405 49.765 ;
        RECT 55.655 49.760 56.405 49.815 ;
        RECT 57.520 49.760 58.330 49.785 ;
        RECT 61.455 49.760 62.205 49.815 ;
        RECT 30.280 46.660 32.280 49.760 ;
        RECT 33.280 48.865 34.730 49.760 ;
        RECT 35.280 48.920 36.750 49.760 ;
        RECT 33.280 48.760 34.280 48.865 ;
        RECT 35.280 48.760 36.280 48.920 ;
        RECT 37.280 48.760 38.280 49.760 ;
        RECT 38.965 48.945 40.280 49.760 ;
        RECT 40.930 48.955 42.280 49.760 ;
        RECT 39.280 48.760 40.280 48.945 ;
        RECT 41.280 48.760 42.280 48.955 ;
        RECT 43.280 49.035 44.385 49.760 ;
        RECT 45.280 49.685 46.280 49.760 ;
        RECT 47.280 49.685 48.280 49.760 ;
        RECT 49.280 49.735 50.280 49.760 ;
        RECT 43.280 48.760 44.280 49.035 ;
        RECT 45.280 48.935 46.610 49.685 ;
        RECT 47.280 48.935 48.760 49.685 ;
        RECT 49.280 48.985 50.610 49.735 ;
        RECT 45.280 48.760 46.280 48.935 ;
        RECT 47.280 48.760 48.280 48.935 ;
        RECT 49.280 48.760 50.280 48.985 ;
        RECT 51.280 48.955 52.405 49.760 ;
        RECT 53.280 49.735 54.280 49.760 ;
        RECT 53.280 48.985 54.485 49.735 ;
        RECT 55.280 49.005 56.405 49.760 ;
        RECT 57.280 49.035 58.330 49.760 ;
        RECT 59.280 49.715 60.280 49.760 ;
        RECT 51.280 48.760 52.280 48.955 ;
        RECT 53.280 48.760 54.280 48.985 ;
        RECT 55.280 48.760 56.280 49.005 ;
        RECT 57.280 48.760 58.280 49.035 ;
        RECT 59.280 48.905 60.455 49.715 ;
        RECT 59.280 48.760 60.280 48.905 ;
        RECT 61.280 48.760 62.280 49.760 ;
        RECT 33.850 47.100 34.760 47.725 ;
        RECT 33.820 46.870 34.780 47.100 ;
        RECT 63.280 46.760 66.280 49.810 ;
        RECT 71.500 47.500 73.500 50.600 ;
        RECT 74.500 49.705 75.950 50.600 ;
        RECT 76.500 49.760 77.970 50.600 ;
        RECT 74.500 49.600 75.500 49.705 ;
        RECT 76.500 49.600 77.500 49.760 ;
        RECT 78.500 49.600 79.500 50.600 ;
        RECT 80.185 49.785 81.500 50.600 ;
        RECT 82.150 49.795 83.500 50.600 ;
        RECT 80.500 49.600 81.500 49.785 ;
        RECT 82.500 49.600 83.500 49.795 ;
        RECT 84.500 49.875 85.605 50.600 ;
        RECT 86.500 50.525 87.500 50.600 ;
        RECT 88.500 50.525 89.500 50.600 ;
        RECT 90.500 50.575 91.500 50.600 ;
        RECT 84.500 49.600 85.500 49.875 ;
        RECT 86.500 49.775 87.830 50.525 ;
        RECT 88.500 49.775 89.980 50.525 ;
        RECT 90.500 49.825 91.830 50.575 ;
        RECT 86.500 49.600 87.500 49.775 ;
        RECT 88.500 49.600 89.500 49.775 ;
        RECT 90.500 49.600 91.500 49.825 ;
        RECT 92.500 49.795 93.625 50.600 ;
        RECT 94.500 50.575 95.500 50.600 ;
        RECT 94.500 49.825 95.705 50.575 ;
        RECT 96.500 49.845 97.625 50.600 ;
        RECT 98.500 49.875 99.550 50.600 ;
        RECT 100.500 50.555 101.500 50.600 ;
        RECT 92.500 49.600 93.500 49.795 ;
        RECT 94.500 49.600 95.500 49.825 ;
        RECT 96.500 49.600 97.500 49.845 ;
        RECT 98.500 49.600 99.500 49.875 ;
        RECT 100.500 49.745 101.675 50.555 ;
        RECT 100.500 49.600 101.500 49.745 ;
        RECT 102.500 49.600 103.500 50.600 ;
        RECT 75.070 47.940 75.980 48.565 ;
        RECT 75.040 47.710 76.000 47.940 ;
        RECT 104.500 47.600 107.500 50.650 ;
        RECT 111.380 48.900 113.380 52.000 ;
        RECT 114.380 51.105 115.830 52.000 ;
        RECT 116.380 51.160 117.850 52.000 ;
        RECT 114.380 51.000 115.380 51.105 ;
        RECT 116.380 51.000 117.380 51.160 ;
        RECT 118.380 51.000 119.380 52.000 ;
        RECT 120.065 51.185 121.380 52.000 ;
        RECT 122.030 51.195 123.380 52.000 ;
        RECT 120.380 51.000 121.380 51.185 ;
        RECT 122.380 51.000 123.380 51.195 ;
        RECT 124.380 51.275 125.485 52.000 ;
        RECT 126.380 51.925 127.380 52.000 ;
        RECT 128.380 51.925 129.380 52.000 ;
        RECT 130.380 51.975 131.380 52.000 ;
        RECT 124.380 51.000 125.380 51.275 ;
        RECT 126.380 51.175 127.710 51.925 ;
        RECT 128.380 51.175 129.860 51.925 ;
        RECT 130.380 51.225 131.710 51.975 ;
        RECT 126.380 51.000 127.380 51.175 ;
        RECT 128.380 51.000 129.380 51.175 ;
        RECT 130.380 51.000 131.380 51.225 ;
        RECT 132.380 51.195 133.505 52.000 ;
        RECT 134.380 51.975 135.380 52.000 ;
        RECT 134.380 51.225 135.585 51.975 ;
        RECT 136.380 51.245 137.505 52.000 ;
        RECT 138.380 51.275 139.430 52.000 ;
        RECT 140.380 51.955 141.380 52.000 ;
        RECT 132.380 51.000 133.380 51.195 ;
        RECT 134.380 51.000 135.380 51.225 ;
        RECT 136.380 51.000 137.380 51.245 ;
        RECT 138.380 51.000 139.380 51.275 ;
        RECT 140.380 51.145 141.555 51.955 ;
        RECT 140.380 51.000 141.380 51.145 ;
        RECT 142.380 51.000 143.380 52.000 ;
        RECT 114.950 49.340 115.860 49.965 ;
        RECT 114.920 49.110 115.880 49.340 ;
        RECT 144.380 49.000 147.380 52.050 ;
        RECT 30.250 44.660 33.280 46.660 ;
        RECT 33.540 46.650 33.770 46.710 ;
        RECT 33.465 44.360 33.770 46.650 ;
        RECT 31.280 34.760 33.770 44.360 ;
        RECT 31.280 32.360 33.280 34.760 ;
        RECT 33.540 34.710 33.770 34.760 ;
        RECT 34.830 46.650 35.060 46.710 ;
        RECT 36.780 46.650 66.280 46.760 ;
        RECT 34.830 43.760 66.280 46.650 ;
        RECT 71.470 45.500 74.500 47.500 ;
        RECT 74.760 47.490 74.990 47.550 ;
        RECT 74.685 45.200 74.990 47.490 ;
        RECT 34.830 37.700 37.760 43.760 ;
        RECT 40.900 38.100 41.710 38.635 ;
        RECT 40.820 37.870 41.780 38.100 ;
        RECT 40.540 37.700 40.770 37.710 ;
        RECT 34.830 34.770 40.770 37.700 ;
        RECT 34.830 34.710 35.060 34.770 ;
        RECT 33.820 34.320 34.780 34.550 ;
        RECT 33.850 33.675 34.760 34.320 ;
        RECT 35.850 32.600 36.750 33.230 ;
        RECT 35.820 32.370 36.780 32.600 ;
        RECT 31.280 29.660 33.080 32.360 ;
        RECT 35.540 32.150 35.770 32.210 ;
        RECT 33.280 30.030 35.280 32.090 ;
        RECT 35.480 29.660 35.770 32.150 ;
        RECT 31.280 24.260 35.770 29.660 ;
        RECT 31.280 23.260 32.780 24.260 ;
        RECT 33.780 23.800 35.770 24.260 ;
        RECT 33.780 23.260 34.880 23.800 ;
        RECT 35.540 23.730 35.770 23.800 ;
        RECT 36.830 32.150 37.060 32.210 ;
        RECT 37.880 32.150 39.680 34.770 ;
        RECT 40.540 34.710 40.770 34.770 ;
        RECT 41.830 36.260 42.060 37.710 ;
        RECT 42.280 36.410 43.980 38.160 ;
        RECT 44.680 37.680 45.325 37.710 ;
        RECT 44.650 37.650 45.355 37.680 ;
        RECT 44.520 37.420 45.480 37.650 ;
        RECT 44.240 36.260 44.470 37.260 ;
        RECT 44.650 37.035 45.355 37.420 ;
        RECT 45.530 37.210 45.760 37.260 ;
        RECT 46.530 37.210 48.530 43.760 ;
        RECT 44.680 37.005 45.325 37.035 ;
        RECT 41.830 35.210 44.470 36.260 ;
        RECT 41.830 35.030 43.580 35.210 ;
        RECT 44.240 35.140 44.470 35.210 ;
        RECT 41.830 34.760 43.600 35.030 ;
        RECT 44.650 34.980 45.355 35.385 ;
        RECT 45.530 35.210 52.180 37.210 ;
        RECT 45.530 35.140 45.760 35.210 ;
        RECT 41.830 34.710 42.060 34.760 ;
        RECT 40.820 34.320 41.780 34.550 ;
        RECT 40.900 33.735 41.710 34.320 ;
        RECT 36.830 25.660 39.680 32.150 ;
        RECT 42.230 29.010 43.600 34.760 ;
        RECT 44.520 34.750 45.480 34.980 ;
        RECT 44.650 34.740 45.355 34.750 ;
        RECT 47.680 34.390 48.980 35.210 ;
        RECT 47.580 34.160 49.080 34.390 ;
        RECT 47.190 34.010 47.420 34.110 ;
        RECT 49.240 34.010 49.470 34.110 ;
        RECT 45.580 33.890 46.930 34.010 ;
        RECT 44.480 33.860 46.930 33.890 ;
        RECT 44.430 32.760 46.930 33.860 ;
        RECT 47.160 33.980 47.800 34.010 ;
        RECT 48.910 33.980 49.550 34.010 ;
        RECT 47.160 33.340 49.550 33.980 ;
        RECT 47.160 33.310 47.800 33.340 ;
        RECT 48.910 33.310 49.550 33.340 ;
        RECT 47.190 33.150 47.420 33.310 ;
        RECT 49.240 33.150 49.470 33.310 ;
        RECT 47.580 32.870 49.080 33.100 ;
        RECT 44.480 32.730 45.580 32.760 ;
        RECT 47.680 32.560 48.980 32.870 ;
        RECT 49.730 32.760 50.630 34.510 ;
        RECT 51.380 34.390 52.180 35.210 ;
        RECT 51.280 34.160 52.280 34.390 ;
        RECT 50.890 33.965 51.120 34.110 ;
        RECT 52.440 33.965 52.670 34.110 ;
        RECT 50.855 33.250 51.510 33.965 ;
        RECT 52.050 33.250 52.705 33.965 ;
        RECT 50.890 33.150 51.120 33.250 ;
        RECT 52.440 33.150 52.670 33.250 ;
        RECT 51.280 32.870 52.280 33.100 ;
        RECT 51.380 32.560 52.230 32.870 ;
        RECT 47.680 31.785 52.230 32.560 ;
        RECT 47.680 29.010 48.980 31.785 ;
        RECT 51.380 31.440 52.230 31.785 ;
        RECT 51.280 31.210 52.280 31.440 ;
        RECT 50.890 30.585 51.120 31.160 ;
        RECT 51.380 31.060 52.230 31.210 ;
        RECT 52.440 30.865 52.670 31.160 ;
        RECT 50.180 30.490 50.630 30.510 ;
        RECT 49.130 29.330 50.630 30.490 ;
        RECT 50.875 29.835 51.685 30.585 ;
        RECT 52.055 30.055 52.805 30.865 ;
        RECT 50.890 29.700 51.120 29.835 ;
        RECT 52.440 29.700 52.670 30.055 ;
        RECT 42.230 27.160 48.980 29.010 ;
        RECT 49.280 29.310 50.630 29.330 ;
        RECT 51.280 29.560 52.280 29.650 ;
        RECT 51.280 29.410 52.330 29.560 ;
        RECT 63.280 29.420 66.280 43.760 ;
        RECT 54.070 29.410 66.280 29.420 ;
        RECT 49.280 28.410 50.280 29.310 ;
        RECT 51.280 28.510 66.280 29.410 ;
        RECT 54.070 28.420 66.280 28.510 ;
        RECT 49.280 27.960 50.880 28.410 ;
        RECT 51.055 28.285 51.805 28.315 ;
        RECT 49.280 27.310 50.280 27.960 ;
        RECT 51.055 27.750 52.885 28.285 ;
        RECT 50.800 27.520 52.885 27.750 ;
        RECT 51.055 27.505 52.885 27.520 ;
        RECT 63.280 27.360 66.280 28.420 ;
        RECT 50.520 27.160 50.830 27.360 ;
        RECT 42.230 26.360 50.830 27.160 ;
        RECT 36.830 23.860 40.680 25.660 ;
        RECT 36.830 23.800 38.630 23.860 ;
        RECT 36.830 23.730 37.060 23.800 ;
        RECT 35.850 23.570 36.750 23.600 ;
        RECT 35.820 23.340 36.780 23.570 ;
        RECT 31.280 21.360 34.880 23.260 ;
        RECT 35.850 22.760 36.750 23.340 ;
        RECT 37.360 21.600 38.240 22.150 ;
        RECT 37.320 21.370 38.280 21.600 ;
        RECT 31.280 18.760 34.280 21.360 ;
        RECT 37.360 21.330 38.240 21.370 ;
        RECT 37.040 21.130 37.270 21.210 ;
        RECT 34.780 19.030 36.780 21.090 ;
        RECT 36.980 18.760 37.270 21.130 ;
        RECT 31.280 15.760 37.270 18.760 ;
        RECT 31.280 14.760 34.280 15.760 ;
        RECT 35.280 15.300 37.270 15.760 ;
        RECT 37.040 15.210 37.270 15.300 ;
        RECT 38.330 21.130 38.560 21.210 ;
        RECT 38.880 21.130 40.680 23.860 ;
        RECT 38.330 20.140 40.680 21.130 ;
        RECT 42.230 23.840 48.980 26.360 ;
        RECT 51.025 26.200 52.780 26.685 ;
        RECT 52.930 26.360 66.280 27.360 ;
        RECT 50.800 25.970 52.880 26.200 ;
        RECT 51.025 25.950 52.780 25.970 ;
        RECT 50.370 25.700 53.420 25.730 ;
        RECT 50.360 25.660 53.420 25.700 ;
        RECT 50.350 24.510 53.420 25.660 ;
        RECT 50.360 24.460 53.420 24.510 ;
        RECT 51.175 24.200 51.925 24.275 ;
        RECT 50.970 23.970 53.930 24.200 ;
        RECT 42.230 23.810 50.890 23.840 ;
        RECT 42.230 22.810 50.920 23.810 ;
        RECT 51.175 23.465 51.925 23.970 ;
        RECT 63.280 23.810 66.280 26.360 ;
        RECT 42.230 22.800 50.890 22.810 ;
        RECT 42.230 21.560 48.980 22.800 ;
        RECT 51.145 22.650 51.955 23.145 ;
        RECT 53.980 22.810 66.280 23.810 ;
        RECT 54.030 22.800 66.280 22.810 ;
        RECT 50.970 22.420 53.930 22.650 ;
        RECT 51.145 22.395 51.955 22.420 ;
        RECT 50.370 22.120 53.420 22.150 ;
        RECT 50.360 22.080 53.420 22.120 ;
        RECT 42.230 21.110 49.000 21.560 ;
        RECT 43.480 20.230 49.000 21.110 ;
        RECT 50.350 20.930 53.420 22.080 ;
        RECT 50.360 20.880 53.420 20.930 ;
        RECT 51.115 20.620 51.865 20.670 ;
        RECT 54.215 20.620 54.965 20.665 ;
        RECT 50.940 20.390 55.140 20.620 ;
        RECT 38.330 15.880 43.080 20.140 ;
        RECT 38.330 15.360 40.680 15.880 ;
        RECT 38.330 15.300 40.440 15.360 ;
        RECT 38.330 15.210 38.560 15.300 ;
        RECT 37.320 14.820 38.280 15.050 ;
        RECT 31.280 10.560 36.180 14.760 ;
        RECT 37.360 14.200 38.240 14.820 ;
        RECT 39.370 13.100 40.240 13.705 ;
        RECT 36.780 10.830 38.780 12.890 ;
        RECT 39.320 12.870 40.280 13.100 ;
        RECT 39.040 12.630 39.270 12.710 ;
        RECT 38.980 10.560 39.270 12.630 ;
        RECT 31.280 8.560 39.270 10.560 ;
        RECT 31.280 7.160 36.180 8.560 ;
        RECT 36.490 8.550 39.270 8.560 ;
        RECT 39.040 8.470 39.270 8.550 ;
        RECT 40.330 12.630 40.560 12.710 ;
        RECT 41.090 12.630 43.080 15.880 ;
        RECT 40.330 8.550 43.080 12.630 ;
        RECT 43.480 19.230 50.890 20.230 ;
        RECT 51.115 19.860 51.865 20.390 ;
        RECT 54.215 19.855 54.965 20.390 ;
        RECT 55.190 20.220 55.420 20.230 ;
        RECT 63.280 20.220 66.280 22.800 ;
        RECT 43.480 16.660 48.980 19.230 ;
        RECT 51.085 19.070 51.895 19.535 ;
        RECT 54.295 19.070 55.045 19.565 ;
        RECT 55.190 19.290 66.280 20.220 ;
        RECT 55.190 19.230 55.420 19.290 ;
        RECT 50.940 18.840 55.140 19.070 ;
        RECT 51.085 18.785 51.895 18.840 ;
        RECT 54.295 18.755 55.045 18.840 ;
        RECT 50.370 18.540 53.420 18.570 ;
        RECT 50.360 18.500 53.420 18.540 ;
        RECT 50.350 17.350 53.420 18.500 ;
        RECT 50.360 17.300 53.420 17.350 ;
        RECT 50.985 17.040 51.735 17.110 ;
        RECT 55.825 17.040 56.635 17.075 ;
        RECT 50.810 16.810 56.770 17.040 ;
        RECT 43.480 16.650 50.730 16.660 ;
        RECT 43.480 15.660 50.760 16.650 ;
        RECT 50.985 16.300 51.735 16.810 ;
        RECT 55.825 16.325 56.635 16.810 ;
        RECT 56.820 16.640 57.050 16.650 ;
        RECT 63.280 16.640 66.280 19.290 ;
        RECT 43.480 13.060 48.980 15.660 ;
        RECT 50.530 15.650 50.760 15.660 ;
        RECT 50.955 15.490 51.765 15.955 ;
        RECT 55.855 15.490 56.605 15.985 ;
        RECT 56.800 15.710 66.280 16.640 ;
        RECT 56.820 15.650 57.050 15.710 ;
        RECT 50.810 15.260 56.770 15.490 ;
        RECT 50.955 15.205 51.765 15.260 ;
        RECT 55.855 15.175 56.605 15.260 ;
        RECT 50.370 14.960 53.420 14.990 ;
        RECT 50.360 14.920 53.420 14.960 ;
        RECT 50.350 13.770 53.420 14.920 ;
        RECT 50.360 13.720 53.420 13.770 ;
        RECT 50.965 13.460 51.715 13.550 ;
        RECT 58.355 13.460 59.165 13.505 ;
        RECT 50.830 13.230 59.270 13.460 ;
        RECT 50.550 13.060 50.780 13.070 ;
        RECT 43.480 12.070 50.780 13.060 ;
        RECT 50.965 12.740 51.715 13.230 ;
        RECT 58.355 12.755 59.165 13.230 ;
        RECT 59.320 13.060 59.550 13.070 ;
        RECT 63.280 13.060 66.280 15.710 ;
        RECT 43.480 12.060 50.740 12.070 ;
        RECT 43.480 9.500 48.980 12.060 ;
        RECT 50.935 11.910 51.745 12.385 ;
        RECT 58.385 11.910 59.135 12.415 ;
        RECT 59.320 12.130 66.280 13.060 ;
        RECT 59.320 12.070 59.550 12.130 ;
        RECT 50.830 11.680 59.270 11.910 ;
        RECT 50.935 11.635 51.745 11.680 ;
        RECT 58.385 11.605 59.135 11.680 ;
        RECT 50.370 11.380 53.420 11.410 ;
        RECT 50.360 11.340 53.420 11.380 ;
        RECT 50.350 10.190 53.420 11.340 ;
        RECT 63.280 10.760 66.280 12.130 ;
        RECT 72.500 35.600 74.990 45.200 ;
        RECT 72.500 33.200 74.500 35.600 ;
        RECT 74.760 35.550 74.990 35.600 ;
        RECT 76.050 47.490 76.280 47.550 ;
        RECT 78.000 47.490 107.500 47.600 ;
        RECT 76.050 45.950 107.500 47.490 ;
        RECT 111.350 46.900 114.380 48.900 ;
        RECT 114.640 48.890 114.870 48.950 ;
        RECT 114.565 46.600 114.870 48.890 ;
        RECT 76.050 44.600 107.530 45.950 ;
        RECT 76.050 38.540 78.980 44.600 ;
        RECT 82.120 38.940 82.930 39.475 ;
        RECT 82.040 38.710 83.000 38.940 ;
        RECT 81.760 38.540 81.990 38.550 ;
        RECT 76.050 35.610 81.990 38.540 ;
        RECT 76.050 35.550 76.280 35.610 ;
        RECT 75.040 35.160 76.000 35.390 ;
        RECT 75.070 34.515 75.980 35.160 ;
        RECT 77.070 33.440 77.970 34.070 ;
        RECT 77.040 33.210 78.000 33.440 ;
        RECT 72.500 30.500 74.300 33.200 ;
        RECT 76.760 32.990 76.990 33.050 ;
        RECT 74.500 30.870 76.500 32.930 ;
        RECT 76.700 30.500 76.990 32.990 ;
        RECT 72.500 25.100 76.990 30.500 ;
        RECT 72.500 24.100 74.000 25.100 ;
        RECT 75.000 24.640 76.990 25.100 ;
        RECT 75.000 24.100 76.100 24.640 ;
        RECT 76.760 24.570 76.990 24.640 ;
        RECT 78.050 32.990 78.280 33.050 ;
        RECT 79.100 32.990 80.900 35.610 ;
        RECT 81.760 35.550 81.990 35.610 ;
        RECT 83.050 37.100 83.280 38.550 ;
        RECT 83.500 37.250 85.200 39.000 ;
        RECT 85.900 38.520 86.545 38.550 ;
        RECT 85.870 38.490 86.575 38.520 ;
        RECT 85.740 38.260 86.700 38.490 ;
        RECT 85.460 37.100 85.690 38.100 ;
        RECT 85.870 37.875 86.575 38.260 ;
        RECT 86.750 38.050 86.980 38.100 ;
        RECT 87.750 38.050 89.750 44.600 ;
        RECT 85.900 37.845 86.545 37.875 ;
        RECT 83.050 36.050 85.690 37.100 ;
        RECT 83.050 35.870 84.800 36.050 ;
        RECT 85.460 35.980 85.690 36.050 ;
        RECT 83.050 35.600 84.820 35.870 ;
        RECT 85.870 35.820 86.575 36.225 ;
        RECT 86.750 36.050 93.400 38.050 ;
        RECT 86.750 35.980 86.980 36.050 ;
        RECT 83.050 35.550 83.280 35.600 ;
        RECT 82.040 35.160 83.000 35.390 ;
        RECT 82.120 34.575 82.930 35.160 ;
        RECT 78.050 26.500 80.900 32.990 ;
        RECT 83.450 29.850 84.820 35.600 ;
        RECT 85.740 35.590 86.700 35.820 ;
        RECT 85.870 35.580 86.575 35.590 ;
        RECT 88.900 35.230 90.200 36.050 ;
        RECT 88.800 35.000 90.300 35.230 ;
        RECT 88.410 34.850 88.640 34.950 ;
        RECT 90.460 34.850 90.690 34.950 ;
        RECT 86.800 34.730 88.150 34.850 ;
        RECT 85.700 34.700 88.150 34.730 ;
        RECT 85.650 33.600 88.150 34.700 ;
        RECT 88.380 34.820 89.020 34.850 ;
        RECT 90.130 34.820 90.770 34.850 ;
        RECT 88.380 34.180 90.770 34.820 ;
        RECT 88.380 34.150 89.020 34.180 ;
        RECT 90.130 34.150 90.770 34.180 ;
        RECT 88.410 33.990 88.640 34.150 ;
        RECT 90.460 33.990 90.690 34.150 ;
        RECT 88.800 33.710 90.300 33.940 ;
        RECT 85.700 33.570 86.800 33.600 ;
        RECT 88.900 33.400 90.200 33.710 ;
        RECT 90.950 33.600 91.850 35.350 ;
        RECT 92.600 35.230 93.400 36.050 ;
        RECT 92.500 35.000 93.500 35.230 ;
        RECT 92.110 34.805 92.340 34.950 ;
        RECT 93.660 34.805 93.890 34.950 ;
        RECT 92.075 34.090 92.730 34.805 ;
        RECT 93.270 34.090 93.925 34.805 ;
        RECT 92.110 33.990 92.340 34.090 ;
        RECT 93.660 33.990 93.890 34.090 ;
        RECT 92.500 33.710 93.500 33.940 ;
        RECT 92.600 33.400 93.450 33.710 ;
        RECT 88.900 32.625 93.450 33.400 ;
        RECT 88.900 29.850 90.200 32.625 ;
        RECT 92.600 32.280 93.450 32.625 ;
        RECT 92.500 32.050 93.500 32.280 ;
        RECT 92.110 31.425 92.340 32.000 ;
        RECT 92.600 31.900 93.450 32.050 ;
        RECT 93.660 31.705 93.890 32.000 ;
        RECT 91.400 31.330 91.850 31.350 ;
        RECT 90.350 30.170 91.850 31.330 ;
        RECT 92.095 30.675 92.905 31.425 ;
        RECT 93.275 30.895 94.025 31.705 ;
        RECT 92.110 30.540 92.340 30.675 ;
        RECT 93.660 30.540 93.890 30.895 ;
        RECT 83.450 28.000 90.200 29.850 ;
        RECT 90.500 30.150 91.850 30.170 ;
        RECT 92.500 30.400 93.500 30.490 ;
        RECT 92.500 30.250 93.550 30.400 ;
        RECT 104.500 30.260 107.530 44.600 ;
        RECT 95.290 30.250 107.530 30.260 ;
        RECT 90.500 29.250 91.500 30.150 ;
        RECT 92.500 29.350 107.530 30.250 ;
        RECT 95.290 29.260 107.530 29.350 ;
        RECT 90.500 28.800 92.100 29.250 ;
        RECT 92.275 29.125 93.025 29.155 ;
        RECT 90.500 28.150 91.500 28.800 ;
        RECT 92.275 28.590 94.105 29.125 ;
        RECT 92.020 28.360 94.105 28.590 ;
        RECT 92.275 28.345 94.105 28.360 ;
        RECT 104.500 28.200 107.530 29.260 ;
        RECT 91.740 28.000 92.050 28.200 ;
        RECT 83.450 27.200 92.050 28.000 ;
        RECT 78.050 24.700 81.900 26.500 ;
        RECT 78.050 24.640 79.850 24.700 ;
        RECT 78.050 24.570 78.280 24.640 ;
        RECT 77.070 24.410 77.970 24.440 ;
        RECT 77.040 24.180 78.000 24.410 ;
        RECT 72.500 22.200 76.100 24.100 ;
        RECT 77.070 23.600 77.970 24.180 ;
        RECT 78.580 22.440 79.460 22.990 ;
        RECT 78.540 22.210 79.500 22.440 ;
        RECT 72.500 19.600 75.500 22.200 ;
        RECT 78.580 22.170 79.460 22.210 ;
        RECT 78.260 21.970 78.490 22.050 ;
        RECT 76.000 19.870 78.000 21.930 ;
        RECT 78.200 19.600 78.490 21.970 ;
        RECT 72.500 16.600 78.490 19.600 ;
        RECT 72.500 15.600 75.500 16.600 ;
        RECT 76.500 16.140 78.490 16.600 ;
        RECT 78.260 16.050 78.490 16.140 ;
        RECT 79.550 21.970 79.780 22.050 ;
        RECT 80.100 21.970 81.900 24.700 ;
        RECT 79.550 20.980 81.900 21.970 ;
        RECT 83.450 24.680 90.200 27.200 ;
        RECT 92.245 27.040 94.000 27.525 ;
        RECT 94.150 27.200 107.530 28.200 ;
        RECT 92.020 26.810 94.100 27.040 ;
        RECT 92.245 26.790 94.000 26.810 ;
        RECT 91.590 26.540 94.640 26.570 ;
        RECT 91.580 26.500 94.640 26.540 ;
        RECT 91.570 25.350 94.640 26.500 ;
        RECT 91.580 25.300 94.640 25.350 ;
        RECT 92.395 25.040 93.145 25.115 ;
        RECT 92.190 24.810 95.150 25.040 ;
        RECT 83.450 24.650 92.110 24.680 ;
        RECT 83.450 23.650 92.140 24.650 ;
        RECT 92.395 24.305 93.145 24.810 ;
        RECT 104.500 24.650 107.530 27.200 ;
        RECT 83.450 23.640 92.110 23.650 ;
        RECT 83.450 22.400 90.200 23.640 ;
        RECT 92.365 23.490 93.175 23.985 ;
        RECT 95.200 23.650 107.530 24.650 ;
        RECT 95.250 23.640 107.530 23.650 ;
        RECT 92.190 23.260 95.150 23.490 ;
        RECT 92.365 23.235 93.175 23.260 ;
        RECT 91.590 22.960 94.640 22.990 ;
        RECT 91.580 22.920 94.640 22.960 ;
        RECT 83.450 21.950 90.220 22.400 ;
        RECT 84.700 21.070 90.220 21.950 ;
        RECT 91.570 21.770 94.640 22.920 ;
        RECT 91.580 21.720 94.640 21.770 ;
        RECT 92.335 21.460 93.085 21.510 ;
        RECT 95.435 21.460 96.185 21.505 ;
        RECT 92.160 21.230 96.360 21.460 ;
        RECT 79.550 16.720 84.300 20.980 ;
        RECT 79.550 16.200 81.900 16.720 ;
        RECT 79.550 16.140 81.660 16.200 ;
        RECT 79.550 16.050 79.780 16.140 ;
        RECT 78.540 15.660 79.500 15.890 ;
        RECT 72.500 11.400 77.400 15.600 ;
        RECT 78.580 15.040 79.460 15.660 ;
        RECT 80.590 13.940 81.460 14.545 ;
        RECT 78.000 11.670 80.000 13.730 ;
        RECT 80.540 13.710 81.500 13.940 ;
        RECT 80.260 13.470 80.490 13.550 ;
        RECT 80.200 11.400 80.490 13.470 ;
        RECT 50.360 10.140 53.420 10.190 ;
        RECT 50.995 9.880 51.745 9.950 ;
        RECT 61.875 9.880 62.685 9.915 ;
        RECT 50.840 9.650 62.800 9.880 ;
        RECT 43.480 9.490 50.770 9.500 ;
        RECT 40.330 8.470 40.560 8.550 ;
        RECT 43.480 8.500 50.790 9.490 ;
        RECT 50.995 9.140 51.745 9.650 ;
        RECT 61.875 9.165 62.685 9.650 ;
        RECT 62.850 9.480 63.080 9.490 ;
        RECT 64.000 9.480 65.020 10.760 ;
        RECT 39.320 8.080 40.280 8.310 ;
        RECT 39.370 7.495 40.240 8.080 ;
        RECT 43.480 7.240 48.980 8.500 ;
        RECT 50.560 8.490 50.790 8.500 ;
        RECT 50.965 8.330 51.775 8.785 ;
        RECT 61.905 8.330 62.655 8.815 ;
        RECT 62.850 8.500 65.020 9.480 ;
        RECT 72.500 9.400 80.490 11.400 ;
        RECT 62.850 8.490 63.080 8.500 ;
        RECT 50.840 8.100 62.800 8.330 ;
        RECT 50.965 8.035 51.775 8.100 ;
        RECT 61.905 8.005 62.655 8.100 ;
        RECT 72.500 8.000 77.400 9.400 ;
        RECT 77.710 9.390 80.490 9.400 ;
        RECT 80.260 9.310 80.490 9.390 ;
        RECT 81.550 13.470 81.780 13.550 ;
        RECT 82.310 13.470 84.300 16.720 ;
        RECT 81.550 9.390 84.300 13.470 ;
        RECT 84.700 20.070 92.110 21.070 ;
        RECT 92.335 20.700 93.085 21.230 ;
        RECT 95.435 20.695 96.185 21.230 ;
        RECT 96.410 21.060 96.640 21.070 ;
        RECT 104.500 21.060 107.530 23.640 ;
        RECT 84.700 17.500 90.200 20.070 ;
        RECT 92.305 19.910 93.115 20.375 ;
        RECT 95.515 19.910 96.265 20.405 ;
        RECT 96.410 20.130 107.530 21.060 ;
        RECT 96.410 20.070 96.640 20.130 ;
        RECT 92.160 19.680 96.360 19.910 ;
        RECT 92.305 19.625 93.115 19.680 ;
        RECT 95.515 19.595 96.265 19.680 ;
        RECT 91.590 19.380 94.640 19.410 ;
        RECT 91.580 19.340 94.640 19.380 ;
        RECT 91.570 18.190 94.640 19.340 ;
        RECT 91.580 18.140 94.640 18.190 ;
        RECT 92.205 17.880 92.955 17.950 ;
        RECT 97.045 17.880 97.855 17.915 ;
        RECT 92.030 17.650 97.990 17.880 ;
        RECT 84.700 17.490 91.950 17.500 ;
        RECT 84.700 16.500 91.980 17.490 ;
        RECT 92.205 17.140 92.955 17.650 ;
        RECT 97.045 17.165 97.855 17.650 ;
        RECT 98.040 17.480 98.270 17.490 ;
        RECT 104.500 17.480 107.530 20.130 ;
        RECT 84.700 13.900 90.200 16.500 ;
        RECT 91.750 16.490 91.980 16.500 ;
        RECT 92.175 16.330 92.985 16.795 ;
        RECT 97.075 16.330 97.825 16.825 ;
        RECT 98.020 16.550 107.530 17.480 ;
        RECT 98.040 16.490 98.270 16.550 ;
        RECT 92.030 16.100 97.990 16.330 ;
        RECT 92.175 16.045 92.985 16.100 ;
        RECT 97.075 16.015 97.825 16.100 ;
        RECT 91.590 15.800 94.640 15.830 ;
        RECT 91.580 15.760 94.640 15.800 ;
        RECT 91.570 14.610 94.640 15.760 ;
        RECT 91.580 14.560 94.640 14.610 ;
        RECT 92.185 14.300 92.935 14.390 ;
        RECT 99.575 14.300 100.385 14.345 ;
        RECT 92.050 14.070 100.490 14.300 ;
        RECT 91.770 13.900 92.000 13.910 ;
        RECT 84.700 12.910 92.000 13.900 ;
        RECT 92.185 13.580 92.935 14.070 ;
        RECT 99.575 13.595 100.385 14.070 ;
        RECT 100.540 13.900 100.770 13.910 ;
        RECT 104.500 13.900 107.530 16.550 ;
        RECT 84.700 12.900 91.960 12.910 ;
        RECT 84.700 10.340 90.200 12.900 ;
        RECT 92.155 12.750 92.965 13.225 ;
        RECT 99.605 12.750 100.355 13.255 ;
        RECT 100.540 12.970 107.530 13.900 ;
        RECT 100.540 12.910 100.770 12.970 ;
        RECT 92.050 12.520 100.490 12.750 ;
        RECT 92.155 12.475 92.965 12.520 ;
        RECT 99.605 12.445 100.355 12.520 ;
        RECT 91.590 12.220 94.640 12.250 ;
        RECT 91.580 12.180 94.640 12.220 ;
        RECT 91.570 11.030 94.640 12.180 ;
        RECT 104.500 11.600 107.530 12.970 ;
        RECT 91.580 10.980 94.640 11.030 ;
        RECT 105.220 10.850 107.530 11.600 ;
        RECT 112.380 37.000 114.870 46.600 ;
        RECT 112.380 34.600 114.380 37.000 ;
        RECT 114.640 36.950 114.870 37.000 ;
        RECT 115.930 48.890 116.160 48.950 ;
        RECT 117.880 48.890 147.380 49.000 ;
        RECT 115.930 46.000 147.380 48.890 ;
        RECT 115.930 39.940 118.860 46.000 ;
        RECT 122.000 40.340 122.810 40.875 ;
        RECT 121.920 40.110 122.880 40.340 ;
        RECT 121.640 39.940 121.870 39.950 ;
        RECT 115.930 37.010 121.870 39.940 ;
        RECT 115.930 36.950 116.160 37.010 ;
        RECT 114.920 36.560 115.880 36.790 ;
        RECT 114.950 35.915 115.860 36.560 ;
        RECT 116.950 34.840 117.850 35.470 ;
        RECT 116.920 34.610 117.880 34.840 ;
        RECT 112.380 31.900 114.180 34.600 ;
        RECT 116.640 34.390 116.870 34.450 ;
        RECT 114.380 32.270 116.380 34.330 ;
        RECT 116.580 31.900 116.870 34.390 ;
        RECT 112.380 26.500 116.870 31.900 ;
        RECT 112.380 25.500 113.880 26.500 ;
        RECT 114.880 26.040 116.870 26.500 ;
        RECT 114.880 25.500 115.980 26.040 ;
        RECT 116.640 25.970 116.870 26.040 ;
        RECT 117.930 34.390 118.160 34.450 ;
        RECT 118.980 34.390 120.780 37.010 ;
        RECT 121.640 36.950 121.870 37.010 ;
        RECT 122.930 38.500 123.160 39.950 ;
        RECT 123.380 38.650 125.080 40.400 ;
        RECT 125.780 39.920 126.425 39.950 ;
        RECT 125.750 39.890 126.455 39.920 ;
        RECT 125.620 39.660 126.580 39.890 ;
        RECT 125.340 38.500 125.570 39.500 ;
        RECT 125.750 39.275 126.455 39.660 ;
        RECT 126.630 39.450 126.860 39.500 ;
        RECT 127.630 39.450 129.630 46.000 ;
        RECT 144.380 45.850 147.380 46.000 ;
        RECT 125.780 39.245 126.425 39.275 ;
        RECT 122.930 37.450 125.570 38.500 ;
        RECT 122.930 37.270 124.680 37.450 ;
        RECT 125.340 37.380 125.570 37.450 ;
        RECT 122.930 37.000 124.700 37.270 ;
        RECT 125.750 37.220 126.455 37.625 ;
        RECT 126.630 37.450 133.280 39.450 ;
        RECT 126.630 37.380 126.860 37.450 ;
        RECT 122.930 36.950 123.160 37.000 ;
        RECT 121.920 36.560 122.880 36.790 ;
        RECT 122.000 35.975 122.810 36.560 ;
        RECT 117.930 27.900 120.780 34.390 ;
        RECT 123.330 31.250 124.700 37.000 ;
        RECT 125.620 36.990 126.580 37.220 ;
        RECT 125.750 36.980 126.455 36.990 ;
        RECT 128.780 36.630 130.080 37.450 ;
        RECT 128.680 36.400 130.180 36.630 ;
        RECT 128.290 36.250 128.520 36.350 ;
        RECT 130.340 36.250 130.570 36.350 ;
        RECT 126.680 36.130 128.030 36.250 ;
        RECT 125.580 36.100 128.030 36.130 ;
        RECT 125.530 35.000 128.030 36.100 ;
        RECT 128.260 36.220 128.900 36.250 ;
        RECT 130.010 36.220 130.650 36.250 ;
        RECT 128.260 35.580 130.650 36.220 ;
        RECT 128.260 35.550 128.900 35.580 ;
        RECT 130.010 35.550 130.650 35.580 ;
        RECT 128.290 35.390 128.520 35.550 ;
        RECT 130.340 35.390 130.570 35.550 ;
        RECT 128.680 35.110 130.180 35.340 ;
        RECT 125.580 34.970 126.680 35.000 ;
        RECT 128.780 34.800 130.080 35.110 ;
        RECT 130.830 35.000 131.730 36.750 ;
        RECT 132.480 36.630 133.280 37.450 ;
        RECT 132.380 36.400 133.380 36.630 ;
        RECT 131.990 36.205 132.220 36.350 ;
        RECT 133.540 36.205 133.770 36.350 ;
        RECT 131.955 35.490 132.610 36.205 ;
        RECT 133.150 35.490 133.805 36.205 ;
        RECT 131.990 35.390 132.220 35.490 ;
        RECT 133.540 35.390 133.770 35.490 ;
        RECT 132.380 35.110 133.380 35.340 ;
        RECT 132.480 34.800 133.330 35.110 ;
        RECT 128.780 34.025 133.330 34.800 ;
        RECT 128.780 31.250 130.080 34.025 ;
        RECT 132.480 33.680 133.330 34.025 ;
        RECT 132.380 33.450 133.380 33.680 ;
        RECT 131.990 32.825 132.220 33.400 ;
        RECT 132.480 33.300 133.330 33.450 ;
        RECT 133.540 33.105 133.770 33.400 ;
        RECT 131.280 32.730 131.730 32.750 ;
        RECT 130.230 31.570 131.730 32.730 ;
        RECT 131.975 32.075 132.785 32.825 ;
        RECT 133.155 32.295 133.905 33.105 ;
        RECT 131.990 31.940 132.220 32.075 ;
        RECT 133.540 31.940 133.770 32.295 ;
        RECT 123.330 29.400 130.080 31.250 ;
        RECT 130.380 31.550 131.730 31.570 ;
        RECT 132.380 31.800 133.380 31.890 ;
        RECT 132.380 31.650 133.430 31.800 ;
        RECT 144.380 31.660 147.400 45.850 ;
        RECT 135.170 31.650 147.400 31.660 ;
        RECT 130.380 30.650 131.380 31.550 ;
        RECT 132.380 30.750 147.400 31.650 ;
        RECT 135.170 30.660 147.400 30.750 ;
        RECT 130.380 30.200 131.980 30.650 ;
        RECT 132.155 30.525 132.905 30.555 ;
        RECT 130.380 29.550 131.380 30.200 ;
        RECT 132.155 29.990 133.985 30.525 ;
        RECT 131.900 29.760 133.985 29.990 ;
        RECT 132.155 29.745 133.985 29.760 ;
        RECT 144.380 29.600 147.400 30.660 ;
        RECT 131.620 29.400 131.930 29.600 ;
        RECT 123.330 28.600 131.930 29.400 ;
        RECT 117.930 26.100 121.780 27.900 ;
        RECT 117.930 26.040 119.730 26.100 ;
        RECT 117.930 25.970 118.160 26.040 ;
        RECT 116.950 25.810 117.850 25.840 ;
        RECT 116.920 25.580 117.880 25.810 ;
        RECT 112.380 23.600 115.980 25.500 ;
        RECT 116.950 25.000 117.850 25.580 ;
        RECT 118.460 23.840 119.340 24.390 ;
        RECT 118.420 23.610 119.380 23.840 ;
        RECT 112.380 21.000 115.380 23.600 ;
        RECT 118.460 23.570 119.340 23.610 ;
        RECT 118.140 23.370 118.370 23.450 ;
        RECT 115.880 21.270 117.880 23.330 ;
        RECT 118.080 21.000 118.370 23.370 ;
        RECT 112.380 18.000 118.370 21.000 ;
        RECT 112.380 17.000 115.380 18.000 ;
        RECT 116.380 17.540 118.370 18.000 ;
        RECT 118.140 17.450 118.370 17.540 ;
        RECT 119.430 23.370 119.660 23.450 ;
        RECT 119.980 23.370 121.780 26.100 ;
        RECT 119.430 22.380 121.780 23.370 ;
        RECT 123.330 26.080 130.080 28.600 ;
        RECT 132.125 28.440 133.880 28.925 ;
        RECT 134.030 28.600 147.400 29.600 ;
        RECT 131.900 28.210 133.980 28.440 ;
        RECT 132.125 28.190 133.880 28.210 ;
        RECT 131.470 27.940 134.520 27.970 ;
        RECT 131.460 27.900 134.520 27.940 ;
        RECT 131.450 26.750 134.520 27.900 ;
        RECT 131.460 26.700 134.520 26.750 ;
        RECT 132.275 26.440 133.025 26.515 ;
        RECT 132.070 26.210 135.030 26.440 ;
        RECT 123.330 26.050 131.990 26.080 ;
        RECT 123.330 25.050 132.020 26.050 ;
        RECT 132.275 25.705 133.025 26.210 ;
        RECT 144.380 26.050 147.400 28.600 ;
        RECT 123.330 25.040 131.990 25.050 ;
        RECT 123.330 23.800 130.080 25.040 ;
        RECT 132.245 24.890 133.055 25.385 ;
        RECT 135.080 25.050 147.400 26.050 ;
        RECT 135.130 25.040 147.400 25.050 ;
        RECT 132.070 24.660 135.030 24.890 ;
        RECT 132.245 24.635 133.055 24.660 ;
        RECT 131.470 24.360 134.520 24.390 ;
        RECT 131.460 24.320 134.520 24.360 ;
        RECT 123.330 23.350 130.100 23.800 ;
        RECT 124.580 22.470 130.100 23.350 ;
        RECT 131.450 23.170 134.520 24.320 ;
        RECT 131.460 23.120 134.520 23.170 ;
        RECT 132.215 22.860 132.965 22.910 ;
        RECT 135.315 22.860 136.065 22.905 ;
        RECT 132.040 22.630 136.240 22.860 ;
        RECT 119.430 18.120 124.180 22.380 ;
        RECT 119.430 17.600 121.780 18.120 ;
        RECT 119.430 17.540 121.540 17.600 ;
        RECT 119.430 17.450 119.660 17.540 ;
        RECT 118.420 17.060 119.380 17.290 ;
        RECT 112.380 12.800 117.280 17.000 ;
        RECT 118.460 16.440 119.340 17.060 ;
        RECT 120.470 15.340 121.340 15.945 ;
        RECT 117.880 13.070 119.880 15.130 ;
        RECT 120.420 15.110 121.380 15.340 ;
        RECT 120.140 14.870 120.370 14.950 ;
        RECT 120.080 12.800 120.370 14.870 ;
        RECT 92.215 10.720 92.965 10.790 ;
        RECT 103.095 10.720 103.905 10.755 ;
        RECT 92.060 10.490 104.020 10.720 ;
        RECT 84.700 10.330 91.990 10.340 ;
        RECT 81.550 9.310 81.780 9.390 ;
        RECT 84.700 9.340 92.010 10.330 ;
        RECT 92.215 9.980 92.965 10.490 ;
        RECT 103.095 10.005 103.905 10.490 ;
        RECT 104.070 10.320 104.300 10.330 ;
        RECT 105.220 10.320 106.240 10.850 ;
        RECT 80.540 8.920 81.500 9.150 ;
        RECT 80.590 8.335 81.460 8.920 ;
        RECT 84.700 8.080 90.200 9.340 ;
        RECT 91.780 9.330 92.010 9.340 ;
        RECT 92.185 9.170 92.995 9.625 ;
        RECT 103.125 9.170 103.875 9.655 ;
        RECT 104.070 9.340 106.240 10.320 ;
        RECT 112.380 10.800 120.370 12.800 ;
        RECT 112.380 9.400 117.280 10.800 ;
        RECT 117.590 10.790 120.370 10.800 ;
        RECT 120.140 10.710 120.370 10.790 ;
        RECT 121.430 14.870 121.660 14.950 ;
        RECT 122.190 14.870 124.180 18.120 ;
        RECT 121.430 10.790 124.180 14.870 ;
        RECT 124.580 21.470 131.990 22.470 ;
        RECT 132.215 22.100 132.965 22.630 ;
        RECT 135.315 22.095 136.065 22.630 ;
        RECT 136.290 22.460 136.520 22.470 ;
        RECT 144.380 22.460 147.400 25.040 ;
        RECT 124.580 18.900 130.080 21.470 ;
        RECT 132.185 21.310 132.995 21.775 ;
        RECT 135.395 21.310 136.145 21.805 ;
        RECT 136.290 21.530 147.400 22.460 ;
        RECT 136.290 21.470 136.520 21.530 ;
        RECT 132.040 21.080 136.240 21.310 ;
        RECT 132.185 21.025 132.995 21.080 ;
        RECT 135.395 20.995 136.145 21.080 ;
        RECT 131.470 20.780 134.520 20.810 ;
        RECT 131.460 20.740 134.520 20.780 ;
        RECT 131.450 19.590 134.520 20.740 ;
        RECT 131.460 19.540 134.520 19.590 ;
        RECT 132.085 19.280 132.835 19.350 ;
        RECT 136.925 19.280 137.735 19.315 ;
        RECT 131.910 19.050 137.870 19.280 ;
        RECT 124.580 18.890 131.830 18.900 ;
        RECT 124.580 17.900 131.860 18.890 ;
        RECT 132.085 18.540 132.835 19.050 ;
        RECT 136.925 18.565 137.735 19.050 ;
        RECT 137.920 18.880 138.150 18.890 ;
        RECT 144.380 18.880 147.400 21.530 ;
        RECT 124.580 15.300 130.080 17.900 ;
        RECT 131.630 17.890 131.860 17.900 ;
        RECT 132.055 17.730 132.865 18.195 ;
        RECT 136.955 17.730 137.705 18.225 ;
        RECT 137.900 17.950 147.400 18.880 ;
        RECT 137.920 17.890 138.150 17.950 ;
        RECT 131.910 17.500 137.870 17.730 ;
        RECT 132.055 17.445 132.865 17.500 ;
        RECT 136.955 17.415 137.705 17.500 ;
        RECT 131.470 17.200 134.520 17.230 ;
        RECT 131.460 17.160 134.520 17.200 ;
        RECT 131.450 16.010 134.520 17.160 ;
        RECT 131.460 15.960 134.520 16.010 ;
        RECT 132.065 15.700 132.815 15.790 ;
        RECT 139.455 15.700 140.265 15.745 ;
        RECT 131.930 15.470 140.370 15.700 ;
        RECT 131.650 15.300 131.880 15.310 ;
        RECT 124.580 14.310 131.880 15.300 ;
        RECT 132.065 14.980 132.815 15.470 ;
        RECT 139.455 14.995 140.265 15.470 ;
        RECT 140.420 15.300 140.650 15.310 ;
        RECT 144.380 15.300 147.400 17.950 ;
        RECT 124.580 14.300 131.840 14.310 ;
        RECT 124.580 11.740 130.080 14.300 ;
        RECT 132.035 14.150 132.845 14.625 ;
        RECT 139.485 14.150 140.235 14.655 ;
        RECT 140.420 14.370 147.400 15.300 ;
        RECT 140.420 14.310 140.650 14.370 ;
        RECT 131.930 13.920 140.370 14.150 ;
        RECT 132.035 13.875 132.845 13.920 ;
        RECT 139.485 13.845 140.235 13.920 ;
        RECT 131.470 13.620 134.520 13.650 ;
        RECT 131.460 13.580 134.520 13.620 ;
        RECT 131.450 12.430 134.520 13.580 ;
        RECT 144.380 13.000 147.400 14.370 ;
        RECT 131.460 12.380 134.520 12.430 ;
        RECT 132.095 12.120 132.845 12.190 ;
        RECT 142.975 12.120 143.785 12.155 ;
        RECT 131.940 11.890 143.900 12.120 ;
        RECT 124.580 11.730 131.870 11.740 ;
        RECT 121.430 10.710 121.660 10.790 ;
        RECT 124.580 10.740 131.890 11.730 ;
        RECT 132.095 11.380 132.845 11.890 ;
        RECT 142.975 11.405 143.785 11.890 ;
        RECT 143.950 11.720 144.180 11.730 ;
        RECT 145.100 11.720 147.400 13.000 ;
        RECT 120.420 10.320 121.380 10.550 ;
        RECT 120.470 9.735 121.340 10.320 ;
        RECT 124.580 9.480 130.080 10.740 ;
        RECT 131.660 10.730 131.890 10.740 ;
        RECT 132.065 10.570 132.875 11.025 ;
        RECT 143.005 10.570 143.755 11.055 ;
        RECT 143.950 10.900 147.400 11.720 ;
        RECT 143.950 10.740 146.120 10.900 ;
        RECT 143.950 10.730 144.180 10.740 ;
        RECT 131.940 10.340 143.900 10.570 ;
        RECT 132.065 10.275 132.875 10.340 ;
        RECT 143.005 10.245 143.755 10.340 ;
        RECT 141.380 9.850 144.530 10.100 ;
        RECT 124.580 9.400 130.070 9.480 ;
        RECT 104.070 9.330 104.300 9.340 ;
        RECT 92.060 8.940 104.020 9.170 ;
        RECT 92.185 8.875 92.995 8.940 ;
        RECT 103.125 8.845 103.875 8.940 ;
        RECT 101.500 8.450 104.650 8.700 ;
        RECT 84.700 8.000 90.190 8.080 ;
        RECT 60.280 7.610 63.430 7.860 ;
        RECT 43.480 7.160 48.970 7.240 ;
        RECT 31.280 2.260 48.970 7.160 ;
        RECT 60.280 6.210 63.580 7.610 ;
        RECT 72.500 3.100 90.190 8.000 ;
        RECT 101.500 7.050 104.800 8.450 ;
        RECT 112.380 4.500 130.070 9.400 ;
        RECT 141.380 8.450 144.680 9.850 ;
        RECT 124.155 4.475 126.245 4.500 ;
        RECT 41.640 2.255 43.860 2.260 ;
      LAYER met2 ;
        RECT 78.460 220.900 78.740 220.935 ;
        RECT 26.950 217.940 27.250 217.950 ;
        RECT 26.915 217.660 27.285 217.940 ;
        RECT 26.950 215.690 27.250 217.660 ;
        RECT 34.300 217.240 34.600 217.250 ;
        RECT 34.265 216.960 34.635 217.240 ;
        RECT 26.930 215.100 27.250 215.690 ;
        RECT 34.300 215.290 34.600 216.960 ;
        RECT 41.650 216.540 41.950 216.550 ;
        RECT 41.615 216.260 41.985 216.540 ;
        RECT 26.930 214.200 27.210 215.100 ;
        RECT 34.290 214.650 34.600 215.290 ;
        RECT 41.650 214.700 41.950 216.260 ;
        RECT 63.700 214.940 64.000 214.950 ;
        RECT 49.010 214.900 49.290 214.935 ;
        RECT 34.290 214.200 34.570 214.650 ;
        RECT 41.650 214.200 41.930 214.700 ;
        RECT 26.920 213.760 27.210 214.200 ;
        RECT 26.920 212.200 27.200 213.760 ;
        RECT 34.280 213.360 34.570 214.200 ;
        RECT 41.640 213.510 41.930 214.200 ;
        RECT 49.000 213.700 49.300 214.900 ;
        RECT 56.350 214.890 56.650 214.900 ;
        RECT 56.315 214.610 56.685 214.890 ;
        RECT 63.665 214.660 64.035 214.940 ;
        RECT 71.050 214.890 71.350 214.900 ;
        RECT 56.350 213.700 56.650 214.610 ;
        RECT 63.700 214.090 64.000 214.660 ;
        RECT 71.015 214.610 71.385 214.890 ;
        RECT 71.050 214.200 71.350 214.610 ;
        RECT 78.450 214.600 78.750 220.900 ;
        RECT 85.800 220.190 86.100 220.200 ;
        RECT 85.765 219.910 86.135 220.190 ;
        RECT 78.450 214.200 78.730 214.600 ;
        RECT 63.700 213.800 64.010 214.090 ;
        RECT 63.720 213.700 64.010 213.800 ;
        RECT 71.050 214.040 71.360 214.200 ;
        RECT 71.050 213.700 71.370 214.040 ;
        RECT 78.440 213.700 78.730 214.200 ;
        RECT 85.800 213.700 86.100 219.910 ;
        RECT 93.160 219.550 93.440 219.585 ;
        RECT 93.150 213.700 93.450 219.550 ;
        RECT 100.560 218.850 100.840 218.885 ;
        RECT 100.550 214.200 100.850 218.850 ;
        RECT 107.910 218.150 108.190 218.185 ;
        RECT 107.900 214.200 108.200 218.150 ;
        RECT 115.260 217.400 115.540 217.435 ;
        RECT 115.250 214.200 115.550 217.400 ;
        RECT 122.610 216.750 122.890 216.785 ;
        RECT 100.520 213.700 100.850 214.200 ;
        RECT 107.880 213.700 108.200 214.200 ;
        RECT 115.240 213.700 115.550 214.200 ;
        RECT 122.600 213.700 122.900 216.750 ;
        RECT 129.950 216.090 130.250 216.100 ;
        RECT 129.915 215.810 130.285 216.090 ;
        RECT 129.950 213.700 130.250 215.810 ;
        RECT 137.300 215.460 137.580 215.495 ;
        RECT 137.290 214.200 137.590 215.460 ;
        RECT 144.690 214.790 144.970 214.825 ;
        RECT 137.290 213.700 137.600 214.200 ;
        RECT 34.280 212.200 34.560 213.360 ;
        RECT 41.640 212.200 41.920 213.510 ;
        RECT 49.000 212.200 49.280 213.700 ;
        RECT 56.360 212.200 56.640 213.700 ;
        RECT 63.720 212.200 64.000 213.700 ;
        RECT 71.080 212.200 71.360 213.700 ;
        RECT 78.440 212.200 78.720 213.700 ;
        RECT 85.800 212.200 86.080 213.700 ;
        RECT 93.160 212.200 93.440 213.700 ;
        RECT 100.520 212.200 100.800 213.700 ;
        RECT 107.880 212.200 108.160 213.700 ;
        RECT 115.240 212.200 115.520 213.700 ;
        RECT 122.600 213.610 122.890 213.700 ;
        RECT 122.600 212.200 122.880 213.610 ;
        RECT 129.960 212.200 130.240 213.700 ;
        RECT 137.320 212.200 137.600 213.700 ;
        RECT 144.680 213.700 144.980 214.790 ;
        RECT 152.040 214.140 152.320 214.200 ;
        RECT 152.570 214.140 152.850 214.175 ;
        RECT 152.040 213.840 152.860 214.140 ;
        RECT 152.040 213.700 152.340 213.840 ;
        RECT 152.570 213.805 152.850 213.840 ;
        RECT 144.680 212.200 144.960 213.700 ;
        RECT 152.040 212.200 152.320 213.700 ;
        RECT 26.990 208.890 27.130 212.200 ;
        RECT 26.930 208.570 27.190 208.890 ;
        RECT 30.150 207.890 30.410 208.210 ;
        RECT 30.210 206.365 30.350 207.890 ;
        RECT 31.530 207.550 31.790 207.870 ;
        RECT 30.140 205.995 30.420 206.365 ;
        RECT 31.590 205.150 31.730 207.550 ;
        RECT 34.350 205.830 34.490 212.200 ;
        RECT 37.510 207.890 37.770 208.210 ;
        RECT 34.290 205.510 34.550 205.830 ;
        RECT 31.530 204.830 31.790 205.150 ;
        RECT 29.230 204.490 29.490 204.810 ;
        RECT 28.770 204.150 29.030 204.470 ;
        RECT 28.830 202.170 28.970 204.150 ;
        RECT 29.290 202.965 29.430 204.490 ;
        RECT 37.570 203.450 37.710 207.890 ;
        RECT 37.970 206.870 38.230 207.190 ;
        RECT 38.030 204.810 38.170 206.870 ;
        RECT 38.710 206.335 40.250 206.705 ;
        RECT 37.970 204.490 38.230 204.810 ;
        RECT 37.510 203.130 37.770 203.450 ;
        RECT 29.220 202.595 29.500 202.965 ;
        RECT 40.730 202.790 40.990 203.110 ;
        RECT 30.150 202.450 30.410 202.770 ;
        RECT 37.970 202.450 38.230 202.770 ;
        RECT 29.230 202.170 29.490 202.430 ;
        RECT 28.830 202.110 29.490 202.170 ;
        RECT 28.830 202.030 29.430 202.110 ;
        RECT 29.290 196.990 29.430 202.030 ;
        RECT 29.230 196.670 29.490 196.990 ;
        RECT 26.010 186.130 26.270 186.450 ;
        RECT 26.070 184.410 26.210 186.130 ;
        RECT 26.010 184.090 26.270 184.410 ;
        RECT 26.010 180.690 26.270 181.010 ;
        RECT 25.550 179.670 25.810 179.990 ;
        RECT 25.610 177.610 25.750 179.670 ;
        RECT 26.070 177.610 26.210 180.690 ;
        RECT 25.550 177.290 25.810 177.610 ;
        RECT 26.010 177.290 26.270 177.610 ;
        RECT 29.230 177.290 29.490 177.610 ;
        RECT 29.290 175.570 29.430 177.290 ;
        RECT 29.230 175.250 29.490 175.570 ;
        RECT 25.550 174.230 25.810 174.550 ;
        RECT 25.610 172.510 25.750 174.230 ;
        RECT 24.170 172.190 24.430 172.510 ;
        RECT 25.550 172.190 25.810 172.510 ;
        RECT 24.230 167.410 24.370 172.190 ;
        RECT 24.170 167.090 24.430 167.410 ;
        RECT 24.230 159.250 24.370 167.090 ;
        RECT 26.010 166.410 26.270 166.730 ;
        RECT 26.070 165.370 26.210 166.410 ;
        RECT 26.010 165.050 26.270 165.370 ;
        RECT 30.210 164.670 30.350 202.450 ;
        RECT 38.030 200.730 38.170 202.450 ;
        RECT 38.710 200.895 40.250 201.265 ;
        RECT 40.790 200.730 40.930 202.790 ;
        RECT 41.710 201.750 41.850 212.200 ;
        RECT 49.070 208.890 49.210 212.200 ;
        RECT 56.430 210.330 56.570 212.200 ;
        RECT 56.430 210.190 57.490 210.330 ;
        RECT 55.500 209.055 57.040 209.425 ;
        RECT 57.350 208.890 57.490 210.190 ;
        RECT 63.790 208.890 63.930 212.200 ;
        RECT 49.010 208.570 49.270 208.890 ;
        RECT 57.290 208.570 57.550 208.890 ;
        RECT 63.730 208.570 63.990 208.890 ;
        RECT 71.150 208.290 71.290 212.200 ;
        RECT 71.150 208.210 71.750 208.290 ;
        RECT 78.510 208.210 78.650 212.200 ;
        RECT 85.870 208.210 86.010 212.200 ;
        RECT 87.190 209.930 87.450 210.250 ;
        RECT 68.330 207.890 68.590 208.210 ;
        RECT 69.250 207.890 69.510 208.210 ;
        RECT 71.150 208.150 71.810 208.210 ;
        RECT 71.550 207.890 71.810 208.150 ;
        RECT 78.450 207.890 78.710 208.210 ;
        RECT 83.510 207.890 83.770 208.210 ;
        RECT 85.810 207.890 86.070 208.210 ;
        RECT 49.470 206.870 49.730 207.190 ;
        RECT 56.830 206.870 57.090 207.190 ;
        RECT 62.350 206.870 62.610 207.190 ;
        RECT 63.730 206.870 63.990 207.190 ;
        RECT 49.530 206.170 49.670 206.870 ;
        RECT 49.470 205.850 49.730 206.170 ;
        RECT 56.890 205.830 57.030 206.870 ;
        RECT 56.830 205.510 57.090 205.830 ;
        RECT 42.570 204.830 42.830 205.150 ;
        RECT 49.470 204.830 49.730 205.150 ;
        RECT 54.070 204.830 54.330 205.150 ;
        RECT 41.190 201.430 41.450 201.750 ;
        RECT 41.650 201.430 41.910 201.750 ;
        RECT 41.250 200.810 41.390 201.430 ;
        RECT 37.970 200.410 38.230 200.730 ;
        RECT 40.730 200.410 40.990 200.730 ;
        RECT 41.250 200.670 42.310 200.810 ;
        RECT 35.210 199.390 35.470 199.710 ;
        RECT 30.610 197.010 30.870 197.330 ;
        RECT 30.670 195.290 30.810 197.010 ;
        RECT 31.070 195.990 31.330 196.310 ;
        RECT 33.830 195.990 34.090 196.310 ;
        RECT 30.610 194.970 30.870 195.290 ;
        RECT 31.130 191.550 31.270 195.990 ;
        RECT 33.890 193.930 34.030 195.990 ;
        RECT 35.270 194.950 35.410 199.390 ;
        RECT 39.810 199.280 40.070 199.370 ;
        RECT 40.720 199.280 41.000 199.565 ;
        RECT 39.810 199.140 41.390 199.280 ;
        RECT 39.810 199.050 40.070 199.140 ;
        RECT 36.130 197.690 36.390 198.010 ;
        RECT 36.190 194.950 36.330 197.690 ;
        RECT 41.250 197.670 41.390 199.140 ;
        RECT 42.170 197.670 42.310 200.670 ;
        RECT 41.190 197.350 41.450 197.670 ;
        RECT 42.110 197.350 42.370 197.670 ;
        RECT 37.970 197.010 38.230 197.330 ;
        RECT 37.050 195.990 37.310 196.310 ;
        RECT 37.110 195.290 37.250 195.990 ;
        RECT 37.050 194.970 37.310 195.290 ;
        RECT 35.210 194.630 35.470 194.950 ;
        RECT 36.130 194.630 36.390 194.950 ;
        RECT 34.290 193.950 34.550 194.270 ;
        RECT 33.830 193.610 34.090 193.930 ;
        RECT 32.450 193.270 32.710 193.590 ;
        RECT 32.510 192.230 32.650 193.270 ;
        RECT 34.350 192.570 34.490 193.950 ;
        RECT 38.030 193.930 38.170 197.010 ;
        RECT 41.190 196.670 41.450 196.990 ;
        RECT 38.710 195.455 40.250 195.825 ;
        RECT 36.130 193.610 36.390 193.930 ;
        RECT 37.970 193.610 38.230 193.930 ;
        RECT 34.290 192.250 34.550 192.570 ;
        RECT 32.450 191.910 32.710 192.230 ;
        RECT 31.070 191.230 31.330 191.550 ;
        RECT 31.130 187.130 31.270 191.230 ;
        RECT 32.450 188.510 32.710 188.830 ;
        RECT 31.530 188.170 31.790 188.490 ;
        RECT 31.070 186.810 31.330 187.130 ;
        RECT 31.590 185.770 31.730 188.170 ;
        RECT 31.530 185.450 31.790 185.770 ;
        RECT 31.590 183.390 31.730 185.450 ;
        RECT 31.990 185.110 32.250 185.430 ;
        RECT 32.050 184.410 32.190 185.110 ;
        RECT 31.990 184.090 32.250 184.410 ;
        RECT 31.530 183.070 31.790 183.390 ;
        RECT 31.990 183.300 32.250 183.390 ;
        RECT 32.510 183.300 32.650 188.510 ;
        RECT 32.910 187.830 33.170 188.150 ;
        RECT 33.370 187.830 33.630 188.150 ;
        RECT 32.970 185.430 33.110 187.830 ;
        RECT 33.430 186.450 33.570 187.830 ;
        RECT 33.370 186.130 33.630 186.450 ;
        RECT 32.910 185.110 33.170 185.430 ;
        RECT 31.990 183.160 32.650 183.300 ;
        RECT 31.990 183.070 32.250 183.160 ;
        RECT 32.510 182.710 32.650 183.160 ;
        RECT 32.450 182.390 32.710 182.710 ;
        RECT 31.070 180.690 31.330 181.010 ;
        RECT 31.990 180.690 32.250 181.010 ;
        RECT 31.130 175.910 31.270 180.690 ;
        RECT 32.050 178.970 32.190 180.690 ;
        RECT 32.910 179.670 33.170 179.990 ;
        RECT 32.970 178.970 33.110 179.670 ;
        RECT 31.990 178.650 32.250 178.970 ;
        RECT 32.910 178.650 33.170 178.970 ;
        RECT 33.430 177.270 33.570 186.130 ;
        RECT 34.750 185.450 35.010 185.770 ;
        RECT 34.810 184.070 34.950 185.450 ;
        RECT 35.670 185.110 35.930 185.430 ;
        RECT 34.750 183.750 35.010 184.070 ;
        RECT 35.730 183.390 35.870 185.110 ;
        RECT 35.670 183.070 35.930 183.390 ;
        RECT 34.290 182.390 34.550 182.710 ;
        RECT 35.210 182.390 35.470 182.710 ;
        RECT 34.350 178.630 34.490 182.390 ;
        RECT 35.270 181.690 35.410 182.390 ;
        RECT 35.210 181.370 35.470 181.690 ;
        RECT 35.210 178.650 35.470 178.970 ;
        RECT 34.290 178.310 34.550 178.630 ;
        RECT 33.370 176.950 33.630 177.270 ;
        RECT 31.070 175.590 31.330 175.910 ;
        RECT 33.430 175.820 33.570 176.950 ;
        RECT 35.270 176.250 35.410 178.650 ;
        RECT 35.730 177.610 35.870 183.070 ;
        RECT 35.670 177.290 35.930 177.610 ;
        RECT 35.730 176.250 35.870 177.290 ;
        RECT 35.210 175.930 35.470 176.250 ;
        RECT 35.670 175.930 35.930 176.250 ;
        RECT 33.830 175.820 34.090 175.910 ;
        RECT 33.430 175.680 34.090 175.820 ;
        RECT 33.430 172.930 33.570 175.680 ;
        RECT 33.830 175.590 34.090 175.680 ;
        RECT 35.270 173.530 35.410 175.930 ;
        RECT 35.210 173.210 35.470 173.530 ;
        RECT 33.430 172.790 34.030 172.930 ;
        RECT 33.370 171.850 33.630 172.170 ;
        RECT 33.430 170.810 33.570 171.850 ;
        RECT 33.890 170.810 34.030 172.790 ;
        RECT 35.210 171.510 35.470 171.830 ;
        RECT 33.370 170.490 33.630 170.810 ;
        RECT 33.830 170.490 34.090 170.810 ;
        RECT 31.070 169.470 31.330 169.790 ;
        RECT 31.130 168.090 31.270 169.470 ;
        RECT 31.070 167.770 31.330 168.090 ;
        RECT 32.450 167.770 32.710 168.090 ;
        RECT 31.530 166.070 31.790 166.390 ;
        RECT 31.590 165.370 31.730 166.070 ;
        RECT 32.510 165.370 32.650 167.770 ;
        RECT 33.430 167.750 33.570 170.490 ;
        RECT 33.370 167.430 33.630 167.750 ;
        RECT 33.890 166.390 34.030 170.490 ;
        RECT 34.290 169.810 34.550 170.130 ;
        RECT 33.830 166.070 34.090 166.390 ;
        RECT 31.530 165.050 31.790 165.370 ;
        RECT 32.450 165.050 32.710 165.370 ;
        RECT 34.350 165.030 34.490 169.810 ;
        RECT 35.270 169.110 35.410 171.510 ;
        RECT 35.210 168.790 35.470 169.110 ;
        RECT 34.750 167.770 35.010 168.090 ;
        RECT 34.810 165.370 34.950 167.770 ;
        RECT 35.670 166.070 35.930 166.390 ;
        RECT 35.730 165.370 35.870 166.070 ;
        RECT 34.750 165.050 35.010 165.370 ;
        RECT 35.670 165.050 35.930 165.370 ;
        RECT 34.290 164.710 34.550 165.030 ;
        RECT 29.290 164.530 30.350 164.670 ;
        RECT 27.850 161.310 28.110 161.630 ;
        RECT 25.090 160.630 25.350 160.950 ;
        RECT 24.170 158.930 24.430 159.250 ;
        RECT 24.230 156.190 24.370 158.930 ;
        RECT 24.170 155.870 24.430 156.190 ;
        RECT 24.230 150.750 24.370 155.870 ;
        RECT 24.170 150.430 24.430 150.750 ;
        RECT 24.230 148.370 24.370 150.430 ;
        RECT 25.150 150.070 25.290 160.630 ;
        RECT 27.910 158.910 28.050 161.310 ;
        RECT 27.850 158.590 28.110 158.910 ;
        RECT 25.550 157.910 25.810 158.230 ;
        RECT 25.610 156.190 25.750 157.910 ;
        RECT 25.550 155.870 25.810 156.190 ;
        RECT 26.930 153.490 27.190 153.810 ;
        RECT 25.550 152.470 25.810 152.790 ;
        RECT 25.610 150.750 25.750 152.470 ;
        RECT 25.550 150.430 25.810 150.750 ;
        RECT 25.090 149.750 25.350 150.070 ;
        RECT 25.150 148.370 25.290 149.750 ;
        RECT 26.990 149.050 27.130 153.490 ;
        RECT 26.930 148.730 27.190 149.050 ;
        RECT 24.170 148.050 24.430 148.370 ;
        RECT 25.090 148.050 25.350 148.370 ;
        RECT 24.230 142.930 24.370 148.050 ;
        RECT 26.930 147.370 27.190 147.690 ;
        RECT 26.990 145.310 27.130 147.370 ;
        RECT 26.930 144.990 27.190 145.310 ;
        RECT 28.310 144.310 28.570 144.630 ;
        RECT 28.770 144.310 29.030 144.630 ;
        RECT 24.170 142.610 24.430 142.930 ;
        RECT 26.930 142.610 27.190 142.930 ;
        RECT 26.990 140.890 27.130 142.610 ;
        RECT 26.930 140.570 27.190 140.890 ;
        RECT 28.370 139.870 28.510 144.310 ;
        RECT 28.830 143.610 28.970 144.310 ;
        RECT 28.770 143.290 29.030 143.610 ;
        RECT 28.830 140.890 28.970 143.290 ;
        RECT 28.770 140.570 29.030 140.890 ;
        RECT 28.310 139.550 28.570 139.870 ;
        RECT 25.090 137.170 25.350 137.490 ;
        RECT 24.630 131.730 24.890 132.050 ;
        RECT 24.690 130.010 24.830 131.730 ;
        RECT 24.630 129.690 24.890 130.010 ;
        RECT 25.150 129.330 25.290 137.170 ;
        RECT 28.310 133.770 28.570 134.090 ;
        RECT 28.370 132.730 28.510 133.770 ;
        RECT 28.770 133.430 29.030 133.750 ;
        RECT 28.830 132.730 28.970 133.430 ;
        RECT 28.310 132.410 28.570 132.730 ;
        RECT 28.770 132.410 29.030 132.730 ;
        RECT 25.550 130.710 25.810 131.030 ;
        RECT 27.850 130.710 28.110 131.030 ;
        RECT 25.090 129.010 25.350 129.330 ;
        RECT 25.150 127.290 25.290 129.010 ;
        RECT 25.090 126.970 25.350 127.290 ;
        RECT 25.610 126.950 25.750 130.710 ;
        RECT 25.550 126.630 25.810 126.950 ;
        RECT 26.470 122.890 26.730 123.210 ;
        RECT 25.550 122.550 25.810 122.870 ;
        RECT 26.530 122.610 26.670 122.890 ;
        RECT 25.610 118.110 25.750 122.550 ;
        RECT 26.070 122.470 26.670 122.610 ;
        RECT 26.070 120.150 26.210 122.470 ;
        RECT 26.010 119.830 26.270 120.150 ;
        RECT 25.550 117.790 25.810 118.110 ;
        RECT 25.610 116.370 25.750 117.790 ;
        RECT 25.150 116.230 25.750 116.370 ;
        RECT 25.150 115.730 25.290 116.230 ;
        RECT 25.090 115.410 25.350 115.730 ;
        RECT 25.150 107.230 25.290 115.410 ;
        RECT 26.070 115.130 26.210 119.830 ;
        RECT 26.470 117.110 26.730 117.430 ;
        RECT 25.610 114.990 26.210 115.130 ;
        RECT 25.610 114.710 25.750 114.990 ;
        RECT 25.550 114.390 25.810 114.710 ;
        RECT 26.530 114.450 26.670 117.110 ;
        RECT 25.610 111.900 25.750 114.390 ;
        RECT 26.070 114.310 26.670 114.450 ;
        RECT 26.070 112.670 26.210 114.310 ;
        RECT 26.010 112.350 26.270 112.670 ;
        RECT 25.610 111.760 26.210 111.900 ;
        RECT 25.550 109.970 25.810 110.290 ;
        RECT 25.610 108.250 25.750 109.970 ;
        RECT 25.550 107.930 25.810 108.250 ;
        RECT 26.070 107.230 26.210 111.760 ;
        RECT 27.390 111.670 27.650 111.990 ;
        RECT 27.450 107.570 27.590 111.670 ;
        RECT 27.390 107.250 27.650 107.570 ;
        RECT 25.090 106.910 25.350 107.230 ;
        RECT 26.010 106.910 26.270 107.230 ;
        RECT 26.470 104.190 26.730 104.510 ;
        RECT 24.170 100.790 24.430 101.110 ;
        RECT 24.230 99.410 24.370 100.790 ;
        RECT 26.530 100.090 26.670 104.190 ;
        RECT 26.470 99.770 26.730 100.090 ;
        RECT 24.170 99.090 24.430 99.410 ;
        RECT 27.910 96.690 28.050 130.710 ;
        RECT 28.770 126.630 29.030 126.950 ;
        RECT 28.830 115.730 28.970 126.630 ;
        RECT 28.310 115.410 28.570 115.730 ;
        RECT 28.770 115.410 29.030 115.730 ;
        RECT 28.370 108.250 28.510 115.410 ;
        RECT 28.770 112.350 29.030 112.670 ;
        RECT 28.830 110.970 28.970 112.350 ;
        RECT 28.770 110.650 29.030 110.970 ;
        RECT 28.310 107.930 28.570 108.250 ;
        RECT 29.290 105.530 29.430 164.530 ;
        RECT 31.070 161.310 31.330 161.630 ;
        RECT 31.990 161.310 32.250 161.630 ;
        RECT 33.830 161.310 34.090 161.630 ;
        RECT 31.130 157.210 31.270 161.310 ;
        RECT 31.070 156.890 31.330 157.210 ;
        RECT 31.530 155.870 31.790 156.190 ;
        RECT 31.590 150.870 31.730 155.870 ;
        RECT 31.130 150.730 31.730 150.870 ;
        RECT 29.690 148.730 29.950 149.050 ;
        RECT 29.750 145.650 29.890 148.730 ;
        RECT 31.130 148.370 31.270 150.730 ;
        RECT 31.070 148.050 31.330 148.370 ;
        RECT 29.690 145.330 29.950 145.650 ;
        RECT 29.750 140.210 29.890 145.330 ;
        RECT 31.130 145.310 31.270 148.050 ;
        RECT 32.050 145.990 32.190 161.310 ;
        RECT 33.370 160.630 33.630 160.950 ;
        RECT 33.430 159.930 33.570 160.630 ;
        RECT 33.370 159.610 33.630 159.930 ;
        RECT 33.890 157.210 34.030 161.310 ;
        RECT 33.830 156.890 34.090 157.210 ;
        RECT 34.290 155.190 34.550 155.510 ;
        RECT 34.350 154.150 34.490 155.190 ;
        RECT 34.290 153.830 34.550 154.150 ;
        RECT 35.730 150.750 35.870 165.050 ;
        RECT 36.190 159.590 36.330 193.610 ;
        RECT 38.030 191.210 38.170 193.610 ;
        RECT 41.250 192.230 41.390 196.670 ;
        RECT 42.170 192.570 42.310 197.350 ;
        RECT 42.630 195.290 42.770 204.830 ;
        RECT 47.170 204.490 47.430 204.810 ;
        RECT 45.790 204.150 46.050 204.470 ;
        RECT 45.330 202.110 45.590 202.430 ;
        RECT 43.950 201.430 44.210 201.750 ;
        RECT 44.410 201.430 44.670 201.750 ;
        RECT 43.030 199.565 43.290 199.710 ;
        RECT 43.020 199.195 43.300 199.565 ;
        RECT 44.010 199.370 44.150 201.430 ;
        RECT 44.470 200.730 44.610 201.430 ;
        RECT 45.390 200.730 45.530 202.110 ;
        RECT 44.410 200.410 44.670 200.730 ;
        RECT 45.330 200.410 45.590 200.730 ;
        RECT 43.950 199.050 44.210 199.370 ;
        RECT 44.010 197.670 44.150 199.050 ;
        RECT 43.950 197.350 44.210 197.670 ;
        RECT 42.570 194.970 42.830 195.290 ;
        RECT 42.110 192.250 42.370 192.570 ;
        RECT 41.190 191.910 41.450 192.230 ;
        RECT 37.970 190.890 38.230 191.210 ;
        RECT 38.710 190.015 40.250 190.385 ;
        RECT 41.250 189.850 41.390 191.910 ;
        RECT 41.190 189.530 41.450 189.850 ;
        RECT 36.590 186.130 36.850 186.450 ;
        RECT 37.510 186.130 37.770 186.450 ;
        RECT 36.650 183.050 36.790 186.130 ;
        RECT 37.050 185.110 37.310 185.430 ;
        RECT 36.590 182.730 36.850 183.050 ;
        RECT 37.110 181.690 37.250 185.110 ;
        RECT 37.570 181.690 37.710 186.130 ;
        RECT 37.970 185.110 38.230 185.430 ;
        RECT 38.030 183.050 38.170 185.110 ;
        RECT 38.710 184.575 40.250 184.945 ;
        RECT 37.970 182.730 38.230 183.050 ;
        RECT 37.050 181.370 37.310 181.690 ;
        RECT 37.510 181.370 37.770 181.690 ;
        RECT 42.170 181.010 42.310 192.250 ;
        RECT 43.030 191.570 43.290 191.890 ;
        RECT 43.090 190.870 43.230 191.570 ;
        RECT 43.030 190.550 43.290 190.870 ;
        RECT 45.330 188.510 45.590 188.830 ;
        RECT 44.870 186.130 45.130 186.450 ;
        RECT 42.570 184.090 42.830 184.410 ;
        RECT 42.110 180.690 42.370 181.010 ;
        RECT 42.170 179.990 42.310 180.690 ;
        RECT 42.110 179.670 42.370 179.990 ;
        RECT 38.710 179.135 40.250 179.505 ;
        RECT 37.050 177.630 37.310 177.950 ;
        RECT 37.110 174.550 37.250 177.630 ;
        RECT 37.510 175.250 37.770 175.570 ;
        RECT 37.050 174.230 37.310 174.550 ;
        RECT 36.590 172.190 36.850 172.510 ;
        RECT 36.650 170.810 36.790 172.190 ;
        RECT 36.590 170.490 36.850 170.810 ;
        RECT 37.110 169.790 37.250 174.230 ;
        RECT 37.570 173.530 37.710 175.250 ;
        RECT 37.970 174.230 38.230 174.550 ;
        RECT 37.510 173.210 37.770 173.530 ;
        RECT 38.030 172.510 38.170 174.230 ;
        RECT 38.710 173.695 40.250 174.065 ;
        RECT 37.970 172.190 38.230 172.510 ;
        RECT 37.510 171.510 37.770 171.830 ;
        RECT 37.570 170.810 37.710 171.510 ;
        RECT 37.510 170.490 37.770 170.810 ;
        RECT 38.030 170.470 38.170 172.190 ;
        RECT 37.970 170.150 38.230 170.470 ;
        RECT 40.270 169.810 40.530 170.130 ;
        RECT 37.050 169.470 37.310 169.790 ;
        RECT 40.330 169.530 40.470 169.810 ;
        RECT 40.330 169.390 40.930 169.530 ;
        RECT 37.970 168.790 38.230 169.110 ;
        RECT 37.050 166.750 37.310 167.070 ;
        RECT 37.110 164.670 37.250 166.750 ;
        RECT 38.030 166.390 38.170 168.790 ;
        RECT 38.710 168.255 40.250 168.625 ;
        RECT 40.790 168.000 40.930 169.390 ;
        RECT 40.330 167.860 40.930 168.000 ;
        RECT 37.970 166.070 38.230 166.390 ;
        RECT 40.330 165.370 40.470 167.860 ;
        RECT 40.270 165.050 40.530 165.370 ;
        RECT 37.110 164.530 38.170 164.670 ;
        RECT 37.510 161.990 37.770 162.310 ;
        RECT 37.050 161.310 37.310 161.630 ;
        RECT 36.590 160.630 36.850 160.950 ;
        RECT 36.130 159.270 36.390 159.590 ;
        RECT 36.650 157.210 36.790 160.630 ;
        RECT 37.110 159.930 37.250 161.310 ;
        RECT 37.050 159.610 37.310 159.930 ;
        RECT 36.590 156.890 36.850 157.210 ;
        RECT 36.590 156.210 36.850 156.530 ;
        RECT 32.910 150.430 33.170 150.750 ;
        RECT 34.290 150.430 34.550 150.750 ;
        RECT 35.670 150.430 35.930 150.750 ;
        RECT 32.970 149.050 33.110 150.430 ;
        RECT 33.830 149.750 34.090 150.070 ;
        RECT 32.910 148.730 33.170 149.050 ;
        RECT 33.890 148.710 34.030 149.750 ;
        RECT 33.830 148.390 34.090 148.710 ;
        RECT 34.350 146.330 34.490 150.430 ;
        RECT 34.290 146.010 34.550 146.330 ;
        RECT 35.730 145.990 35.870 150.430 ;
        RECT 36.650 150.410 36.790 156.210 ;
        RECT 37.110 155.850 37.250 159.610 ;
        RECT 37.570 157.210 37.710 161.990 ;
        RECT 38.030 158.910 38.170 164.530 ;
        RECT 38.710 162.815 40.250 163.185 ;
        RECT 38.890 162.330 39.150 162.650 ;
        RECT 38.950 161.630 39.090 162.330 ;
        RECT 38.890 161.310 39.150 161.630 ;
        RECT 37.970 158.590 38.230 158.910 ;
        RECT 38.030 157.210 38.170 158.590 ;
        RECT 38.710 157.375 40.250 157.745 ;
        RECT 37.510 156.890 37.770 157.210 ;
        RECT 37.970 156.890 38.230 157.210 ;
        RECT 42.170 156.190 42.310 179.670 ;
        RECT 42.630 178.630 42.770 184.090 ;
        RECT 43.950 178.650 44.210 178.970 ;
        RECT 42.570 178.310 42.830 178.630 ;
        RECT 44.010 177.270 44.150 178.650 ;
        RECT 43.950 176.950 44.210 177.270 ;
        RECT 44.410 176.950 44.670 177.270 ;
        RECT 44.010 175.910 44.150 176.950 ;
        RECT 43.950 175.590 44.210 175.910 ;
        RECT 44.470 174.890 44.610 176.950 ;
        RECT 44.410 174.570 44.670 174.890 ;
        RECT 43.490 172.870 43.750 173.190 ;
        RECT 43.550 170.130 43.690 172.870 ;
        RECT 44.930 172.250 45.070 186.130 ;
        RECT 45.390 185.770 45.530 188.510 ;
        RECT 45.330 185.450 45.590 185.770 ;
        RECT 45.390 178.290 45.530 185.450 ;
        RECT 45.330 177.970 45.590 178.290 ;
        RECT 44.930 172.110 45.530 172.250 ;
        RECT 45.850 172.170 45.990 204.150 ;
        RECT 47.230 199.710 47.370 204.490 ;
        RECT 47.630 204.150 47.890 204.470 ;
        RECT 49.010 204.150 49.270 204.470 ;
        RECT 47.170 199.390 47.430 199.710 ;
        RECT 46.250 191.570 46.510 191.890 ;
        RECT 46.310 189.850 46.450 191.570 ;
        RECT 46.250 189.530 46.510 189.850 ;
        RECT 46.710 189.530 46.970 189.850 ;
        RECT 46.250 189.080 46.510 189.170 ;
        RECT 46.770 189.080 46.910 189.530 ;
        RECT 46.250 188.940 46.910 189.080 ;
        RECT 46.250 188.850 46.510 188.940 ;
        RECT 47.170 185.110 47.430 185.430 ;
        RECT 46.250 182.730 46.510 183.050 ;
        RECT 46.310 181.690 46.450 182.730 ;
        RECT 47.230 181.690 47.370 185.110 ;
        RECT 46.250 181.370 46.510 181.690 ;
        RECT 47.170 181.370 47.430 181.690 ;
        RECT 47.170 176.950 47.430 177.270 ;
        RECT 46.250 175.250 46.510 175.570 ;
        RECT 46.310 173.530 46.450 175.250 ;
        RECT 46.250 173.210 46.510 173.530 ;
        RECT 44.410 171.510 44.670 171.830 ;
        RECT 44.870 171.510 45.130 171.830 ;
        RECT 44.470 170.810 44.610 171.510 ;
        RECT 44.410 170.490 44.670 170.810 ;
        RECT 44.930 170.130 45.070 171.510 ;
        RECT 43.490 169.810 43.750 170.130 ;
        RECT 44.870 169.810 45.130 170.130 ;
        RECT 42.570 169.130 42.830 169.450 ;
        RECT 42.630 168.090 42.770 169.130 ;
        RECT 42.570 167.770 42.830 168.090 ;
        RECT 43.550 167.750 43.690 169.810 ;
        RECT 43.490 167.430 43.750 167.750 ;
        RECT 44.930 167.070 45.070 169.810 ;
        RECT 45.390 167.070 45.530 172.110 ;
        RECT 45.790 171.850 46.050 172.170 ;
        RECT 46.710 171.850 46.970 172.170 ;
        RECT 46.250 171.510 46.510 171.830 ;
        RECT 45.790 169.810 46.050 170.130 ;
        RECT 44.870 166.750 45.130 167.070 ;
        RECT 45.330 166.750 45.590 167.070 ;
        RECT 44.410 166.070 44.670 166.390 ;
        RECT 44.470 163.670 44.610 166.070 ;
        RECT 44.410 163.350 44.670 163.670 ;
        RECT 44.930 161.630 45.070 166.750 ;
        RECT 45.850 166.730 45.990 169.810 ;
        RECT 45.790 166.410 46.050 166.730 ;
        RECT 45.850 161.970 45.990 166.410 ;
        RECT 46.310 162.650 46.450 171.510 ;
        RECT 46.250 162.330 46.510 162.650 ;
        RECT 45.790 161.650 46.050 161.970 ;
        RECT 44.870 161.540 45.130 161.630 ;
        RECT 44.870 161.400 45.530 161.540 ;
        RECT 44.870 161.310 45.130 161.400 ;
        RECT 44.410 160.630 44.670 160.950 ;
        RECT 42.110 155.870 42.370 156.190 ;
        RECT 37.050 155.530 37.310 155.850 ;
        RECT 39.810 155.530 40.070 155.850 ;
        RECT 39.870 154.490 40.010 155.530 ;
        RECT 39.810 154.170 40.070 154.490 ;
        RECT 42.170 154.150 42.310 155.870 ;
        RECT 42.110 153.830 42.370 154.150 ;
        RECT 38.710 151.935 40.250 152.305 ;
        RECT 42.170 151.770 42.310 153.830 ;
        RECT 44.470 152.790 44.610 160.630 ;
        RECT 45.390 159.930 45.530 161.400 ;
        RECT 45.330 159.840 45.590 159.930 ;
        RECT 44.930 159.700 45.590 159.840 ;
        RECT 44.930 157.210 45.070 159.700 ;
        RECT 45.330 159.610 45.590 159.700 ;
        RECT 45.330 157.910 45.590 158.230 ;
        RECT 44.870 156.890 45.130 157.210 ;
        RECT 44.930 153.810 45.070 156.890 ;
        RECT 45.390 154.490 45.530 157.910 ;
        RECT 46.250 155.190 46.510 155.510 ;
        RECT 46.310 154.490 46.450 155.190 ;
        RECT 45.330 154.170 45.590 154.490 ;
        RECT 46.250 154.170 46.510 154.490 ;
        RECT 44.870 153.490 45.130 153.810 ;
        RECT 44.410 152.470 44.670 152.790 ;
        RECT 42.110 151.450 42.370 151.770 ;
        RECT 40.730 150.430 40.990 150.750 ;
        RECT 43.030 150.430 43.290 150.750 ;
        RECT 36.590 150.090 36.850 150.410 ;
        RECT 40.790 147.350 40.930 150.430 ;
        RECT 41.190 149.750 41.450 150.070 ;
        RECT 41.250 148.370 41.390 149.750 ;
        RECT 41.190 148.050 41.450 148.370 ;
        RECT 37.970 147.030 38.230 147.350 ;
        RECT 40.730 147.030 40.990 147.350 ;
        RECT 38.030 145.990 38.170 147.030 ;
        RECT 38.710 146.495 40.250 146.865 ;
        RECT 31.990 145.670 32.250 145.990 ;
        RECT 35.210 145.670 35.470 145.990 ;
        RECT 35.670 145.670 35.930 145.990 ;
        RECT 37.050 145.670 37.310 145.990 ;
        RECT 37.970 145.670 38.230 145.990 ;
        RECT 31.070 144.990 31.330 145.310 ;
        RECT 31.530 144.310 31.790 144.630 ;
        RECT 29.690 139.890 29.950 140.210 ;
        RECT 30.610 134.110 30.870 134.430 ;
        RECT 29.690 133.770 29.950 134.090 ;
        RECT 29.750 116.410 29.890 133.770 ;
        RECT 30.670 131.370 30.810 134.110 ;
        RECT 31.590 134.090 31.730 144.310 ;
        RECT 33.830 141.930 34.090 142.250 ;
        RECT 33.890 140.890 34.030 141.930 ;
        RECT 33.830 140.570 34.090 140.890 ;
        RECT 34.750 140.230 35.010 140.550 ;
        RECT 32.450 139.890 32.710 140.210 ;
        RECT 32.510 139.190 32.650 139.890 ;
        RECT 31.990 138.870 32.250 139.190 ;
        RECT 32.450 138.870 32.710 139.190 ;
        RECT 32.050 138.170 32.190 138.870 ;
        RECT 31.990 137.850 32.250 138.170 ;
        RECT 33.370 137.170 33.630 137.490 ;
        RECT 34.290 137.170 34.550 137.490 ;
        RECT 33.430 135.450 33.570 137.170 ;
        RECT 33.370 135.130 33.630 135.450 ;
        RECT 32.910 134.450 33.170 134.770 ;
        RECT 31.990 134.110 32.250 134.430 ;
        RECT 31.530 133.770 31.790 134.090 ;
        RECT 30.610 131.050 30.870 131.370 ;
        RECT 30.150 129.690 30.410 130.010 ;
        RECT 30.210 120.570 30.350 129.690 ;
        RECT 30.670 126.950 30.810 131.050 ;
        RECT 31.590 131.030 31.730 133.770 ;
        RECT 32.050 132.050 32.190 134.110 ;
        RECT 32.970 132.730 33.110 134.450 ;
        RECT 34.350 134.430 34.490 137.170 ;
        RECT 34.810 136.810 34.950 140.230 ;
        RECT 34.750 136.490 35.010 136.810 ;
        RECT 34.810 134.430 34.950 136.490 ;
        RECT 34.290 134.110 34.550 134.430 ;
        RECT 34.750 134.110 35.010 134.430 ;
        RECT 32.910 132.410 33.170 132.730 ;
        RECT 31.990 131.730 32.250 132.050 ;
        RECT 32.050 131.450 32.190 131.730 ;
        RECT 32.050 131.310 32.650 131.450 ;
        RECT 31.530 130.710 31.790 131.030 ;
        RECT 31.990 130.710 32.250 131.030 ;
        RECT 32.050 128.990 32.190 130.710 ;
        RECT 32.510 128.990 32.650 131.310 ;
        RECT 33.830 130.710 34.090 131.030 ;
        RECT 33.890 130.090 34.030 130.710 ;
        RECT 33.430 130.010 34.030 130.090 ;
        RECT 33.370 129.950 34.030 130.010 ;
        RECT 33.370 129.690 33.630 129.950 ;
        RECT 31.990 128.670 32.250 128.990 ;
        RECT 32.450 128.670 32.710 128.990 ;
        RECT 31.530 127.990 31.790 128.310 ;
        RECT 30.610 126.630 30.870 126.950 ;
        RECT 31.590 125.590 31.730 127.990 ;
        RECT 32.510 126.610 32.650 128.670 ;
        RECT 33.370 126.630 33.630 126.950 ;
        RECT 32.450 126.290 32.710 126.610 ;
        RECT 31.530 125.270 31.790 125.590 ;
        RECT 30.610 122.550 30.870 122.870 ;
        RECT 31.070 122.550 31.330 122.870 ;
        RECT 30.670 121.170 30.810 122.550 ;
        RECT 31.130 121.850 31.270 122.550 ;
        RECT 31.070 121.530 31.330 121.850 ;
        RECT 30.610 120.850 30.870 121.170 ;
        RECT 31.070 120.850 31.330 121.170 ;
        RECT 31.130 120.570 31.270 120.850 ;
        RECT 30.210 120.430 31.270 120.570 ;
        RECT 31.130 118.110 31.270 120.430 ;
        RECT 31.070 117.790 31.330 118.110 ;
        RECT 31.590 117.770 31.730 125.270 ;
        RECT 32.510 121.850 32.650 126.290 ;
        RECT 33.430 121.850 33.570 126.630 ;
        RECT 33.830 126.290 34.090 126.610 ;
        RECT 33.890 124.570 34.030 126.290 ;
        RECT 33.830 124.250 34.090 124.570 ;
        RECT 34.290 123.230 34.550 123.550 ;
        RECT 34.350 121.850 34.490 123.230 ;
        RECT 35.270 122.870 35.410 145.670 ;
        RECT 37.110 143.270 37.250 145.670 ;
        RECT 37.970 144.990 38.230 145.310 ;
        RECT 37.050 142.950 37.310 143.270 ;
        RECT 37.510 142.950 37.770 143.270 ;
        RECT 37.110 142.590 37.250 142.950 ;
        RECT 37.050 142.270 37.310 142.590 ;
        RECT 36.590 141.590 36.850 141.910 ;
        RECT 36.650 139.530 36.790 141.590 ;
        RECT 37.570 139.870 37.710 142.950 ;
        RECT 38.030 142.930 38.170 144.990 ;
        RECT 43.090 143.610 43.230 150.430 ;
        RECT 44.870 150.090 45.130 150.410 ;
        RECT 45.330 150.090 45.590 150.410 ;
        RECT 43.030 143.290 43.290 143.610 ;
        RECT 44.410 143.290 44.670 143.610 ;
        RECT 37.970 142.610 38.230 142.930 ;
        RECT 43.030 142.610 43.290 142.930 ;
        RECT 40.730 141.930 40.990 142.250 ;
        RECT 38.710 141.055 40.250 141.425 ;
        RECT 40.790 140.890 40.930 141.930 ;
        RECT 42.110 141.590 42.370 141.910 ;
        RECT 40.730 140.570 40.990 140.890 ;
        RECT 41.190 140.570 41.450 140.890 ;
        RECT 37.510 139.550 37.770 139.870 ;
        RECT 36.590 139.210 36.850 139.530 ;
        RECT 36.130 138.870 36.390 139.190 ;
        RECT 36.190 137.490 36.330 138.870 ;
        RECT 36.650 138.170 36.790 139.210 ;
        RECT 36.590 137.850 36.850 138.170 ;
        RECT 36.130 137.170 36.390 137.490 ;
        RECT 38.710 135.615 40.250 135.985 ;
        RECT 36.590 133.770 36.850 134.090 ;
        RECT 35.670 131.390 35.930 131.710 ;
        RECT 35.730 128.310 35.870 131.390 ;
        RECT 35.670 127.990 35.930 128.310 ;
        RECT 36.650 126.950 36.790 133.770 ;
        RECT 41.250 132.050 41.390 140.570 ;
        RECT 42.170 138.170 42.310 141.590 ;
        RECT 43.090 140.890 43.230 142.610 ;
        RECT 43.030 140.570 43.290 140.890 ;
        RECT 44.470 139.530 44.610 143.290 ;
        RECT 44.930 142.930 45.070 150.090 ;
        RECT 45.390 149.050 45.530 150.090 ;
        RECT 45.330 148.730 45.590 149.050 ;
        RECT 45.330 144.990 45.590 145.310 ;
        RECT 45.390 143.270 45.530 144.990 ;
        RECT 45.330 142.950 45.590 143.270 ;
        RECT 44.870 142.610 45.130 142.930 ;
        RECT 46.770 142.250 46.910 171.850 ;
        RECT 47.230 170.810 47.370 176.950 ;
        RECT 47.690 172.510 47.830 204.150 ;
        RECT 49.070 203.450 49.210 204.150 ;
        RECT 49.530 203.450 49.670 204.830 ;
        RECT 53.610 204.150 53.870 204.470 ;
        RECT 49.010 203.130 49.270 203.450 ;
        RECT 49.470 203.130 49.730 203.450 ;
        RECT 53.670 203.110 53.810 204.150 ;
        RECT 53.610 202.790 53.870 203.110 ;
        RECT 51.770 202.110 52.030 202.430 ;
        RECT 49.470 200.070 49.730 200.390 ;
        RECT 49.530 197.330 49.670 200.070 ;
        RECT 51.830 199.710 51.970 202.110 ;
        RECT 52.220 201.235 52.500 201.605 ;
        RECT 52.290 200.730 52.430 201.235 ;
        RECT 52.230 200.410 52.490 200.730 ;
        RECT 51.770 199.390 52.030 199.710 ;
        RECT 53.150 199.390 53.410 199.710 ;
        RECT 53.210 198.010 53.350 199.390 ;
        RECT 53.150 197.690 53.410 198.010 ;
        RECT 49.470 197.010 49.730 197.330 ;
        RECT 54.130 196.990 54.270 204.830 ;
        RECT 57.290 204.490 57.550 204.810 ;
        RECT 60.050 204.490 60.310 204.810 ;
        RECT 55.500 203.615 57.040 203.985 ;
        RECT 57.350 203.450 57.490 204.490 ;
        RECT 58.210 204.150 58.470 204.470 ;
        RECT 57.290 203.130 57.550 203.450 ;
        RECT 54.530 202.450 54.790 202.770 ;
        RECT 55.450 202.450 55.710 202.770 ;
        RECT 54.590 200.730 54.730 202.450 ;
        RECT 54.990 202.110 55.250 202.430 ;
        RECT 54.530 200.410 54.790 200.730 ;
        RECT 55.050 199.450 55.190 202.110 ;
        RECT 55.510 201.750 55.650 202.450 ;
        RECT 58.270 202.430 58.410 204.150 ;
        RECT 59.590 203.130 59.850 203.450 ;
        RECT 59.130 202.790 59.390 203.110 ;
        RECT 58.670 202.450 58.930 202.770 ;
        RECT 55.910 202.110 56.170 202.430 ;
        RECT 58.210 202.110 58.470 202.430 ;
        RECT 55.450 201.430 55.710 201.750 ;
        RECT 55.970 200.730 56.110 202.110 ;
        RECT 57.750 201.430 58.010 201.750 ;
        RECT 55.910 200.410 56.170 200.730 ;
        RECT 54.590 199.310 55.190 199.450 ;
        RECT 54.070 196.670 54.330 196.990 ;
        RECT 52.690 194.630 52.950 194.950 ;
        RECT 50.390 189.530 50.650 189.850 ;
        RECT 49.010 188.170 49.270 188.490 ;
        RECT 49.070 187.130 49.210 188.170 ;
        RECT 49.010 186.810 49.270 187.130 ;
        RECT 48.090 185.110 48.350 185.430 ;
        RECT 48.150 182.710 48.290 185.110 ;
        RECT 48.090 182.390 48.350 182.710 ;
        RECT 48.550 182.390 48.810 182.710 ;
        RECT 48.150 177.610 48.290 182.390 ;
        RECT 48.610 178.630 48.750 182.390 ;
        RECT 48.550 178.310 48.810 178.630 ;
        RECT 50.450 178.370 50.590 189.530 ;
        RECT 50.850 185.790 51.110 186.110 ;
        RECT 50.910 182.710 51.050 185.790 ;
        RECT 50.850 182.390 51.110 182.710 ;
        RECT 52.230 182.390 52.490 182.710 ;
        RECT 52.290 181.690 52.430 182.390 ;
        RECT 52.230 181.370 52.490 181.690 ;
        RECT 51.760 178.370 52.040 178.485 ;
        RECT 50.450 178.230 52.040 178.370 ;
        RECT 52.230 178.310 52.490 178.630 ;
        RECT 48.090 177.290 48.350 177.610 ;
        RECT 50.450 175.910 50.590 178.230 ;
        RECT 51.760 178.115 52.040 178.230 ;
        RECT 51.760 177.690 52.040 177.805 ;
        RECT 50.910 177.550 52.040 177.690 ;
        RECT 50.390 175.590 50.650 175.910 ;
        RECT 50.910 175.570 51.050 177.550 ;
        RECT 51.760 177.435 52.040 177.550 ;
        RECT 50.850 175.250 51.110 175.570 ;
        RECT 51.760 175.395 52.040 175.765 ;
        RECT 52.290 175.570 52.430 178.310 ;
        RECT 52.750 175.650 52.890 194.630 ;
        RECT 53.610 193.950 53.870 194.270 ;
        RECT 53.670 189.850 53.810 193.950 ;
        RECT 54.130 191.890 54.270 196.670 ;
        RECT 54.590 196.650 54.730 199.310 ;
        RECT 57.290 199.050 57.550 199.370 ;
        RECT 54.990 198.710 55.250 199.030 ;
        RECT 54.530 196.330 54.790 196.650 ;
        RECT 55.050 195.290 55.190 198.710 ;
        RECT 55.500 198.175 57.040 198.545 ;
        RECT 57.350 198.010 57.490 199.050 ;
        RECT 57.810 198.010 57.950 201.430 ;
        RECT 58.270 200.730 58.410 202.110 ;
        RECT 58.730 202.090 58.870 202.450 ;
        RECT 58.670 201.770 58.930 202.090 ;
        RECT 58.730 201.605 58.870 201.770 ;
        RECT 58.660 201.235 58.940 201.605 ;
        RECT 58.210 200.410 58.470 200.730 ;
        RECT 58.210 199.050 58.470 199.370 ;
        RECT 56.370 197.690 56.630 198.010 ;
        RECT 57.290 197.690 57.550 198.010 ;
        RECT 57.750 197.690 58.010 198.010 ;
        RECT 56.430 197.410 56.570 197.690 ;
        RECT 56.430 197.330 57.950 197.410 ;
        RECT 55.910 197.010 56.170 197.330 ;
        RECT 56.430 197.270 58.010 197.330 ;
        RECT 57.750 197.010 58.010 197.270 ;
        RECT 55.970 196.730 56.110 197.010 ;
        RECT 58.270 196.730 58.410 199.050 ;
        RECT 58.670 198.710 58.930 199.030 ;
        RECT 58.730 197.330 58.870 198.710 ;
        RECT 58.670 197.010 58.930 197.330 ;
        RECT 55.970 196.590 58.410 196.730 ;
        RECT 54.990 194.970 55.250 195.290 ;
        RECT 59.190 193.930 59.330 202.790 ;
        RECT 59.650 199.710 59.790 203.130 ;
        RECT 60.110 199.710 60.250 204.490 ;
        RECT 61.430 202.450 61.690 202.770 ;
        RECT 61.490 200.390 61.630 202.450 ;
        RECT 62.410 200.730 62.550 206.870 ;
        RECT 63.270 204.490 63.530 204.810 ;
        RECT 63.330 200.730 63.470 204.490 ;
        RECT 63.790 204.470 63.930 206.870 ;
        RECT 63.730 204.150 63.990 204.470 ;
        RECT 67.870 204.150 68.130 204.470 ;
        RECT 63.790 202.770 63.930 204.150 ;
        RECT 67.930 203.110 68.070 204.150 ;
        RECT 67.870 202.790 68.130 203.110 ;
        RECT 63.730 202.450 63.990 202.770 ;
        RECT 63.730 201.430 63.990 201.750 ;
        RECT 66.950 201.430 67.210 201.750 ;
        RECT 62.350 200.410 62.610 200.730 ;
        RECT 63.270 200.410 63.530 200.730 ;
        RECT 61.430 200.070 61.690 200.390 ;
        RECT 63.790 199.710 63.930 201.430 ;
        RECT 67.010 200.730 67.150 201.430 ;
        RECT 68.390 200.730 68.530 207.890 ;
        RECT 69.310 203.110 69.450 207.890 ;
        RECT 71.090 207.550 71.350 207.870 ;
        RECT 76.150 207.550 76.410 207.870 ;
        RECT 78.910 207.550 79.170 207.870 ;
        RECT 82.130 207.550 82.390 207.870 ;
        RECT 71.150 204.470 71.290 207.550 ;
        RECT 75.230 207.210 75.490 207.530 ;
        RECT 72.290 206.335 73.830 206.705 ;
        RECT 74.770 204.830 75.030 205.150 ;
        RECT 71.090 204.150 71.350 204.470 ;
        RECT 69.250 202.790 69.510 203.110 ;
        RECT 71.090 202.450 71.350 202.770 ;
        RECT 71.550 202.450 71.810 202.770 ;
        RECT 71.150 200.730 71.290 202.450 ;
        RECT 71.610 200.730 71.750 202.450 ;
        RECT 74.830 202.430 74.970 204.830 ;
        RECT 75.290 204.810 75.430 207.210 ;
        RECT 75.230 204.490 75.490 204.810 ;
        RECT 75.690 204.150 75.950 204.470 ;
        RECT 74.770 202.110 75.030 202.430 ;
        RECT 72.290 200.895 73.830 201.265 ;
        RECT 66.950 200.410 67.210 200.730 ;
        RECT 67.410 200.410 67.670 200.730 ;
        RECT 68.330 200.410 68.590 200.730 ;
        RECT 71.090 200.410 71.350 200.730 ;
        RECT 71.550 200.410 71.810 200.730 ;
        RECT 59.590 199.390 59.850 199.710 ;
        RECT 60.050 199.390 60.310 199.710 ;
        RECT 63.730 199.390 63.990 199.710 ;
        RECT 59.650 196.650 59.790 199.390 ;
        RECT 61.890 199.050 62.150 199.370 ;
        RECT 59.590 196.330 59.850 196.650 ;
        RECT 60.050 193.950 60.310 194.270 ;
        RECT 57.750 193.610 58.010 193.930 ;
        RECT 59.130 193.610 59.390 193.930 ;
        RECT 55.500 192.735 57.040 193.105 ;
        RECT 54.070 191.570 54.330 191.890 ;
        RECT 53.610 189.530 53.870 189.850 ;
        RECT 54.130 180.670 54.270 191.570 ;
        RECT 56.370 190.550 56.630 190.870 ;
        RECT 56.430 189.170 56.570 190.550 ;
        RECT 57.290 189.190 57.550 189.510 ;
        RECT 56.370 188.850 56.630 189.170 ;
        RECT 54.530 187.830 54.790 188.150 ;
        RECT 54.990 187.830 55.250 188.150 ;
        RECT 54.590 185.430 54.730 187.830 ;
        RECT 55.050 187.130 55.190 187.830 ;
        RECT 55.500 187.295 57.040 187.665 ;
        RECT 57.350 187.130 57.490 189.190 ;
        RECT 54.990 186.810 55.250 187.130 ;
        RECT 57.290 186.810 57.550 187.130 ;
        RECT 57.810 186.450 57.950 193.610 ;
        RECT 58.670 193.270 58.930 193.590 ;
        RECT 59.590 193.270 59.850 193.590 ;
        RECT 58.730 189.170 58.870 193.270 ;
        RECT 59.130 191.570 59.390 191.890 ;
        RECT 59.190 189.170 59.330 191.570 ;
        RECT 59.650 190.870 59.790 193.270 ;
        RECT 60.110 191.890 60.250 193.950 ;
        RECT 61.950 193.930 62.090 199.050 ;
        RECT 63.790 194.610 63.930 199.390 ;
        RECT 64.650 199.050 64.910 199.370 ;
        RECT 64.710 198.090 64.850 199.050 ;
        RECT 67.470 199.030 67.610 200.410 ;
        RECT 67.410 198.710 67.670 199.030 ;
        RECT 68.330 198.710 68.590 199.030 ;
        RECT 64.710 197.950 65.310 198.090 ;
        RECT 64.650 197.010 64.910 197.330 ;
        RECT 63.730 194.290 63.990 194.610 ;
        RECT 61.890 193.610 62.150 193.930 ;
        RECT 61.950 191.890 62.090 193.610 ;
        RECT 62.810 193.270 63.070 193.590 ;
        RECT 60.050 191.570 60.310 191.890 ;
        RECT 61.890 191.570 62.150 191.890 ;
        RECT 60.110 191.210 60.250 191.570 ;
        RECT 60.050 190.890 60.310 191.210 ;
        RECT 59.590 190.550 59.850 190.870 ;
        RECT 58.670 188.850 58.930 189.170 ;
        RECT 59.130 188.850 59.390 189.170 ;
        RECT 58.210 187.830 58.470 188.150 ;
        RECT 55.450 186.130 55.710 186.450 ;
        RECT 57.750 186.130 58.010 186.450 ;
        RECT 54.990 185.790 55.250 186.110 ;
        RECT 54.530 185.110 54.790 185.430 ;
        RECT 55.050 184.070 55.190 185.790 ;
        RECT 55.510 184.410 55.650 186.130 ;
        RECT 55.450 184.090 55.710 184.410 ;
        RECT 54.990 183.750 55.250 184.070 ;
        RECT 58.270 183.730 58.410 187.830 ;
        RECT 61.950 186.450 62.090 191.570 ;
        RECT 62.870 191.210 63.010 193.270 ;
        RECT 63.790 191.890 63.930 194.290 ;
        RECT 64.190 193.950 64.450 194.270 ;
        RECT 63.730 191.570 63.990 191.890 ;
        RECT 64.250 191.550 64.390 193.950 ;
        RECT 64.710 192.570 64.850 197.010 ;
        RECT 64.650 192.250 64.910 192.570 ;
        RECT 65.170 191.970 65.310 197.950 ;
        RECT 68.390 196.310 68.530 198.710 ;
        RECT 74.830 196.990 74.970 202.110 ;
        RECT 75.750 200.730 75.890 204.150 ;
        RECT 76.210 201.750 76.350 207.550 ;
        RECT 78.970 203.450 79.110 207.550 ;
        RECT 80.750 206.870 81.010 207.190 ;
        RECT 78.910 203.130 79.170 203.450 ;
        RECT 80.810 202.430 80.950 206.870 ;
        RECT 82.190 203.110 82.330 207.550 ;
        RECT 83.050 206.870 83.310 207.190 ;
        RECT 83.110 205.490 83.250 206.870 ;
        RECT 83.050 205.170 83.310 205.490 ;
        RECT 83.570 203.450 83.710 207.890 ;
        RECT 86.270 205.850 86.530 206.170 ;
        RECT 84.890 205.510 85.150 205.830 ;
        RECT 83.970 205.170 84.230 205.490 ;
        RECT 83.510 203.130 83.770 203.450 ;
        RECT 82.130 202.790 82.390 203.110 ;
        RECT 79.820 201.915 80.100 202.285 ;
        RECT 80.750 202.110 81.010 202.430 ;
        RECT 82.130 202.110 82.390 202.430 ;
        RECT 76.150 201.430 76.410 201.750 ;
        RECT 75.690 200.410 75.950 200.730 ;
        RECT 74.770 196.670 75.030 196.990 ;
        RECT 68.330 195.990 68.590 196.310 ;
        RECT 70.630 195.990 70.890 196.310 ;
        RECT 68.390 195.290 68.530 195.990 ;
        RECT 68.330 194.970 68.590 195.290 ;
        RECT 66.030 194.290 66.290 194.610 ;
        RECT 64.710 191.830 65.310 191.970 ;
        RECT 64.190 191.230 64.450 191.550 ;
        RECT 62.810 190.890 63.070 191.210 ;
        RECT 62.870 188.830 63.010 190.890 ;
        RECT 64.250 189.850 64.390 191.230 ;
        RECT 64.190 189.530 64.450 189.850 ;
        RECT 62.810 188.510 63.070 188.830 ;
        RECT 61.890 186.130 62.150 186.450 ;
        RECT 61.950 185.770 62.090 186.130 ;
        RECT 62.350 185.790 62.610 186.110 ;
        RECT 58.670 185.450 58.930 185.770 ;
        RECT 61.890 185.450 62.150 185.770 ;
        RECT 58.210 183.410 58.470 183.730 ;
        RECT 55.500 181.855 57.040 182.225 ;
        RECT 54.070 180.350 54.330 180.670 ;
        RECT 54.530 179.670 54.790 179.990 ;
        RECT 54.590 178.970 54.730 179.670 ;
        RECT 54.530 178.650 54.790 178.970 ;
        RECT 54.530 177.690 54.790 177.950 ;
        RECT 54.530 177.630 55.190 177.690 ;
        RECT 57.750 177.630 58.010 177.950 ;
        RECT 54.590 177.550 55.190 177.630 ;
        RECT 54.070 176.950 54.330 177.270 ;
        RECT 51.830 174.550 51.970 175.395 ;
        RECT 52.230 175.250 52.490 175.570 ;
        RECT 52.750 175.510 53.810 175.650 ;
        RECT 54.130 175.570 54.270 176.950 ;
        RECT 55.050 176.250 55.190 177.550 ;
        RECT 57.290 176.950 57.550 177.270 ;
        RECT 55.500 176.415 57.040 176.785 ;
        RECT 54.990 175.930 55.250 176.250 ;
        RECT 55.050 175.570 55.190 175.930 ;
        RECT 52.690 174.570 52.950 174.890 ;
        RECT 51.770 174.230 52.030 174.550 ;
        RECT 52.230 174.230 52.490 174.550 ;
        RECT 52.290 173.530 52.430 174.230 ;
        RECT 52.750 173.530 52.890 174.570 ;
        RECT 52.230 173.210 52.490 173.530 ;
        RECT 52.690 173.210 52.950 173.530 ;
        RECT 47.630 172.190 47.890 172.510 ;
        RECT 47.170 170.490 47.430 170.810 ;
        RECT 50.390 169.810 50.650 170.130 ;
        RECT 47.630 168.790 47.890 169.110 ;
        RECT 47.170 167.770 47.430 168.090 ;
        RECT 47.230 164.010 47.370 167.770 ;
        RECT 47.690 167.070 47.830 168.790 ;
        RECT 47.630 166.750 47.890 167.070 ;
        RECT 49.010 166.750 49.270 167.070 ;
        RECT 47.690 164.690 47.830 166.750 ;
        RECT 48.090 166.070 48.350 166.390 ;
        RECT 47.630 164.370 47.890 164.690 ;
        RECT 48.150 164.670 48.290 166.070 ;
        RECT 49.070 165.370 49.210 166.750 ;
        RECT 49.010 165.050 49.270 165.370 ;
        RECT 48.150 164.530 49.210 164.670 ;
        RECT 47.170 163.690 47.430 164.010 ;
        RECT 47.630 161.650 47.890 161.970 ;
        RECT 47.170 160.970 47.430 161.290 ;
        RECT 47.230 153.470 47.370 160.970 ;
        RECT 47.690 158.230 47.830 161.650 ;
        RECT 49.070 159.250 49.210 164.530 ;
        RECT 49.930 164.030 50.190 164.350 ;
        RECT 49.990 162.650 50.130 164.030 ;
        RECT 50.450 163.670 50.590 169.810 ;
        RECT 51.310 168.790 51.570 169.110 ;
        RECT 51.370 167.410 51.510 168.790 ;
        RECT 53.150 167.430 53.410 167.750 ;
        RECT 51.310 167.320 51.570 167.410 ;
        RECT 51.310 167.180 51.970 167.320 ;
        RECT 51.310 167.090 51.570 167.180 ;
        RECT 51.310 166.410 51.570 166.730 ;
        RECT 51.370 165.370 51.510 166.410 ;
        RECT 51.830 165.370 51.970 167.180 ;
        RECT 52.690 166.070 52.950 166.390 ;
        RECT 52.750 165.370 52.890 166.070 ;
        RECT 51.310 165.050 51.570 165.370 ;
        RECT 51.770 165.050 52.030 165.370 ;
        RECT 52.690 165.050 52.950 165.370 ;
        RECT 53.210 164.670 53.350 167.430 ;
        RECT 53.670 164.690 53.810 175.510 ;
        RECT 54.070 175.250 54.330 175.570 ;
        RECT 54.990 175.250 55.250 175.570 ;
        RECT 57.350 175.230 57.490 176.950 ;
        RECT 57.290 174.910 57.550 175.230 ;
        RECT 54.530 174.405 54.790 174.550 ;
        RECT 54.520 174.035 54.800 174.405 ;
        RECT 56.830 174.230 57.090 174.550 ;
        RECT 54.530 173.210 54.790 173.530 ;
        RECT 54.590 170.810 54.730 173.210 ;
        RECT 56.890 172.510 57.030 174.230 ;
        RECT 56.830 172.190 57.090 172.510 ;
        RECT 57.350 172.420 57.490 174.910 ;
        RECT 57.810 173.190 57.950 177.630 ;
        RECT 58.200 177.435 58.480 177.805 ;
        RECT 58.210 177.290 58.470 177.435 ;
        RECT 58.210 175.930 58.470 176.250 ;
        RECT 58.270 174.550 58.410 175.930 ;
        RECT 58.210 174.230 58.470 174.550 ;
        RECT 57.750 172.870 58.010 173.190 ;
        RECT 57.750 172.420 58.010 172.510 ;
        RECT 57.350 172.280 58.010 172.420 ;
        RECT 57.750 172.190 58.010 172.280 ;
        RECT 54.990 171.510 55.250 171.830 ;
        RECT 54.530 170.490 54.790 170.810 ;
        RECT 55.050 170.130 55.190 171.510 ;
        RECT 55.500 170.975 57.040 171.345 ;
        RECT 58.730 170.470 58.870 185.450 ;
        RECT 60.050 185.110 60.310 185.430 ;
        RECT 60.110 181.350 60.250 185.110 ;
        RECT 60.050 181.030 60.310 181.350 ;
        RECT 60.500 178.370 60.780 178.485 ;
        RECT 60.110 178.230 60.780 178.370 ;
        RECT 59.130 177.630 59.390 177.950 ;
        RECT 59.190 174.405 59.330 177.630 ;
        RECT 59.580 175.395 59.860 175.765 ;
        RECT 59.590 175.250 59.850 175.395 ;
        RECT 59.590 174.570 59.850 174.890 ;
        RECT 59.120 174.035 59.400 174.405 ;
        RECT 59.190 172.510 59.330 174.035 ;
        RECT 59.650 172.510 59.790 174.570 ;
        RECT 59.130 172.190 59.390 172.510 ;
        RECT 59.590 172.190 59.850 172.510 ;
        RECT 58.670 170.150 58.930 170.470 ;
        RECT 54.070 169.810 54.330 170.130 ;
        RECT 54.990 169.810 55.250 170.130 ;
        RECT 52.750 164.530 53.350 164.670 ;
        RECT 50.390 163.350 50.650 163.670 ;
        RECT 49.930 162.330 50.190 162.650 ;
        RECT 49.010 158.930 49.270 159.250 ;
        RECT 49.470 158.930 49.730 159.250 ;
        RECT 47.630 157.910 47.890 158.230 ;
        RECT 47.690 156.870 47.830 157.910 ;
        RECT 47.630 156.550 47.890 156.870 ;
        RECT 47.170 153.150 47.430 153.470 ;
        RECT 47.230 148.370 47.370 153.150 ;
        RECT 47.170 148.050 47.430 148.370 ;
        RECT 49.070 147.690 49.210 158.930 ;
        RECT 49.530 150.410 49.670 158.930 ;
        RECT 51.310 155.870 51.570 156.190 ;
        RECT 51.370 150.750 51.510 155.870 ;
        RECT 52.750 154.150 52.890 164.530 ;
        RECT 53.610 164.370 53.870 164.690 ;
        RECT 54.130 164.090 54.270 169.810 ;
        RECT 55.050 167.490 55.190 169.810 ;
        RECT 58.210 169.130 58.470 169.450 ;
        RECT 57.290 168.790 57.550 169.110 ;
        RECT 55.050 167.350 55.650 167.490 ;
        RECT 55.510 167.070 55.650 167.350 ;
        RECT 54.990 166.750 55.250 167.070 ;
        RECT 55.450 166.750 55.710 167.070 ;
        RECT 57.350 166.810 57.490 168.790 ;
        RECT 55.050 164.350 55.190 166.750 ;
        RECT 57.350 166.670 57.950 166.810 ;
        RECT 57.290 166.070 57.550 166.390 ;
        RECT 55.500 165.535 57.040 165.905 ;
        RECT 57.350 165.370 57.490 166.070 ;
        RECT 57.290 165.050 57.550 165.370 ;
        RECT 57.810 164.690 57.950 166.670 ;
        RECT 58.270 165.370 58.410 169.130 ;
        RECT 58.730 167.070 58.870 170.150 ;
        RECT 59.590 167.090 59.850 167.410 ;
        RECT 58.670 166.750 58.930 167.070 ;
        RECT 59.130 166.410 59.390 166.730 ;
        RECT 58.210 165.050 58.470 165.370 ;
        RECT 57.750 164.370 58.010 164.690 ;
        RECT 58.670 164.370 58.930 164.690 ;
        RECT 53.210 164.010 54.270 164.090 ;
        RECT 54.990 164.030 55.250 164.350 ;
        RECT 53.150 163.950 54.270 164.010 ;
        RECT 53.150 163.690 53.410 163.950 ;
        RECT 54.530 163.690 54.790 164.010 ;
        RECT 52.690 153.830 52.950 154.150 ;
        RECT 51.770 152.470 52.030 152.790 ;
        RECT 50.390 150.430 50.650 150.750 ;
        RECT 51.310 150.430 51.570 150.750 ;
        RECT 49.470 150.090 49.730 150.410 ;
        RECT 49.010 147.370 49.270 147.690 ;
        RECT 49.070 145.310 49.210 147.370 ;
        RECT 50.450 147.350 50.590 150.430 ;
        RECT 51.370 148.370 51.510 150.430 ;
        RECT 51.310 148.050 51.570 148.370 ;
        RECT 50.390 147.030 50.650 147.350 ;
        RECT 49.010 144.990 49.270 145.310 ;
        RECT 46.710 141.930 46.970 142.250 ;
        RECT 50.450 139.870 50.590 147.030 ;
        RECT 51.370 142.930 51.510 148.050 ;
        RECT 51.830 145.310 51.970 152.470 ;
        RECT 52.230 148.050 52.490 148.370 ;
        RECT 52.290 146.330 52.430 148.050 ;
        RECT 52.230 146.010 52.490 146.330 ;
        RECT 51.770 144.990 52.030 145.310 ;
        RECT 51.310 142.610 51.570 142.930 ;
        RECT 51.370 140.210 51.510 142.610 ;
        RECT 51.310 139.890 51.570 140.210 ;
        RECT 50.390 139.550 50.650 139.870 ;
        RECT 44.410 139.210 44.670 139.530 ;
        RECT 42.110 137.850 42.370 138.170 ;
        RECT 52.750 137.150 52.890 153.830 ;
        RECT 54.590 147.350 54.730 163.690 ;
        RECT 55.050 162.650 55.190 164.030 ;
        RECT 58.730 162.650 58.870 164.370 ;
        RECT 54.990 162.330 55.250 162.650 ;
        RECT 58.670 162.330 58.930 162.650 ;
        RECT 58.670 161.650 58.930 161.970 ;
        RECT 54.990 161.310 55.250 161.630 ;
        RECT 55.050 159.930 55.190 161.310 ;
        RECT 57.750 160.970 58.010 161.290 ;
        RECT 57.290 160.630 57.550 160.950 ;
        RECT 55.500 160.095 57.040 160.465 ;
        RECT 57.350 159.930 57.490 160.630 ;
        RECT 54.990 159.610 55.250 159.930 ;
        RECT 57.290 159.610 57.550 159.930 ;
        RECT 57.810 159.330 57.950 160.970 ;
        RECT 58.210 160.630 58.470 160.950 ;
        RECT 57.350 159.250 57.950 159.330 ;
        RECT 57.290 159.190 57.950 159.250 ;
        RECT 57.290 158.930 57.550 159.190 ;
        RECT 54.990 158.250 55.250 158.570 ;
        RECT 55.050 152.790 55.190 158.250 ;
        RECT 57.350 157.210 57.490 158.930 ;
        RECT 58.270 158.910 58.410 160.630 ;
        RECT 58.210 158.590 58.470 158.910 ;
        RECT 57.290 156.890 57.550 157.210 ;
        RECT 55.500 154.655 57.040 155.025 ;
        RECT 58.270 154.490 58.410 158.590 ;
        RECT 58.730 156.190 58.870 161.650 ;
        RECT 59.190 159.930 59.330 166.410 ;
        RECT 59.650 164.690 59.790 167.090 ;
        RECT 59.590 164.370 59.850 164.690 ;
        RECT 60.110 164.670 60.250 178.230 ;
        RECT 60.500 178.115 60.780 178.230 ;
        RECT 60.510 174.910 60.770 175.230 ;
        RECT 60.570 173.530 60.710 174.910 ;
        RECT 60.510 173.210 60.770 173.530 ;
        RECT 60.970 172.190 61.230 172.510 ;
        RECT 61.030 170.810 61.170 172.190 ;
        RECT 60.970 170.490 61.230 170.810 ;
        RECT 61.950 168.090 62.090 185.450 ;
        RECT 61.890 167.770 62.150 168.090 ;
        RECT 60.110 164.530 60.710 164.670 ;
        RECT 60.050 164.030 60.310 164.350 ;
        RECT 59.590 160.630 59.850 160.950 ;
        RECT 59.130 159.610 59.390 159.930 ;
        RECT 59.650 158.230 59.790 160.630 ;
        RECT 59.130 157.910 59.390 158.230 ;
        RECT 59.590 157.910 59.850 158.230 ;
        RECT 58.670 155.870 58.930 156.190 ;
        RECT 58.210 154.170 58.470 154.490 ;
        RECT 59.190 153.810 59.330 157.910 ;
        RECT 59.650 157.210 59.790 157.910 ;
        RECT 59.590 156.890 59.850 157.210 ;
        RECT 59.130 153.490 59.390 153.810 ;
        RECT 57.750 153.150 58.010 153.470 ;
        RECT 54.990 152.470 55.250 152.790 ;
        RECT 55.500 149.215 57.040 149.585 ;
        RECT 57.810 149.050 57.950 153.150 ;
        RECT 60.110 150.750 60.250 164.030 ;
        RECT 60.570 151.170 60.710 164.530 ;
        RECT 60.970 163.690 61.230 164.010 ;
        RECT 61.030 162.650 61.170 163.690 ;
        RECT 60.970 162.330 61.230 162.650 ;
        RECT 62.410 154.490 62.550 185.790 ;
        RECT 63.730 185.110 63.990 185.430 ;
        RECT 63.790 183.050 63.930 185.110 ;
        RECT 63.730 182.730 63.990 183.050 ;
        RECT 63.270 177.290 63.530 177.610 ;
        RECT 63.330 176.250 63.470 177.290 ;
        RECT 64.190 176.950 64.450 177.270 ;
        RECT 63.270 175.930 63.530 176.250 ;
        RECT 64.250 175.570 64.390 176.950 ;
        RECT 64.710 175.570 64.850 191.830 ;
        RECT 65.110 189.530 65.370 189.850 ;
        RECT 65.170 186.450 65.310 189.530 ;
        RECT 65.110 186.130 65.370 186.450 ;
        RECT 65.170 185.770 65.310 186.130 ;
        RECT 65.110 185.450 65.370 185.770 ;
        RECT 65.110 180.350 65.370 180.670 ;
        RECT 65.170 178.970 65.310 180.350 ;
        RECT 65.110 178.650 65.370 178.970 ;
        RECT 64.190 175.250 64.450 175.570 ;
        RECT 64.650 175.250 64.910 175.570 ;
        RECT 62.810 174.910 63.070 175.230 ;
        RECT 62.870 172.510 63.010 174.910 ;
        RECT 64.250 172.510 64.390 175.250 ;
        RECT 62.810 172.190 63.070 172.510 ;
        RECT 64.190 172.190 64.450 172.510 ;
        RECT 63.730 164.370 63.990 164.690 ;
        RECT 63.790 162.650 63.930 164.370 ;
        RECT 63.730 162.330 63.990 162.650 ;
        RECT 64.250 161.630 64.390 172.190 ;
        RECT 65.110 171.510 65.370 171.830 ;
        RECT 65.170 170.470 65.310 171.510 ;
        RECT 65.110 170.150 65.370 170.470 ;
        RECT 64.190 161.310 64.450 161.630 ;
        RECT 62.810 156.890 63.070 157.210 ;
        RECT 62.350 154.170 62.610 154.490 ;
        RECT 62.870 153.470 63.010 156.890 ;
        RECT 62.810 153.150 63.070 153.470 ;
        RECT 60.570 151.030 61.170 151.170 ;
        RECT 60.050 150.430 60.310 150.750 ;
        RECT 61.030 150.070 61.170 151.030 ;
        RECT 62.350 150.430 62.610 150.750 ;
        RECT 60.970 149.750 61.230 150.070 ;
        RECT 61.890 149.750 62.150 150.070 ;
        RECT 57.750 148.730 58.010 149.050 ;
        RECT 61.030 147.690 61.170 149.750 ;
        RECT 60.970 147.370 61.230 147.690 ;
        RECT 61.430 147.370 61.690 147.690 ;
        RECT 54.530 147.030 54.790 147.350 ;
        RECT 59.130 147.030 59.390 147.350 ;
        RECT 54.590 145.650 54.730 147.030 ;
        RECT 59.190 145.990 59.330 147.030 ;
        RECT 59.130 145.670 59.390 145.990 ;
        RECT 54.530 145.330 54.790 145.650 ;
        RECT 53.610 145.050 53.870 145.310 ;
        RECT 53.610 144.990 54.730 145.050 ;
        RECT 53.670 144.910 54.730 144.990 ;
        RECT 54.590 144.630 54.730 144.910 ;
        RECT 54.530 144.310 54.790 144.630 ;
        RECT 54.990 144.310 55.250 144.630 ;
        RECT 53.150 142.610 53.410 142.930 ;
        RECT 53.210 140.890 53.350 142.610 ;
        RECT 53.150 140.570 53.410 140.890 ;
        RECT 54.590 139.530 54.730 144.310 ;
        RECT 55.050 139.870 55.190 144.310 ;
        RECT 55.500 143.775 57.040 144.145 ;
        RECT 54.990 139.550 55.250 139.870 ;
        RECT 54.530 139.210 54.790 139.530 ;
        RECT 57.750 139.210 58.010 139.530 ;
        RECT 54.590 137.490 54.730 139.210 ;
        RECT 55.500 138.335 57.040 138.705 ;
        RECT 57.810 137.490 57.950 139.210 ;
        RECT 59.190 138.170 59.330 145.670 ;
        RECT 61.490 143.610 61.630 147.370 ;
        RECT 61.950 146.330 62.090 149.750 ;
        RECT 61.890 146.010 62.150 146.330 ;
        RECT 62.410 145.310 62.550 150.430 ;
        RECT 62.870 148.370 63.010 153.150 ;
        RECT 64.250 153.130 64.390 161.310 ;
        RECT 66.090 161.290 66.230 194.290 ;
        RECT 66.950 193.950 67.210 194.270 ;
        RECT 67.010 192.570 67.150 193.950 ;
        RECT 66.950 192.250 67.210 192.570 ;
        RECT 67.870 191.570 68.130 191.890 ;
        RECT 66.490 190.890 66.750 191.210 ;
        RECT 66.550 172.170 66.690 190.890 ;
        RECT 67.930 187.130 68.070 191.570 ;
        RECT 68.390 188.830 68.530 194.970 ;
        RECT 68.790 193.610 69.050 193.930 ;
        RECT 68.850 192.570 68.990 193.610 ;
        RECT 69.250 193.270 69.510 193.590 ;
        RECT 68.790 192.250 69.050 192.570 ;
        RECT 68.330 188.510 68.590 188.830 ;
        RECT 69.310 188.490 69.450 193.270 ;
        RECT 70.690 191.890 70.830 195.990 ;
        RECT 72.290 195.455 73.830 195.825 ;
        RECT 74.310 194.630 74.570 194.950 ;
        RECT 74.370 192.230 74.510 194.630 ;
        RECT 74.770 193.270 75.030 193.590 ;
        RECT 74.830 192.570 74.970 193.270 ;
        RECT 74.770 192.250 75.030 192.570 ;
        RECT 74.310 191.910 74.570 192.230 ;
        RECT 69.710 191.570 69.970 191.890 ;
        RECT 70.630 191.570 70.890 191.890 ;
        RECT 74.770 191.570 75.030 191.890 ;
        RECT 75.230 191.570 75.490 191.890 ;
        RECT 69.250 188.170 69.510 188.490 ;
        RECT 67.870 186.810 68.130 187.130 ;
        RECT 68.330 186.810 68.590 187.130 ;
        RECT 66.950 179.670 67.210 179.990 ;
        RECT 67.010 175.570 67.150 179.670 ;
        RECT 66.950 175.250 67.210 175.570 ;
        RECT 66.490 171.850 66.750 172.170 ;
        RECT 66.030 160.970 66.290 161.290 ;
        RECT 66.030 158.930 66.290 159.250 ;
        RECT 65.110 155.190 65.370 155.510 ;
        RECT 65.170 154.490 65.310 155.190 ;
        RECT 66.090 154.490 66.230 158.930 ;
        RECT 64.650 154.170 64.910 154.490 ;
        RECT 65.110 154.170 65.370 154.490 ;
        RECT 66.030 154.170 66.290 154.490 ;
        RECT 64.710 153.810 64.850 154.170 ;
        RECT 64.650 153.490 64.910 153.810 ;
        RECT 64.190 152.810 64.450 153.130 ;
        RECT 64.710 151.430 64.850 153.490 ;
        RECT 66.030 151.450 66.290 151.770 ;
        RECT 64.650 151.110 64.910 151.430 ;
        RECT 63.270 150.430 63.530 150.750 ;
        RECT 63.730 150.430 63.990 150.750 ;
        RECT 64.650 150.660 64.910 150.750 ;
        RECT 64.650 150.520 65.310 150.660 ;
        RECT 64.650 150.430 64.910 150.520 ;
        RECT 63.330 148.710 63.470 150.430 ;
        RECT 63.270 148.390 63.530 148.710 ;
        RECT 62.810 148.050 63.070 148.370 ;
        RECT 62.350 144.990 62.610 145.310 ;
        RECT 61.430 143.290 61.690 143.610 ;
        RECT 62.410 142.930 62.550 144.990 ;
        RECT 63.330 144.630 63.470 148.390 ;
        RECT 63.790 148.370 63.930 150.430 ;
        RECT 64.190 149.750 64.450 150.070 ;
        RECT 64.650 149.750 64.910 150.070 ;
        RECT 63.730 148.050 63.990 148.370 ;
        RECT 63.270 144.310 63.530 144.630 ;
        RECT 63.330 143.610 63.470 144.310 ;
        RECT 63.270 143.290 63.530 143.610 ;
        RECT 63.790 142.930 63.930 148.050 ;
        RECT 64.250 144.970 64.390 149.750 ;
        RECT 64.710 145.990 64.850 149.750 ;
        RECT 65.170 147.690 65.310 150.520 ;
        RECT 65.570 149.750 65.830 150.070 ;
        RECT 65.110 147.370 65.370 147.690 ;
        RECT 65.170 145.990 65.310 147.370 ;
        RECT 64.650 145.670 64.910 145.990 ;
        RECT 65.110 145.670 65.370 145.990 ;
        RECT 65.170 145.310 65.310 145.670 ;
        RECT 64.650 144.990 64.910 145.310 ;
        RECT 65.110 144.990 65.370 145.310 ;
        RECT 64.190 144.650 64.450 144.970 ;
        RECT 62.350 142.610 62.610 142.930 ;
        RECT 63.730 142.610 63.990 142.930 ;
        RECT 59.590 141.590 59.850 141.910 ;
        RECT 59.650 140.210 59.790 141.590 ;
        RECT 62.410 140.405 62.550 142.610 ;
        RECT 59.590 139.890 59.850 140.210 ;
        RECT 60.110 140.150 61.170 140.290 ;
        RECT 60.110 139.870 60.250 140.150 ;
        RECT 61.030 140.120 61.170 140.150 ;
        RECT 61.030 139.980 62.090 140.120 ;
        RECT 62.340 140.035 62.620 140.405 ;
        RECT 60.050 139.550 60.310 139.870 ;
        RECT 61.430 139.210 61.690 139.530 ;
        RECT 60.050 138.870 60.310 139.190 ;
        RECT 60.110 138.170 60.250 138.870 ;
        RECT 59.130 137.850 59.390 138.170 ;
        RECT 60.050 137.850 60.310 138.170 ;
        RECT 54.070 137.170 54.330 137.490 ;
        RECT 54.530 137.170 54.790 137.490 ;
        RECT 54.990 137.170 55.250 137.490 ;
        RECT 57.750 137.170 58.010 137.490 ;
        RECT 60.970 137.170 61.230 137.490 ;
        RECT 52.690 136.830 52.950 137.150 ;
        RECT 53.150 136.830 53.410 137.150 ;
        RECT 42.110 136.150 42.370 136.470 ;
        RECT 52.230 136.150 52.490 136.470 ;
        RECT 42.170 134.430 42.310 136.150 ;
        RECT 50.850 135.130 51.110 135.450 ;
        RECT 42.110 134.110 42.370 134.430 ;
        RECT 50.390 134.110 50.650 134.430 ;
        RECT 42.170 132.390 42.310 134.110 ;
        RECT 42.110 132.070 42.370 132.390 ;
        RECT 37.510 131.730 37.770 132.050 ;
        RECT 41.190 131.730 41.450 132.050 ;
        RECT 37.570 130.010 37.710 131.730 ;
        RECT 40.730 130.710 40.990 131.030 ;
        RECT 38.710 130.175 40.250 130.545 ;
        RECT 37.510 129.690 37.770 130.010 ;
        RECT 38.430 128.900 38.690 128.990 ;
        RECT 38.030 128.760 38.690 128.900 ;
        RECT 37.050 127.990 37.310 128.310 ;
        RECT 36.590 126.630 36.850 126.950 ;
        RECT 36.650 123.210 36.790 126.630 ;
        RECT 36.590 122.890 36.850 123.210 ;
        RECT 35.210 122.550 35.470 122.870 ;
        RECT 32.450 121.530 32.710 121.850 ;
        RECT 33.370 121.530 33.630 121.850 ;
        RECT 34.290 121.530 34.550 121.850 ;
        RECT 31.990 120.850 32.250 121.170 ;
        RECT 32.050 119.130 32.190 120.850 ;
        RECT 31.990 118.810 32.250 119.130 ;
        RECT 31.530 117.450 31.790 117.770 ;
        RECT 29.690 116.090 29.950 116.410 ;
        RECT 32.510 115.730 32.650 121.530 ;
        RECT 36.650 121.510 36.790 122.890 ;
        RECT 37.110 121.510 37.250 127.990 ;
        RECT 37.510 125.950 37.770 126.270 ;
        RECT 37.570 124.570 37.710 125.950 ;
        RECT 37.510 124.250 37.770 124.570 ;
        RECT 36.590 121.190 36.850 121.510 ;
        RECT 37.050 121.190 37.310 121.510 ;
        RECT 37.570 121.170 37.710 124.250 ;
        RECT 37.510 120.850 37.770 121.170 ;
        RECT 35.670 119.830 35.930 120.150 ;
        RECT 35.730 118.020 35.870 119.830 ;
        RECT 35.730 117.880 36.790 118.020 ;
        RECT 33.370 117.450 33.630 117.770 ;
        RECT 33.830 117.450 34.090 117.770 ;
        RECT 33.430 115.810 33.570 117.450 ;
        RECT 33.890 116.410 34.030 117.450 ;
        RECT 35.670 117.110 35.930 117.430 ;
        RECT 36.130 117.110 36.390 117.430 ;
        RECT 33.830 116.090 34.090 116.410 ;
        RECT 32.450 115.410 32.710 115.730 ;
        RECT 33.430 115.670 34.030 115.810 ;
        RECT 35.730 115.730 35.870 117.110 ;
        RECT 36.190 116.410 36.330 117.110 ;
        RECT 36.130 116.090 36.390 116.410 ;
        RECT 32.510 112.670 32.650 115.410 ;
        RECT 33.890 115.390 34.030 115.670 ;
        RECT 34.750 115.410 35.010 115.730 ;
        RECT 35.670 115.410 35.930 115.730 ;
        RECT 33.830 115.070 34.090 115.390 ;
        RECT 34.810 113.350 34.950 115.410 ;
        RECT 36.650 113.690 36.790 117.880 ;
        RECT 37.570 116.070 37.710 120.850 ;
        RECT 37.510 115.750 37.770 116.070 ;
        RECT 36.590 113.600 36.850 113.690 ;
        RECT 36.590 113.460 37.250 113.600 ;
        RECT 36.590 113.370 36.850 113.460 ;
        RECT 33.370 113.030 33.630 113.350 ;
        RECT 34.750 113.030 35.010 113.350 ;
        RECT 33.430 112.670 33.570 113.030 ;
        RECT 32.450 112.350 32.710 112.670 ;
        RECT 33.370 112.350 33.630 112.670 ;
        RECT 30.610 111.670 30.870 111.990 ;
        RECT 30.670 110.970 30.810 111.670 ;
        RECT 30.610 110.650 30.870 110.970 ;
        RECT 32.510 109.610 32.650 112.350 ;
        RECT 32.450 109.290 32.710 109.610 ;
        RECT 30.610 108.950 30.870 109.270 ;
        RECT 29.230 105.210 29.490 105.530 ;
        RECT 29.230 104.530 29.490 104.850 ;
        RECT 29.290 99.410 29.430 104.530 ;
        RECT 30.670 104.510 30.810 108.950 ;
        RECT 31.530 106.230 31.790 106.550 ;
        RECT 30.610 104.190 30.870 104.510 ;
        RECT 30.150 103.510 30.410 103.830 ;
        RECT 29.690 101.130 29.950 101.450 ;
        RECT 28.310 99.090 28.570 99.410 ;
        RECT 29.230 99.090 29.490 99.410 ;
        RECT 28.370 96.690 28.510 99.090 ;
        RECT 27.850 96.370 28.110 96.690 ;
        RECT 28.310 96.370 28.570 96.690 ;
        RECT 27.910 91.250 28.050 96.370 ;
        RECT 29.290 96.350 29.430 99.090 ;
        RECT 29.750 96.690 29.890 101.130 ;
        RECT 30.210 99.410 30.350 103.510 ;
        RECT 30.670 101.790 30.810 104.190 ;
        RECT 31.070 102.490 31.330 102.810 ;
        RECT 30.610 101.470 30.870 101.790 ;
        RECT 31.130 99.410 31.270 102.490 ;
        RECT 31.590 101.110 31.730 106.230 ;
        RECT 31.990 104.530 32.250 104.850 ;
        RECT 31.530 100.790 31.790 101.110 ;
        RECT 30.150 99.090 30.410 99.410 ;
        RECT 30.610 99.090 30.870 99.410 ;
        RECT 31.070 99.090 31.330 99.410 ;
        RECT 29.690 96.370 29.950 96.690 ;
        RECT 29.230 96.090 29.490 96.350 ;
        RECT 29.230 96.030 29.890 96.090 ;
        RECT 29.290 95.950 29.890 96.030 ;
        RECT 27.850 90.930 28.110 91.250 ;
        RECT 29.230 90.590 29.490 90.910 ;
        RECT 28.770 90.250 29.030 90.570 ;
        RECT 28.310 89.910 28.570 90.230 ;
        RECT 25.550 88.210 25.810 88.530 ;
        RECT 25.610 86.490 25.750 88.210 ;
        RECT 25.550 86.170 25.810 86.490 ;
        RECT 28.370 85.470 28.510 89.910 ;
        RECT 28.830 85.810 28.970 90.250 ;
        RECT 29.290 89.210 29.430 90.590 ;
        RECT 29.230 88.890 29.490 89.210 ;
        RECT 29.290 86.490 29.430 88.890 ;
        RECT 29.230 86.170 29.490 86.490 ;
        RECT 28.770 85.490 29.030 85.810 ;
        RECT 28.310 85.150 28.570 85.470 ;
        RECT 26.010 81.750 26.270 82.070 ;
        RECT 26.070 80.030 26.210 81.750 ;
        RECT 25.550 79.710 25.810 80.030 ;
        RECT 26.010 79.710 26.270 80.030 ;
        RECT 25.610 78.330 25.750 79.710 ;
        RECT 29.750 78.330 29.890 95.950 ;
        RECT 30.670 94.650 30.810 99.090 ;
        RECT 32.050 99.070 32.190 104.530 ;
        RECT 32.510 103.830 32.650 109.290 ;
        RECT 33.430 105.530 33.570 112.350 ;
        RECT 33.830 111.670 34.090 111.990 ;
        RECT 33.370 105.210 33.630 105.530 ;
        RECT 32.450 103.510 32.710 103.830 ;
        RECT 32.510 101.790 32.650 103.510 ;
        RECT 33.430 102.810 33.570 105.210 ;
        RECT 33.370 102.490 33.630 102.810 ;
        RECT 33.430 101.790 33.570 102.490 ;
        RECT 32.450 101.470 32.710 101.790 ;
        RECT 32.910 101.470 33.170 101.790 ;
        RECT 33.370 101.470 33.630 101.790 ;
        RECT 32.450 100.790 32.710 101.110 ;
        RECT 32.510 99.750 32.650 100.790 ;
        RECT 32.450 99.430 32.710 99.750 ;
        RECT 31.990 98.750 32.250 99.070 ;
        RECT 32.970 97.370 33.110 101.470 ;
        RECT 32.910 97.050 33.170 97.370 ;
        RECT 31.990 96.710 32.250 97.030 ;
        RECT 32.050 96.350 32.190 96.710 ;
        RECT 31.990 96.030 32.250 96.350 ;
        RECT 32.050 95.670 32.190 96.030 ;
        RECT 33.890 96.010 34.030 111.670 ;
        RECT 34.810 110.970 34.950 113.030 ;
        RECT 36.130 111.670 36.390 111.990 ;
        RECT 34.750 110.650 35.010 110.970 ;
        RECT 34.750 109.970 35.010 110.290 ;
        RECT 34.810 102.470 34.950 109.970 ;
        RECT 35.210 106.230 35.470 106.550 ;
        RECT 35.270 103.830 35.410 106.230 ;
        RECT 35.670 104.870 35.930 105.190 ;
        RECT 35.210 103.510 35.470 103.830 ;
        RECT 34.750 102.150 35.010 102.470 ;
        RECT 34.750 100.790 35.010 101.110 ;
        RECT 34.290 98.750 34.550 99.070 ;
        RECT 34.350 97.030 34.490 98.750 ;
        RECT 34.810 98.730 34.950 100.790 ;
        RECT 35.730 100.090 35.870 104.870 ;
        RECT 36.190 101.790 36.330 111.670 ;
        RECT 36.590 107.250 36.850 107.570 ;
        RECT 36.130 101.470 36.390 101.790 ;
        RECT 35.670 99.770 35.930 100.090 ;
        RECT 35.210 99.090 35.470 99.410 ;
        RECT 34.750 98.410 35.010 98.730 ;
        RECT 34.290 96.710 34.550 97.030 ;
        RECT 34.290 96.260 34.550 96.350 ;
        RECT 34.810 96.260 34.950 98.410 ;
        RECT 34.290 96.120 34.950 96.260 ;
        RECT 34.290 96.030 34.550 96.120 ;
        RECT 33.830 95.690 34.090 96.010 ;
        RECT 31.990 95.350 32.250 95.670 ;
        RECT 30.610 94.330 30.870 94.650 ;
        RECT 32.050 91.930 32.190 95.350 ;
        RECT 31.990 91.610 32.250 91.930 ;
        RECT 30.610 90.590 30.870 90.910 ;
        RECT 30.670 87.510 30.810 90.590 ;
        RECT 32.450 90.250 32.710 90.570 ;
        RECT 32.510 88.530 32.650 90.250 ;
        RECT 34.350 88.870 34.490 96.030 ;
        RECT 35.270 96.010 35.410 99.090 ;
        RECT 36.190 98.810 36.330 101.470 ;
        RECT 36.650 100.090 36.790 107.250 ;
        RECT 37.110 101.790 37.250 113.460 ;
        RECT 37.510 106.570 37.770 106.890 ;
        RECT 37.570 102.810 37.710 106.570 ;
        RECT 38.030 105.190 38.170 128.760 ;
        RECT 38.430 128.670 38.690 128.760 ;
        RECT 38.710 124.735 40.250 125.105 ;
        RECT 40.270 123.290 40.530 123.550 ;
        RECT 40.790 123.290 40.930 130.710 ;
        RECT 40.270 123.230 40.930 123.290 ;
        RECT 40.330 123.150 40.930 123.230 ;
        RECT 40.330 120.150 40.470 123.150 ;
        RECT 40.730 120.850 40.990 121.170 ;
        RECT 40.270 119.830 40.530 120.150 ;
        RECT 38.710 119.295 40.250 119.665 ;
        RECT 39.810 117.110 40.070 117.430 ;
        RECT 39.870 116.070 40.010 117.110 ;
        RECT 40.790 116.410 40.930 120.850 ;
        RECT 40.730 116.090 40.990 116.410 ;
        RECT 39.810 115.750 40.070 116.070 ;
        RECT 38.710 113.855 40.250 114.225 ;
        RECT 40.270 113.370 40.530 113.690 ;
        RECT 40.330 110.290 40.470 113.370 ;
        RECT 40.730 111.670 40.990 111.990 ;
        RECT 40.270 109.970 40.530 110.290 ;
        RECT 40.790 109.610 40.930 111.670 ;
        RECT 41.250 110.290 41.390 131.730 ;
        RECT 42.170 130.010 42.310 132.070 ;
        RECT 50.450 132.050 50.590 134.110 ;
        RECT 50.910 132.050 51.050 135.130 ;
        RECT 52.290 133.750 52.430 136.150 ;
        RECT 52.690 133.770 52.950 134.090 ;
        RECT 52.230 133.430 52.490 133.750 ;
        RECT 50.390 131.730 50.650 132.050 ;
        RECT 50.850 131.730 51.110 132.050 ;
        RECT 48.550 131.050 48.810 131.370 ;
        RECT 43.490 130.710 43.750 131.030 ;
        RECT 47.630 130.710 47.890 131.030 ;
        RECT 42.110 129.690 42.370 130.010 ;
        RECT 41.650 125.610 41.910 125.930 ;
        RECT 41.710 123.550 41.850 125.610 ;
        RECT 42.170 124.570 42.310 129.690 ;
        RECT 43.550 129.670 43.690 130.710 ;
        RECT 42.570 129.350 42.830 129.670 ;
        RECT 43.490 129.350 43.750 129.670 ;
        RECT 42.630 127.290 42.770 129.350 ;
        RECT 47.690 128.650 47.830 130.710 ;
        RECT 45.330 128.330 45.590 128.650 ;
        RECT 47.630 128.330 47.890 128.650 ;
        RECT 42.570 126.970 42.830 127.290 ;
        RECT 42.630 126.610 42.770 126.970 ;
        RECT 42.570 126.290 42.830 126.610 ;
        RECT 42.110 124.250 42.370 124.570 ;
        RECT 41.650 123.230 41.910 123.550 ;
        RECT 42.110 117.790 42.370 118.110 ;
        RECT 42.170 115.130 42.310 117.790 ;
        RECT 41.710 114.990 42.310 115.130 ;
        RECT 41.190 109.970 41.450 110.290 ;
        RECT 40.730 109.290 40.990 109.610 ;
        RECT 38.710 108.415 40.250 108.785 ;
        RECT 38.430 106.910 38.690 107.230 ;
        RECT 38.490 105.530 38.630 106.910 ;
        RECT 40.730 106.230 40.990 106.550 ;
        RECT 38.430 105.210 38.690 105.530 ;
        RECT 37.970 104.870 38.230 105.190 ;
        RECT 38.710 102.975 40.250 103.345 ;
        RECT 37.510 102.490 37.770 102.810 ;
        RECT 37.050 101.470 37.310 101.790 ;
        RECT 39.350 101.470 39.610 101.790 ;
        RECT 36.590 99.770 36.850 100.090 ;
        RECT 37.110 99.410 37.250 101.470 ;
        RECT 37.050 99.090 37.310 99.410 ;
        RECT 36.190 98.670 36.790 98.810 ;
        RECT 35.210 95.690 35.470 96.010 ;
        RECT 35.670 95.690 35.930 96.010 ;
        RECT 35.210 93.990 35.470 94.310 ;
        RECT 34.750 93.310 35.010 93.630 ;
        RECT 34.810 89.210 34.950 93.310 ;
        RECT 35.270 90.570 35.410 93.990 ;
        RECT 35.730 93.290 35.870 95.690 ;
        RECT 36.650 94.310 36.790 98.670 ;
        RECT 36.590 93.990 36.850 94.310 ;
        RECT 37.110 94.220 37.250 99.090 ;
        RECT 39.410 99.070 39.550 101.470 ;
        RECT 40.790 99.410 40.930 106.230 ;
        RECT 41.710 102.470 41.850 114.990 ;
        RECT 42.110 114.390 42.370 114.710 ;
        RECT 42.170 113.010 42.310 114.390 ;
        RECT 42.110 112.690 42.370 113.010 ;
        RECT 42.630 112.670 42.770 126.290 ;
        RECT 43.950 125.950 44.210 126.270 ;
        RECT 44.010 122.870 44.150 125.950 ;
        RECT 45.390 124.570 45.530 128.330 ;
        RECT 45.330 124.250 45.590 124.570 ;
        RECT 43.950 122.550 44.210 122.870 ;
        RECT 44.010 121.850 44.150 122.550 ;
        RECT 43.950 121.530 44.210 121.850 ;
        RECT 43.950 120.510 44.210 120.830 ;
        RECT 44.010 118.110 44.150 120.510 ;
        RECT 45.330 118.470 45.590 118.790 ;
        RECT 43.950 117.790 44.210 118.110 ;
        RECT 44.010 114.710 44.150 117.790 ;
        RECT 44.870 117.450 45.130 117.770 ;
        RECT 44.930 115.730 45.070 117.450 ;
        RECT 45.390 117.430 45.530 118.470 ;
        RECT 48.610 118.110 48.750 131.050 ;
        RECT 50.910 128.650 51.050 131.730 ;
        RECT 52.290 129.330 52.430 133.430 ;
        RECT 52.750 130.010 52.890 133.770 ;
        RECT 53.210 132.050 53.350 136.830 ;
        RECT 54.130 132.730 54.270 137.170 ;
        RECT 54.070 132.410 54.330 132.730 ;
        RECT 53.150 131.730 53.410 132.050 ;
        RECT 53.610 131.730 53.870 132.050 ;
        RECT 52.690 129.690 52.950 130.010 ;
        RECT 51.310 129.010 51.570 129.330 ;
        RECT 52.230 129.010 52.490 129.330 ;
        RECT 50.850 128.330 51.110 128.650 ;
        RECT 51.370 126.950 51.510 129.010 ;
        RECT 53.670 128.990 53.810 131.730 ;
        RECT 54.070 129.010 54.330 129.330 ;
        RECT 53.610 128.670 53.870 128.990 ;
        RECT 51.770 128.330 52.030 128.650 ;
        RECT 51.830 127.290 51.970 128.330 ;
        RECT 53.670 128.310 53.810 128.670 ;
        RECT 53.610 127.990 53.870 128.310 ;
        RECT 51.770 126.970 52.030 127.290 ;
        RECT 51.310 126.630 51.570 126.950 ;
        RECT 49.470 125.270 49.730 125.590 ;
        RECT 49.530 123.550 49.670 125.270 ;
        RECT 49.990 123.890 51.050 123.970 ;
        RECT 49.990 123.830 51.110 123.890 ;
        RECT 49.470 123.230 49.730 123.550 ;
        RECT 49.990 121.510 50.130 123.830 ;
        RECT 50.850 123.570 51.110 123.830 ;
        RECT 50.390 123.230 50.650 123.550 ;
        RECT 50.450 121.850 50.590 123.230 ;
        RECT 51.370 123.210 51.510 126.630 ;
        RECT 54.130 126.610 54.270 129.010 ;
        RECT 54.590 127.290 54.730 137.170 ;
        RECT 55.050 130.010 55.190 137.170 ;
        RECT 57.750 136.150 58.010 136.470 ;
        RECT 57.290 133.430 57.550 133.750 ;
        RECT 55.500 132.895 57.040 133.265 ;
        RECT 57.350 132.730 57.490 133.430 ;
        RECT 57.810 132.730 57.950 136.150 ;
        RECT 61.030 134.770 61.170 137.170 ;
        RECT 61.490 136.470 61.630 139.210 ;
        RECT 61.950 138.080 62.090 139.980 ;
        RECT 62.350 138.080 62.610 138.170 ;
        RECT 61.950 137.940 62.610 138.080 ;
        RECT 62.350 137.850 62.610 137.940 ;
        RECT 61.890 137.400 62.150 137.490 ;
        RECT 62.810 137.400 63.070 137.490 ;
        RECT 61.890 137.260 63.070 137.400 ;
        RECT 61.890 137.170 62.150 137.260 ;
        RECT 62.810 137.170 63.070 137.260 ;
        RECT 61.430 136.150 61.690 136.470 ;
        RECT 64.250 135.450 64.390 144.650 ;
        RECT 64.710 142.930 64.850 144.990 ;
        RECT 65.630 143.610 65.770 149.750 ;
        RECT 66.090 149.050 66.230 151.450 ;
        RECT 66.030 148.730 66.290 149.050 ;
        RECT 66.550 147.770 66.690 171.850 ;
        RECT 68.390 170.470 68.530 186.810 ;
        RECT 69.250 185.790 69.510 186.110 ;
        RECT 69.310 184.410 69.450 185.790 ;
        RECT 69.250 184.090 69.510 184.410 ;
        RECT 69.310 181.690 69.450 184.090 ;
        RECT 69.250 181.370 69.510 181.690 ;
        RECT 69.770 181.350 69.910 191.570 ;
        RECT 70.170 190.890 70.430 191.210 ;
        RECT 70.230 189.850 70.370 190.890 ;
        RECT 72.290 190.015 73.830 190.385 ;
        RECT 70.170 189.530 70.430 189.850 ;
        RECT 70.630 186.130 70.890 186.450 ;
        RECT 70.690 182.710 70.830 186.130 ;
        RECT 72.290 184.575 73.830 184.945 ;
        RECT 74.830 183.390 74.970 191.570 ;
        RECT 75.290 189.850 75.430 191.570 ;
        RECT 75.230 189.530 75.490 189.850 ;
        RECT 75.230 188.400 75.490 188.490 ;
        RECT 75.750 188.400 75.890 200.410 ;
        RECT 79.890 199.370 80.030 201.915 ;
        RECT 82.190 200.390 82.330 202.110 ;
        RECT 82.130 200.070 82.390 200.390 ;
        RECT 77.990 199.050 78.250 199.370 ;
        RECT 79.830 199.050 80.090 199.370 ;
        RECT 80.290 199.050 80.550 199.370 ;
        RECT 77.530 193.270 77.790 193.590 ;
        RECT 77.590 188.830 77.730 193.270 ;
        RECT 78.050 188.830 78.190 199.050 ;
        RECT 78.450 198.710 78.710 199.030 ;
        RECT 78.510 197.670 78.650 198.710 ;
        RECT 78.450 197.350 78.710 197.670 ;
        RECT 78.450 193.950 78.710 194.270 ;
        RECT 77.070 188.510 77.330 188.830 ;
        RECT 77.530 188.510 77.790 188.830 ;
        RECT 77.990 188.510 78.250 188.830 ;
        RECT 75.230 188.260 75.890 188.400 ;
        RECT 75.230 188.170 75.490 188.260 ;
        RECT 76.610 188.170 76.870 188.490 ;
        RECT 74.770 183.070 75.030 183.390 ;
        RECT 70.630 182.390 70.890 182.710 ;
        RECT 69.710 181.030 69.970 181.350 ;
        RECT 69.250 176.950 69.510 177.270 ;
        RECT 69.310 173.530 69.450 176.950 ;
        RECT 69.250 173.210 69.510 173.530 ;
        RECT 69.770 170.810 69.910 181.030 ;
        RECT 70.630 179.670 70.890 179.990 ;
        RECT 70.690 177.950 70.830 179.670 ;
        RECT 72.290 179.135 73.830 179.505 ;
        RECT 74.830 178.970 74.970 183.070 ;
        RECT 75.290 179.990 75.430 188.170 ;
        RECT 76.670 186.790 76.810 188.170 ;
        RECT 75.690 186.470 75.950 186.790 ;
        RECT 76.610 186.470 76.870 186.790 ;
        RECT 75.230 179.670 75.490 179.990 ;
        RECT 74.770 178.650 75.030 178.970 ;
        RECT 70.170 177.630 70.430 177.950 ;
        RECT 70.630 177.630 70.890 177.950 ;
        RECT 72.010 177.630 72.270 177.950 ;
        RECT 70.230 175.570 70.370 177.630 ;
        RECT 71.090 177.290 71.350 177.610 ;
        RECT 71.550 177.290 71.810 177.610 ;
        RECT 71.150 175.910 71.290 177.290 ;
        RECT 71.610 176.250 71.750 177.290 ;
        RECT 72.070 176.250 72.210 177.630 ;
        RECT 71.550 175.930 71.810 176.250 ;
        RECT 72.010 175.930 72.270 176.250 ;
        RECT 71.090 175.590 71.350 175.910 ;
        RECT 70.170 175.250 70.430 175.570 ;
        RECT 69.710 170.490 69.970 170.810 ;
        RECT 68.330 170.150 68.590 170.470 ;
        RECT 70.230 170.130 70.370 175.250 ;
        RECT 71.150 173.530 71.290 175.590 ;
        RECT 74.830 175.570 74.970 178.650 ;
        RECT 75.230 177.630 75.490 177.950 ;
        RECT 74.770 175.250 75.030 175.570 ;
        RECT 72.290 173.695 73.830 174.065 ;
        RECT 71.090 173.210 71.350 173.530 ;
        RECT 71.150 170.130 71.290 173.210 ;
        RECT 75.290 172.510 75.430 177.630 ;
        RECT 75.230 172.190 75.490 172.510 ;
        RECT 72.010 170.490 72.270 170.810 ;
        RECT 72.070 170.130 72.210 170.490 ;
        RECT 75.290 170.130 75.430 172.190 ;
        RECT 75.750 170.470 75.890 186.470 ;
        RECT 77.130 186.450 77.270 188.510 ;
        RECT 77.070 186.130 77.330 186.450 ;
        RECT 76.150 185.110 76.410 185.430 ;
        RECT 76.210 183.050 76.350 185.110 ;
        RECT 76.150 182.730 76.410 183.050 ;
        RECT 76.610 174.230 76.870 174.550 ;
        RECT 76.670 173.530 76.810 174.230 ;
        RECT 76.610 173.210 76.870 173.530 ;
        RECT 75.690 170.150 75.950 170.470 ;
        RECT 77.530 170.150 77.790 170.470 ;
        RECT 69.250 169.810 69.510 170.130 ;
        RECT 69.710 169.810 69.970 170.130 ;
        RECT 70.170 169.810 70.430 170.130 ;
        RECT 70.630 169.810 70.890 170.130 ;
        RECT 71.090 169.810 71.350 170.130 ;
        RECT 72.010 169.810 72.270 170.130 ;
        RECT 75.230 169.810 75.490 170.130 ;
        RECT 69.310 167.410 69.450 169.810 ;
        RECT 69.250 167.090 69.510 167.410 ;
        RECT 69.770 166.730 69.910 169.810 ;
        RECT 70.170 166.750 70.430 167.070 ;
        RECT 69.710 166.410 69.970 166.730 ;
        RECT 68.330 166.070 68.590 166.390 ;
        RECT 67.870 161.650 68.130 161.970 ;
        RECT 66.950 157.910 67.210 158.230 ;
        RECT 67.010 156.530 67.150 157.910 ;
        RECT 66.950 156.210 67.210 156.530 ;
        RECT 66.950 155.530 67.210 155.850 ;
        RECT 67.010 151.090 67.150 155.530 ;
        RECT 67.930 153.720 68.070 161.650 ;
        RECT 68.390 161.630 68.530 166.070 ;
        RECT 70.230 164.010 70.370 166.750 ;
        RECT 70.690 165.370 70.830 169.810 ;
        RECT 70.630 165.050 70.890 165.370 ;
        RECT 70.170 163.690 70.430 164.010 ;
        RECT 70.630 163.350 70.890 163.670 ;
        RECT 70.690 162.310 70.830 163.350 ;
        RECT 70.630 161.990 70.890 162.310 ;
        RECT 71.150 161.970 71.290 169.810 ;
        RECT 72.070 169.530 72.210 169.810 ;
        RECT 71.610 169.390 72.210 169.530 ;
        RECT 71.610 166.390 71.750 169.390 ;
        RECT 72.290 168.255 73.830 168.625 ;
        RECT 74.310 166.750 74.570 167.070 ;
        RECT 71.550 166.070 71.810 166.390 ;
        RECT 72.290 162.815 73.830 163.185 ;
        RECT 71.090 161.650 71.350 161.970 ;
        RECT 72.010 161.650 72.270 161.970 ;
        RECT 68.330 161.310 68.590 161.630 ;
        RECT 69.250 160.970 69.510 161.290 ;
        RECT 68.790 158.590 69.050 158.910 ;
        RECT 68.850 156.530 68.990 158.590 ;
        RECT 68.790 156.210 69.050 156.530 ;
        RECT 68.330 153.720 68.590 153.810 ;
        RECT 67.930 153.580 68.590 153.720 ;
        RECT 67.930 153.130 68.070 153.580 ;
        RECT 68.330 153.490 68.590 153.580 ;
        RECT 67.870 152.810 68.130 153.130 ;
        RECT 66.950 150.770 67.210 151.090 ;
        RECT 69.310 150.410 69.450 160.970 ;
        RECT 72.070 159.930 72.210 161.650 ;
        RECT 72.010 159.610 72.270 159.930 ;
        RECT 69.710 158.930 69.970 159.250 ;
        RECT 69.770 154.490 69.910 158.930 ;
        RECT 72.290 157.375 73.830 157.745 ;
        RECT 71.090 156.210 71.350 156.530 ;
        RECT 70.170 155.190 70.430 155.510 ;
        RECT 69.710 154.170 69.970 154.490 ;
        RECT 70.230 153.810 70.370 155.190 ;
        RECT 70.170 153.490 70.430 153.810 ;
        RECT 69.250 150.090 69.510 150.410 ;
        RECT 66.950 149.750 67.210 150.070 ;
        RECT 67.010 149.050 67.150 149.750 ;
        RECT 66.950 148.730 67.210 149.050 ;
        RECT 66.550 147.630 67.150 147.770 ;
        RECT 66.490 147.030 66.750 147.350 ;
        RECT 66.030 144.310 66.290 144.630 ;
        RECT 65.570 143.290 65.830 143.610 ;
        RECT 66.090 142.930 66.230 144.310 ;
        RECT 66.550 142.930 66.690 147.030 ;
        RECT 64.650 142.610 64.910 142.930 ;
        RECT 65.570 142.610 65.830 142.930 ;
        RECT 66.030 142.610 66.290 142.930 ;
        RECT 66.490 142.610 66.750 142.930 ;
        RECT 65.630 142.330 65.770 142.610 ;
        RECT 65.630 142.250 66.230 142.330 ;
        RECT 65.630 142.190 66.290 142.250 ;
        RECT 66.030 141.930 66.290 142.190 ;
        RECT 65.570 141.590 65.830 141.910 ;
        RECT 65.630 140.890 65.770 141.590 ;
        RECT 65.110 140.570 65.370 140.890 ;
        RECT 65.570 140.570 65.830 140.890 ;
        RECT 65.170 140.120 65.310 140.570 ;
        RECT 64.710 139.980 65.310 140.120 ;
        RECT 64.190 135.130 64.450 135.450 ;
        RECT 60.970 134.450 61.230 134.770 ;
        RECT 58.210 133.770 58.470 134.090 ;
        RECT 57.290 132.410 57.550 132.730 ;
        RECT 57.750 132.410 58.010 132.730 ;
        RECT 57.290 131.390 57.550 131.710 ;
        RECT 54.990 129.690 55.250 130.010 ;
        RECT 55.500 127.455 57.040 127.825 ;
        RECT 57.350 127.290 57.490 131.390 ;
        RECT 54.530 126.970 54.790 127.290 ;
        RECT 57.290 126.970 57.550 127.290 ;
        RECT 54.070 126.290 54.330 126.610 ;
        RECT 51.770 125.610 52.030 125.930 ;
        RECT 51.830 123.210 51.970 125.610 ;
        RECT 54.130 124.570 54.270 126.290 ;
        RECT 54.990 125.270 55.250 125.590 ;
        RECT 55.050 124.570 55.190 125.270 ;
        RECT 57.350 124.570 57.490 126.970 ;
        RECT 54.070 124.250 54.330 124.570 ;
        RECT 54.990 124.250 55.250 124.570 ;
        RECT 57.290 124.250 57.550 124.570 ;
        RECT 58.270 123.890 58.410 133.770 ;
        RECT 62.350 132.410 62.610 132.730 ;
        RECT 60.050 132.070 60.310 132.390 ;
        RECT 60.110 127.290 60.250 132.070 ;
        RECT 61.890 131.390 62.150 131.710 ;
        RECT 61.950 130.010 62.090 131.390 ;
        RECT 61.890 129.690 62.150 130.010 ;
        RECT 61.430 128.220 61.690 128.310 ;
        RECT 61.030 128.080 61.690 128.220 ;
        RECT 60.050 126.970 60.310 127.290 ;
        RECT 60.510 126.970 60.770 127.290 ;
        RECT 58.210 123.570 58.470 123.890 ;
        RECT 51.310 122.890 51.570 123.210 ;
        RECT 51.770 122.890 52.030 123.210 ;
        RECT 55.500 122.015 57.040 122.385 ;
        RECT 50.390 121.530 50.650 121.850 ;
        RECT 49.930 121.190 50.190 121.510 ;
        RECT 51.310 121.190 51.570 121.510 ;
        RECT 49.470 120.170 49.730 120.490 ;
        RECT 48.550 117.790 48.810 118.110 ;
        RECT 49.530 117.430 49.670 120.170 ;
        RECT 51.370 119.130 51.510 121.190 ;
        RECT 60.570 121.170 60.710 126.970 ;
        RECT 61.030 123.210 61.170 128.080 ;
        RECT 61.430 127.990 61.690 128.080 ;
        RECT 60.970 122.890 61.230 123.210 ;
        RECT 60.510 120.850 60.770 121.170 ;
        RECT 58.210 120.510 58.470 120.830 ;
        RECT 54.530 119.830 54.790 120.150 ;
        RECT 56.830 119.830 57.090 120.150 ;
        RECT 51.310 118.810 51.570 119.130 ;
        RECT 52.230 117.790 52.490 118.110 ;
        RECT 45.330 117.110 45.590 117.430 ;
        RECT 49.470 117.110 49.730 117.430 ;
        RECT 45.390 115.730 45.530 117.110 ;
        RECT 44.870 115.410 45.130 115.730 ;
        RECT 45.330 115.410 45.590 115.730 ;
        RECT 43.950 114.390 44.210 114.710 ;
        RECT 42.570 112.350 42.830 112.670 ;
        RECT 43.030 112.350 43.290 112.670 ;
        RECT 43.090 110.970 43.230 112.350 ;
        RECT 43.030 110.650 43.290 110.970 ;
        RECT 44.010 110.630 44.150 114.390 ;
        RECT 44.870 113.260 45.130 113.350 ;
        RECT 45.390 113.260 45.530 115.410 ;
        RECT 52.290 114.710 52.430 117.790 ;
        RECT 52.690 115.070 52.950 115.390 ;
        RECT 47.170 114.390 47.430 114.710 ;
        RECT 52.230 114.390 52.490 114.710 ;
        RECT 44.870 113.120 45.530 113.260 ;
        RECT 44.870 113.030 45.130 113.120 ;
        RECT 44.410 112.690 44.670 113.010 ;
        RECT 43.950 110.310 44.210 110.630 ;
        RECT 43.950 106.230 44.210 106.550 ;
        RECT 41.650 102.150 41.910 102.470 ;
        RECT 44.010 101.790 44.150 106.230 ;
        RECT 44.470 105.530 44.610 112.690 ;
        RECT 44.930 110.290 45.070 113.030 ;
        RECT 47.230 110.290 47.370 114.390 ;
        RECT 52.750 112.410 52.890 115.070 ;
        RECT 54.070 114.390 54.330 114.710 ;
        RECT 52.750 112.270 53.350 112.410 ;
        RECT 52.690 111.670 52.950 111.990 ;
        RECT 52.750 110.290 52.890 111.670 ;
        RECT 53.210 111.050 53.350 112.270 ;
        RECT 53.210 110.910 53.810 111.050 ;
        RECT 53.670 110.290 53.810 110.910 ;
        RECT 54.130 110.290 54.270 114.390 ;
        RECT 54.590 110.970 54.730 119.830 ;
        RECT 56.890 119.130 57.030 119.830 ;
        RECT 56.830 118.810 57.090 119.130 ;
        RECT 54.990 117.450 55.250 117.770 ;
        RECT 57.290 117.450 57.550 117.770 ;
        RECT 55.050 115.730 55.190 117.450 ;
        RECT 55.500 116.575 57.040 116.945 ;
        RECT 54.990 115.410 55.250 115.730 ;
        RECT 57.350 113.690 57.490 117.450 ;
        RECT 58.270 115.730 58.410 120.510 ;
        RECT 58.670 120.170 58.930 120.490 ;
        RECT 58.730 118.450 58.870 120.170 ;
        RECT 60.570 119.130 60.710 120.850 ;
        RECT 60.510 118.810 60.770 119.130 ;
        RECT 58.670 118.130 58.930 118.450 ;
        RECT 58.730 116.410 58.870 118.130 ;
        RECT 58.670 116.090 58.930 116.410 ;
        RECT 61.030 115.730 61.170 122.890 ;
        RECT 61.950 120.830 62.090 129.690 ;
        RECT 62.410 125.590 62.550 132.410 ;
        RECT 63.270 130.710 63.530 131.030 ;
        RECT 63.330 128.990 63.470 130.710 ;
        RECT 64.250 128.990 64.390 135.130 ;
        RECT 63.270 128.670 63.530 128.990 ;
        RECT 64.190 128.670 64.450 128.990 ;
        RECT 63.270 126.290 63.530 126.610 ;
        RECT 62.350 125.270 62.610 125.590 ;
        RECT 63.330 124.570 63.470 126.290 ;
        RECT 63.270 124.250 63.530 124.570 ;
        RECT 64.250 123.550 64.390 128.670 ;
        RECT 64.190 123.230 64.450 123.550 ;
        RECT 61.890 120.510 62.150 120.830 ;
        RECT 62.810 119.830 63.070 120.150 ;
        RECT 62.870 119.130 63.010 119.830 ;
        RECT 62.810 118.810 63.070 119.130 ;
        RECT 61.430 117.110 61.690 117.430 ;
        RECT 61.490 115.730 61.630 117.110 ;
        RECT 64.710 116.370 64.850 139.980 ;
        RECT 65.110 139.210 65.370 139.530 ;
        RECT 65.170 138.170 65.310 139.210 ;
        RECT 65.110 137.850 65.370 138.170 ;
        RECT 65.110 136.830 65.370 137.150 ;
        RECT 65.170 134.770 65.310 136.830 ;
        RECT 67.010 135.450 67.150 147.630 ;
        RECT 67.870 145.670 68.130 145.990 ;
        RECT 67.410 144.310 67.670 144.630 ;
        RECT 67.470 143.610 67.610 144.310 ;
        RECT 67.410 143.290 67.670 143.610 ;
        RECT 67.930 142.840 68.070 145.670 ;
        RECT 68.330 145.330 68.590 145.650 ;
        RECT 68.390 143.610 68.530 145.330 ;
        RECT 68.330 143.290 68.590 143.610 ;
        RECT 68.790 142.840 69.050 142.930 ;
        RECT 67.930 142.700 69.050 142.840 ;
        RECT 68.790 142.610 69.050 142.700 ;
        RECT 68.330 140.570 68.590 140.890 ;
        RECT 66.950 135.130 67.210 135.450 ;
        RECT 65.110 134.450 65.370 134.770 ;
        RECT 65.170 132.730 65.310 134.450 ;
        RECT 65.110 132.410 65.370 132.730 ;
        RECT 68.390 128.990 68.530 140.570 ;
        RECT 68.330 128.670 68.590 128.990 ;
        RECT 65.570 128.330 65.830 128.650 ;
        RECT 66.950 128.330 67.210 128.650 ;
        RECT 65.110 126.630 65.370 126.950 ;
        RECT 65.170 125.500 65.310 126.630 ;
        RECT 65.630 126.270 65.770 128.330 ;
        RECT 67.010 127.290 67.150 128.330 ;
        RECT 66.950 126.970 67.210 127.290 ;
        RECT 67.410 126.970 67.670 127.290 ;
        RECT 65.570 125.950 65.830 126.270 ;
        RECT 67.470 125.500 67.610 126.970 ;
        RECT 67.870 126.290 68.130 126.610 ;
        RECT 67.930 125.930 68.070 126.290 ;
        RECT 67.870 125.610 68.130 125.930 ;
        RECT 65.170 125.360 67.610 125.500 ;
        RECT 66.030 117.110 66.290 117.430 ;
        RECT 63.330 116.230 64.850 116.370 ;
        RECT 66.090 116.370 66.230 117.110 ;
        RECT 66.090 116.230 66.690 116.370 ;
        RECT 63.330 115.730 63.470 116.230 ;
        RECT 64.650 115.750 64.910 116.070 ;
        RECT 58.210 115.410 58.470 115.730 ;
        RECT 60.970 115.410 61.230 115.730 ;
        RECT 61.430 115.410 61.690 115.730 ;
        RECT 62.350 115.410 62.610 115.730 ;
        RECT 63.270 115.410 63.530 115.730 ;
        RECT 57.750 115.070 58.010 115.390 ;
        RECT 57.290 113.370 57.550 113.690 ;
        RECT 55.500 111.135 57.040 111.505 ;
        RECT 54.530 110.650 54.790 110.970 ;
        RECT 57.350 110.630 57.490 113.370 ;
        RECT 57.810 112.670 57.950 115.070 ;
        RECT 62.410 113.690 62.550 115.410 ;
        RECT 62.350 113.370 62.610 113.690 ;
        RECT 57.750 112.350 58.010 112.670 ;
        RECT 57.290 110.310 57.550 110.630 ;
        RECT 44.870 109.970 45.130 110.290 ;
        RECT 47.170 109.970 47.430 110.290 ;
        RECT 52.690 109.970 52.950 110.290 ;
        RECT 53.150 109.970 53.410 110.290 ;
        RECT 53.610 109.970 53.870 110.290 ;
        RECT 54.070 109.970 54.330 110.290 ;
        RECT 54.530 109.970 54.790 110.290 ;
        RECT 44.930 108.250 45.070 109.970 ;
        RECT 47.230 109.690 47.370 109.970 ;
        RECT 47.230 109.550 47.830 109.690 ;
        RECT 44.870 107.930 45.130 108.250 ;
        RECT 44.930 107.230 45.070 107.930 ;
        RECT 47.690 107.910 47.830 109.550 ;
        RECT 50.390 108.950 50.650 109.270 ;
        RECT 47.630 107.590 47.890 107.910 ;
        RECT 49.010 107.590 49.270 107.910 ;
        RECT 47.690 107.230 47.830 107.590 ;
        RECT 44.870 106.910 45.130 107.230 ;
        RECT 45.790 106.910 46.050 107.230 ;
        RECT 47.630 106.910 47.890 107.230 ;
        RECT 45.850 106.550 45.990 106.910 ;
        RECT 45.790 106.230 46.050 106.550 ;
        RECT 44.410 105.210 44.670 105.530 ;
        RECT 44.470 102.810 44.610 105.210 ;
        RECT 49.070 105.190 49.210 107.590 ;
        RECT 49.010 104.870 49.270 105.190 ;
        RECT 49.070 102.810 49.210 104.870 ;
        RECT 50.450 104.850 50.590 108.950 ;
        RECT 51.310 107.590 51.570 107.910 ;
        RECT 51.370 106.550 51.510 107.590 ;
        RECT 52.690 106.910 52.950 107.230 ;
        RECT 51.310 106.230 51.570 106.550 ;
        RECT 51.770 106.230 52.030 106.550 ;
        RECT 52.230 106.230 52.490 106.550 ;
        RECT 50.390 104.530 50.650 104.850 ;
        RECT 49.930 104.190 50.190 104.510 ;
        RECT 44.410 102.490 44.670 102.810 ;
        RECT 49.010 102.490 49.270 102.810 ;
        RECT 43.950 101.470 44.210 101.790 ;
        RECT 49.990 101.450 50.130 104.190 ;
        RECT 51.830 101.450 51.970 106.230 ;
        RECT 52.290 104.850 52.430 106.230 ;
        RECT 52.230 104.530 52.490 104.850 ;
        RECT 52.230 103.740 52.490 103.830 ;
        RECT 52.750 103.740 52.890 106.910 ;
        RECT 53.210 105.530 53.350 109.970 ;
        RECT 53.610 107.930 53.870 108.250 ;
        RECT 54.070 107.930 54.330 108.250 ;
        RECT 53.670 107.230 53.810 107.930 ;
        RECT 54.130 107.230 54.270 107.930 ;
        RECT 53.610 106.910 53.870 107.230 ;
        RECT 54.070 106.910 54.330 107.230 ;
        RECT 53.150 105.210 53.410 105.530 ;
        RECT 54.590 104.850 54.730 109.970 ;
        RECT 57.350 107.230 57.490 110.310 ;
        RECT 57.290 106.910 57.550 107.230 ;
        RECT 55.500 105.695 57.040 106.065 ;
        RECT 57.810 105.530 57.950 112.350 ;
        RECT 58.670 112.010 58.930 112.330 ;
        RECT 58.730 110.970 58.870 112.010 ;
        RECT 61.890 111.670 62.150 111.990 ;
        RECT 61.950 110.970 62.090 111.670 ;
        RECT 58.670 110.650 58.930 110.970 ;
        RECT 61.890 110.650 62.150 110.970 ;
        RECT 62.410 109.270 62.550 113.370 ;
        RECT 63.330 110.290 63.470 115.410 ;
        RECT 63.730 112.350 63.990 112.670 ;
        RECT 64.190 112.350 64.450 112.670 ;
        RECT 63.790 110.970 63.930 112.350 ;
        RECT 64.250 110.970 64.390 112.350 ;
        RECT 63.730 110.650 63.990 110.970 ;
        RECT 64.190 110.650 64.450 110.970 ;
        RECT 64.710 110.290 64.850 115.750 ;
        RECT 66.550 115.730 66.690 116.230 ;
        RECT 68.390 116.070 68.530 128.670 ;
        RECT 68.790 126.520 69.050 126.610 ;
        RECT 69.310 126.520 69.450 150.090 ;
        RECT 69.710 149.750 69.970 150.070 ;
        RECT 69.770 146.330 69.910 149.750 ;
        RECT 71.150 148.370 71.290 156.210 ;
        RECT 72.290 151.935 73.830 152.305 ;
        RECT 72.010 150.430 72.270 150.750 ;
        RECT 72.470 150.430 72.730 150.750 ;
        RECT 71.550 149.750 71.810 150.070 ;
        RECT 71.090 148.280 71.350 148.370 ;
        RECT 70.690 148.140 71.350 148.280 ;
        RECT 69.710 146.010 69.970 146.330 ;
        RECT 70.690 145.730 70.830 148.140 ;
        RECT 71.090 148.050 71.350 148.140 ;
        RECT 71.090 147.370 71.350 147.690 ;
        RECT 69.770 145.590 70.830 145.730 ;
        RECT 69.770 139.870 69.910 145.590 ;
        RECT 70.170 144.990 70.430 145.310 ;
        RECT 70.230 139.870 70.370 144.990 ;
        RECT 70.630 142.270 70.890 142.590 ;
        RECT 69.710 139.550 69.970 139.870 ;
        RECT 70.170 139.550 70.430 139.870 ;
        RECT 70.230 137.490 70.370 139.550 ;
        RECT 70.690 139.190 70.830 142.270 ;
        RECT 71.150 141.910 71.290 147.370 ;
        RECT 71.610 142.930 71.750 149.750 ;
        RECT 72.070 147.690 72.210 150.430 ;
        RECT 72.010 147.370 72.270 147.690 ;
        RECT 72.530 147.350 72.670 150.430 ;
        RECT 72.470 147.030 72.730 147.350 ;
        RECT 72.290 146.495 73.830 146.865 ;
        RECT 74.370 142.930 74.510 166.750 ;
        RECT 75.290 166.390 75.430 169.810 ;
        RECT 75.690 168.790 75.950 169.110 ;
        RECT 76.150 168.790 76.410 169.110 ;
        RECT 75.230 166.070 75.490 166.390 ;
        RECT 75.290 164.690 75.430 166.070 ;
        RECT 75.230 164.370 75.490 164.690 ;
        RECT 74.760 163.835 75.040 164.205 ;
        RECT 74.830 161.290 74.970 163.835 ;
        RECT 75.750 161.630 75.890 168.790 ;
        RECT 76.210 165.030 76.350 168.790 ;
        RECT 76.150 164.710 76.410 165.030 ;
        RECT 77.070 164.370 77.330 164.690 ;
        RECT 77.130 161.630 77.270 164.370 ;
        RECT 75.690 161.310 75.950 161.630 ;
        RECT 77.070 161.310 77.330 161.630 ;
        RECT 74.770 160.970 75.030 161.290 ;
        RECT 74.770 158.930 75.030 159.250 ;
        RECT 74.830 154.490 74.970 158.930 ;
        RECT 77.590 157.290 77.730 170.150 ;
        RECT 78.050 167.070 78.190 188.510 ;
        RECT 78.510 186.450 78.650 193.950 ;
        RECT 80.350 187.130 80.490 199.050 ;
        RECT 83.050 198.710 83.310 199.030 ;
        RECT 83.110 194.270 83.250 198.710 ;
        RECT 83.510 197.010 83.770 197.330 ;
        RECT 83.570 195.290 83.710 197.010 ;
        RECT 84.030 196.990 84.170 205.170 ;
        RECT 84.950 203.450 85.090 205.510 ;
        RECT 85.350 204.830 85.610 205.150 ;
        RECT 84.890 203.130 85.150 203.450 ;
        RECT 85.410 202.770 85.550 204.830 ;
        RECT 85.350 202.450 85.610 202.770 ;
        RECT 84.890 201.430 85.150 201.750 ;
        RECT 85.350 201.660 85.610 201.750 ;
        RECT 85.350 201.520 86.010 201.660 ;
        RECT 85.350 201.430 85.610 201.520 ;
        RECT 83.970 196.670 84.230 196.990 ;
        RECT 83.510 194.970 83.770 195.290 ;
        RECT 82.590 193.950 82.850 194.270 ;
        RECT 83.050 193.950 83.310 194.270 ;
        RECT 82.650 191.210 82.790 193.950 ;
        RECT 82.590 190.890 82.850 191.210 ;
        RECT 80.290 186.810 80.550 187.130 ;
        RECT 81.210 186.470 81.470 186.790 ;
        RECT 78.450 186.130 78.710 186.450 ;
        RECT 80.290 186.130 80.550 186.450 ;
        RECT 79.370 182.730 79.630 183.050 ;
        RECT 79.430 181.690 79.570 182.730 ;
        RECT 79.370 181.370 79.630 181.690 ;
        RECT 80.350 179.990 80.490 186.130 ;
        RECT 81.270 181.010 81.410 186.470 ;
        RECT 83.110 186.450 83.250 193.950 ;
        RECT 84.030 191.890 84.170 196.670 ;
        RECT 83.970 191.570 84.230 191.890 ;
        RECT 84.430 191.570 84.690 191.890 ;
        RECT 84.030 189.850 84.170 191.570 ;
        RECT 83.970 189.530 84.230 189.850 ;
        RECT 83.970 188.510 84.230 188.830 ;
        RECT 83.050 186.130 83.310 186.450 ;
        RECT 84.030 186.360 84.170 188.510 ;
        RECT 84.490 187.130 84.630 191.570 ;
        RECT 84.430 186.810 84.690 187.130 ;
        RECT 84.430 186.360 84.690 186.450 ;
        RECT 84.030 186.220 84.690 186.360 ;
        RECT 82.590 185.790 82.850 186.110 ;
        RECT 82.650 184.410 82.790 185.790 ;
        RECT 82.590 184.090 82.850 184.410 ;
        RECT 81.210 180.690 81.470 181.010 ;
        RECT 80.290 179.670 80.550 179.990 ;
        RECT 78.910 176.950 79.170 177.270 ;
        RECT 78.970 176.250 79.110 176.950 ;
        RECT 78.910 175.930 79.170 176.250 ;
        RECT 79.370 171.850 79.630 172.170 ;
        RECT 79.430 169.110 79.570 171.850 ;
        RECT 80.350 170.130 80.490 179.670 ;
        RECT 80.750 175.250 81.010 175.570 ;
        RECT 80.810 173.530 80.950 175.250 ;
        RECT 80.750 173.210 81.010 173.530 ;
        RECT 81.270 170.130 81.410 180.690 ;
        RECT 84.030 174.890 84.170 186.220 ;
        RECT 84.430 186.130 84.690 186.220 ;
        RECT 84.430 177.290 84.690 177.610 ;
        RECT 83.970 174.570 84.230 174.890 ;
        RECT 84.490 173.530 84.630 177.290 ;
        RECT 84.430 173.210 84.690 173.530 ;
        RECT 79.830 169.810 80.090 170.130 ;
        RECT 80.290 169.810 80.550 170.130 ;
        RECT 81.210 169.810 81.470 170.130 ;
        RECT 79.370 168.790 79.630 169.110 ;
        RECT 79.890 168.090 80.030 169.810 ;
        RECT 80.350 169.450 80.490 169.810 ;
        RECT 80.290 169.130 80.550 169.450 ;
        RECT 79.830 167.770 80.090 168.090 ;
        RECT 77.990 166.750 78.250 167.070 ;
        RECT 76.670 157.150 77.730 157.290 ;
        RECT 76.670 155.850 76.810 157.150 ;
        RECT 75.230 155.530 75.490 155.850 ;
        RECT 76.610 155.530 76.870 155.850 ;
        RECT 75.290 154.490 75.430 155.530 ;
        RECT 75.690 155.190 75.950 155.510 ;
        RECT 74.770 154.170 75.030 154.490 ;
        RECT 75.230 154.170 75.490 154.490 ;
        RECT 75.750 152.790 75.890 155.190 ;
        RECT 76.670 154.150 76.810 155.530 ;
        RECT 76.610 153.830 76.870 154.150 ;
        RECT 76.150 153.490 76.410 153.810 ;
        RECT 77.070 153.490 77.330 153.810 ;
        RECT 74.770 152.470 75.030 152.790 ;
        RECT 75.690 152.470 75.950 152.790 ;
        RECT 71.550 142.610 71.810 142.930 ;
        RECT 74.310 142.610 74.570 142.930 ;
        RECT 74.310 141.930 74.570 142.250 ;
        RECT 71.090 141.590 71.350 141.910 ;
        RECT 71.550 141.590 71.810 141.910 ;
        RECT 71.610 140.800 71.750 141.590 ;
        RECT 72.290 141.055 73.830 141.425 ;
        RECT 71.610 140.660 72.210 140.800 ;
        RECT 71.090 139.890 71.350 140.210 ;
        RECT 71.550 139.890 71.810 140.210 ;
        RECT 70.630 138.870 70.890 139.190 ;
        RECT 70.170 137.170 70.430 137.490 ;
        RECT 70.690 137.400 70.830 138.870 ;
        RECT 71.150 138.170 71.290 139.890 ;
        RECT 71.610 138.170 71.750 139.890 ;
        RECT 72.070 139.870 72.210 140.660 ;
        RECT 72.930 140.570 73.190 140.890 ;
        RECT 72.460 140.035 72.740 140.405 ;
        RECT 72.530 139.870 72.670 140.035 ;
        RECT 72.010 139.550 72.270 139.870 ;
        RECT 72.470 139.550 72.730 139.870 ;
        RECT 71.090 137.850 71.350 138.170 ;
        RECT 71.550 137.850 71.810 138.170 ;
        RECT 71.550 137.400 71.810 137.490 ;
        RECT 70.690 137.260 71.810 137.400 ;
        RECT 71.550 137.170 71.810 137.260 ;
        RECT 72.990 136.810 73.130 140.570 ;
        RECT 74.370 138.170 74.510 141.930 ;
        RECT 74.830 140.890 74.970 152.470 ;
        RECT 75.230 151.450 75.490 151.770 ;
        RECT 75.290 151.170 75.430 151.450 ;
        RECT 75.290 151.030 75.890 151.170 ;
        RECT 76.210 151.090 76.350 153.490 ;
        RECT 77.130 151.770 77.270 153.490 ;
        RECT 77.070 151.450 77.330 151.770 ;
        RECT 75.230 150.430 75.490 150.750 ;
        RECT 75.290 149.050 75.430 150.430 ;
        RECT 75.750 150.070 75.890 151.030 ;
        RECT 76.150 150.770 76.410 151.090 ;
        RECT 75.690 149.750 75.950 150.070 ;
        RECT 75.230 148.730 75.490 149.050 ;
        RECT 75.230 145.330 75.490 145.650 ;
        RECT 75.290 143.610 75.430 145.330 ;
        RECT 78.050 145.310 78.190 166.750 ;
        RECT 78.910 161.310 79.170 161.630 ;
        RECT 78.970 159.250 79.110 161.310 ;
        RECT 78.910 158.930 79.170 159.250 ;
        RECT 78.970 156.530 79.110 158.930 ;
        RECT 78.910 156.210 79.170 156.530 ;
        RECT 79.890 150.070 80.030 167.770 ;
        RECT 80.350 167.750 80.490 169.130 ;
        RECT 80.290 167.430 80.550 167.750 ;
        RECT 81.270 162.650 81.410 169.810 ;
        RECT 83.970 169.470 84.230 169.790 ;
        RECT 82.130 167.090 82.390 167.410 ;
        RECT 82.190 166.730 82.330 167.090 ;
        RECT 82.130 166.410 82.390 166.730 ;
        RECT 81.210 162.330 81.470 162.650 ;
        RECT 82.190 161.630 82.330 166.410 ;
        RECT 84.030 165.370 84.170 169.470 ;
        RECT 84.430 166.750 84.690 167.070 ;
        RECT 83.970 165.050 84.230 165.370 ;
        RECT 84.490 161.970 84.630 166.750 ;
        RECT 84.430 161.650 84.690 161.970 ;
        RECT 82.130 161.310 82.390 161.630 ;
        RECT 82.190 159.930 82.330 161.310 ;
        RECT 83.970 160.970 84.230 161.290 ;
        RECT 82.130 159.610 82.390 159.930 ;
        RECT 83.050 158.590 83.310 158.910 ;
        RECT 81.670 157.910 81.930 158.230 ;
        RECT 81.730 156.190 81.870 157.910 ;
        RECT 81.670 155.870 81.930 156.190 ;
        RECT 82.590 155.190 82.850 155.510 ;
        RECT 82.650 153.810 82.790 155.190 ;
        RECT 83.110 154.490 83.250 158.590 ;
        RECT 83.050 154.170 83.310 154.490 ;
        RECT 82.590 153.490 82.850 153.810 ;
        RECT 80.290 151.450 80.550 151.770 ;
        RECT 80.350 150.410 80.490 151.450 ;
        RECT 81.210 151.110 81.470 151.430 ;
        RECT 81.270 150.750 81.410 151.110 ;
        RECT 81.210 150.660 81.470 150.750 ;
        RECT 81.210 150.520 81.870 150.660 ;
        RECT 81.210 150.430 81.470 150.520 ;
        RECT 80.290 150.090 80.550 150.410 ;
        RECT 79.830 149.750 80.090 150.070 ;
        RECT 81.210 149.810 81.470 150.070 ;
        RECT 80.810 149.750 81.470 149.810 ;
        RECT 77.990 144.990 78.250 145.310 ;
        RECT 75.230 143.290 75.490 143.610 ;
        RECT 75.690 141.590 75.950 141.910 ;
        RECT 74.770 140.570 75.030 140.890 ;
        RECT 75.750 139.870 75.890 141.590 ;
        RECT 74.770 139.550 75.030 139.870 ;
        RECT 75.690 139.550 75.950 139.870 ;
        RECT 74.830 138.170 74.970 139.550 ;
        RECT 79.370 138.870 79.630 139.190 ;
        RECT 74.310 137.850 74.570 138.170 ;
        RECT 74.770 137.850 75.030 138.170 ;
        RECT 75.230 137.170 75.490 137.490 ;
        RECT 72.930 136.490 73.190 136.810 ;
        RECT 74.310 136.150 74.570 136.470 ;
        RECT 72.290 135.615 73.830 135.985 ;
        RECT 69.710 133.770 69.970 134.090 ;
        RECT 73.380 133.915 73.660 134.285 ;
        RECT 73.390 133.770 73.650 133.915 ;
        RECT 68.790 126.380 69.450 126.520 ;
        RECT 68.790 126.290 69.050 126.380 ;
        RECT 69.240 125.755 69.520 126.125 ;
        RECT 69.310 125.590 69.450 125.755 ;
        RECT 69.250 125.270 69.510 125.590 ;
        RECT 68.790 121.530 69.050 121.850 ;
        RECT 68.850 118.450 68.990 121.530 ;
        RECT 68.790 118.130 69.050 118.450 ;
        RECT 68.330 115.750 68.590 116.070 ;
        RECT 65.570 115.410 65.830 115.730 ;
        RECT 66.490 115.410 66.750 115.730 ;
        RECT 65.630 112.670 65.770 115.410 ;
        RECT 66.490 114.390 66.750 114.710 ;
        RECT 67.870 114.390 68.130 114.710 ;
        RECT 66.550 112.670 66.690 114.390 ;
        RECT 65.570 112.350 65.830 112.670 ;
        RECT 66.490 112.350 66.750 112.670 ;
        RECT 63.270 109.970 63.530 110.290 ;
        RECT 64.650 109.970 64.910 110.290 ;
        RECT 62.350 108.950 62.610 109.270 ;
        RECT 60.970 106.910 61.230 107.230 ;
        RECT 60.050 106.230 60.310 106.550 ;
        RECT 60.110 105.530 60.250 106.230 ;
        RECT 57.750 105.210 58.010 105.530 ;
        RECT 60.050 105.210 60.310 105.530 ;
        RECT 54.530 104.530 54.790 104.850 ;
        RECT 52.230 103.600 52.890 103.740 ;
        RECT 52.230 103.510 52.490 103.600 ;
        RECT 49.930 101.130 50.190 101.450 ;
        RECT 51.770 101.130 52.030 101.450 ;
        RECT 49.990 100.090 50.130 101.130 ;
        RECT 52.290 101.110 52.430 103.510 ;
        RECT 54.590 102.810 54.730 104.530 ;
        RECT 61.030 102.810 61.170 106.910 ;
        RECT 64.710 105.530 64.850 109.970 ;
        RECT 65.630 107.230 65.770 112.350 ;
        RECT 65.570 106.910 65.830 107.230 ;
        RECT 64.650 105.440 64.910 105.530 ;
        RECT 64.650 105.300 65.310 105.440 ;
        RECT 64.650 105.210 64.910 105.300 ;
        RECT 63.270 103.510 63.530 103.830 ;
        RECT 54.530 102.490 54.790 102.810 ;
        RECT 57.290 102.490 57.550 102.810 ;
        RECT 60.970 102.490 61.230 102.810 ;
        RECT 52.230 100.790 52.490 101.110 ;
        RECT 55.500 100.255 57.040 100.625 ;
        RECT 49.930 99.770 50.190 100.090 ;
        RECT 57.350 99.410 57.490 102.490 ;
        RECT 59.590 101.470 59.850 101.790 ;
        RECT 59.650 99.410 59.790 101.470 ;
        RECT 63.330 101.450 63.470 103.510 ;
        RECT 65.170 102.130 65.310 105.300 ;
        RECT 64.190 101.810 64.450 102.130 ;
        RECT 65.110 101.810 65.370 102.130 ;
        RECT 63.270 101.130 63.530 101.450 ;
        RECT 64.250 100.090 64.390 101.810 ;
        RECT 65.170 100.090 65.310 101.810 ;
        RECT 64.190 99.770 64.450 100.090 ;
        RECT 65.110 99.770 65.370 100.090 ;
        RECT 40.730 99.090 40.990 99.410 ;
        RECT 57.290 99.090 57.550 99.410 ;
        RECT 59.590 99.090 59.850 99.410 ;
        RECT 39.350 98.750 39.610 99.070 ;
        RECT 60.050 98.070 60.310 98.390 ;
        RECT 38.710 97.535 40.250 97.905 ;
        RECT 50.390 96.030 50.650 96.350 ;
        RECT 40.730 95.350 40.990 95.670 ;
        RECT 43.030 95.350 43.290 95.670 ;
        RECT 37.510 94.220 37.770 94.310 ;
        RECT 37.110 94.080 37.770 94.220 ;
        RECT 37.510 93.990 37.770 94.080 ;
        RECT 40.790 93.970 40.930 95.350 ;
        RECT 36.130 93.650 36.390 93.970 ;
        RECT 40.730 93.650 40.990 93.970 ;
        RECT 35.670 92.970 35.930 93.290 ;
        RECT 36.190 91.930 36.330 93.650 ;
        RECT 37.970 93.310 38.230 93.630 ;
        RECT 41.650 93.310 41.910 93.630 ;
        RECT 36.130 91.610 36.390 91.930 ;
        RECT 38.030 91.590 38.170 93.310 ;
        RECT 41.190 92.630 41.450 92.950 ;
        RECT 38.710 92.095 40.250 92.465 ;
        RECT 37.970 91.500 38.230 91.590 ;
        RECT 37.570 91.360 38.230 91.500 ;
        RECT 35.210 90.250 35.470 90.570 ;
        RECT 34.750 88.890 35.010 89.210 ;
        RECT 34.290 88.550 34.550 88.870 ;
        RECT 32.450 88.210 32.710 88.530 ;
        RECT 30.610 87.190 30.870 87.510 ;
        RECT 31.070 87.190 31.330 87.510 ;
        RECT 30.670 86.490 30.810 87.190 ;
        RECT 31.130 86.490 31.270 87.190 ;
        RECT 32.510 86.490 32.650 88.210 ;
        RECT 30.610 86.170 30.870 86.490 ;
        RECT 31.070 86.170 31.330 86.490 ;
        RECT 32.450 86.170 32.710 86.490 ;
        RECT 37.570 85.470 37.710 91.360 ;
        RECT 37.970 91.270 38.230 91.360 ;
        RECT 40.730 91.270 40.990 91.590 ;
        RECT 40.790 90.910 40.930 91.270 ;
        RECT 41.250 91.250 41.390 92.630 ;
        RECT 41.710 91.930 41.850 93.310 ;
        RECT 42.110 92.970 42.370 93.290 ;
        RECT 41.650 91.610 41.910 91.930 ;
        RECT 41.190 90.930 41.450 91.250 ;
        RECT 38.430 90.590 38.690 90.910 ;
        RECT 40.730 90.590 40.990 90.910 ;
        RECT 42.170 90.820 42.310 92.970 ;
        RECT 43.090 91.590 43.230 95.350 ;
        RECT 45.330 93.650 45.590 93.970 ;
        RECT 44.870 92.630 45.130 92.950 ;
        RECT 43.030 91.270 43.290 91.590 ;
        RECT 42.570 90.820 42.830 90.910 ;
        RECT 42.170 90.680 42.830 90.820 ;
        RECT 42.570 90.590 42.830 90.680 ;
        RECT 37.970 88.210 38.230 88.530 ;
        RECT 38.030 86.490 38.170 88.210 ;
        RECT 38.490 88.190 38.630 90.590 ;
        RECT 40.790 90.230 40.930 90.590 ;
        RECT 40.730 89.910 40.990 90.230 ;
        RECT 42.630 88.870 42.770 90.590 ;
        RECT 42.570 88.550 42.830 88.870 ;
        RECT 38.430 87.870 38.690 88.190 ;
        RECT 41.190 87.530 41.450 87.850 ;
        RECT 38.710 86.655 40.250 87.025 ;
        RECT 41.250 86.490 41.390 87.530 ;
        RECT 37.970 86.170 38.230 86.490 ;
        RECT 41.190 86.170 41.450 86.490 ;
        RECT 33.370 85.150 33.630 85.470 ;
        RECT 37.510 85.150 37.770 85.470 ;
        RECT 31.070 84.470 31.330 84.790 ;
        RECT 30.610 81.750 30.870 82.070 ;
        RECT 30.670 80.030 30.810 81.750 ;
        RECT 31.130 81.050 31.270 84.470 ;
        RECT 33.430 83.770 33.570 85.150 ;
        RECT 38.030 83.770 38.170 86.170 ;
        RECT 42.630 83.770 42.770 88.550 ;
        RECT 43.090 88.530 43.230 91.270 ;
        RECT 44.930 90.230 45.070 92.630 ;
        RECT 45.390 91.930 45.530 93.650 ;
        RECT 45.790 92.630 46.050 92.950 ;
        RECT 45.850 91.930 45.990 92.630 ;
        RECT 45.330 91.610 45.590 91.930 ;
        RECT 45.790 91.610 46.050 91.930 ;
        RECT 44.870 89.910 45.130 90.230 ;
        RECT 46.710 89.910 46.970 90.230 ;
        RECT 46.770 88.870 46.910 89.910 ;
        RECT 46.710 88.550 46.970 88.870 ;
        RECT 50.450 88.530 50.590 96.030 ;
        RECT 60.110 96.010 60.250 98.070 ;
        RECT 64.250 97.370 64.390 99.770 ;
        RECT 65.630 98.390 65.770 106.910 ;
        RECT 66.550 102.470 66.690 112.350 ;
        RECT 67.930 110.970 68.070 114.390 ;
        RECT 67.870 110.650 68.130 110.970 ;
        RECT 68.330 110.310 68.590 110.630 ;
        RECT 66.950 108.950 67.210 109.270 ;
        RECT 67.010 107.230 67.150 108.950 ;
        RECT 66.950 106.910 67.210 107.230 ;
        RECT 66.490 102.150 66.750 102.470 ;
        RECT 66.030 100.790 66.290 101.110 ;
        RECT 66.090 100.090 66.230 100.790 ;
        RECT 66.030 99.770 66.290 100.090 ;
        RECT 67.010 99.410 67.150 106.910 ;
        RECT 68.390 106.890 68.530 110.310 ;
        RECT 68.790 109.970 69.050 110.290 ;
        RECT 68.850 109.270 68.990 109.970 ;
        RECT 68.790 108.950 69.050 109.270 ;
        RECT 68.330 106.570 68.590 106.890 ;
        RECT 67.410 104.530 67.670 104.850 ;
        RECT 67.470 101.790 67.610 104.530 ;
        RECT 67.410 101.470 67.670 101.790 ;
        RECT 69.770 101.530 69.910 133.770 ;
        RECT 74.370 132.730 74.510 136.150 ;
        RECT 75.290 135.450 75.430 137.170 ;
        RECT 76.150 136.150 76.410 136.470 ;
        RECT 75.230 135.130 75.490 135.450 ;
        RECT 75.690 135.130 75.950 135.450 ;
        RECT 75.230 134.000 75.490 134.090 ;
        RECT 75.750 134.000 75.890 135.130 ;
        RECT 76.210 134.430 76.350 136.150 ;
        RECT 77.070 135.130 77.330 135.450 ;
        RECT 76.610 134.790 76.870 135.110 ;
        RECT 76.670 134.430 76.810 134.790 ;
        RECT 76.150 134.110 76.410 134.430 ;
        RECT 76.610 134.110 76.870 134.430 ;
        RECT 75.230 133.860 75.890 134.000 ;
        RECT 75.230 133.770 75.490 133.860 ;
        RECT 74.310 132.410 74.570 132.730 ;
        RECT 71.550 131.730 71.810 132.050 ;
        RECT 76.150 131.730 76.410 132.050 ;
        RECT 71.090 129.690 71.350 130.010 ;
        RECT 71.150 128.310 71.290 129.690 ;
        RECT 71.090 127.990 71.350 128.310 ;
        RECT 71.090 126.630 71.350 126.950 ;
        RECT 71.150 126.125 71.290 126.630 ;
        RECT 71.080 125.755 71.360 126.125 ;
        RECT 71.610 122.870 71.750 131.730 ;
        RECT 72.290 130.175 73.830 130.545 ;
        RECT 74.310 128.670 74.570 128.990 ;
        RECT 72.470 127.990 72.730 128.310 ;
        RECT 72.530 126.010 72.670 127.990 ;
        RECT 72.070 125.930 72.670 126.010 ;
        RECT 72.010 125.870 72.670 125.930 ;
        RECT 72.010 125.610 72.270 125.870 ;
        RECT 72.290 124.735 73.830 125.105 ;
        RECT 71.550 122.550 71.810 122.870 ;
        RECT 73.850 122.550 74.110 122.870 ;
        RECT 73.910 120.830 74.050 122.550 ;
        RECT 74.370 120.830 74.510 128.670 ;
        RECT 75.230 126.630 75.490 126.950 ;
        RECT 74.770 125.950 75.030 126.270 ;
        RECT 74.830 121.850 74.970 125.950 ;
        RECT 75.290 124.570 75.430 126.630 ;
        RECT 76.210 125.930 76.350 131.730 ;
        RECT 77.130 128.050 77.270 135.130 ;
        RECT 79.430 134.430 79.570 138.870 ;
        RECT 79.370 134.110 79.630 134.430 ;
        RECT 78.450 133.430 78.710 133.750 ;
        RECT 78.510 128.650 78.650 133.430 ;
        RECT 78.450 128.330 78.710 128.650 ;
        RECT 76.670 127.910 77.270 128.050 ;
        RECT 76.150 125.610 76.410 125.930 ;
        RECT 75.230 124.250 75.490 124.570 ;
        RECT 76.670 123.970 76.810 127.910 ;
        RECT 77.990 125.270 78.250 125.590 ;
        RECT 76.210 123.830 76.810 123.970 ;
        RECT 75.230 122.550 75.490 122.870 ;
        RECT 74.770 121.530 75.030 121.850 ;
        RECT 75.290 121.170 75.430 122.550 ;
        RECT 75.230 120.850 75.490 121.170 ;
        RECT 73.850 120.510 74.110 120.830 ;
        RECT 74.310 120.510 74.570 120.830 ;
        RECT 72.290 119.295 73.830 119.665 ;
        RECT 74.370 117.770 74.510 120.510 ;
        RECT 74.770 119.830 75.030 120.150 ;
        RECT 74.830 119.130 74.970 119.830 ;
        RECT 74.770 118.810 75.030 119.130 ;
        RECT 74.310 117.450 74.570 117.770 ;
        RECT 70.630 117.110 70.890 117.430 ;
        RECT 70.690 116.410 70.830 117.110 ;
        RECT 70.630 116.090 70.890 116.410 ;
        RECT 76.210 116.370 76.350 123.830 ;
        RECT 76.610 123.460 76.870 123.550 ;
        RECT 76.610 123.320 77.730 123.460 ;
        RECT 76.610 123.230 76.870 123.320 ;
        RECT 76.210 116.230 76.810 116.370 ;
        RECT 75.230 115.410 75.490 115.730 ;
        RECT 70.170 115.070 70.430 115.390 ;
        RECT 70.230 110.970 70.370 115.070 ;
        RECT 71.550 114.390 71.810 114.710 ;
        RECT 71.610 112.330 71.750 114.390 ;
        RECT 72.290 113.855 73.830 114.225 ;
        RECT 75.290 113.010 75.430 115.410 ;
        RECT 75.230 112.920 75.490 113.010 ;
        RECT 74.830 112.780 75.490 112.920 ;
        RECT 71.550 112.010 71.810 112.330 ;
        RECT 70.170 110.650 70.430 110.970 ;
        RECT 70.170 109.970 70.430 110.290 ;
        RECT 70.230 108.250 70.370 109.970 ;
        RECT 71.090 108.950 71.350 109.270 ;
        RECT 70.170 107.930 70.430 108.250 ;
        RECT 71.150 107.570 71.290 108.950 ;
        RECT 72.290 108.415 73.830 108.785 ;
        RECT 71.090 107.250 71.350 107.570 ;
        RECT 70.630 106.910 70.890 107.230 ;
        RECT 74.310 106.910 74.570 107.230 ;
        RECT 70.690 105.530 70.830 106.910 ;
        RECT 73.850 106.230 74.110 106.550 ;
        RECT 73.910 105.530 74.050 106.230 ;
        RECT 70.630 105.210 70.890 105.530 ;
        RECT 73.850 105.210 74.110 105.530 ;
        RECT 70.690 102.130 70.830 105.210 ;
        RECT 74.370 105.190 74.510 106.910 ;
        RECT 74.310 104.870 74.570 105.190 ;
        RECT 74.830 104.850 74.970 112.780 ;
        RECT 75.230 112.690 75.490 112.780 ;
        RECT 76.150 111.670 76.410 111.990 ;
        RECT 76.210 110.290 76.350 111.670 ;
        RECT 76.150 109.970 76.410 110.290 ;
        RECT 75.230 109.290 75.490 109.610 ;
        RECT 75.290 104.850 75.430 109.290 ;
        RECT 74.770 104.530 75.030 104.850 ;
        RECT 75.230 104.530 75.490 104.850 ;
        RECT 72.290 102.975 73.830 103.345 ;
        RECT 75.290 102.810 75.430 104.530 ;
        RECT 74.770 102.490 75.030 102.810 ;
        RECT 75.230 102.490 75.490 102.810 ;
        RECT 70.630 101.810 70.890 102.130 ;
        RECT 67.470 101.110 67.610 101.470 ;
        RECT 69.770 101.390 70.370 101.530 ;
        RECT 67.410 100.790 67.670 101.110 ;
        RECT 69.710 100.790 69.970 101.110 ;
        RECT 67.470 99.750 67.610 100.790 ;
        RECT 67.410 99.430 67.670 99.750 ;
        RECT 66.950 99.090 67.210 99.410 ;
        RECT 67.470 99.070 67.610 99.430 ;
        RECT 69.770 99.410 69.910 100.790 ;
        RECT 69.710 99.090 69.970 99.410 ;
        RECT 67.410 98.750 67.670 99.070 ;
        RECT 65.570 98.070 65.830 98.390 ;
        RECT 68.330 98.070 68.590 98.390 ;
        RECT 64.190 97.050 64.450 97.370 ;
        RECT 66.030 96.030 66.290 96.350 ;
        RECT 51.770 95.690 52.030 96.010 ;
        RECT 60.050 95.690 60.310 96.010 ;
        RECT 51.830 94.650 51.970 95.690 ;
        RECT 53.150 95.350 53.410 95.670 ;
        RECT 51.770 94.330 52.030 94.650 ;
        RECT 53.210 88.530 53.350 95.350 ;
        RECT 55.500 94.815 57.040 95.185 ;
        RECT 54.070 93.650 54.330 93.970 ;
        RECT 54.130 91.930 54.270 93.650 ;
        RECT 64.190 93.310 64.450 93.630 ;
        RECT 54.070 91.610 54.330 91.930 ;
        RECT 64.250 91.250 64.390 93.310 ;
        RECT 54.990 90.930 55.250 91.250 ;
        RECT 64.190 90.930 64.450 91.250 ;
        RECT 54.530 90.590 54.790 90.910 ;
        RECT 54.590 88.530 54.730 90.590 ;
        RECT 55.050 89.210 55.190 90.930 ;
        RECT 63.270 90.590 63.530 90.910 ;
        RECT 57.290 90.250 57.550 90.570 ;
        RECT 55.500 89.375 57.040 89.745 ;
        RECT 57.350 89.210 57.490 90.250 ;
        RECT 62.350 89.910 62.610 90.230 ;
        RECT 54.990 88.890 55.250 89.210 ;
        RECT 57.290 88.890 57.550 89.210 ;
        RECT 62.410 88.530 62.550 89.910 ;
        RECT 43.030 88.210 43.290 88.530 ;
        RECT 50.390 88.210 50.650 88.530 ;
        RECT 50.850 88.210 51.110 88.530 ;
        RECT 53.150 88.440 53.410 88.530 ;
        RECT 52.750 88.300 53.410 88.440 ;
        RECT 50.910 86.490 51.050 88.210 ;
        RECT 50.850 86.170 51.110 86.490 ;
        RECT 52.750 85.470 52.890 88.300 ;
        RECT 53.150 88.210 53.410 88.300 ;
        RECT 54.530 88.210 54.790 88.530 ;
        RECT 62.350 88.210 62.610 88.530 ;
        RECT 62.810 88.210 63.070 88.530 ;
        RECT 53.150 87.190 53.410 87.510 ;
        RECT 53.210 86.490 53.350 87.190 ;
        RECT 54.590 86.490 54.730 88.210 ;
        RECT 62.870 87.510 63.010 88.210 ;
        RECT 59.590 87.190 59.850 87.510 ;
        RECT 62.810 87.190 63.070 87.510 ;
        RECT 53.150 86.170 53.410 86.490 ;
        RECT 54.530 86.170 54.790 86.490 ;
        RECT 58.670 85.490 58.930 85.810 ;
        RECT 43.950 85.150 44.210 85.470 ;
        RECT 49.010 85.150 49.270 85.470 ;
        RECT 52.690 85.150 52.950 85.470 ;
        RECT 53.610 85.150 53.870 85.470 ;
        RECT 44.010 83.770 44.150 85.150 ;
        RECT 49.070 83.770 49.210 85.150 ;
        RECT 53.670 83.770 53.810 85.150 ;
        RECT 55.500 83.935 57.040 84.305 ;
        RECT 58.730 83.770 58.870 85.490 ;
        RECT 33.370 83.450 33.630 83.770 ;
        RECT 37.970 83.450 38.230 83.770 ;
        RECT 42.570 83.450 42.830 83.770 ;
        RECT 43.950 83.450 44.210 83.770 ;
        RECT 49.010 83.450 49.270 83.770 ;
        RECT 53.610 83.450 53.870 83.770 ;
        RECT 58.670 83.450 58.930 83.770 ;
        RECT 59.650 83.090 59.790 87.190 ;
        RECT 63.330 86.490 63.470 90.590 ;
        RECT 66.090 88.530 66.230 96.030 ;
        RECT 67.410 95.690 67.670 96.010 ;
        RECT 67.470 94.650 67.610 95.690 ;
        RECT 68.390 94.650 68.530 98.070 ;
        RECT 67.410 94.330 67.670 94.650 ;
        RECT 68.330 94.330 68.590 94.650 ;
        RECT 69.240 90.395 69.520 90.765 ;
        RECT 69.250 90.250 69.510 90.395 ;
        RECT 68.330 89.910 68.590 90.230 ;
        RECT 66.030 88.210 66.290 88.530 ;
        RECT 66.090 86.490 66.230 88.210 ;
        RECT 68.390 88.190 68.530 89.910 ;
        RECT 70.230 89.210 70.370 101.390 ;
        RECT 71.550 101.130 71.810 101.450 ;
        RECT 70.630 100.790 70.890 101.110 ;
        RECT 70.690 99.410 70.830 100.790 ;
        RECT 70.630 99.090 70.890 99.410 ;
        RECT 71.610 97.370 71.750 101.130 ;
        RECT 72.290 97.535 73.830 97.905 ;
        RECT 71.550 97.050 71.810 97.370 ;
        RECT 74.830 96.350 74.970 102.490 ;
        RECT 75.290 99.410 75.430 102.490 ;
        RECT 75.230 99.090 75.490 99.410 ;
        RECT 75.290 96.690 75.430 99.090 ;
        RECT 75.230 96.370 75.490 96.690 ;
        RECT 74.770 96.030 75.030 96.350 ;
        RECT 72.290 92.095 73.830 92.465 ;
        RECT 70.630 90.590 70.890 90.910 ;
        RECT 71.550 90.590 71.810 90.910 ;
        RECT 72.470 90.590 72.730 90.910 ;
        RECT 70.170 88.890 70.430 89.210 ;
        RECT 70.690 88.530 70.830 90.590 ;
        RECT 71.610 89.210 71.750 90.590 ;
        RECT 71.550 88.890 71.810 89.210 ;
        RECT 72.530 88.870 72.670 90.590 ;
        RECT 75.230 89.910 75.490 90.230 ;
        RECT 75.290 88.870 75.430 89.910 ;
        RECT 72.470 88.550 72.730 88.870 ;
        RECT 75.230 88.550 75.490 88.870 ;
        RECT 70.630 88.210 70.890 88.530 ;
        RECT 71.090 88.210 71.350 88.530 ;
        RECT 68.330 87.870 68.590 88.190 ;
        RECT 63.270 86.170 63.530 86.490 ;
        RECT 66.030 86.170 66.290 86.490 ;
        RECT 60.510 85.830 60.770 86.150 ;
        RECT 61.430 85.830 61.690 86.150 ;
        RECT 60.570 83.770 60.710 85.830 ;
        RECT 60.970 84.470 61.230 84.790 ;
        RECT 60.510 83.450 60.770 83.770 ;
        RECT 31.530 82.770 31.790 83.090 ;
        RECT 34.750 82.770 35.010 83.090 ;
        RECT 46.250 82.770 46.510 83.090 ;
        RECT 50.390 82.770 50.650 83.090 ;
        RECT 58.210 82.770 58.470 83.090 ;
        RECT 59.590 82.770 59.850 83.090 ;
        RECT 31.070 80.730 31.330 81.050 ;
        RECT 30.610 79.710 30.870 80.030 ;
        RECT 25.550 78.010 25.810 78.330 ;
        RECT 29.690 78.010 29.950 78.330 ;
        RECT 30.610 77.330 30.870 77.650 ;
        RECT 30.670 73.910 30.810 77.330 ;
        RECT 31.070 74.270 31.330 74.590 ;
        RECT 30.610 73.590 30.870 73.910 ;
        RECT 30.150 71.210 30.410 71.530 ;
        RECT 30.210 69.150 30.350 71.210 ;
        RECT 31.130 70.170 31.270 74.270 ;
        RECT 31.590 74.250 31.730 82.770 ;
        RECT 32.910 82.430 33.170 82.750 ;
        RECT 32.970 77.990 33.110 82.430 ;
        RECT 34.810 81.050 34.950 82.770 ;
        RECT 36.130 81.750 36.390 82.070 ;
        RECT 34.750 80.730 35.010 81.050 ;
        RECT 32.910 77.670 33.170 77.990 ;
        RECT 35.210 77.330 35.470 77.650 ;
        RECT 32.910 76.990 33.170 77.310 ;
        RECT 32.970 74.590 33.110 76.990 ;
        RECT 35.270 75.270 35.410 77.330 ;
        RECT 35.210 74.950 35.470 75.270 ;
        RECT 32.910 74.270 33.170 74.590 ;
        RECT 31.530 73.930 31.790 74.250 ;
        RECT 33.830 73.930 34.090 74.250 ;
        RECT 34.740 74.075 35.020 74.445 ;
        RECT 31.070 69.850 31.330 70.170 ;
        RECT 33.890 69.490 34.030 73.930 ;
        RECT 34.810 72.890 34.950 74.075 ;
        RECT 34.750 72.570 35.010 72.890 ;
        RECT 35.210 72.570 35.470 72.890 ;
        RECT 35.270 69.490 35.410 72.570 ;
        RECT 36.190 71.530 36.330 81.750 ;
        RECT 38.710 81.215 40.250 81.585 ;
        RECT 46.310 81.050 46.450 82.770 ;
        RECT 50.450 81.050 50.590 82.770 ;
        RECT 54.530 81.750 54.790 82.070 ;
        RECT 54.590 81.050 54.730 81.750 ;
        RECT 58.270 81.050 58.410 82.770 ;
        RECT 46.250 80.730 46.510 81.050 ;
        RECT 50.390 80.730 50.650 81.050 ;
        RECT 54.530 80.730 54.790 81.050 ;
        RECT 58.210 80.730 58.470 81.050 ;
        RECT 36.590 79.710 36.850 80.030 ;
        RECT 45.330 79.710 45.590 80.030 ;
        RECT 48.550 79.710 48.810 80.030 ;
        RECT 51.770 79.710 52.030 80.030 ;
        RECT 36.650 77.650 36.790 79.710 ;
        RECT 37.050 79.030 37.310 79.350 ;
        RECT 36.590 77.330 36.850 77.650 ;
        RECT 36.650 74.930 36.790 77.330 ;
        RECT 37.110 76.970 37.250 79.030 ;
        RECT 40.730 77.670 40.990 77.990 ;
        RECT 37.510 77.560 37.770 77.650 ;
        RECT 37.510 77.420 38.170 77.560 ;
        RECT 37.510 77.330 37.770 77.420 ;
        RECT 37.050 76.650 37.310 76.970 ;
        RECT 37.050 74.950 37.310 75.270 ;
        RECT 36.590 74.610 36.850 74.930 ;
        RECT 36.650 72.210 36.790 74.610 ;
        RECT 37.110 72.210 37.250 74.950 ;
        RECT 37.510 74.270 37.770 74.590 ;
        RECT 38.030 74.445 38.170 77.420 ;
        RECT 38.710 75.775 40.250 76.145 ;
        RECT 40.790 74.590 40.930 77.670 ;
        RECT 41.650 77.330 41.910 77.650 ;
        RECT 43.950 77.330 44.210 77.650 ;
        RECT 41.190 76.990 41.450 77.310 ;
        RECT 41.250 75.610 41.390 76.990 ;
        RECT 41.190 75.290 41.450 75.610 ;
        RECT 36.590 71.890 36.850 72.210 ;
        RECT 37.050 71.890 37.310 72.210 ;
        RECT 36.130 71.210 36.390 71.530 ;
        RECT 33.830 69.170 34.090 69.490 ;
        RECT 35.210 69.170 35.470 69.490 ;
        RECT 36.190 69.150 36.330 71.210 ;
        RECT 30.150 68.830 30.410 69.150 ;
        RECT 31.990 68.830 32.250 69.150 ;
        RECT 36.130 68.830 36.390 69.150 ;
        RECT 26.470 68.150 26.730 68.470 ;
        RECT 30.150 68.150 30.410 68.470 ;
        RECT 24.630 63.390 24.890 63.710 ;
        RECT 25.550 63.390 25.810 63.710 ;
        RECT 24.690 58.610 24.830 63.390 ;
        RECT 25.610 61.330 25.750 63.390 ;
        RECT 26.530 62.010 26.670 68.150 ;
        RECT 30.210 62.010 30.350 68.150 ;
        RECT 32.050 66.770 32.190 68.830 ;
        RECT 32.450 68.490 32.710 68.810 ;
        RECT 31.990 66.450 32.250 66.770 ;
        RECT 26.470 61.690 26.730 62.010 ;
        RECT 30.150 61.690 30.410 62.010 ;
        RECT 25.550 61.010 25.810 61.330 ;
        RECT 31.530 61.010 31.790 61.330 ;
        RECT 30.610 60.670 30.870 60.990 ;
        RECT 30.670 59.290 30.810 60.670 ;
        RECT 30.610 58.970 30.870 59.290 ;
        RECT 24.630 58.290 24.890 58.610 ;
        RECT 28.770 57.950 29.030 58.270 ;
        RECT 28.830 56.200 28.970 57.950 ;
        RECT 31.590 56.200 31.730 61.010 ;
        RECT 32.510 58.270 32.650 68.490 ;
        RECT 33.370 68.150 33.630 68.470 ;
        RECT 33.430 66.770 33.570 68.150 ;
        RECT 33.370 66.450 33.630 66.770 ;
        RECT 33.370 65.770 33.630 66.090 ;
        RECT 33.430 63.710 33.570 65.770 ;
        RECT 37.570 63.710 37.710 74.270 ;
        RECT 37.960 74.075 38.240 74.445 ;
        RECT 40.730 74.270 40.990 74.590 ;
        RECT 41.250 74.250 41.390 75.290 ;
        RECT 41.710 75.010 41.850 77.330 ;
        RECT 42.110 76.650 42.370 76.970 ;
        RECT 42.170 75.610 42.310 76.650 ;
        RECT 42.110 75.290 42.370 75.610 ;
        RECT 41.710 74.870 42.310 75.010 ;
        RECT 40.270 73.930 40.530 74.250 ;
        RECT 41.190 73.930 41.450 74.250 ;
        RECT 41.650 73.930 41.910 74.250 ;
        RECT 40.330 72.120 40.470 73.930 ;
        RECT 40.730 72.120 40.990 72.210 ;
        RECT 40.330 71.980 40.990 72.120 ;
        RECT 40.730 71.890 40.990 71.980 ;
        RECT 38.710 70.335 40.250 70.705 ;
        RECT 38.890 69.170 39.150 69.490 ;
        RECT 38.950 66.430 39.090 69.170 ;
        RECT 41.250 68.470 41.390 73.930 ;
        RECT 41.710 72.210 41.850 73.930 ;
        RECT 41.650 71.890 41.910 72.210 ;
        RECT 42.170 71.870 42.310 74.870 ;
        RECT 44.010 74.590 44.150 77.330 ;
        RECT 44.410 75.290 44.670 75.610 ;
        RECT 44.470 74.590 44.610 75.290 ;
        RECT 44.870 74.950 45.130 75.270 ;
        RECT 43.950 74.270 44.210 74.590 ;
        RECT 44.410 74.270 44.670 74.590 ;
        RECT 44.410 73.590 44.670 73.910 ;
        RECT 42.570 71.890 42.830 72.210 ;
        RECT 43.490 71.890 43.750 72.210 ;
        RECT 42.110 71.610 42.370 71.870 ;
        RECT 41.710 71.550 42.370 71.610 ;
        RECT 41.710 71.470 42.310 71.550 ;
        RECT 41.710 68.810 41.850 71.470 ;
        RECT 42.110 70.870 42.370 71.190 ;
        RECT 41.650 68.490 41.910 68.810 ;
        RECT 41.190 68.150 41.450 68.470 ;
        RECT 42.170 66.965 42.310 70.870 ;
        RECT 42.100 66.850 42.380 66.965 ;
        RECT 41.710 66.770 42.380 66.850 ;
        RECT 42.630 66.770 42.770 71.890 ;
        RECT 43.550 67.450 43.690 71.890 ;
        RECT 44.470 68.380 44.610 73.590 ;
        RECT 44.930 71.725 45.070 74.950 ;
        RECT 45.390 72.890 45.530 79.710 ;
        RECT 48.610 78.330 48.750 79.710 ;
        RECT 48.550 78.010 48.810 78.330 ;
        RECT 47.630 77.330 47.890 77.650 ;
        RECT 47.170 76.310 47.430 76.630 ;
        RECT 47.230 74.590 47.370 76.310 ;
        RECT 47.170 74.270 47.430 74.590 ;
        RECT 46.250 73.590 46.510 73.910 ;
        RECT 47.170 73.590 47.430 73.910 ;
        RECT 45.330 72.570 45.590 72.890 ;
        RECT 44.860 71.355 45.140 71.725 ;
        RECT 46.310 69.830 46.450 73.590 ;
        RECT 46.250 69.510 46.510 69.830 ;
        RECT 46.310 68.810 46.450 69.510 ;
        RECT 46.250 68.490 46.510 68.810 ;
        RECT 44.470 68.240 45.530 68.380 ;
        RECT 43.490 67.130 43.750 67.450 ;
        RECT 41.650 66.710 42.380 66.770 ;
        RECT 41.650 66.450 41.910 66.710 ;
        RECT 42.100 66.595 42.380 66.710 ;
        RECT 42.570 66.450 42.830 66.770 ;
        RECT 38.890 66.110 39.150 66.430 ;
        RECT 37.970 65.430 38.230 65.750 ;
        RECT 40.730 65.430 40.990 65.750 ;
        RECT 43.030 65.430 43.290 65.750 ;
        RECT 33.370 63.390 33.630 63.710 ;
        RECT 34.750 63.620 35.010 63.710 ;
        RECT 34.350 63.480 35.010 63.620 ;
        RECT 32.450 57.950 32.710 58.270 ;
        RECT 34.350 56.200 34.490 63.480 ;
        RECT 34.750 63.390 35.010 63.480 ;
        RECT 36.590 63.390 36.850 63.710 ;
        RECT 37.510 63.390 37.770 63.710 ;
        RECT 36.130 61.010 36.390 61.330 ;
        RECT 36.190 58.010 36.330 61.010 ;
        RECT 36.650 60.990 36.790 63.390 ;
        RECT 37.510 62.710 37.770 63.030 ;
        RECT 37.570 62.010 37.710 62.710 ;
        RECT 37.510 61.690 37.770 62.010 ;
        RECT 36.590 60.670 36.850 60.990 ;
        RECT 38.030 58.270 38.170 65.430 ;
        RECT 38.710 64.895 40.250 65.265 ;
        RECT 40.270 64.640 40.530 64.730 ;
        RECT 40.790 64.640 40.930 65.430 ;
        RECT 40.270 64.500 40.930 64.640 ;
        RECT 40.270 64.410 40.530 64.500 ;
        RECT 40.270 63.050 40.530 63.370 ;
        RECT 40.330 60.730 40.470 63.050 ;
        RECT 42.110 61.240 42.370 61.330 ;
        RECT 42.110 61.100 42.770 61.240 ;
        RECT 42.110 61.010 42.370 61.100 ;
        RECT 40.330 60.590 40.930 60.730 ;
        RECT 38.710 59.455 40.250 59.825 ;
        RECT 40.790 59.290 40.930 60.590 ;
        RECT 40.730 58.970 40.990 59.290 ;
        RECT 36.190 57.870 37.250 58.010 ;
        RECT 37.970 57.950 38.230 58.270 ;
        RECT 40.270 58.180 40.530 58.270 ;
        RECT 39.870 58.040 40.530 58.180 ;
        RECT 37.110 56.200 37.250 57.870 ;
        RECT 39.870 56.200 40.010 58.040 ;
        RECT 40.270 57.950 40.530 58.040 ;
        RECT 42.630 56.200 42.770 61.100 ;
        RECT 43.090 58.270 43.230 65.430 ;
        RECT 43.550 61.330 43.690 67.130 ;
        RECT 45.390 66.770 45.530 68.240 ;
        RECT 47.230 66.965 47.370 73.590 ;
        RECT 44.410 66.450 44.670 66.770 ;
        RECT 45.330 66.450 45.590 66.770 ;
        RECT 47.160 66.595 47.440 66.965 ;
        RECT 43.950 65.430 44.210 65.750 ;
        RECT 44.010 64.730 44.150 65.430 ;
        RECT 44.470 64.730 44.610 66.450 ;
        RECT 47.690 65.750 47.830 77.330 ;
        RECT 49.930 76.990 50.190 77.310 ;
        RECT 49.010 74.270 49.270 74.590 ;
        RECT 49.070 71.870 49.210 74.270 ;
        RECT 49.990 73.910 50.130 76.990 ;
        RECT 51.830 75.610 51.970 79.710 ;
        RECT 55.500 78.495 57.040 78.865 ;
        RECT 61.030 78.330 61.170 84.470 ;
        RECT 61.490 83.090 61.630 85.830 ;
        RECT 68.390 83.770 68.530 87.870 ;
        RECT 68.330 83.450 68.590 83.770 ;
        RECT 67.410 83.110 67.670 83.430 ;
        RECT 61.430 82.770 61.690 83.090 ;
        RECT 64.190 80.050 64.450 80.370 ;
        RECT 62.810 79.710 63.070 80.030 ;
        RECT 62.350 79.030 62.610 79.350 ;
        RECT 60.970 78.010 61.230 78.330 ;
        RECT 61.430 77.670 61.690 77.990 ;
        RECT 60.050 76.990 60.310 77.310 ;
        RECT 54.990 76.310 55.250 76.630 ;
        RECT 51.770 75.290 52.030 75.610 ;
        RECT 52.230 74.950 52.490 75.270 ;
        RECT 50.850 73.930 51.110 74.250 ;
        RECT 49.930 73.590 50.190 73.910 ;
        RECT 49.010 71.550 49.270 71.870 ;
        RECT 48.090 66.450 48.350 66.770 ;
        RECT 47.630 65.430 47.890 65.750 ;
        RECT 48.150 64.730 48.290 66.450 ;
        RECT 43.950 64.410 44.210 64.730 ;
        RECT 44.410 64.410 44.670 64.730 ;
        RECT 48.090 64.410 48.350 64.730 ;
        RECT 49.070 63.710 49.210 71.550 ;
        RECT 50.910 68.380 51.050 73.930 ;
        RECT 51.310 71.550 51.570 71.870 ;
        RECT 51.370 70.170 51.510 71.550 ;
        RECT 52.290 71.190 52.430 74.950 ;
        RECT 55.050 74.590 55.190 76.310 ;
        RECT 60.110 75.610 60.250 76.990 ;
        RECT 60.050 75.290 60.310 75.610 ;
        RECT 53.610 74.270 53.870 74.590 ;
        RECT 54.990 74.270 55.250 74.590 ;
        RECT 53.150 73.590 53.410 73.910 ;
        RECT 53.210 72.210 53.350 73.590 ;
        RECT 53.670 72.890 53.810 74.270 ;
        RECT 58.200 74.075 58.480 74.445 ;
        RECT 55.500 73.055 57.040 73.425 ;
        RECT 53.610 72.570 53.870 72.890 ;
        RECT 53.150 71.890 53.410 72.210 ;
        RECT 54.070 71.890 54.330 72.210 ;
        RECT 51.770 70.870 52.030 71.190 ;
        RECT 52.230 70.870 52.490 71.190 ;
        RECT 51.310 69.850 51.570 70.170 ;
        RECT 51.830 68.470 51.970 70.870 ;
        RECT 51.310 68.380 51.570 68.470 ;
        RECT 50.910 68.240 51.570 68.380 ;
        RECT 51.310 68.150 51.570 68.240 ;
        RECT 51.770 68.150 52.030 68.470 ;
        RECT 50.390 65.430 50.650 65.750 ;
        RECT 45.790 63.620 46.050 63.710 ;
        RECT 45.390 63.480 46.050 63.620 ;
        RECT 43.490 61.010 43.750 61.330 ;
        RECT 43.030 57.950 43.290 58.270 ;
        RECT 45.390 56.200 45.530 63.480 ;
        RECT 45.790 63.390 46.050 63.480 ;
        RECT 46.250 63.390 46.510 63.710 ;
        RECT 48.550 63.390 48.810 63.710 ;
        RECT 49.010 63.390 49.270 63.710 ;
        RECT 46.310 61.330 46.450 63.390 ;
        RECT 48.610 61.330 48.750 63.390 ;
        RECT 46.250 61.010 46.510 61.330 ;
        RECT 48.550 61.010 48.810 61.330 ;
        RECT 50.450 58.270 50.590 65.430 ;
        RECT 51.370 62.010 51.510 68.150 ;
        RECT 52.290 67.450 52.430 70.870 ;
        RECT 53.150 68.830 53.410 69.150 ;
        RECT 53.210 67.450 53.350 68.830 ;
        RECT 52.230 67.130 52.490 67.450 ;
        RECT 53.150 67.130 53.410 67.450 ;
        RECT 52.220 66.595 52.500 66.965 ;
        RECT 52.230 66.450 52.490 66.595 ;
        RECT 53.210 64.730 53.350 67.130 ;
        RECT 54.130 66.430 54.270 71.890 ;
        RECT 55.900 71.355 56.180 71.725 ;
        RECT 54.530 70.870 54.790 71.190 ;
        RECT 54.590 69.830 54.730 70.870 ;
        RECT 54.990 69.850 55.250 70.170 ;
        RECT 54.530 69.510 54.790 69.830 ;
        RECT 55.050 68.070 55.190 69.850 ;
        RECT 55.970 68.810 56.110 71.355 ;
        RECT 56.830 70.870 57.090 71.190 ;
        RECT 57.290 70.870 57.550 71.190 ;
        RECT 56.890 69.150 57.030 70.870 ;
        RECT 57.350 70.170 57.490 70.870 ;
        RECT 57.290 69.850 57.550 70.170 ;
        RECT 56.830 68.830 57.090 69.150 ;
        RECT 55.910 68.490 56.170 68.810 ;
        RECT 54.590 67.930 55.190 68.070 ;
        RECT 54.070 66.110 54.330 66.430 ;
        RECT 53.150 64.410 53.410 64.730 ;
        RECT 53.150 63.390 53.410 63.710 ;
        RECT 51.310 61.690 51.570 62.010 ;
        RECT 50.850 61.350 51.110 61.670 ;
        RECT 47.630 58.180 47.890 58.270 ;
        RECT 47.630 58.040 48.290 58.180 ;
        RECT 47.630 57.950 47.890 58.040 ;
        RECT 48.150 56.200 48.290 58.040 ;
        RECT 50.390 57.950 50.650 58.270 ;
        RECT 50.910 56.200 51.050 61.350 ;
        RECT 51.310 59.990 51.570 60.310 ;
        RECT 51.370 59.290 51.510 59.990 ;
        RECT 51.310 58.970 51.570 59.290 ;
        RECT 53.210 56.650 53.350 63.390 ;
        RECT 54.590 61.240 54.730 67.930 ;
        RECT 55.500 67.615 57.040 67.985 ;
        RECT 58.270 66.770 58.410 74.075 ;
        RECT 61.490 73.910 61.630 77.670 ;
        RECT 62.410 76.970 62.550 79.030 ;
        RECT 62.870 77.990 63.010 79.710 ;
        RECT 63.730 79.030 63.990 79.350 ;
        RECT 63.790 78.330 63.930 79.030 ;
        RECT 63.730 78.010 63.990 78.330 ;
        RECT 62.810 77.670 63.070 77.990 ;
        RECT 62.350 76.650 62.610 76.970 ;
        RECT 62.410 75.610 62.550 76.650 ;
        RECT 62.350 75.290 62.610 75.610 ;
        RECT 62.870 74.590 63.010 77.670 ;
        RECT 64.250 77.650 64.390 80.050 ;
        RECT 65.110 77.670 65.370 77.990 ;
        RECT 64.190 77.330 64.450 77.650 ;
        RECT 64.250 74.590 64.390 77.330 ;
        RECT 62.810 74.270 63.070 74.590 ;
        RECT 64.190 74.270 64.450 74.590 ;
        RECT 61.430 73.590 61.690 73.910 ;
        RECT 62.810 71.890 63.070 72.210 ;
        RECT 60.970 71.550 61.230 71.870 ;
        RECT 61.030 70.170 61.170 71.550 ;
        RECT 62.870 70.170 63.010 71.890 ;
        RECT 64.190 70.870 64.450 71.190 ;
        RECT 60.970 69.850 61.230 70.170 ;
        RECT 62.810 69.850 63.070 70.170 ;
        RECT 61.430 68.150 61.690 68.470 ;
        RECT 58.210 66.450 58.470 66.770 ;
        RECT 54.990 65.430 55.250 65.750 ;
        RECT 55.450 65.430 55.710 65.750 ;
        RECT 55.050 64.730 55.190 65.430 ;
        RECT 54.990 64.410 55.250 64.730 ;
        RECT 55.510 63.710 55.650 65.430 ;
        RECT 55.450 63.390 55.710 63.710 ;
        RECT 59.130 63.390 59.390 63.710 ;
        RECT 59.590 63.390 59.850 63.710 ;
        RECT 55.500 62.175 57.040 62.545 ;
        RECT 56.830 61.690 57.090 62.010 ;
        RECT 55.450 61.240 55.710 61.330 ;
        RECT 54.590 61.100 55.710 61.240 ;
        RECT 55.450 61.010 55.710 61.100 ;
        RECT 53.610 59.990 53.870 60.310 ;
        RECT 53.670 59.290 53.810 59.990 ;
        RECT 53.610 58.970 53.870 59.290 ;
        RECT 56.890 58.270 57.030 61.690 ;
        RECT 54.990 57.950 55.250 58.270 ;
        RECT 56.830 57.950 57.090 58.270 ;
        RECT 53.210 56.510 53.810 56.650 ;
        RECT 53.670 56.200 53.810 56.510 ;
        RECT 28.760 54.700 29.040 56.200 ;
        RECT 31.520 54.870 31.800 56.200 ;
        RECT 28.760 54.200 29.050 54.700 ;
        RECT 31.520 54.200 31.810 54.870 ;
        RECT 34.280 54.610 34.560 56.200 ;
        RECT 37.040 54.700 37.320 56.200 ;
        RECT 39.800 54.760 40.080 56.200 ;
        RECT 42.560 54.780 42.840 56.200 ;
        RECT 45.320 54.980 45.600 56.200 ;
        RECT 48.080 55.070 48.360 56.200 ;
        RECT 34.280 54.200 34.570 54.610 ;
        RECT 37.040 54.200 37.330 54.700 ;
        RECT 39.800 54.200 40.090 54.760 ;
        RECT 42.560 54.200 42.850 54.780 ;
        RECT 45.320 54.200 45.610 54.980 ;
        RECT 48.080 54.200 48.370 55.070 ;
        RECT 50.840 54.830 51.120 56.200 ;
        RECT 53.600 55.000 53.880 56.200 ;
        RECT 55.050 55.970 55.190 57.950 ;
        RECT 55.500 56.735 57.040 57.105 ;
        RECT 55.970 56.340 56.570 56.480 ;
        RECT 55.970 55.970 56.110 56.340 ;
        RECT 56.430 56.200 56.570 56.340 ;
        RECT 59.190 56.200 59.330 63.390 ;
        RECT 59.650 62.010 59.790 63.390 ;
        RECT 59.590 61.690 59.850 62.010 ;
        RECT 61.490 61.330 61.630 68.150 ;
        RECT 64.250 67.450 64.390 70.870 ;
        RECT 64.190 67.130 64.450 67.450 ;
        RECT 65.170 66.430 65.310 77.670 ;
        RECT 65.570 76.310 65.830 76.630 ;
        RECT 65.630 75.610 65.770 76.310 ;
        RECT 65.570 75.290 65.830 75.610 ;
        RECT 65.570 74.270 65.830 74.590 ;
        RECT 65.630 71.190 65.770 74.270 ;
        RECT 65.570 70.870 65.830 71.190 ;
        RECT 65.110 66.110 65.370 66.430 ;
        RECT 65.630 65.750 65.770 70.870 ;
        RECT 67.470 66.430 67.610 83.110 ;
        RECT 68.390 83.090 68.530 83.450 ;
        RECT 68.330 82.770 68.590 83.090 ;
        RECT 70.690 82.070 70.830 88.210 ;
        RECT 68.790 81.750 69.050 82.070 ;
        RECT 70.630 81.750 70.890 82.070 ;
        RECT 67.870 79.030 68.130 79.350 ;
        RECT 67.930 77.990 68.070 79.030 ;
        RECT 68.850 78.330 68.990 81.750 ;
        RECT 71.150 80.030 71.290 88.210 ;
        RECT 76.150 87.870 76.410 88.190 ;
        RECT 71.550 87.530 71.810 87.850 ;
        RECT 71.610 86.490 71.750 87.530 ;
        RECT 72.290 86.655 73.830 87.025 ;
        RECT 71.550 86.170 71.810 86.490 ;
        RECT 71.610 84.790 71.750 86.170 ;
        RECT 76.210 85.470 76.350 87.870 ;
        RECT 76.150 85.150 76.410 85.470 ;
        RECT 71.550 84.470 71.810 84.790 ;
        RECT 71.610 82.660 71.750 84.470 ;
        RECT 72.470 82.660 72.730 82.750 ;
        RECT 71.610 82.520 72.730 82.660 ;
        RECT 71.090 79.710 71.350 80.030 ;
        RECT 68.790 78.010 69.050 78.330 ;
        RECT 67.870 77.670 68.130 77.990 ;
        RECT 68.330 76.310 68.590 76.630 ;
        RECT 68.390 74.590 68.530 76.310 ;
        RECT 68.330 74.270 68.590 74.590 ;
        RECT 71.610 74.250 71.750 82.520 ;
        RECT 72.470 82.430 72.730 82.520 ;
        RECT 72.290 81.215 73.830 81.585 ;
        RECT 76.210 80.710 76.350 85.150 ;
        RECT 76.150 80.390 76.410 80.710 ;
        RECT 73.850 79.710 74.110 80.030 ;
        RECT 73.910 78.330 74.050 79.710 ;
        RECT 76.670 79.350 76.810 116.230 ;
        RECT 77.590 116.070 77.730 123.320 ;
        RECT 78.050 117.770 78.190 125.270 ;
        RECT 78.510 119.130 78.650 128.330 ;
        RECT 79.370 126.970 79.630 127.290 ;
        RECT 78.910 125.270 79.170 125.590 ;
        RECT 78.970 121.510 79.110 125.270 ;
        RECT 79.430 121.760 79.570 126.970 ;
        RECT 79.890 126.950 80.030 149.750 ;
        RECT 80.810 149.670 81.410 149.750 ;
        RECT 80.810 148.370 80.950 149.670 ;
        RECT 81.730 149.050 81.870 150.520 ;
        RECT 81.670 148.730 81.930 149.050 ;
        RECT 82.650 148.370 82.790 153.490 ;
        RECT 84.030 150.750 84.170 160.970 ;
        RECT 84.950 154.490 85.090 201.430 ;
        RECT 85.870 199.170 86.010 201.520 ;
        RECT 86.330 200.730 86.470 205.850 ;
        RECT 87.250 202.090 87.390 209.930 ;
        RECT 89.080 209.055 90.620 209.425 ;
        RECT 93.230 208.210 93.370 212.200 ;
        RECT 100.590 208.890 100.730 212.200 ;
        RECT 100.530 208.570 100.790 208.890 ;
        RECT 107.950 208.550 108.090 212.200 ;
        RECT 107.890 208.230 108.150 208.550 ;
        RECT 93.170 207.890 93.430 208.210 ;
        RECT 96.390 207.890 96.650 208.210 ;
        RECT 103.750 207.890 104.010 208.210 ;
        RECT 110.190 207.890 110.450 208.210 ;
        RECT 90.410 207.550 90.670 207.870 ;
        RECT 88.110 207.210 88.370 207.530 ;
        RECT 87.650 206.870 87.910 207.190 ;
        RECT 87.710 205.150 87.850 206.870 ;
        RECT 87.650 204.830 87.910 205.150 ;
        RECT 87.650 202.110 87.910 202.430 ;
        RECT 86.730 201.770 86.990 202.090 ;
        RECT 87.190 201.770 87.450 202.090 ;
        RECT 86.270 200.410 86.530 200.730 ;
        RECT 86.790 200.050 86.930 201.770 ;
        RECT 86.730 199.730 86.990 200.050 ;
        RECT 85.870 199.030 86.470 199.170 ;
        RECT 87.250 199.030 87.390 201.770 ;
        RECT 87.710 200.730 87.850 202.110 ;
        RECT 88.170 201.750 88.310 207.210 ;
        RECT 90.470 206.170 90.610 207.550 ;
        RECT 92.710 207.210 92.970 207.530 ;
        RECT 90.410 205.850 90.670 206.170 ;
        RECT 92.770 205.150 92.910 207.210 ;
        RECT 93.170 206.870 93.430 207.190 ;
        RECT 93.230 205.150 93.370 206.870 ;
        RECT 92.710 204.830 92.970 205.150 ;
        RECT 93.170 204.830 93.430 205.150 ;
        RECT 88.570 204.490 88.830 204.810 ;
        RECT 91.330 204.490 91.590 204.810 ;
        RECT 88.110 201.430 88.370 201.750 ;
        RECT 87.650 200.410 87.910 200.730 ;
        RECT 85.350 193.610 85.610 193.930 ;
        RECT 85.410 186.790 85.550 193.610 ;
        RECT 85.350 186.470 85.610 186.790 ;
        RECT 85.810 183.750 86.070 184.070 ;
        RECT 85.870 181.010 86.010 183.750 ;
        RECT 85.810 180.690 86.070 181.010 ;
        RECT 85.350 176.950 85.610 177.270 ;
        RECT 85.410 176.250 85.550 176.950 ;
        RECT 85.350 175.930 85.610 176.250 ;
        RECT 85.350 174.230 85.610 174.550 ;
        RECT 85.810 174.230 86.070 174.550 ;
        RECT 85.410 173.530 85.550 174.230 ;
        RECT 85.350 173.210 85.610 173.530 ;
        RECT 85.870 172.850 86.010 174.230 ;
        RECT 85.810 172.530 86.070 172.850 ;
        RECT 85.810 166.070 86.070 166.390 ;
        RECT 85.350 155.190 85.610 155.510 ;
        RECT 85.410 154.490 85.550 155.190 ;
        RECT 84.890 154.170 85.150 154.490 ;
        RECT 85.350 154.170 85.610 154.490 ;
        RECT 84.890 153.490 85.150 153.810 ;
        RECT 84.950 153.325 85.090 153.490 ;
        RECT 84.880 152.955 85.160 153.325 ;
        RECT 83.050 150.430 83.310 150.750 ;
        RECT 83.970 150.430 84.230 150.750 ;
        RECT 80.750 148.050 81.010 148.370 ;
        RECT 82.130 148.050 82.390 148.370 ;
        RECT 82.590 148.050 82.850 148.370 ;
        RECT 82.190 146.330 82.330 148.050 ;
        RECT 82.130 146.010 82.390 146.330 ;
        RECT 82.190 139.530 82.330 146.010 ;
        RECT 83.110 142.930 83.250 150.430 ;
        RECT 83.050 142.610 83.310 142.930 ;
        RECT 82.130 139.210 82.390 139.530 ;
        RECT 82.190 137.490 82.330 139.210 ;
        RECT 82.130 137.170 82.390 137.490 ;
        RECT 83.050 137.170 83.310 137.490 ;
        RECT 82.190 132.050 82.330 137.170 ;
        RECT 82.130 131.730 82.390 132.050 ;
        RECT 81.670 130.710 81.930 131.030 ;
        RECT 81.730 128.990 81.870 130.710 ;
        RECT 83.110 129.670 83.250 137.170 ;
        RECT 83.510 131.730 83.770 132.050 ;
        RECT 83.570 129.670 83.710 131.730 ;
        RECT 83.050 129.350 83.310 129.670 ;
        RECT 83.510 129.350 83.770 129.670 ;
        RECT 81.670 128.670 81.930 128.990 ;
        RECT 80.290 127.990 80.550 128.310 ;
        RECT 79.830 126.630 80.090 126.950 ;
        RECT 80.350 126.270 80.490 127.990 ;
        RECT 80.290 125.950 80.550 126.270 ;
        RECT 80.750 125.950 81.010 126.270 ;
        RECT 83.500 126.010 83.780 126.125 ;
        RECT 84.030 126.010 84.170 150.430 ;
        RECT 85.870 143.610 86.010 166.070 ;
        RECT 86.330 159.590 86.470 199.030 ;
        RECT 87.190 198.710 87.450 199.030 ;
        RECT 87.650 198.710 87.910 199.030 ;
        RECT 87.250 195.290 87.390 198.710 ;
        RECT 87.710 196.310 87.850 198.710 ;
        RECT 87.650 195.990 87.910 196.310 ;
        RECT 87.190 194.970 87.450 195.290 ;
        RECT 87.710 194.270 87.850 195.990 ;
        RECT 87.650 193.950 87.910 194.270 ;
        RECT 88.170 188.830 88.310 201.430 ;
        RECT 88.630 200.730 88.770 204.490 ;
        RECT 89.080 203.615 90.620 203.985 ;
        RECT 91.390 203.450 91.530 204.490 ;
        RECT 93.230 204.470 93.370 204.830 ;
        RECT 95.470 204.490 95.730 204.810 ;
        RECT 93.170 204.150 93.430 204.470 ;
        RECT 91.330 203.130 91.590 203.450 ;
        RECT 95.010 203.130 95.270 203.450 ;
        RECT 92.250 202.790 92.510 203.110 ;
        RECT 92.310 202.090 92.450 202.790 ;
        RECT 92.250 201.770 92.510 202.090 ;
        RECT 93.170 201.770 93.430 202.090 ;
        RECT 88.570 200.410 88.830 200.730 ;
        RECT 92.250 199.390 92.510 199.710 ;
        RECT 89.080 198.175 90.620 198.545 ;
        RECT 91.330 195.990 91.590 196.310 ;
        RECT 91.390 195.290 91.530 195.990 ;
        RECT 91.330 194.970 91.590 195.290 ;
        RECT 89.080 192.735 90.620 193.105 ;
        RECT 90.870 190.890 91.130 191.210 ;
        RECT 90.930 189.170 91.070 190.890 ;
        RECT 90.870 188.850 91.130 189.170 ;
        RECT 88.110 188.510 88.370 188.830 ;
        RECT 87.650 187.830 87.910 188.150 ;
        RECT 87.710 187.130 87.850 187.830 ;
        RECT 89.080 187.295 90.620 187.665 ;
        RECT 87.650 186.810 87.910 187.130 ;
        RECT 87.190 186.130 87.450 186.450 ;
        RECT 91.330 186.130 91.590 186.450 ;
        RECT 87.250 179.990 87.390 186.130 ;
        RECT 90.870 185.450 91.130 185.770 ;
        RECT 88.570 185.110 88.830 185.430 ;
        RECT 89.030 185.110 89.290 185.430 ;
        RECT 88.630 184.070 88.770 185.110 ;
        RECT 88.570 183.750 88.830 184.070 ;
        RECT 88.630 183.390 88.770 183.750 ;
        RECT 88.110 183.070 88.370 183.390 ;
        RECT 88.570 183.070 88.830 183.390 ;
        RECT 87.650 182.390 87.910 182.710 ;
        RECT 87.710 181.690 87.850 182.390 ;
        RECT 88.170 181.690 88.310 183.070 ;
        RECT 89.090 182.710 89.230 185.110 ;
        RECT 90.930 183.390 91.070 185.450 ;
        RECT 90.870 183.070 91.130 183.390 ;
        RECT 89.030 182.620 89.290 182.710 ;
        RECT 88.630 182.480 89.290 182.620 ;
        RECT 87.650 181.370 87.910 181.690 ;
        RECT 88.110 181.370 88.370 181.690 ;
        RECT 88.630 181.350 88.770 182.480 ;
        RECT 89.030 182.390 89.290 182.480 ;
        RECT 89.080 181.855 90.620 182.225 ;
        RECT 90.930 181.690 91.070 183.070 ;
        RECT 90.870 181.370 91.130 181.690 ;
        RECT 88.570 181.030 88.830 181.350 ;
        RECT 90.410 180.690 90.670 181.010 ;
        RECT 89.030 180.010 89.290 180.330 ;
        RECT 87.190 179.670 87.450 179.990 ;
        RECT 88.570 179.670 88.830 179.990 ;
        RECT 87.190 177.970 87.450 178.290 ;
        RECT 87.250 174.550 87.390 177.970 ;
        RECT 88.630 175.910 88.770 179.670 ;
        RECT 89.090 178.290 89.230 180.010 ;
        RECT 89.950 179.670 90.210 179.990 ;
        RECT 89.030 177.970 89.290 178.290 ;
        RECT 90.010 177.950 90.150 179.670 ;
        RECT 90.470 178.970 90.610 180.690 ;
        RECT 90.410 178.650 90.670 178.970 ;
        RECT 91.390 178.630 91.530 186.130 ;
        RECT 91.790 183.070 92.050 183.390 ;
        RECT 91.850 180.670 91.990 183.070 ;
        RECT 91.790 180.350 92.050 180.670 ;
        RECT 92.310 178.630 92.450 199.390 ;
        RECT 92.710 197.350 92.970 197.670 ;
        RECT 92.770 194.270 92.910 197.350 ;
        RECT 92.710 193.950 92.970 194.270 ;
        RECT 92.770 191.890 92.910 193.950 ;
        RECT 92.710 191.570 92.970 191.890 ;
        RECT 92.710 185.110 92.970 185.430 ;
        RECT 91.330 178.310 91.590 178.630 ;
        RECT 92.250 178.310 92.510 178.630 ;
        RECT 92.770 178.290 92.910 185.110 ;
        RECT 93.230 180.330 93.370 201.770 ;
        RECT 95.070 200.050 95.210 203.130 ;
        RECT 95.010 199.730 95.270 200.050 ;
        RECT 95.530 199.710 95.670 204.490 ;
        RECT 96.450 203.450 96.590 207.890 ;
        RECT 101.910 206.870 102.170 207.190 ;
        RECT 101.970 206.170 102.110 206.870 ;
        RECT 98.230 205.850 98.490 206.170 ;
        RECT 101.910 205.850 102.170 206.170 ;
        RECT 97.770 204.490 98.030 204.810 ;
        RECT 96.390 203.130 96.650 203.450 ;
        RECT 97.830 203.110 97.970 204.490 ;
        RECT 96.850 202.790 97.110 203.110 ;
        RECT 97.770 202.790 98.030 203.110 ;
        RECT 95.470 199.390 95.730 199.710 ;
        RECT 95.010 193.950 95.270 194.270 ;
        RECT 94.090 193.270 94.350 193.590 ;
        RECT 94.150 192.570 94.290 193.270 ;
        RECT 94.090 192.250 94.350 192.570 ;
        RECT 95.070 191.210 95.210 193.950 ;
        RECT 95.530 193.930 95.670 199.390 ;
        RECT 96.910 198.010 97.050 202.790 ;
        RECT 97.770 202.340 98.030 202.430 ;
        RECT 98.290 202.340 98.430 205.850 ;
        RECT 101.970 205.150 102.110 205.850 ;
        RECT 101.910 204.830 102.170 205.150 ;
        RECT 102.830 204.490 103.090 204.810 ;
        RECT 100.530 204.150 100.790 204.470 ;
        RECT 100.590 203.450 100.730 204.150 ;
        RECT 100.530 203.130 100.790 203.450 ;
        RECT 100.990 203.020 101.250 203.110 ;
        RECT 102.370 203.020 102.630 203.110 ;
        RECT 100.990 202.880 102.630 203.020 ;
        RECT 100.990 202.790 101.250 202.880 ;
        RECT 102.370 202.790 102.630 202.880 ;
        RECT 97.770 202.200 98.430 202.340 ;
        RECT 102.890 202.285 103.030 204.490 ;
        RECT 103.810 203.450 103.950 207.890 ;
        RECT 108.810 207.100 109.070 207.190 ;
        RECT 108.410 206.960 109.070 207.100 ;
        RECT 105.870 206.335 107.410 206.705 ;
        RECT 105.130 205.510 105.390 205.830 ;
        RECT 104.670 205.400 104.930 205.490 ;
        RECT 104.270 205.260 104.930 205.400 ;
        RECT 103.750 203.130 104.010 203.450 ;
        RECT 97.770 202.110 98.030 202.200 ;
        RECT 98.290 201.750 98.430 202.200 ;
        RECT 100.530 201.770 100.790 202.090 ;
        RECT 102.820 201.915 103.100 202.285 ;
        RECT 98.230 201.430 98.490 201.750 ;
        RECT 99.610 201.430 99.870 201.750 ;
        RECT 97.770 198.710 98.030 199.030 ;
        RECT 96.850 197.690 97.110 198.010 ;
        RECT 96.390 195.990 96.650 196.310 ;
        RECT 96.450 194.950 96.590 195.990 ;
        RECT 96.390 194.630 96.650 194.950 ;
        RECT 95.470 193.610 95.730 193.930 ;
        RECT 95.530 191.890 95.670 193.610 ;
        RECT 95.470 191.570 95.730 191.890 ;
        RECT 95.010 190.890 95.270 191.210 ;
        RECT 95.930 190.890 96.190 191.210 ;
        RECT 95.990 189.850 96.130 190.890 ;
        RECT 95.930 189.530 96.190 189.850 ;
        RECT 96.450 189.510 96.590 194.630 ;
        RECT 97.830 193.590 97.970 198.710 ;
        RECT 98.290 197.330 98.430 201.430 ;
        RECT 98.690 199.390 98.950 199.710 ;
        RECT 98.230 197.010 98.490 197.330 ;
        RECT 98.750 196.310 98.890 199.390 ;
        RECT 99.670 199.370 99.810 201.430 ;
        RECT 100.590 200.390 100.730 201.770 ;
        RECT 103.290 201.430 103.550 201.750 ;
        RECT 103.750 201.430 104.010 201.750 ;
        RECT 102.830 200.410 103.090 200.730 ;
        RECT 100.530 200.070 100.790 200.390 ;
        RECT 99.610 199.050 99.870 199.370 ;
        RECT 99.150 198.710 99.410 199.030 ;
        RECT 98.230 195.990 98.490 196.310 ;
        RECT 98.690 195.990 98.950 196.310 ;
        RECT 96.850 193.270 97.110 193.590 ;
        RECT 97.310 193.270 97.570 193.590 ;
        RECT 97.770 193.270 98.030 193.590 ;
        RECT 96.910 190.870 97.050 193.270 ;
        RECT 97.370 192.650 97.510 193.270 ;
        RECT 97.370 192.510 97.970 192.650 ;
        RECT 97.830 192.230 97.970 192.510 ;
        RECT 97.770 191.910 98.030 192.230 ;
        RECT 96.850 190.550 97.110 190.870 ;
        RECT 96.390 189.190 96.650 189.510 ;
        RECT 96.910 188.150 97.050 190.550 ;
        RECT 97.830 188.490 97.970 191.910 ;
        RECT 98.290 188.830 98.430 195.990 ;
        RECT 99.210 195.290 99.350 198.710 ;
        RECT 99.670 198.010 99.810 199.050 ;
        RECT 99.610 197.690 99.870 198.010 ;
        RECT 99.610 197.010 99.870 197.330 ;
        RECT 99.150 194.970 99.410 195.290 ;
        RECT 99.670 191.210 99.810 197.010 ;
        RECT 100.590 196.310 100.730 200.070 ;
        RECT 101.910 198.710 102.170 199.030 ;
        RECT 101.970 197.330 102.110 198.710 ;
        RECT 102.890 197.410 103.030 200.410 ;
        RECT 103.350 200.390 103.490 201.430 ;
        RECT 103.290 200.070 103.550 200.390 ;
        RECT 103.350 197.670 103.490 200.070 ;
        RECT 103.810 199.030 103.950 201.430 ;
        RECT 104.270 199.170 104.410 205.260 ;
        RECT 104.670 205.170 104.930 205.260 ;
        RECT 105.190 203.450 105.330 205.510 ;
        RECT 106.510 205.170 106.770 205.490 ;
        RECT 105.130 203.130 105.390 203.450 ;
        RECT 104.670 202.790 104.930 203.110 ;
        RECT 104.730 200.730 104.870 202.790 ;
        RECT 106.570 202.770 106.710 205.170 ;
        RECT 106.510 202.450 106.770 202.770 ;
        RECT 105.130 201.770 105.390 202.090 ;
        RECT 104.670 200.410 104.930 200.730 ;
        RECT 105.190 199.710 105.330 201.770 ;
        RECT 107.890 201.430 108.150 201.750 ;
        RECT 105.870 200.895 107.410 201.265 ;
        RECT 105.590 200.410 105.850 200.730 ;
        RECT 105.130 199.390 105.390 199.710 ;
        RECT 104.270 199.030 105.330 199.170 ;
        RECT 103.750 198.710 104.010 199.030 ;
        RECT 101.910 197.010 102.170 197.330 ;
        RECT 102.430 197.270 103.030 197.410 ;
        RECT 103.290 197.350 103.550 197.670 ;
        RECT 100.530 195.990 100.790 196.310 ;
        RECT 101.970 193.590 102.110 197.010 ;
        RECT 101.910 193.270 102.170 193.590 ;
        RECT 101.970 192.570 102.110 193.270 ;
        RECT 101.910 192.250 102.170 192.570 ;
        RECT 99.610 190.890 99.870 191.210 ;
        RECT 102.430 190.870 102.570 197.270 ;
        RECT 102.830 196.670 103.090 196.990 ;
        RECT 102.890 195.290 103.030 196.670 ;
        RECT 103.290 196.330 103.550 196.650 ;
        RECT 103.350 195.290 103.490 196.330 ;
        RECT 103.750 195.990 104.010 196.310 ;
        RECT 102.830 194.970 103.090 195.290 ;
        RECT 103.290 194.970 103.550 195.290 ;
        RECT 102.890 190.870 103.030 194.970 ;
        RECT 103.290 193.445 103.550 193.590 ;
        RECT 103.280 193.075 103.560 193.445 ;
        RECT 103.810 193.330 103.950 195.990 ;
        RECT 104.670 194.290 104.930 194.610 ;
        RECT 104.730 193.500 104.870 194.290 ;
        RECT 104.270 193.360 104.870 193.500 ;
        RECT 103.810 193.190 104.030 193.330 ;
        RECT 103.290 192.250 103.550 192.570 ;
        RECT 103.890 192.270 104.030 193.190 ;
        RECT 99.150 190.550 99.410 190.870 ;
        RECT 102.370 190.550 102.630 190.870 ;
        RECT 102.830 190.550 103.090 190.870 ;
        RECT 98.230 188.510 98.490 188.830 ;
        RECT 97.770 188.170 98.030 188.490 ;
        RECT 96.850 187.830 97.110 188.150 ;
        RECT 98.230 187.830 98.490 188.150 ;
        RECT 98.690 187.830 98.950 188.150 ;
        RECT 98.290 186.790 98.430 187.830 ;
        RECT 98.750 187.130 98.890 187.830 ;
        RECT 99.210 187.130 99.350 190.550 ;
        RECT 102.430 189.930 102.570 190.550 ;
        RECT 102.430 189.790 103.030 189.930 ;
        RECT 98.690 186.810 98.950 187.130 ;
        RECT 99.150 186.810 99.410 187.130 ;
        RECT 98.230 186.470 98.490 186.790 ;
        RECT 97.770 186.130 98.030 186.450 ;
        RECT 96.390 185.450 96.650 185.770 ;
        RECT 95.930 182.390 96.190 182.710 ;
        RECT 94.090 181.370 94.350 181.690 ;
        RECT 93.170 180.010 93.430 180.330 ;
        RECT 94.150 179.990 94.290 181.370 ;
        RECT 94.550 181.030 94.810 181.350 ;
        RECT 94.090 179.670 94.350 179.990 ;
        RECT 94.610 178.970 94.750 181.030 ;
        RECT 95.990 180.410 96.130 182.390 ;
        RECT 95.010 180.010 95.270 180.330 ;
        RECT 95.530 180.270 96.130 180.410 ;
        RECT 95.070 178.970 95.210 180.010 ;
        RECT 94.550 178.650 94.810 178.970 ;
        RECT 95.010 178.650 95.270 178.970 ;
        RECT 94.090 178.310 94.350 178.630 ;
        RECT 90.870 177.970 91.130 178.290 ;
        RECT 92.710 177.970 92.970 178.290 ;
        RECT 89.950 177.630 90.210 177.950 ;
        RECT 89.080 176.415 90.620 176.785 ;
        RECT 88.570 175.590 88.830 175.910 ;
        RECT 89.030 175.250 89.290 175.570 ;
        RECT 87.190 174.230 87.450 174.550 ;
        RECT 87.250 166.730 87.390 174.230 ;
        RECT 89.090 173.190 89.230 175.250 ;
        RECT 90.930 174.550 91.070 177.970 ;
        RECT 94.150 177.860 94.290 178.310 ;
        RECT 95.530 178.290 95.670 180.270 ;
        RECT 95.930 179.670 96.190 179.990 ;
        RECT 95.990 178.290 96.130 179.670 ;
        RECT 95.470 177.970 95.730 178.290 ;
        RECT 95.930 177.970 96.190 178.290 ;
        RECT 94.150 177.720 94.750 177.860 ;
        RECT 92.250 177.290 92.510 177.610 ;
        RECT 91.330 174.910 91.590 175.230 ;
        RECT 90.870 174.230 91.130 174.550 ;
        RECT 89.030 172.870 89.290 173.190 ;
        RECT 87.650 171.510 87.910 171.830 ;
        RECT 89.090 171.740 89.230 172.870 ;
        RECT 88.630 171.600 89.230 171.740 ;
        RECT 87.710 170.130 87.850 171.510 ;
        RECT 87.650 169.810 87.910 170.130 ;
        RECT 88.630 168.090 88.770 171.600 ;
        RECT 89.080 170.975 90.620 171.345 ;
        RECT 91.390 170.130 91.530 174.910 ;
        RECT 92.310 174.890 92.450 177.290 ;
        RECT 93.630 176.950 93.890 177.270 ;
        RECT 93.690 175.230 93.830 176.950 ;
        RECT 93.630 174.910 93.890 175.230 ;
        RECT 92.250 174.570 92.510 174.890 ;
        RECT 92.310 173.530 92.450 174.570 ;
        RECT 92.250 173.210 92.510 173.530 ;
        RECT 93.690 173.190 93.830 174.910 ;
        RECT 93.630 173.100 93.890 173.190 ;
        RECT 93.230 172.960 93.890 173.100 ;
        RECT 91.330 169.810 91.590 170.130 ;
        RECT 89.030 169.130 89.290 169.450 ;
        RECT 88.570 167.770 88.830 168.090 ;
        RECT 89.090 167.070 89.230 169.130 ;
        RECT 91.330 167.430 91.590 167.750 ;
        RECT 89.030 166.810 89.290 167.070 ;
        RECT 88.630 166.750 89.290 166.810 ;
        RECT 87.190 166.410 87.450 166.730 ;
        RECT 88.630 166.670 89.230 166.750 ;
        RECT 88.110 166.070 88.370 166.390 ;
        RECT 88.170 162.650 88.310 166.070 ;
        RECT 88.630 164.770 88.770 166.670 ;
        RECT 89.080 165.535 90.620 165.905 ;
        RECT 88.630 164.630 89.230 164.770 ;
        RECT 89.090 163.670 89.230 164.630 ;
        RECT 90.870 164.370 91.130 164.690 ;
        RECT 89.030 163.350 89.290 163.670 ;
        RECT 88.110 162.330 88.370 162.650 ;
        RECT 89.090 161.630 89.230 163.350 ;
        RECT 90.930 162.650 91.070 164.370 ;
        RECT 91.390 163.410 91.530 167.430 ;
        RECT 93.230 167.070 93.370 172.960 ;
        RECT 93.630 172.870 93.890 172.960 ;
        RECT 93.630 171.510 93.890 171.830 ;
        RECT 93.690 170.810 93.830 171.510 ;
        RECT 93.630 170.490 93.890 170.810 ;
        RECT 93.170 166.750 93.430 167.070 ;
        RECT 92.710 166.410 92.970 166.730 ;
        RECT 91.390 163.270 91.990 163.410 ;
        RECT 90.870 162.330 91.130 162.650 ;
        RECT 91.850 161.630 91.990 163.270 ;
        RECT 89.030 161.310 89.290 161.630 ;
        RECT 91.790 161.310 92.050 161.630 ;
        RECT 90.870 160.970 91.130 161.290 ;
        RECT 89.080 160.095 90.620 160.465 ;
        RECT 86.270 159.270 86.530 159.590 ;
        RECT 86.330 156.530 86.470 159.270 ;
        RECT 88.110 158.590 88.370 158.910 ;
        RECT 86.270 156.210 86.530 156.530 ;
        RECT 88.170 156.190 88.310 158.590 ;
        RECT 90.410 157.910 90.670 158.230 ;
        RECT 90.470 156.190 90.610 157.910 ;
        RECT 90.930 157.210 91.070 160.970 ;
        RECT 91.330 160.630 91.590 160.950 ;
        RECT 91.790 160.630 92.050 160.950 ;
        RECT 91.390 159.930 91.530 160.630 ;
        RECT 91.330 159.610 91.590 159.930 ;
        RECT 90.870 156.890 91.130 157.210 ;
        RECT 91.850 156.530 91.990 160.630 ;
        RECT 92.250 156.550 92.510 156.870 ;
        RECT 90.870 156.210 91.130 156.530 ;
        RECT 91.790 156.210 92.050 156.530 ;
        RECT 88.110 155.870 88.370 156.190 ;
        RECT 90.410 155.870 90.670 156.190 ;
        RECT 88.170 153.810 88.310 155.870 ;
        RECT 89.080 154.655 90.620 155.025 ;
        RECT 90.930 154.490 91.070 156.210 ;
        RECT 90.870 154.170 91.130 154.490 ;
        RECT 90.930 153.810 91.070 154.170 ;
        RECT 88.110 153.490 88.370 153.810 ;
        RECT 90.870 153.490 91.130 153.810 ;
        RECT 90.410 152.810 90.670 153.130 ;
        RECT 90.470 151.770 90.610 152.810 ;
        RECT 87.190 151.450 87.450 151.770 ;
        RECT 90.410 151.450 90.670 151.770 ;
        RECT 86.270 144.990 86.530 145.310 ;
        RECT 85.810 143.290 86.070 143.610 ;
        RECT 86.330 142.930 86.470 144.990 ;
        RECT 87.250 142.930 87.390 151.450 ;
        RECT 87.650 150.430 87.910 150.750 ;
        RECT 87.710 150.070 87.850 150.430 ;
        RECT 87.650 149.750 87.910 150.070 ;
        RECT 88.570 149.750 88.830 150.070 ;
        RECT 91.330 149.750 91.590 150.070 ;
        RECT 88.630 149.050 88.770 149.750 ;
        RECT 89.080 149.215 90.620 149.585 ;
        RECT 91.390 149.050 91.530 149.750 ;
        RECT 88.570 148.730 88.830 149.050 ;
        RECT 91.330 148.730 91.590 149.050 ;
        RECT 88.630 142.930 88.770 148.730 ;
        RECT 91.330 147.030 91.590 147.350 ;
        RECT 90.870 144.650 91.130 144.970 ;
        RECT 89.080 143.775 90.620 144.145 ;
        RECT 89.950 142.950 90.210 143.270 ;
        RECT 86.270 142.610 86.530 142.930 ;
        RECT 87.190 142.610 87.450 142.930 ;
        RECT 88.570 142.610 88.830 142.930 ;
        RECT 89.030 142.610 89.290 142.930 ;
        RECT 85.350 137.850 85.610 138.170 ;
        RECT 84.430 134.790 84.690 135.110 ;
        RECT 80.810 124.570 80.950 125.950 ;
        RECT 83.500 125.870 84.170 126.010 ;
        RECT 83.500 125.755 83.780 125.870 ;
        RECT 83.050 125.270 83.310 125.590 ;
        RECT 80.750 124.250 81.010 124.570 ;
        RECT 81.210 122.890 81.470 123.210 ;
        RECT 81.270 121.850 81.410 122.890 ;
        RECT 83.110 121.850 83.250 125.270 ;
        RECT 83.510 123.230 83.770 123.550 ;
        RECT 83.570 122.870 83.710 123.230 ;
        RECT 83.510 122.550 83.770 122.870 ;
        RECT 79.430 121.620 80.030 121.760 ;
        RECT 78.910 121.190 79.170 121.510 ;
        RECT 79.370 120.850 79.630 121.170 ;
        RECT 79.430 119.130 79.570 120.850 ;
        RECT 78.450 118.810 78.710 119.130 ;
        RECT 79.370 118.810 79.630 119.130 ;
        RECT 79.890 118.110 80.030 121.620 ;
        RECT 81.210 121.530 81.470 121.850 ;
        RECT 83.050 121.530 83.310 121.850 ;
        RECT 80.290 118.470 80.550 118.790 ;
        RECT 79.830 117.790 80.090 118.110 ;
        RECT 77.990 117.450 78.250 117.770 ;
        RECT 79.830 117.110 80.090 117.430 ;
        RECT 79.890 116.410 80.030 117.110 ;
        RECT 79.830 116.090 80.090 116.410 ;
        RECT 77.530 115.750 77.790 116.070 ;
        RECT 77.590 85.470 77.730 115.750 ;
        RECT 79.370 115.410 79.630 115.730 ;
        RECT 77.990 111.670 78.250 111.990 ;
        RECT 78.050 110.630 78.190 111.670 ;
        RECT 77.990 110.310 78.250 110.630 ;
        RECT 79.430 110.290 79.570 115.410 ;
        RECT 80.350 112.670 80.490 118.470 ;
        RECT 82.130 117.790 82.390 118.110 ;
        RECT 81.670 117.110 81.930 117.430 ;
        RECT 81.730 113.010 81.870 117.110 ;
        RECT 82.190 113.690 82.330 117.790 ;
        RECT 82.590 117.110 82.850 117.430 ;
        RECT 82.650 114.710 82.790 117.110 ;
        RECT 82.590 114.390 82.850 114.710 ;
        RECT 82.130 113.370 82.390 113.690 ;
        RECT 81.670 112.690 81.930 113.010 ;
        RECT 80.290 112.350 80.550 112.670 ;
        RECT 79.370 109.970 79.630 110.290 ;
        RECT 80.750 106.910 81.010 107.230 ;
        RECT 79.830 106.230 80.090 106.550 ;
        RECT 79.370 93.650 79.630 93.970 ;
        RECT 78.450 92.630 78.710 92.950 ;
        RECT 78.510 91.930 78.650 92.630 ;
        RECT 78.450 91.610 78.710 91.930 ;
        RECT 79.430 90.085 79.570 93.650 ;
        RECT 79.360 89.715 79.640 90.085 ;
        RECT 79.430 89.210 79.570 89.715 ;
        RECT 79.370 88.890 79.630 89.210 ;
        RECT 78.910 88.210 79.170 88.530 ;
        RECT 78.450 87.190 78.710 87.510 ;
        RECT 78.510 86.490 78.650 87.190 ;
        RECT 78.450 86.170 78.710 86.490 ;
        RECT 78.970 85.470 79.110 88.210 ;
        RECT 77.530 85.150 77.790 85.470 ;
        RECT 78.910 85.150 79.170 85.470 ;
        RECT 79.370 85.150 79.630 85.470 ;
        RECT 77.530 84.470 77.790 84.790 ;
        RECT 77.990 84.470 78.250 84.790 ;
        RECT 77.590 82.070 77.730 84.470 ;
        RECT 78.050 83.430 78.190 84.470 ;
        RECT 77.990 83.110 78.250 83.430 ;
        RECT 78.910 82.770 79.170 83.090 ;
        RECT 77.530 81.750 77.790 82.070 ;
        RECT 77.590 79.690 77.730 81.750 ;
        RECT 77.530 79.370 77.790 79.690 ;
        RECT 76.610 79.030 76.870 79.350 ;
        RECT 73.850 78.010 74.110 78.330 ;
        RECT 73.390 77.730 73.650 77.990 ;
        RECT 73.390 77.670 74.510 77.730 ;
        RECT 73.450 77.590 74.510 77.670 ;
        RECT 78.970 77.650 79.110 82.770 ;
        RECT 79.430 81.050 79.570 85.150 ;
        RECT 79.890 83.090 80.030 106.230 ;
        RECT 80.810 102.130 80.950 106.910 ;
        RECT 83.570 102.570 83.710 122.550 ;
        RECT 83.970 120.850 84.230 121.170 ;
        RECT 84.030 119.130 84.170 120.850 ;
        RECT 83.970 118.810 84.230 119.130 ;
        RECT 84.490 117.430 84.630 134.790 ;
        RECT 84.890 131.730 85.150 132.050 ;
        RECT 84.950 130.010 85.090 131.730 ;
        RECT 84.890 129.690 85.150 130.010 ;
        RECT 85.410 128.990 85.550 137.850 ;
        RECT 87.250 134.430 87.390 142.610 ;
        RECT 88.110 142.270 88.370 142.590 ;
        RECT 87.650 139.210 87.910 139.530 ;
        RECT 87.190 134.110 87.450 134.430 ;
        RECT 87.710 132.390 87.850 139.210 ;
        RECT 87.650 132.070 87.910 132.390 ;
        RECT 87.190 130.710 87.450 131.030 ;
        RECT 87.250 128.990 87.390 130.710 ;
        RECT 85.350 128.670 85.610 128.990 ;
        RECT 85.810 128.670 86.070 128.990 ;
        RECT 87.190 128.670 87.450 128.990 ;
        RECT 85.410 123.890 85.550 128.670 ;
        RECT 85.350 123.570 85.610 123.890 ;
        RECT 85.410 122.870 85.550 123.570 ;
        RECT 85.350 122.550 85.610 122.870 ;
        RECT 85.410 118.450 85.550 122.550 ;
        RECT 85.350 118.130 85.610 118.450 ;
        RECT 84.430 117.110 84.690 117.430 ;
        RECT 84.490 112.670 84.630 117.110 ;
        RECT 84.430 112.350 84.690 112.670 ;
        RECT 84.890 111.670 85.150 111.990 ;
        RECT 84.950 110.970 85.090 111.670 ;
        RECT 84.890 110.650 85.150 110.970 ;
        RECT 84.890 108.950 85.150 109.270 ;
        RECT 84.950 107.230 85.090 108.950 ;
        RECT 85.350 107.590 85.610 107.910 ;
        RECT 84.890 106.910 85.150 107.230 ;
        RECT 84.430 106.230 84.690 106.550 ;
        RECT 82.650 102.430 83.710 102.570 ;
        RECT 80.750 101.810 81.010 102.130 ;
        RECT 81.670 101.470 81.930 101.790 ;
        RECT 82.650 101.700 82.790 102.430 ;
        RECT 83.970 102.150 84.230 102.470 ;
        RECT 83.050 101.700 83.310 101.790 ;
        RECT 82.650 101.560 83.310 101.700 ;
        RECT 83.050 101.470 83.310 101.560 ;
        RECT 81.730 96.350 81.870 101.470 ;
        RECT 82.590 100.790 82.850 101.110 ;
        RECT 82.130 98.750 82.390 99.070 ;
        RECT 81.670 96.030 81.930 96.350 ;
        RECT 81.730 93.970 81.870 96.030 ;
        RECT 82.190 94.310 82.330 98.750 ;
        RECT 82.650 96.690 82.790 100.790 ;
        RECT 84.030 100.090 84.170 102.150 ;
        RECT 84.490 100.090 84.630 106.230 ;
        RECT 84.950 104.850 85.090 106.910 ;
        RECT 85.410 106.550 85.550 107.590 ;
        RECT 85.350 106.230 85.610 106.550 ;
        RECT 85.410 104.850 85.550 106.230 ;
        RECT 84.890 104.530 85.150 104.850 ;
        RECT 85.350 104.530 85.610 104.850 ;
        RECT 84.950 101.450 85.090 104.530 ;
        RECT 85.350 103.510 85.610 103.830 ;
        RECT 84.890 101.130 85.150 101.450 ;
        RECT 83.970 99.770 84.230 100.090 ;
        RECT 84.430 99.770 84.690 100.090 ;
        RECT 84.490 97.030 84.630 99.770 ;
        RECT 84.430 96.710 84.690 97.030 ;
        RECT 82.590 96.370 82.850 96.690 ;
        RECT 83.050 96.370 83.310 96.690 ;
        RECT 82.650 94.650 82.790 96.370 ;
        RECT 82.590 94.330 82.850 94.650 ;
        RECT 82.130 93.990 82.390 94.310 ;
        RECT 81.670 93.650 81.930 93.970 ;
        RECT 82.590 93.880 82.850 93.970 ;
        RECT 83.110 93.880 83.250 96.370 ;
        RECT 83.970 95.690 84.230 96.010 ;
        RECT 82.590 93.740 83.250 93.880 ;
        RECT 82.590 93.650 82.850 93.740 ;
        RECT 80.750 93.310 81.010 93.630 ;
        RECT 80.810 89.210 80.950 93.310 ;
        RECT 81.670 92.630 81.930 92.950 ;
        RECT 80.750 88.890 81.010 89.210 ;
        RECT 80.290 87.190 80.550 87.510 ;
        RECT 80.350 86.490 80.490 87.190 ;
        RECT 80.290 86.170 80.550 86.490 ;
        RECT 81.730 83.090 81.870 92.630 ;
        RECT 83.050 90.930 83.310 91.250 ;
        RECT 82.130 90.590 82.390 90.910 ;
        RECT 82.190 87.850 82.330 90.590 ;
        RECT 82.590 88.210 82.850 88.530 ;
        RECT 82.130 87.530 82.390 87.850 ;
        RECT 82.650 85.810 82.790 88.210 ;
        RECT 83.110 85.810 83.250 90.930 ;
        RECT 83.510 88.210 83.770 88.530 ;
        RECT 83.570 87.850 83.710 88.210 ;
        RECT 83.510 87.530 83.770 87.850 ;
        RECT 82.590 85.490 82.850 85.810 ;
        RECT 83.050 85.490 83.310 85.810 ;
        RECT 83.570 85.130 83.710 87.530 ;
        RECT 83.510 84.810 83.770 85.130 ;
        RECT 79.830 82.770 80.090 83.090 ;
        RECT 81.210 82.770 81.470 83.090 ;
        RECT 81.670 82.770 81.930 83.090 ;
        RECT 82.590 82.770 82.850 83.090 ;
        RECT 80.290 81.750 80.550 82.070 ;
        RECT 79.370 80.730 79.630 81.050 ;
        RECT 79.830 80.730 80.090 81.050 ;
        RECT 79.890 80.450 80.030 80.730 ;
        RECT 79.430 80.310 80.030 80.450 ;
        RECT 79.430 79.350 79.570 80.310 ;
        RECT 80.350 80.030 80.490 81.750 ;
        RECT 80.290 79.710 80.550 80.030 ;
        RECT 80.750 79.370 81.010 79.690 ;
        RECT 79.370 79.030 79.630 79.350 ;
        RECT 80.290 79.030 80.550 79.350 ;
        RECT 80.350 77.990 80.490 79.030 ;
        RECT 80.290 77.670 80.550 77.990 ;
        RECT 72.290 75.775 73.830 76.145 ;
        RECT 74.370 75.270 74.510 77.590 ;
        RECT 76.150 77.330 76.410 77.650 ;
        RECT 78.910 77.330 79.170 77.650 ;
        RECT 74.770 76.310 75.030 76.630 ;
        RECT 74.310 74.950 74.570 75.270 ;
        RECT 74.830 74.930 74.970 76.310 ;
        RECT 74.770 74.610 75.030 74.930 ;
        RECT 72.930 74.270 73.190 74.590 ;
        RECT 69.710 73.930 69.970 74.250 ;
        RECT 71.550 73.930 71.810 74.250 ;
        RECT 68.790 72.570 69.050 72.890 ;
        RECT 68.330 68.490 68.590 68.810 ;
        RECT 68.390 67.450 68.530 68.490 ;
        RECT 68.330 67.130 68.590 67.450 ;
        RECT 67.410 66.110 67.670 66.430 ;
        RECT 65.570 65.430 65.830 65.750 ;
        RECT 66.030 63.390 66.290 63.710 ;
        RECT 64.650 61.350 64.910 61.670 ;
        RECT 61.430 61.010 61.690 61.330 ;
        RECT 60.050 60.670 60.310 60.990 ;
        RECT 60.110 59.290 60.250 60.670 ;
        RECT 60.050 58.970 60.310 59.290 ;
        RECT 61.430 58.180 61.690 58.270 ;
        RECT 61.430 58.040 62.090 58.180 ;
        RECT 61.430 57.950 61.690 58.040 ;
        RECT 61.950 56.200 62.090 58.040 ;
        RECT 64.710 56.200 64.850 61.350 ;
        RECT 66.090 58.610 66.230 63.390 ;
        RECT 66.490 61.240 66.750 61.330 ;
        RECT 66.490 61.100 67.610 61.240 ;
        RECT 66.490 61.010 66.750 61.100 ;
        RECT 66.030 58.290 66.290 58.610 ;
        RECT 67.470 56.200 67.610 61.100 ;
        RECT 68.330 58.180 68.590 58.270 ;
        RECT 68.850 58.180 68.990 72.570 ;
        RECT 69.770 69.490 69.910 73.930 ;
        RECT 72.990 72.210 73.130 74.270 ;
        RECT 75.230 73.590 75.490 73.910 ;
        RECT 73.850 72.570 74.110 72.890 ;
        RECT 73.910 72.405 74.050 72.570 ;
        RECT 71.090 71.890 71.350 72.210 ;
        RECT 72.930 71.890 73.190 72.210 ;
        RECT 73.840 72.035 74.120 72.405 ;
        RECT 71.150 70.170 71.290 71.890 ;
        RECT 72.290 70.335 73.830 70.705 ;
        RECT 71.090 69.850 71.350 70.170 ;
        RECT 73.390 69.740 73.650 69.830 ;
        RECT 73.390 69.600 74.510 69.740 ;
        RECT 73.390 69.510 73.650 69.600 ;
        RECT 69.710 69.170 69.970 69.490 ;
        RECT 73.850 68.830 74.110 69.150 ;
        RECT 70.170 68.150 70.430 68.470 ;
        RECT 69.250 61.240 69.510 61.330 ;
        RECT 70.230 61.240 70.370 68.150 ;
        RECT 73.910 67.450 74.050 68.830 ;
        RECT 73.850 67.130 74.110 67.450 ;
        RECT 70.630 65.770 70.890 66.090 ;
        RECT 70.690 63.710 70.830 65.770 ;
        RECT 71.550 65.430 71.810 65.750 ;
        RECT 71.610 64.730 71.750 65.430 ;
        RECT 72.290 64.895 73.830 65.265 ;
        RECT 71.550 64.410 71.810 64.730 ;
        RECT 70.630 63.390 70.890 63.710 ;
        RECT 73.850 63.620 74.110 63.710 ;
        RECT 74.370 63.620 74.510 69.600 ;
        RECT 75.290 69.150 75.430 73.590 ;
        RECT 76.210 69.150 76.350 77.330 ;
        RECT 78.970 74.590 79.110 77.330 ;
        RECT 80.290 77.220 80.550 77.310 ;
        RECT 80.810 77.220 80.950 79.370 ;
        RECT 81.270 78.330 81.410 82.770 ;
        RECT 81.210 78.010 81.470 78.330 ;
        RECT 80.290 77.080 80.950 77.220 ;
        RECT 80.290 76.990 80.550 77.080 ;
        RECT 80.350 74.590 80.490 76.990 ;
        RECT 78.910 74.270 79.170 74.590 ;
        RECT 80.290 74.270 80.550 74.590 ;
        RECT 76.610 71.550 76.870 71.870 ;
        RECT 75.230 68.830 75.490 69.150 ;
        RECT 76.150 68.830 76.410 69.150 ;
        RECT 76.670 68.810 76.810 71.550 ;
        RECT 78.970 71.530 79.110 74.270 ;
        RECT 80.350 72.890 80.490 74.270 ;
        RECT 80.290 72.570 80.550 72.890 ;
        RECT 78.910 71.210 79.170 71.530 ;
        RECT 77.070 70.870 77.330 71.190 ;
        RECT 81.210 70.870 81.470 71.190 ;
        RECT 76.610 68.490 76.870 68.810 ;
        RECT 74.770 68.150 75.030 68.470 ;
        RECT 74.830 66.090 74.970 68.150 ;
        RECT 76.670 67.450 76.810 68.490 ;
        RECT 76.610 67.130 76.870 67.450 ;
        RECT 77.130 66.770 77.270 70.870 ;
        RECT 79.370 69.850 79.630 70.170 ;
        RECT 79.430 66.770 79.570 69.850 ;
        RECT 81.270 68.070 81.410 70.870 ;
        RECT 81.730 69.150 81.870 82.770 ;
        RECT 82.650 77.650 82.790 82.770 ;
        RECT 83.510 81.750 83.770 82.070 ;
        RECT 83.570 80.030 83.710 81.750 ;
        RECT 83.510 79.710 83.770 80.030 ;
        RECT 82.590 77.330 82.850 77.650 ;
        RECT 84.030 77.310 84.170 95.690 ;
        RECT 84.430 93.310 84.690 93.630 ;
        RECT 84.490 91.930 84.630 93.310 ;
        RECT 84.430 91.610 84.690 91.930 ;
        RECT 84.890 90.590 85.150 90.910 ;
        RECT 84.950 90.085 85.090 90.590 ;
        RECT 84.880 89.715 85.160 90.085 ;
        RECT 84.430 88.550 84.690 88.870 ;
        RECT 84.490 86.490 84.630 88.550 ;
        RECT 84.430 86.170 84.690 86.490 ;
        RECT 84.430 82.770 84.690 83.090 ;
        RECT 84.490 81.050 84.630 82.770 ;
        RECT 84.890 82.430 85.150 82.750 ;
        RECT 84.950 81.050 85.090 82.430 ;
        RECT 84.430 80.730 84.690 81.050 ;
        RECT 84.890 80.730 85.150 81.050 ;
        RECT 85.410 80.030 85.550 103.510 ;
        RECT 85.870 101.790 86.010 128.670 ;
        RECT 87.710 128.310 87.850 132.070 ;
        RECT 87.650 127.990 87.910 128.310 ;
        RECT 87.710 123.290 87.850 127.990 ;
        RECT 88.170 127.290 88.310 142.270 ;
        RECT 88.630 136.470 88.770 142.610 ;
        RECT 89.090 139.530 89.230 142.610 ;
        RECT 89.490 141.590 89.750 141.910 ;
        RECT 89.550 140.210 89.690 141.590 ;
        RECT 90.010 140.210 90.150 142.950 ;
        RECT 90.930 140.890 91.070 144.650 ;
        RECT 90.870 140.570 91.130 140.890 ;
        RECT 89.490 139.890 89.750 140.210 ;
        RECT 89.950 139.890 90.210 140.210 ;
        RECT 91.390 139.870 91.530 147.030 ;
        RECT 91.850 143.610 91.990 156.210 ;
        RECT 91.790 143.290 92.050 143.610 ;
        RECT 91.330 139.550 91.590 139.870 ;
        RECT 89.030 139.210 89.290 139.530 ;
        RECT 89.080 138.335 90.620 138.705 ;
        RECT 90.410 137.170 90.670 137.490 ;
        RECT 88.570 136.150 88.830 136.470 ;
        RECT 90.470 135.450 90.610 137.170 ;
        RECT 90.410 135.130 90.670 135.450 ;
        RECT 89.080 132.895 90.620 133.265 ;
        RECT 91.330 131.960 91.590 132.050 ;
        RECT 92.310 131.960 92.450 156.550 ;
        RECT 92.770 152.790 92.910 166.410 ;
        RECT 93.230 165.370 93.370 166.750 ;
        RECT 93.170 165.050 93.430 165.370 ;
        RECT 93.230 161.970 93.370 165.050 ;
        RECT 93.170 161.650 93.430 161.970 ;
        RECT 94.090 156.890 94.350 157.210 ;
        RECT 94.150 155.510 94.290 156.890 ;
        RECT 93.170 155.190 93.430 155.510 ;
        RECT 93.630 155.190 93.890 155.510 ;
        RECT 94.090 155.190 94.350 155.510 ;
        RECT 93.230 154.490 93.370 155.190 ;
        RECT 93.170 154.170 93.430 154.490 ;
        RECT 93.170 153.150 93.430 153.470 ;
        RECT 92.710 152.470 92.970 152.790 ;
        RECT 93.230 148.030 93.370 153.150 ;
        RECT 93.690 151.770 93.830 155.190 ;
        RECT 94.610 153.380 94.750 177.720 ;
        RECT 95.930 176.950 96.190 177.270 ;
        RECT 95.990 176.250 96.130 176.950 ;
        RECT 96.450 176.250 96.590 185.450 ;
        RECT 97.830 184.410 97.970 186.130 ;
        RECT 97.770 184.090 98.030 184.410 ;
        RECT 97.310 181.030 97.570 181.350 ;
        RECT 96.850 179.670 97.110 179.990 ;
        RECT 95.930 175.930 96.190 176.250 ;
        RECT 96.390 175.930 96.650 176.250 ;
        RECT 96.910 175.570 97.050 179.670 ;
        RECT 97.370 176.250 97.510 181.030 ;
        RECT 98.290 179.990 98.430 186.470 ;
        RECT 99.610 185.790 99.870 186.110 ;
        RECT 99.150 182.730 99.410 183.050 ;
        RECT 98.230 179.670 98.490 179.990 ;
        RECT 98.690 179.670 98.950 179.990 ;
        RECT 98.750 178.970 98.890 179.670 ;
        RECT 97.770 178.650 98.030 178.970 ;
        RECT 98.690 178.650 98.950 178.970 ;
        RECT 97.830 178.485 97.970 178.650 ;
        RECT 97.760 178.115 98.040 178.485 ;
        RECT 98.230 176.950 98.490 177.270 ;
        RECT 97.310 175.930 97.570 176.250 ;
        RECT 95.010 175.250 95.270 175.570 ;
        RECT 96.850 175.250 97.110 175.570 ;
        RECT 97.770 175.250 98.030 175.570 ;
        RECT 95.070 171.830 95.210 175.250 ;
        RECT 97.310 174.910 97.570 175.230 ;
        RECT 95.930 174.230 96.190 174.550 ;
        RECT 95.990 173.190 96.130 174.230 ;
        RECT 95.930 172.870 96.190 173.190 ;
        RECT 97.370 172.510 97.510 174.910 ;
        RECT 97.830 173.530 97.970 175.250 ;
        RECT 97.770 173.210 98.030 173.530 ;
        RECT 97.310 172.190 97.570 172.510 ;
        RECT 95.010 171.510 95.270 171.830 ;
        RECT 97.370 170.810 97.510 172.190 ;
        RECT 97.310 170.490 97.570 170.810 ;
        RECT 95.010 168.790 95.270 169.110 ;
        RECT 95.070 167.070 95.210 168.790 ;
        RECT 95.010 166.750 95.270 167.070 ;
        RECT 95.930 158.930 96.190 159.250 ;
        RECT 95.470 157.910 95.730 158.230 ;
        RECT 94.150 153.240 94.750 153.380 ;
        RECT 93.630 151.450 93.890 151.770 ;
        RECT 92.710 147.710 92.970 148.030 ;
        RECT 93.170 147.710 93.430 148.030 ;
        RECT 91.330 131.820 92.450 131.960 ;
        RECT 91.330 131.730 91.590 131.820 ;
        RECT 89.030 131.390 89.290 131.710 ;
        RECT 89.090 130.010 89.230 131.390 ;
        RECT 89.490 130.710 89.750 131.030 ;
        RECT 89.030 129.690 89.290 130.010 ;
        RECT 89.550 129.330 89.690 130.710 ;
        RECT 92.770 129.670 92.910 147.710 ;
        RECT 94.150 142.330 94.290 153.240 ;
        RECT 95.010 152.470 95.270 152.790 ;
        RECT 95.530 152.530 95.670 157.910 ;
        RECT 95.990 154.490 96.130 158.930 ;
        RECT 98.290 157.290 98.430 176.950 ;
        RECT 99.210 173.530 99.350 182.730 ;
        RECT 99.670 177.270 99.810 185.790 ;
        RECT 102.890 185.770 103.030 189.790 ;
        RECT 103.350 185.770 103.490 192.250 ;
        RECT 103.810 192.130 104.030 192.270 ;
        RECT 104.270 192.270 104.410 193.360 ;
        RECT 104.270 192.130 104.870 192.270 ;
        RECT 103.810 186.450 103.950 192.130 ;
        RECT 104.730 191.890 104.870 192.130 ;
        RECT 104.670 191.570 104.930 191.890 ;
        RECT 105.190 191.290 105.330 199.030 ;
        RECT 105.650 196.310 105.790 200.410 ;
        RECT 107.950 199.370 108.090 201.430 ;
        RECT 107.890 199.050 108.150 199.370 ;
        RECT 107.890 197.010 108.150 197.330 ;
        RECT 105.590 195.990 105.850 196.310 ;
        RECT 105.870 195.455 107.410 195.825 ;
        RECT 105.590 193.950 105.850 194.270 ;
        RECT 104.270 191.150 105.330 191.290 ;
        RECT 103.750 186.130 104.010 186.450 ;
        RECT 104.270 185.850 104.410 191.150 ;
        RECT 104.670 190.550 104.930 190.870 ;
        RECT 105.650 190.780 105.790 193.950 ;
        RECT 106.050 193.445 106.310 193.590 ;
        RECT 106.040 193.075 106.320 193.445 ;
        RECT 107.950 192.765 108.090 197.010 ;
        RECT 106.040 192.395 106.320 192.765 ;
        RECT 107.880 192.395 108.160 192.765 ;
        RECT 106.050 192.250 106.310 192.395 ;
        RECT 105.190 190.640 105.790 190.780 ;
        RECT 104.730 189.850 104.870 190.550 ;
        RECT 104.670 189.530 104.930 189.850 ;
        RECT 102.830 185.450 103.090 185.770 ;
        RECT 103.290 185.450 103.550 185.770 ;
        RECT 103.810 185.710 104.410 185.850 ;
        RECT 101.450 182.730 101.710 183.050 ;
        RECT 101.510 178.970 101.650 182.730 ;
        RECT 101.910 180.690 102.170 181.010 ;
        RECT 101.970 178.970 102.110 180.690 ;
        RECT 103.290 179.670 103.550 179.990 ;
        RECT 101.450 178.650 101.710 178.970 ;
        RECT 101.910 178.650 102.170 178.970 ;
        RECT 101.450 177.630 101.710 177.950 ;
        RECT 99.610 176.950 99.870 177.270 ;
        RECT 101.510 176.250 101.650 177.630 ;
        RECT 101.450 175.930 101.710 176.250 ;
        RECT 101.970 175.230 102.110 178.650 ;
        RECT 103.350 178.290 103.490 179.670 ;
        RECT 102.830 177.970 103.090 178.290 ;
        RECT 103.290 177.970 103.550 178.290 ;
        RECT 102.890 176.250 103.030 177.970 ;
        RECT 103.810 177.690 103.950 185.710 ;
        RECT 104.210 185.110 104.470 185.430 ;
        RECT 104.270 181.690 104.410 185.110 ;
        RECT 105.190 183.730 105.330 190.640 ;
        RECT 105.870 190.015 107.410 190.385 ;
        RECT 107.430 188.510 107.690 188.830 ;
        RECT 106.970 188.170 107.230 188.490 ;
        RECT 107.030 186.110 107.170 188.170 ;
        RECT 107.490 187.130 107.630 188.510 ;
        RECT 107.430 186.810 107.690 187.130 ;
        RECT 106.970 185.790 107.230 186.110 ;
        RECT 107.890 185.450 108.150 185.770 ;
        RECT 105.870 184.575 107.410 184.945 ;
        RECT 105.130 183.410 105.390 183.730 ;
        RECT 104.210 181.370 104.470 181.690 ;
        RECT 103.350 177.550 103.950 177.690 ;
        RECT 102.830 175.930 103.090 176.250 ;
        RECT 101.910 174.910 102.170 175.230 ;
        RECT 99.150 173.210 99.410 173.530 ;
        RECT 102.830 170.490 103.090 170.810 ;
        RECT 102.890 167.410 103.030 170.490 ;
        RECT 102.830 167.090 103.090 167.410 ;
        RECT 103.350 166.390 103.490 177.550 ;
        RECT 103.750 175.250 104.010 175.570 ;
        RECT 103.290 166.070 103.550 166.390 ;
        RECT 102.830 165.050 103.090 165.370 ;
        RECT 102.890 164.690 103.030 165.050 ;
        RECT 102.830 164.370 103.090 164.690 ;
        RECT 103.290 164.370 103.550 164.690 ;
        RECT 100.530 164.030 100.790 164.350 ;
        RECT 101.450 164.030 101.710 164.350 ;
        RECT 98.690 163.350 98.950 163.670 ;
        RECT 98.750 158.140 98.890 163.350 ;
        RECT 100.590 160.950 100.730 164.030 ;
        RECT 100.990 163.350 101.250 163.670 ;
        RECT 101.050 162.310 101.190 163.350 ;
        RECT 101.510 162.310 101.650 164.030 ;
        RECT 103.350 162.650 103.490 164.370 ;
        RECT 103.290 162.330 103.550 162.650 ;
        RECT 100.990 161.990 101.250 162.310 ;
        RECT 101.450 161.990 101.710 162.310 ;
        RECT 100.530 160.630 100.790 160.950 ;
        RECT 99.610 158.250 99.870 158.570 ;
        RECT 99.150 158.140 99.410 158.230 ;
        RECT 98.750 158.000 99.410 158.140 ;
        RECT 99.150 157.910 99.410 158.000 ;
        RECT 98.290 157.150 98.890 157.290 ;
        RECT 96.390 155.190 96.650 155.510 ;
        RECT 95.930 154.170 96.190 154.490 ;
        RECT 96.450 154.150 96.590 155.190 ;
        RECT 97.770 154.400 98.030 154.490 ;
        RECT 97.770 154.260 98.430 154.400 ;
        RECT 97.770 154.170 98.030 154.260 ;
        RECT 96.390 153.830 96.650 154.150 ;
        RECT 95.070 151.430 95.210 152.470 ;
        RECT 95.530 152.390 97.050 152.530 ;
        RECT 96.390 151.450 96.650 151.770 ;
        RECT 94.540 150.915 94.820 151.285 ;
        RECT 95.010 151.110 95.270 151.430 ;
        RECT 95.930 151.110 96.190 151.430 ;
        RECT 94.610 150.410 94.750 150.915 ;
        RECT 94.550 150.090 94.810 150.410 ;
        RECT 94.550 148.390 94.810 148.710 ;
        RECT 93.230 142.190 94.290 142.330 ;
        RECT 93.230 134.285 93.370 142.190 ;
        RECT 93.630 141.590 93.890 141.910 ;
        RECT 93.690 139.530 93.830 141.590 ;
        RECT 93.630 139.210 93.890 139.530 ;
        RECT 94.090 138.870 94.350 139.190 ;
        RECT 93.160 133.915 93.440 134.285 ;
        RECT 94.150 134.090 94.290 138.870 ;
        RECT 94.610 134.770 94.750 148.390 ;
        RECT 95.070 145.650 95.210 151.110 ;
        RECT 95.470 149.750 95.730 150.070 ;
        RECT 95.530 146.330 95.670 149.750 ;
        RECT 95.470 146.010 95.730 146.330 ;
        RECT 95.010 145.330 95.270 145.650 ;
        RECT 95.530 144.970 95.670 146.010 ;
        RECT 95.990 144.970 96.130 151.110 ;
        RECT 95.470 144.650 95.730 144.970 ;
        RECT 95.930 144.650 96.190 144.970 ;
        RECT 95.530 143.610 95.670 144.650 ;
        RECT 95.470 143.290 95.730 143.610 ;
        RECT 95.990 142.930 96.130 144.650 ;
        RECT 96.450 143.610 96.590 151.450 ;
        RECT 96.910 151.090 97.050 152.390 ;
        RECT 96.850 150.770 97.110 151.090 ;
        RECT 96.910 148.370 97.050 150.770 ;
        RECT 97.310 150.430 97.570 150.750 ;
        RECT 97.770 150.430 98.030 150.750 ;
        RECT 96.850 148.050 97.110 148.370 ;
        RECT 97.370 145.310 97.510 150.430 ;
        RECT 97.830 149.050 97.970 150.430 ;
        RECT 97.770 148.730 98.030 149.050 ;
        RECT 97.310 144.990 97.570 145.310 ;
        RECT 96.390 143.290 96.650 143.610 ;
        RECT 95.930 142.610 96.190 142.930 ;
        RECT 96.390 142.160 96.650 142.250 ;
        RECT 95.530 142.020 96.650 142.160 ;
        RECT 95.010 140.570 95.270 140.890 ;
        RECT 95.070 140.210 95.210 140.570 ;
        RECT 95.010 139.890 95.270 140.210 ;
        RECT 95.070 137.570 95.210 139.890 ;
        RECT 95.530 138.170 95.670 142.020 ;
        RECT 96.390 141.930 96.650 142.020 ;
        RECT 95.470 137.850 95.730 138.170 ;
        RECT 95.070 137.430 95.670 137.570 ;
        RECT 94.550 134.450 94.810 134.770 ;
        RECT 94.090 133.770 94.350 134.090 ;
        RECT 94.090 130.710 94.350 131.030 ;
        RECT 93.630 129.690 93.890 130.010 ;
        RECT 90.410 129.350 90.670 129.670 ;
        RECT 92.710 129.350 92.970 129.670 ;
        RECT 89.490 129.010 89.750 129.330 ;
        RECT 90.470 128.650 90.610 129.350 ;
        RECT 91.790 128.670 92.050 128.990 ;
        RECT 90.410 128.330 90.670 128.650 ;
        RECT 89.080 127.455 90.620 127.825 ;
        RECT 88.110 126.970 88.370 127.290 ;
        RECT 91.850 123.890 91.990 128.670 ;
        RECT 92.770 124.650 92.910 129.350 ;
        RECT 93.690 128.990 93.830 129.690 ;
        RECT 93.630 128.670 93.890 128.990 ;
        RECT 94.150 127.290 94.290 130.710 ;
        RECT 94.550 128.670 94.810 128.990 ;
        RECT 94.090 126.970 94.350 127.290 ;
        RECT 94.610 126.610 94.750 128.670 ;
        RECT 94.550 126.290 94.810 126.610 ;
        RECT 93.170 125.500 93.430 125.590 ;
        RECT 93.170 125.360 93.830 125.500 ;
        RECT 93.170 125.270 93.430 125.360 ;
        RECT 92.770 124.510 93.370 124.650 ;
        RECT 91.790 123.570 92.050 123.890 ;
        RECT 87.710 123.150 88.770 123.290 ;
        RECT 92.710 123.230 92.970 123.550 ;
        RECT 88.110 122.550 88.370 122.870 ;
        RECT 88.170 120.150 88.310 122.550 ;
        RECT 88.630 121.760 88.770 123.150 ;
        RECT 90.870 122.550 91.130 122.870 ;
        RECT 91.330 122.550 91.590 122.870 ;
        RECT 92.250 122.550 92.510 122.870 ;
        RECT 89.080 122.015 90.620 122.385 ;
        RECT 88.630 121.620 89.230 121.760 ;
        RECT 88.110 119.830 88.370 120.150 ;
        RECT 86.730 114.390 86.990 114.710 ;
        RECT 86.270 106.230 86.530 106.550 ;
        RECT 86.330 104.850 86.470 106.230 ;
        RECT 86.790 104.850 86.930 114.390 ;
        RECT 88.170 107.230 88.310 119.830 ;
        RECT 89.090 118.450 89.230 121.620 ;
        RECT 89.490 120.510 89.750 120.830 ;
        RECT 89.030 118.130 89.290 118.450 ;
        RECT 89.090 117.340 89.230 118.130 ;
        RECT 89.550 117.770 89.690 120.510 ;
        RECT 90.930 118.450 91.070 122.550 ;
        RECT 91.390 121.170 91.530 122.550 ;
        RECT 92.310 121.850 92.450 122.550 ;
        RECT 92.250 121.530 92.510 121.850 ;
        RECT 91.330 120.850 91.590 121.170 ;
        RECT 90.870 118.130 91.130 118.450 ;
        RECT 89.490 117.450 89.750 117.770 ;
        RECT 88.630 117.200 89.230 117.340 ;
        RECT 88.630 113.690 88.770 117.200 ;
        RECT 89.080 116.575 90.620 116.945 ;
        RECT 92.310 115.640 92.450 121.530 ;
        RECT 92.770 119.130 92.910 123.230 ;
        RECT 92.710 118.810 92.970 119.130 ;
        RECT 92.710 115.640 92.970 115.730 ;
        RECT 92.310 115.500 92.970 115.640 ;
        RECT 92.710 115.410 92.970 115.500 ;
        RECT 91.790 114.390 92.050 114.710 ;
        RECT 88.570 113.370 88.830 113.690 ;
        RECT 90.870 112.010 91.130 112.330 ;
        RECT 91.330 112.010 91.590 112.330 ;
        RECT 89.080 111.135 90.620 111.505 ;
        RECT 90.930 110.970 91.070 112.010 ;
        RECT 90.870 110.650 91.130 110.970 ;
        RECT 91.390 110.290 91.530 112.010 ;
        RECT 90.870 109.970 91.130 110.290 ;
        RECT 91.330 109.970 91.590 110.290 ;
        RECT 88.110 106.910 88.370 107.230 ;
        RECT 87.190 106.570 87.450 106.890 ;
        RECT 87.250 105.530 87.390 106.570 ;
        RECT 89.080 105.695 90.620 106.065 ;
        RECT 87.190 105.210 87.450 105.530 ;
        RECT 90.930 104.850 91.070 109.970 ;
        RECT 91.330 108.950 91.590 109.270 ;
        RECT 91.390 104.850 91.530 108.950 ;
        RECT 86.270 104.530 86.530 104.850 ;
        RECT 86.730 104.530 86.990 104.850 ;
        RECT 90.870 104.530 91.130 104.850 ;
        RECT 91.330 104.530 91.590 104.850 ;
        RECT 90.930 101.790 91.070 104.530 ;
        RECT 91.850 101.790 91.990 114.390 ;
        RECT 92.250 112.350 92.510 112.670 ;
        RECT 92.310 104.510 92.450 112.350 ;
        RECT 92.770 110.970 92.910 115.410 ;
        RECT 92.710 110.650 92.970 110.970 ;
        RECT 92.710 105.210 92.970 105.530 ;
        RECT 92.250 104.190 92.510 104.510 ;
        RECT 92.250 103.510 92.510 103.830 ;
        RECT 92.310 101.790 92.450 103.510 ;
        RECT 85.810 101.470 86.070 101.790 ;
        RECT 90.870 101.470 91.130 101.790 ;
        RECT 91.790 101.470 92.050 101.790 ;
        RECT 92.250 101.470 92.510 101.790 ;
        RECT 92.770 101.530 92.910 105.210 ;
        RECT 93.230 102.210 93.370 124.510 ;
        RECT 93.690 123.890 93.830 125.360 ;
        RECT 94.090 123.910 94.350 124.230 ;
        RECT 93.630 123.570 93.890 123.890 ;
        RECT 93.690 121.170 93.830 123.570 ;
        RECT 93.630 120.850 93.890 121.170 ;
        RECT 93.690 116.410 93.830 120.850 ;
        RECT 93.630 116.090 93.890 116.410 ;
        RECT 93.690 113.010 93.830 116.090 ;
        RECT 94.150 115.730 94.290 123.910 ;
        RECT 95.010 122.550 95.270 122.870 ;
        RECT 95.070 118.110 95.210 122.550 ;
        RECT 95.010 117.790 95.270 118.110 ;
        RECT 95.530 117.770 95.670 137.430 ;
        RECT 96.850 137.170 97.110 137.490 ;
        RECT 96.390 136.150 96.650 136.470 ;
        RECT 96.450 134.430 96.590 136.150 ;
        RECT 96.390 134.110 96.650 134.430 ;
        RECT 95.930 131.730 96.190 132.050 ;
        RECT 95.990 130.010 96.130 131.730 ;
        RECT 95.930 129.690 96.190 130.010 ;
        RECT 96.910 129.330 97.050 137.170 ;
        RECT 97.770 135.130 98.030 135.450 ;
        RECT 97.310 134.285 97.570 134.430 ;
        RECT 97.300 133.915 97.580 134.285 ;
        RECT 97.310 133.430 97.570 133.750 ;
        RECT 97.370 132.390 97.510 133.430 ;
        RECT 97.310 132.070 97.570 132.390 ;
        RECT 97.830 131.710 97.970 135.130 ;
        RECT 98.290 132.730 98.430 154.260 ;
        RECT 98.750 134.770 98.890 157.150 ;
        RECT 99.210 155.850 99.350 157.910 ;
        RECT 99.670 155.850 99.810 158.250 ;
        RECT 99.150 155.530 99.410 155.850 ;
        RECT 99.610 155.530 99.870 155.850 ;
        RECT 99.210 151.090 99.350 155.530 ;
        RECT 100.070 153.490 100.330 153.810 ;
        RECT 100.130 151.770 100.270 153.490 ;
        RECT 100.530 152.470 100.790 152.790 ;
        RECT 100.070 151.450 100.330 151.770 ;
        RECT 99.150 150.770 99.410 151.090 ;
        RECT 100.590 150.750 100.730 152.470 ;
        RECT 100.530 150.430 100.790 150.750 ;
        RECT 101.050 146.330 101.190 161.990 ;
        RECT 101.510 159.930 101.650 161.990 ;
        RECT 103.810 160.860 103.950 175.250 ;
        RECT 104.270 164.690 104.410 181.370 ;
        RECT 105.130 180.690 105.390 181.010 ;
        RECT 104.670 180.350 104.930 180.670 ;
        RECT 104.730 175.570 104.870 180.350 ;
        RECT 105.190 175.570 105.330 180.690 ;
        RECT 105.870 179.135 107.410 179.505 ;
        RECT 107.950 178.370 108.090 185.450 ;
        RECT 107.490 178.230 108.090 178.370 ;
        RECT 106.970 177.630 107.230 177.950 ;
        RECT 106.050 176.950 106.310 177.270 ;
        RECT 106.510 176.950 106.770 177.270 ;
        RECT 106.110 176.250 106.250 176.950 ;
        RECT 106.570 176.250 106.710 176.950 ;
        RECT 107.030 176.250 107.170 177.630 ;
        RECT 106.050 175.930 106.310 176.250 ;
        RECT 106.510 175.930 106.770 176.250 ;
        RECT 106.970 175.930 107.230 176.250 ;
        RECT 107.490 175.570 107.630 178.230 ;
        RECT 108.410 177.690 108.550 206.960 ;
        RECT 108.810 206.870 109.070 206.960 ;
        RECT 110.250 200.730 110.390 207.890 ;
        RECT 115.310 207.870 115.450 212.200 ;
        RECT 122.670 210.330 122.810 212.200 ;
        RECT 122.210 210.190 122.810 210.330 ;
        RECT 117.090 209.590 117.350 209.910 ;
        RECT 117.150 208.210 117.290 209.590 ;
        RECT 118.010 208.230 118.270 208.550 ;
        RECT 118.470 208.290 118.730 208.550 ;
        RECT 118.470 208.230 119.130 208.290 ;
        RECT 117.090 207.890 117.350 208.210 ;
        RECT 115.250 207.550 115.510 207.870 ;
        RECT 110.650 207.210 110.910 207.530 ;
        RECT 110.710 205.150 110.850 207.210 ;
        RECT 111.110 206.870 111.370 207.190 ;
        RECT 110.650 204.830 110.910 205.150 ;
        RECT 111.170 203.110 111.310 206.870 ;
        RECT 117.150 205.570 117.290 207.890 ;
        RECT 117.550 206.870 117.810 207.190 ;
        RECT 116.690 205.430 117.290 205.570 ;
        RECT 111.110 202.790 111.370 203.110 ;
        RECT 114.790 202.790 115.050 203.110 ;
        RECT 114.850 202.285 114.990 202.790 ;
        RECT 114.780 201.915 115.060 202.285 ;
        RECT 116.170 202.110 116.430 202.430 ;
        RECT 110.650 201.430 110.910 201.750 ;
        RECT 115.710 201.430 115.970 201.750 ;
        RECT 110.190 200.410 110.450 200.730 ;
        RECT 110.710 199.710 110.850 201.430 ;
        RECT 115.770 199.710 115.910 201.430 ;
        RECT 116.230 199.710 116.370 202.110 ;
        RECT 116.690 200.730 116.830 205.430 ;
        RECT 117.090 204.830 117.350 205.150 ;
        RECT 117.150 202.680 117.290 204.830 ;
        RECT 117.610 204.810 117.750 206.870 ;
        RECT 117.550 204.490 117.810 204.810 ;
        RECT 117.550 202.680 117.810 202.770 ;
        RECT 117.150 202.540 117.810 202.680 ;
        RECT 117.550 202.450 117.810 202.540 ;
        RECT 116.630 200.410 116.890 200.730 ;
        RECT 116.690 199.710 116.830 200.410 ;
        RECT 110.650 199.390 110.910 199.710 ;
        RECT 113.410 199.390 113.670 199.710 ;
        RECT 115.710 199.390 115.970 199.710 ;
        RECT 116.170 199.390 116.430 199.710 ;
        RECT 116.630 199.390 116.890 199.710 ;
        RECT 111.110 199.050 111.370 199.370 ;
        RECT 108.810 193.950 109.070 194.270 ;
        RECT 108.870 192.570 109.010 193.950 ;
        RECT 108.810 192.250 109.070 192.570 ;
        RECT 108.810 190.550 109.070 190.870 ;
        RECT 110.190 190.550 110.450 190.870 ;
        RECT 108.870 181.010 109.010 190.550 ;
        RECT 110.250 189.850 110.390 190.550 ;
        RECT 110.190 189.530 110.450 189.850 ;
        RECT 109.270 189.190 109.530 189.510 ;
        RECT 109.330 188.060 109.470 189.190 ;
        RECT 109.730 188.060 109.990 188.150 ;
        RECT 109.330 187.920 109.990 188.060 ;
        RECT 109.330 183.390 109.470 187.920 ;
        RECT 109.730 187.830 109.990 187.920 ;
        RECT 109.730 185.110 109.990 185.430 ;
        RECT 110.650 185.110 110.910 185.430 ;
        RECT 109.790 184.410 109.930 185.110 ;
        RECT 109.730 184.090 109.990 184.410 ;
        RECT 109.270 183.070 109.530 183.390 ;
        RECT 109.790 181.690 109.930 184.090 ;
        RECT 110.710 183.390 110.850 185.110 ;
        RECT 110.650 183.070 110.910 183.390 ;
        RECT 109.730 181.370 109.990 181.690 ;
        RECT 108.810 180.690 109.070 181.010 ;
        RECT 110.650 179.670 110.910 179.990 ;
        RECT 110.710 177.950 110.850 179.670 ;
        RECT 107.950 177.550 108.550 177.690 ;
        RECT 110.650 177.630 110.910 177.950 ;
        RECT 104.670 175.250 104.930 175.570 ;
        RECT 105.130 175.250 105.390 175.570 ;
        RECT 107.430 175.250 107.690 175.570 ;
        RECT 104.730 170.810 104.870 175.250 ;
        RECT 105.870 173.695 107.410 174.065 ;
        RECT 104.670 170.490 104.930 170.810 ;
        RECT 105.130 170.150 105.390 170.470 ;
        RECT 105.190 168.090 105.330 170.150 ;
        RECT 105.870 168.255 107.410 168.625 ;
        RECT 105.130 167.770 105.390 168.090 ;
        RECT 106.970 166.750 107.230 167.070 ;
        RECT 105.130 166.070 105.390 166.390 ;
        RECT 104.210 164.370 104.470 164.690 ;
        RECT 104.210 160.860 104.470 160.950 ;
        RECT 103.810 160.720 104.470 160.860 ;
        RECT 104.210 160.630 104.470 160.720 ;
        RECT 101.450 159.610 101.710 159.930 ;
        RECT 103.290 158.930 103.550 159.250 ;
        RECT 103.350 158.570 103.490 158.930 ;
        RECT 103.290 158.250 103.550 158.570 ;
        RECT 102.370 149.750 102.630 150.070 ;
        RECT 102.430 149.050 102.570 149.750 ;
        RECT 102.370 148.730 102.630 149.050 ;
        RECT 100.990 146.010 101.250 146.330 ;
        RECT 102.830 142.270 103.090 142.590 ;
        RECT 99.610 141.590 99.870 141.910 ;
        RECT 101.450 141.590 101.710 141.910 ;
        RECT 99.670 138.170 99.810 141.590 ;
        RECT 101.510 140.890 101.650 141.590 ;
        RECT 101.450 140.570 101.710 140.890 ;
        RECT 102.370 140.230 102.630 140.550 ;
        RECT 100.520 139.355 100.800 139.725 ;
        RECT 100.530 139.210 100.790 139.355 ;
        RECT 101.450 138.870 101.710 139.190 ;
        RECT 99.610 137.850 99.870 138.170 ;
        RECT 98.690 134.450 98.950 134.770 ;
        RECT 100.990 134.110 101.250 134.430 ;
        RECT 101.050 132.730 101.190 134.110 ;
        RECT 98.230 132.410 98.490 132.730 ;
        RECT 99.610 132.410 99.870 132.730 ;
        RECT 100.990 132.410 101.250 132.730 ;
        RECT 97.770 131.390 98.030 131.710 ;
        RECT 97.770 129.350 98.030 129.670 ;
        RECT 96.850 129.010 97.110 129.330 ;
        RECT 96.390 128.330 96.650 128.650 ;
        RECT 96.450 127.290 96.590 128.330 ;
        RECT 96.390 126.970 96.650 127.290 ;
        RECT 97.310 123.230 97.570 123.550 ;
        RECT 97.370 121.850 97.510 123.230 ;
        RECT 97.310 121.530 97.570 121.850 ;
        RECT 95.930 120.510 96.190 120.830 ;
        RECT 95.470 117.450 95.730 117.770 ;
        RECT 95.990 117.430 96.130 120.510 ;
        RECT 95.930 117.110 96.190 117.430 ;
        RECT 94.090 115.410 94.350 115.730 ;
        RECT 93.630 112.690 93.890 113.010 ;
        RECT 94.150 109.610 94.290 115.410 ;
        RECT 95.010 112.010 95.270 112.330 ;
        RECT 95.070 110.970 95.210 112.010 ;
        RECT 95.470 111.670 95.730 111.990 ;
        RECT 95.530 110.970 95.670 111.670 ;
        RECT 95.010 110.650 95.270 110.970 ;
        RECT 95.470 110.650 95.730 110.970 ;
        RECT 94.090 109.290 94.350 109.610 ;
        RECT 94.550 106.910 94.810 107.230 ;
        RECT 93.630 106.230 93.890 106.550 ;
        RECT 93.690 105.190 93.830 106.230 ;
        RECT 93.630 104.870 93.890 105.190 ;
        RECT 94.610 102.810 94.750 106.910 ;
        RECT 95.930 106.230 96.190 106.550 ;
        RECT 97.310 106.230 97.570 106.550 ;
        RECT 94.550 102.490 94.810 102.810 ;
        RECT 93.230 102.070 95.210 102.210 ;
        RECT 89.080 100.255 90.620 100.625 ;
        RECT 90.410 99.770 90.670 100.090 ;
        RECT 85.810 99.090 86.070 99.410 ;
        RECT 86.730 99.090 86.990 99.410 ;
        RECT 88.570 99.090 88.830 99.410 ;
        RECT 85.870 96.350 86.010 99.090 ;
        RECT 85.810 96.030 86.070 96.350 ;
        RECT 86.790 95.670 86.930 99.090 ;
        RECT 87.650 98.070 87.910 98.390 ;
        RECT 86.730 95.350 86.990 95.670 ;
        RECT 87.710 83.430 87.850 98.070 ;
        RECT 88.630 96.010 88.770 99.090 ;
        RECT 90.470 96.940 90.610 99.770 ;
        RECT 90.930 99.410 91.070 101.470 ;
        RECT 92.310 99.410 92.450 101.470 ;
        RECT 92.770 101.390 94.290 101.530 ;
        RECT 93.170 100.790 93.430 101.110 ;
        RECT 90.870 99.090 91.130 99.410 ;
        RECT 92.250 99.090 92.510 99.410 ;
        RECT 91.330 98.070 91.590 98.390 ;
        RECT 90.470 96.800 91.070 96.940 ;
        RECT 88.570 95.690 88.830 96.010 ;
        RECT 88.110 95.350 88.370 95.670 ;
        RECT 88.170 91.930 88.310 95.350 ;
        RECT 89.080 94.815 90.620 95.185 ;
        RECT 90.930 94.650 91.070 96.800 ;
        RECT 90.870 94.330 91.130 94.650 ;
        RECT 90.870 92.630 91.130 92.950 ;
        RECT 88.110 91.610 88.370 91.930 ;
        RECT 89.080 89.375 90.620 89.745 ;
        RECT 90.410 86.170 90.670 86.490 ;
        RECT 88.570 85.150 88.830 85.470 ;
        RECT 90.470 85.325 90.610 86.170 ;
        RECT 88.630 83.430 88.770 85.150 ;
        RECT 90.400 84.955 90.680 85.325 ;
        RECT 89.080 83.935 90.620 84.305 ;
        RECT 90.930 83.770 91.070 92.630 ;
        RECT 91.390 84.790 91.530 98.070 ;
        RECT 91.790 96.710 92.050 97.030 ;
        RECT 91.850 87.930 91.990 96.710 ;
        RECT 92.310 96.350 92.450 99.090 ;
        RECT 92.250 96.030 92.510 96.350 ;
        RECT 92.310 93.880 92.450 96.030 ;
        RECT 92.710 93.880 92.970 93.970 ;
        RECT 92.310 93.740 92.970 93.880 ;
        RECT 92.710 93.650 92.970 93.740 ;
        RECT 92.710 92.970 92.970 93.290 ;
        RECT 92.770 91.930 92.910 92.970 ;
        RECT 92.710 91.610 92.970 91.930 ;
        RECT 92.250 90.590 92.510 90.910 ;
        RECT 92.310 89.210 92.450 90.590 ;
        RECT 92.250 88.890 92.510 89.210 ;
        RECT 93.230 87.930 93.370 100.790 ;
        RECT 93.630 98.070 93.890 98.390 ;
        RECT 93.690 96.690 93.830 98.070 ;
        RECT 93.630 96.370 93.890 96.690 ;
        RECT 94.150 94.560 94.290 101.390 ;
        RECT 94.550 99.090 94.810 99.410 ;
        RECT 94.610 96.350 94.750 99.090 ;
        RECT 94.550 96.030 94.810 96.350 ;
        RECT 94.610 94.650 94.750 96.030 ;
        RECT 95.070 95.670 95.210 102.070 ;
        RECT 95.990 101.790 96.130 106.230 ;
        RECT 97.370 103.830 97.510 106.230 ;
        RECT 97.830 104.510 97.970 129.350 ;
        RECT 98.690 118.130 98.950 118.450 ;
        RECT 98.230 116.090 98.490 116.410 ;
        RECT 98.290 115.730 98.430 116.090 ;
        RECT 98.230 115.410 98.490 115.730 ;
        RECT 98.750 113.010 98.890 118.130 ;
        RECT 99.150 117.110 99.410 117.430 ;
        RECT 99.210 116.410 99.350 117.110 ;
        RECT 99.150 116.090 99.410 116.410 ;
        RECT 98.690 112.690 98.950 113.010 ;
        RECT 98.230 106.910 98.490 107.230 ;
        RECT 97.770 104.190 98.030 104.510 ;
        RECT 97.310 103.510 97.570 103.830 ;
        RECT 95.930 101.470 96.190 101.790 ;
        RECT 96.850 100.790 97.110 101.110 ;
        RECT 96.910 99.070 97.050 100.790 ;
        RECT 97.370 99.410 97.510 103.510 ;
        RECT 98.290 99.410 98.430 106.910 ;
        RECT 98.750 104.510 98.890 112.690 ;
        RECT 99.670 105.530 99.810 132.410 ;
        RECT 101.050 129.330 101.190 132.410 ;
        RECT 100.990 129.010 101.250 129.330 ;
        RECT 101.510 118.450 101.650 138.870 ;
        RECT 102.430 138.170 102.570 140.230 ;
        RECT 102.370 137.850 102.630 138.170 ;
        RECT 102.430 135.450 102.570 137.850 ;
        RECT 102.370 135.130 102.630 135.450 ;
        RECT 102.370 125.270 102.630 125.590 ;
        RECT 102.430 121.850 102.570 125.270 ;
        RECT 102.370 121.530 102.630 121.850 ;
        RECT 101.450 118.130 101.710 118.450 ;
        RECT 100.990 117.790 101.250 118.110 ;
        RECT 101.050 116.410 101.190 117.790 ;
        RECT 100.990 116.090 101.250 116.410 ;
        RECT 102.890 112.670 103.030 142.270 ;
        RECT 103.350 139.870 103.490 158.250 ;
        RECT 104.270 156.530 104.410 160.630 ;
        RECT 104.210 156.210 104.470 156.530 ;
        RECT 104.670 153.490 104.930 153.810 ;
        RECT 104.730 151.770 104.870 153.490 ;
        RECT 104.670 151.450 104.930 151.770 ;
        RECT 105.190 148.960 105.330 166.070 ;
        RECT 107.030 164.010 107.170 166.750 ;
        RECT 106.970 163.690 107.230 164.010 ;
        RECT 105.870 162.815 107.410 163.185 ;
        RECT 105.870 157.375 107.410 157.745 ;
        RECT 105.870 151.935 107.410 152.305 ;
        RECT 107.950 150.750 108.090 177.550 ;
        RECT 109.270 169.810 109.530 170.130 ;
        RECT 109.330 168.090 109.470 169.810 ;
        RECT 109.730 169.470 109.990 169.790 ;
        RECT 109.270 167.770 109.530 168.090 ;
        RECT 109.270 166.750 109.530 167.070 ;
        RECT 108.350 166.070 108.610 166.390 ;
        RECT 108.410 165.370 108.550 166.070 ;
        RECT 108.350 165.050 108.610 165.370 ;
        RECT 108.410 156.190 108.550 165.050 ;
        RECT 108.810 164.600 109.070 164.690 ;
        RECT 109.330 164.600 109.470 166.750 ;
        RECT 108.810 164.460 109.470 164.600 ;
        RECT 108.810 164.370 109.070 164.460 ;
        RECT 108.350 155.870 108.610 156.190 ;
        RECT 108.870 156.100 109.010 164.370 ;
        RECT 109.270 163.350 109.530 163.670 ;
        RECT 109.330 159.930 109.470 163.350 ;
        RECT 109.790 161.630 109.930 169.470 ;
        RECT 111.170 167.410 111.310 199.050 ;
        RECT 113.470 198.010 113.610 199.390 ;
        RECT 114.330 198.710 114.590 199.030 ;
        RECT 113.410 197.690 113.670 198.010 ;
        RECT 114.390 197.670 114.530 198.710 ;
        RECT 114.330 197.350 114.590 197.670 ;
        RECT 117.610 196.990 117.750 202.450 ;
        RECT 118.070 201.750 118.210 208.230 ;
        RECT 118.530 208.150 119.130 208.230 ;
        RECT 118.470 202.450 118.730 202.770 ;
        RECT 118.010 201.430 118.270 201.750 ;
        RECT 118.530 200.730 118.670 202.450 ;
        RECT 118.470 200.410 118.730 200.730 ;
        RECT 118.010 200.070 118.270 200.390 ;
        RECT 118.990 200.130 119.130 208.150 ;
        RECT 120.310 207.100 120.570 207.190 ;
        RECT 118.070 197.330 118.210 200.070 ;
        RECT 118.530 199.990 119.130 200.130 ;
        RECT 119.450 206.960 120.570 207.100 ;
        RECT 118.010 197.010 118.270 197.330 ;
        RECT 117.550 196.670 117.810 196.990 ;
        RECT 118.530 196.730 118.670 199.990 ;
        RECT 118.930 199.390 119.190 199.710 ;
        RECT 117.610 193.590 117.750 196.670 ;
        RECT 118.070 196.590 118.670 196.730 ;
        RECT 111.570 193.270 111.830 193.590 ;
        RECT 112.490 193.270 112.750 193.590 ;
        RECT 117.550 193.270 117.810 193.590 ;
        RECT 111.630 189.850 111.770 193.270 ;
        RECT 112.550 192.230 112.690 193.270 ;
        RECT 112.490 191.910 112.750 192.230 ;
        RECT 117.610 191.890 117.750 193.270 ;
        RECT 116.630 191.570 116.890 191.890 ;
        RECT 117.550 191.570 117.810 191.890 ;
        RECT 112.030 190.890 112.290 191.210 ;
        RECT 112.090 189.850 112.230 190.890 ;
        RECT 116.690 189.850 116.830 191.570 ;
        RECT 111.570 189.530 111.830 189.850 ;
        RECT 112.030 189.530 112.290 189.850 ;
        RECT 116.630 189.530 116.890 189.850 ;
        RECT 117.610 189.170 117.750 191.570 ;
        RECT 117.550 188.850 117.810 189.170 ;
        RECT 112.490 188.510 112.750 188.830 ;
        RECT 112.030 185.110 112.290 185.430 ;
        RECT 112.090 183.730 112.230 185.110 ;
        RECT 112.550 184.410 112.690 188.510 ;
        RECT 113.410 187.830 113.670 188.150 ;
        RECT 113.470 187.130 113.610 187.830 ;
        RECT 117.610 187.130 117.750 188.850 ;
        RECT 113.410 186.810 113.670 187.130 ;
        RECT 117.550 186.810 117.810 187.130 ;
        RECT 117.550 186.130 117.810 186.450 ;
        RECT 117.610 184.410 117.750 186.130 ;
        RECT 112.490 184.090 112.750 184.410 ;
        RECT 117.550 184.090 117.810 184.410 ;
        RECT 118.070 183.810 118.210 196.590 ;
        RECT 118.990 191.890 119.130 199.390 ;
        RECT 118.930 191.570 119.190 191.890 ;
        RECT 118.990 191.290 119.130 191.570 ;
        RECT 112.030 183.410 112.290 183.730 ;
        RECT 117.610 183.670 118.210 183.810 ;
        RECT 118.530 191.150 119.130 191.290 ;
        RECT 111.570 181.030 111.830 181.350 ;
        RECT 111.630 175.570 111.770 181.030 ;
        RECT 112.090 175.570 112.230 183.410 ;
        RECT 112.490 176.950 112.750 177.270 ;
        RECT 112.550 176.250 112.690 176.950 ;
        RECT 112.490 175.930 112.750 176.250 ;
        RECT 111.570 175.250 111.830 175.570 ;
        RECT 112.030 175.250 112.290 175.570 ;
        RECT 112.030 174.230 112.290 174.550 ;
        RECT 112.090 173.530 112.230 174.230 ;
        RECT 112.030 173.210 112.290 173.530 ;
        RECT 112.550 173.190 112.690 175.930 ;
        RECT 116.630 175.590 116.890 175.910 ;
        RECT 113.870 175.250 114.130 175.570 ;
        RECT 113.410 174.910 113.670 175.230 ;
        RECT 112.490 172.870 112.750 173.190 ;
        RECT 113.470 171.830 113.610 174.910 ;
        RECT 113.930 172.510 114.070 175.250 ;
        RECT 113.870 172.190 114.130 172.510 ;
        RECT 113.410 171.510 113.670 171.830 ;
        RECT 113.470 168.090 113.610 171.510 ;
        RECT 116.690 170.810 116.830 175.590 ;
        RECT 117.090 171.850 117.350 172.170 ;
        RECT 116.630 170.490 116.890 170.810 ;
        RECT 117.150 170.210 117.290 171.850 ;
        RECT 117.610 171.830 117.750 183.670 ;
        RECT 118.530 181.690 118.670 191.150 ;
        RECT 118.930 190.550 119.190 190.870 ;
        RECT 118.990 188.830 119.130 190.550 ;
        RECT 118.930 188.510 119.190 188.830 ;
        RECT 118.930 186.130 119.190 186.450 ;
        RECT 118.990 183.730 119.130 186.130 ;
        RECT 118.930 183.410 119.190 183.730 ;
        RECT 118.470 181.370 118.730 181.690 ;
        RECT 118.990 178.290 119.130 183.410 ;
        RECT 118.930 177.970 119.190 178.290 ;
        RECT 118.470 176.950 118.730 177.270 ;
        RECT 118.530 174.890 118.670 176.950 ;
        RECT 118.990 175.570 119.130 177.970 ;
        RECT 118.930 175.250 119.190 175.570 ;
        RECT 118.470 174.570 118.730 174.890 ;
        RECT 119.450 173.610 119.590 206.960 ;
        RECT 120.310 206.870 120.570 206.960 ;
        RECT 122.210 205.150 122.350 210.190 ;
        RECT 125.370 209.930 125.630 210.250 ;
        RECT 122.660 209.055 124.200 209.425 ;
        RECT 125.430 208.890 125.570 209.930 ;
        RECT 125.370 208.570 125.630 208.890 ;
        RECT 123.990 207.550 124.250 207.870 ;
        RECT 124.050 206.170 124.190 207.550 ;
        RECT 123.990 205.850 124.250 206.170 ;
        RECT 122.150 204.830 122.410 205.150 ;
        RECT 124.050 205.005 124.190 205.850 ;
        RECT 123.980 204.635 124.260 205.005 ;
        RECT 124.910 204.150 125.170 204.470 ;
        RECT 122.660 203.615 124.200 203.985 ;
        RECT 123.070 203.130 123.330 203.450 ;
        RECT 123.130 201.750 123.270 203.130 ;
        RECT 120.310 201.430 120.570 201.750 ;
        RECT 123.070 201.430 123.330 201.750 ;
        RECT 120.370 192.230 120.510 201.430 ;
        RECT 123.130 200.050 123.270 201.430 ;
        RECT 123.070 199.730 123.330 200.050 ;
        RECT 122.660 198.175 124.200 198.545 ;
        RECT 122.660 192.735 124.200 193.105 ;
        RECT 120.310 191.910 120.570 192.230 ;
        RECT 119.850 191.570 120.110 191.890 ;
        RECT 119.910 176.330 120.050 191.570 ;
        RECT 120.370 181.690 120.510 191.910 ;
        RECT 124.450 190.550 124.710 190.870 ;
        RECT 124.510 189.850 124.650 190.550 ;
        RECT 124.450 189.530 124.710 189.850 ;
        RECT 122.660 187.295 124.200 187.665 ;
        RECT 123.530 185.110 123.790 185.430 ;
        RECT 123.590 183.050 123.730 185.110 ;
        RECT 123.530 182.730 123.790 183.050 ;
        RECT 122.660 181.855 124.200 182.225 ;
        RECT 120.310 181.370 120.570 181.690 ;
        RECT 122.610 181.370 122.870 181.690 ;
        RECT 121.690 181.030 121.950 181.350 ;
        RECT 120.310 180.690 120.570 181.010 ;
        RECT 120.370 177.270 120.510 180.690 ;
        RECT 120.310 176.950 120.570 177.270 ;
        RECT 119.910 176.190 121.430 176.330 ;
        RECT 119.850 175.250 120.110 175.570 ;
        RECT 118.530 173.470 119.590 173.610 ;
        RECT 119.910 173.530 120.050 175.250 ;
        RECT 118.010 172.190 118.270 172.510 ;
        RECT 117.550 171.510 117.810 171.830 ;
        RECT 116.690 170.070 117.290 170.210 ;
        RECT 114.790 168.790 115.050 169.110 ;
        RECT 113.410 167.770 113.670 168.090 ;
        RECT 114.850 167.410 114.990 168.790 ;
        RECT 116.690 167.750 116.830 170.070 ;
        RECT 116.630 167.430 116.890 167.750 ;
        RECT 111.110 167.090 111.370 167.410 ;
        RECT 114.790 167.090 115.050 167.410 ;
        RECT 111.170 164.670 111.310 167.090 ;
        RECT 115.250 166.750 115.510 167.070 ;
        RECT 115.710 166.750 115.970 167.070 ;
        RECT 116.630 166.750 116.890 167.070 ;
        RECT 117.090 166.750 117.350 167.070 ;
        RECT 115.310 164.690 115.450 166.750 ;
        RECT 115.770 165.370 115.910 166.750 ;
        RECT 116.170 166.410 116.430 166.730 ;
        RECT 115.710 165.050 115.970 165.370 ;
        RECT 111.170 164.530 112.230 164.670 ;
        RECT 110.190 164.205 110.450 164.350 ;
        RECT 110.180 163.835 110.460 164.205 ;
        RECT 111.570 161.990 111.830 162.310 ;
        RECT 109.730 161.310 109.990 161.630 ;
        RECT 109.270 159.610 109.530 159.930 ;
        RECT 109.790 158.910 109.930 161.310 ;
        RECT 110.650 160.970 110.910 161.290 ;
        RECT 110.190 158.930 110.450 159.250 ;
        RECT 109.730 158.590 109.990 158.910 ;
        RECT 109.730 156.100 109.990 156.190 ;
        RECT 108.870 155.960 109.990 156.100 ;
        RECT 109.730 155.870 109.990 155.960 ;
        RECT 110.250 154.150 110.390 158.930 ;
        RECT 110.710 157.210 110.850 160.970 ;
        RECT 110.650 156.890 110.910 157.210 ;
        RECT 110.190 153.830 110.450 154.150 ;
        RECT 109.730 152.470 109.990 152.790 ;
        RECT 109.270 150.770 109.530 151.090 ;
        RECT 107.890 150.430 108.150 150.750 ;
        RECT 107.950 149.050 108.090 150.430 ;
        RECT 104.730 148.820 105.330 148.960 ;
        RECT 104.210 144.990 104.470 145.310 ;
        RECT 103.750 144.310 104.010 144.630 ;
        RECT 103.810 139.870 103.950 144.310 ;
        RECT 104.270 142.930 104.410 144.990 ;
        RECT 104.210 142.610 104.470 142.930 ;
        RECT 104.730 139.870 104.870 148.820 ;
        RECT 107.890 148.730 108.150 149.050 ;
        RECT 105.130 148.050 105.390 148.370 ;
        RECT 105.190 146.330 105.330 148.050 ;
        RECT 105.870 146.495 107.410 146.865 ;
        RECT 105.130 146.010 105.390 146.330 ;
        RECT 107.950 142.930 108.090 148.730 ;
        RECT 109.330 145.650 109.470 150.770 ;
        RECT 109.790 148.710 109.930 152.470 ;
        RECT 110.250 150.750 110.390 153.830 ;
        RECT 111.630 151.285 111.770 161.990 ;
        RECT 112.090 159.590 112.230 164.530 ;
        RECT 115.250 164.370 115.510 164.690 ;
        RECT 112.490 164.030 112.750 164.350 ;
        RECT 113.410 164.030 113.670 164.350 ;
        RECT 112.030 159.270 112.290 159.590 ;
        RECT 111.560 150.915 111.840 151.285 ;
        RECT 110.190 150.430 110.450 150.750 ;
        RECT 111.570 150.430 111.830 150.750 ;
        RECT 109.730 148.390 109.990 148.710 ;
        RECT 111.110 147.030 111.370 147.350 ;
        RECT 109.270 145.330 109.530 145.650 ;
        RECT 110.650 144.310 110.910 144.630 ;
        RECT 110.710 143.610 110.850 144.310 ;
        RECT 108.350 143.290 108.610 143.610 ;
        RECT 110.650 143.290 110.910 143.610 ;
        RECT 107.890 142.610 108.150 142.930 ;
        RECT 105.870 141.055 107.410 141.425 ;
        RECT 103.290 139.550 103.550 139.870 ;
        RECT 103.750 139.550 104.010 139.870 ;
        RECT 104.670 139.550 104.930 139.870 ;
        RECT 105.590 139.550 105.850 139.870 ;
        RECT 104.670 138.870 104.930 139.190 ;
        RECT 104.210 137.170 104.470 137.490 ;
        RECT 104.270 126.270 104.410 137.170 ;
        RECT 104.210 125.950 104.470 126.270 ;
        RECT 103.290 122.890 103.550 123.210 ;
        RECT 103.350 120.830 103.490 122.890 ;
        RECT 103.290 120.510 103.550 120.830 ;
        RECT 103.290 115.410 103.550 115.730 ;
        RECT 102.830 112.350 103.090 112.670 ;
        RECT 102.830 111.670 103.090 111.990 ;
        RECT 102.890 110.970 103.030 111.670 ;
        RECT 102.830 110.650 103.090 110.970 ;
        RECT 103.350 109.950 103.490 115.410 ;
        RECT 104.730 113.010 104.870 138.870 ;
        RECT 105.650 137.490 105.790 139.550 ;
        RECT 108.410 138.930 108.550 143.290 ;
        RECT 110.190 142.950 110.450 143.270 ;
        RECT 108.810 142.610 109.070 142.930 ;
        RECT 108.870 140.890 109.010 142.610 ;
        RECT 109.730 142.270 109.990 142.590 ;
        RECT 108.810 140.570 109.070 140.890 ;
        RECT 109.790 140.550 109.930 142.270 ;
        RECT 110.250 142.250 110.390 142.950 ;
        RECT 110.190 141.930 110.450 142.250 ;
        RECT 109.730 140.230 109.990 140.550 ;
        RECT 110.190 139.890 110.450 140.210 ;
        RECT 107.950 138.790 108.550 138.930 ;
        RECT 109.270 138.870 109.530 139.190 ;
        RECT 107.950 137.490 108.090 138.790 ;
        RECT 109.330 138.170 109.470 138.870 ;
        RECT 108.350 137.850 108.610 138.170 ;
        RECT 109.270 137.850 109.530 138.170 ;
        RECT 108.410 137.490 108.550 137.850 ;
        RECT 105.590 137.170 105.850 137.490 ;
        RECT 107.890 137.170 108.150 137.490 ;
        RECT 108.350 137.170 108.610 137.490 ;
        RECT 105.870 135.615 107.410 135.985 ;
        RECT 108.810 134.110 109.070 134.430 ;
        RECT 108.350 133.430 108.610 133.750 ;
        RECT 108.410 132.730 108.550 133.430 ;
        RECT 108.350 132.410 108.610 132.730 ;
        RECT 107.890 131.390 108.150 131.710 ;
        RECT 105.870 130.175 107.410 130.545 ;
        RECT 105.130 125.950 105.390 126.270 ;
        RECT 105.190 124.570 105.330 125.950 ;
        RECT 105.870 124.735 107.410 125.105 ;
        RECT 105.130 124.250 105.390 124.570 ;
        RECT 106.510 122.550 106.770 122.870 ;
        RECT 106.570 121.170 106.710 122.550 ;
        RECT 107.950 121.170 108.090 131.390 ;
        RECT 108.870 130.010 109.010 134.110 ;
        RECT 109.730 133.430 109.990 133.750 ;
        RECT 108.810 129.690 109.070 130.010 ;
        RECT 109.790 128.990 109.930 133.430 ;
        RECT 110.250 129.330 110.390 139.890 ;
        RECT 110.190 129.010 110.450 129.330 ;
        RECT 109.730 128.670 109.990 128.990 ;
        RECT 110.250 123.890 110.390 129.010 ;
        RECT 111.170 128.310 111.310 147.030 ;
        RECT 111.630 142.590 111.770 150.430 ;
        RECT 111.570 142.270 111.830 142.590 ;
        RECT 112.090 141.910 112.230 159.270 ;
        RECT 112.550 159.250 112.690 164.030 ;
        RECT 112.490 158.930 112.750 159.250 ;
        RECT 113.470 158.230 113.610 164.030 ;
        RECT 115.310 162.310 115.450 164.370 ;
        RECT 116.230 164.350 116.370 166.410 ;
        RECT 116.170 164.030 116.430 164.350 ;
        RECT 115.710 163.690 115.970 164.010 ;
        RECT 115.250 161.990 115.510 162.310 ;
        RECT 115.770 161.970 115.910 163.690 ;
        RECT 115.710 161.650 115.970 161.970 ;
        RECT 116.230 159.930 116.370 164.030 ;
        RECT 116.690 162.650 116.830 166.750 ;
        RECT 116.630 162.330 116.890 162.650 ;
        RECT 116.690 161.630 116.830 162.330 ;
        RECT 116.630 161.310 116.890 161.630 ;
        RECT 116.170 159.610 116.430 159.930 ;
        RECT 115.710 158.930 115.970 159.250 ;
        RECT 113.410 157.910 113.670 158.230 ;
        RECT 112.490 155.870 112.750 156.190 ;
        RECT 114.790 155.870 115.050 156.190 ;
        RECT 112.550 153.325 112.690 155.870 ;
        RECT 114.850 154.490 114.990 155.870 ;
        RECT 114.790 154.170 115.050 154.490 ;
        RECT 112.480 152.955 112.760 153.325 ;
        RECT 112.550 145.310 112.690 152.955 ;
        RECT 112.950 152.470 113.210 152.790 ;
        RECT 113.010 151.430 113.150 152.470 ;
        RECT 112.950 151.110 113.210 151.430 ;
        RECT 113.410 147.030 113.670 147.350 ;
        RECT 112.490 144.990 112.750 145.310 ;
        RECT 112.030 141.590 112.290 141.910 ;
        RECT 111.570 134.110 111.830 134.430 ;
        RECT 112.030 134.110 112.290 134.430 ;
        RECT 111.630 132.730 111.770 134.110 ;
        RECT 111.570 132.410 111.830 132.730 ;
        RECT 112.090 128.650 112.230 134.110 ;
        RECT 112.550 128.900 112.690 144.990 ;
        RECT 113.470 144.630 113.610 147.030 ;
        RECT 113.410 144.310 113.670 144.630 ;
        RECT 113.470 142.930 113.610 144.310 ;
        RECT 113.410 142.610 113.670 142.930 ;
        RECT 115.250 142.610 115.510 142.930 ;
        RECT 114.330 139.550 114.590 139.870 ;
        RECT 114.390 138.170 114.530 139.550 ;
        RECT 114.790 139.210 115.050 139.530 ;
        RECT 114.850 138.170 114.990 139.210 ;
        RECT 115.310 138.170 115.450 142.610 ;
        RECT 114.330 137.850 114.590 138.170 ;
        RECT 114.790 137.850 115.050 138.170 ;
        RECT 115.250 137.850 115.510 138.170 ;
        RECT 113.870 133.770 114.130 134.090 ;
        RECT 113.930 132.390 114.070 133.770 ;
        RECT 113.870 132.070 114.130 132.390 ;
        RECT 112.550 128.760 113.150 128.900 ;
        RECT 112.030 128.560 112.290 128.650 ;
        RECT 112.030 128.420 112.690 128.560 ;
        RECT 112.030 128.330 112.290 128.420 ;
        RECT 111.110 127.990 111.370 128.310 ;
        RECT 111.570 127.990 111.830 128.310 ;
        RECT 110.650 125.950 110.910 126.270 ;
        RECT 110.190 123.570 110.450 123.890 ;
        RECT 108.810 123.230 109.070 123.550 ;
        RECT 106.510 120.850 106.770 121.170 ;
        RECT 107.890 120.850 108.150 121.170 ;
        RECT 105.870 119.295 107.410 119.665 ;
        RECT 108.870 116.370 109.010 123.230 ;
        RECT 109.270 122.550 109.530 122.870 ;
        RECT 109.330 119.130 109.470 122.550 ;
        RECT 109.270 118.810 109.530 119.130 ;
        RECT 108.870 116.230 109.470 116.370 ;
        RECT 108.350 114.390 108.610 114.710 ;
        RECT 105.870 113.855 107.410 114.225 ;
        RECT 108.410 113.010 108.550 114.390 ;
        RECT 104.670 112.690 104.930 113.010 ;
        RECT 108.350 112.690 108.610 113.010 ;
        RECT 106.970 111.670 107.230 111.990 ;
        RECT 107.030 110.970 107.170 111.670 ;
        RECT 106.970 110.650 107.230 110.970 ;
        RECT 103.290 109.630 103.550 109.950 ;
        RECT 100.070 106.910 100.330 107.230 ;
        RECT 100.130 105.530 100.270 106.910 ;
        RECT 99.610 105.210 99.870 105.530 ;
        RECT 100.070 105.210 100.330 105.530 ;
        RECT 99.670 104.510 99.810 105.210 ;
        RECT 102.830 104.870 103.090 105.190 ;
        RECT 98.690 104.190 98.950 104.510 ;
        RECT 99.610 104.190 99.870 104.510 ;
        RECT 98.750 102.130 98.890 104.190 ;
        RECT 98.690 101.810 98.950 102.130 ;
        RECT 99.150 100.790 99.410 101.110 ;
        RECT 99.210 100.090 99.350 100.790 ;
        RECT 102.890 100.090 103.030 104.870 ;
        RECT 103.350 101.790 103.490 109.630 ;
        RECT 105.870 108.415 107.410 108.785 ;
        RECT 103.750 106.230 104.010 106.550 ;
        RECT 103.290 101.470 103.550 101.790 ;
        RECT 103.810 101.450 103.950 106.230 ;
        RECT 108.410 104.170 108.550 112.690 ;
        RECT 108.810 104.530 109.070 104.850 ;
        RECT 108.350 103.850 108.610 104.170 ;
        RECT 107.890 103.510 108.150 103.830 ;
        RECT 105.870 102.975 107.410 103.345 ;
        RECT 107.950 101.790 108.090 103.510 ;
        RECT 108.870 102.810 109.010 104.530 ;
        RECT 108.810 102.490 109.070 102.810 ;
        RECT 108.350 102.210 108.610 102.470 ;
        RECT 109.330 102.210 109.470 116.230 ;
        RECT 109.730 115.410 109.990 115.730 ;
        RECT 109.790 113.690 109.930 115.410 ;
        RECT 109.730 113.370 109.990 113.690 ;
        RECT 110.710 107.910 110.850 125.950 ;
        RECT 111.170 118.110 111.310 127.990 ;
        RECT 111.630 126.125 111.770 127.990 ;
        RECT 112.030 126.290 112.290 126.610 ;
        RECT 111.560 125.755 111.840 126.125 ;
        RECT 112.090 121.850 112.230 126.290 ;
        RECT 112.030 121.530 112.290 121.850 ;
        RECT 112.090 118.110 112.230 121.530 ;
        RECT 112.550 118.450 112.690 128.420 ;
        RECT 113.010 126.610 113.150 128.760 ;
        RECT 112.950 126.290 113.210 126.610 ;
        RECT 114.330 126.290 114.590 126.610 ;
        RECT 113.010 123.890 113.150 126.290 ;
        RECT 113.410 125.950 113.670 126.270 ;
        RECT 112.950 123.570 113.210 123.890 ;
        RECT 112.490 118.130 112.750 118.450 ;
        RECT 111.110 117.790 111.370 118.110 ;
        RECT 112.030 117.790 112.290 118.110 ;
        RECT 113.470 112.670 113.610 125.950 ;
        RECT 114.390 121.850 114.530 126.290 ;
        RECT 114.330 121.530 114.590 121.850 ;
        RECT 113.870 118.470 114.130 118.790 ;
        RECT 113.930 117.770 114.070 118.470 ;
        RECT 114.390 118.450 114.530 121.530 ;
        RECT 115.770 118.790 115.910 158.930 ;
        RECT 116.630 157.910 116.890 158.230 ;
        RECT 116.690 155.850 116.830 157.910 ;
        RECT 116.630 155.530 116.890 155.850 ;
        RECT 117.150 155.250 117.290 166.750 ;
        RECT 118.070 165.370 118.210 172.190 ;
        RECT 118.010 165.050 118.270 165.370 ;
        RECT 118.010 158.930 118.270 159.250 ;
        RECT 116.690 155.110 117.290 155.250 ;
        RECT 117.550 155.190 117.810 155.510 ;
        RECT 116.690 154.490 116.830 155.110 ;
        RECT 117.610 154.490 117.750 155.190 ;
        RECT 118.070 154.490 118.210 158.930 ;
        RECT 116.630 154.170 116.890 154.490 ;
        RECT 117.550 154.170 117.810 154.490 ;
        RECT 118.010 154.170 118.270 154.490 ;
        RECT 116.690 151.770 116.830 154.170 ;
        RECT 118.010 153.150 118.270 153.470 ;
        RECT 116.630 151.450 116.890 151.770 ;
        RECT 116.690 148.710 116.830 151.450 ;
        RECT 118.070 151.090 118.210 153.150 ;
        RECT 118.010 150.770 118.270 151.090 ;
        RECT 116.630 148.620 116.890 148.710 ;
        RECT 116.630 148.480 117.290 148.620 ;
        RECT 116.630 148.390 116.890 148.480 ;
        RECT 117.150 145.650 117.290 148.480 ;
        RECT 118.070 146.240 118.210 150.770 ;
        RECT 118.530 150.750 118.670 173.470 ;
        RECT 119.850 173.210 120.110 173.530 ;
        RECT 118.930 171.510 119.190 171.830 ;
        RECT 118.990 153.810 119.130 171.510 ;
        RECT 119.390 166.410 119.650 166.730 ;
        RECT 119.450 165.370 119.590 166.410 ;
        RECT 119.390 165.050 119.650 165.370 ;
        RECT 119.390 164.370 119.650 164.690 ;
        RECT 119.450 162.650 119.590 164.370 ;
        RECT 119.850 163.690 120.110 164.010 ;
        RECT 119.390 162.330 119.650 162.650 ;
        RECT 119.910 157.210 120.050 163.690 ;
        RECT 121.290 158.910 121.430 176.190 ;
        RECT 121.750 173.530 121.890 181.030 ;
        RECT 122.150 179.670 122.410 179.990 ;
        RECT 122.210 177.950 122.350 179.670 ;
        RECT 122.150 177.630 122.410 177.950 ;
        RECT 122.670 177.180 122.810 181.370 ;
        RECT 124.450 180.690 124.710 181.010 ;
        RECT 122.210 177.040 122.810 177.180 ;
        RECT 121.690 173.210 121.950 173.530 ;
        RECT 122.210 172.510 122.350 177.040 ;
        RECT 122.660 176.415 124.200 176.785 ;
        RECT 122.150 172.190 122.410 172.510 ;
        RECT 121.690 169.470 121.950 169.790 ;
        RECT 121.750 165.370 121.890 169.470 ;
        RECT 122.210 168.090 122.350 172.190 ;
        RECT 122.660 170.975 124.200 171.345 ;
        RECT 122.150 167.770 122.410 168.090 ;
        RECT 122.660 165.535 124.200 165.905 ;
        RECT 121.690 165.050 121.950 165.370 ;
        RECT 121.750 160.950 121.890 165.050 ;
        RECT 124.510 164.010 124.650 180.690 ;
        RECT 124.450 163.690 124.710 164.010 ;
        RECT 121.690 160.630 121.950 160.950 ;
        RECT 122.150 160.630 122.410 160.950 ;
        RECT 122.210 159.590 122.350 160.630 ;
        RECT 122.660 160.095 124.200 160.465 ;
        RECT 124.970 160.010 125.110 204.150 ;
        RECT 125.430 164.670 125.570 208.570 ;
        RECT 130.030 208.210 130.170 212.200 ;
        RECT 133.650 209.590 133.910 209.910 ;
        RECT 133.710 208.210 133.850 209.590 ;
        RECT 137.390 208.890 137.530 212.200 ;
        RECT 137.330 208.570 137.590 208.890 ;
        RECT 129.970 207.890 130.230 208.210 ;
        RECT 133.650 207.890 133.910 208.210 ;
        RECT 128.590 207.550 128.850 207.870 ;
        RECT 132.270 207.550 132.530 207.870 ;
        RECT 126.750 206.870 127.010 207.190 ;
        RECT 126.290 205.170 126.550 205.490 ;
        RECT 125.830 199.390 126.090 199.710 ;
        RECT 125.890 196.310 126.030 199.390 ;
        RECT 126.350 197.330 126.490 205.170 ;
        RECT 126.290 197.010 126.550 197.330 ;
        RECT 125.830 195.990 126.090 196.310 ;
        RECT 126.350 194.610 126.490 197.010 ;
        RECT 126.290 194.290 126.550 194.610 ;
        RECT 126.290 189.365 126.550 189.510 ;
        RECT 126.280 188.995 126.560 189.365 ;
        RECT 126.290 188.510 126.550 188.830 ;
        RECT 126.350 187.130 126.490 188.510 ;
        RECT 126.290 186.810 126.550 187.130 ;
        RECT 126.810 177.690 126.950 206.870 ;
        RECT 127.670 202.790 127.930 203.110 ;
        RECT 127.730 200.390 127.870 202.790 ;
        RECT 128.650 201.750 128.790 207.550 ;
        RECT 132.330 206.170 132.470 207.550 ;
        RECT 132.270 205.850 132.530 206.170 ;
        RECT 133.190 205.850 133.450 206.170 ;
        RECT 133.250 205.150 133.390 205.850 ;
        RECT 133.710 205.490 133.850 207.890 ;
        RECT 135.950 207.550 136.210 207.870 ;
        RECT 135.030 206.870 135.290 207.190 ;
        RECT 135.490 206.870 135.750 207.190 ;
        RECT 135.090 205.490 135.230 206.870 ;
        RECT 133.650 205.170 133.910 205.490 ;
        RECT 135.030 205.170 135.290 205.490 ;
        RECT 133.190 204.830 133.450 205.150 ;
        RECT 135.030 204.490 135.290 204.810 ;
        RECT 134.100 202.595 134.380 202.965 ;
        RECT 133.190 202.110 133.450 202.430 ;
        RECT 128.590 201.430 128.850 201.750 ;
        RECT 127.670 200.070 127.930 200.390 ;
        RECT 127.730 194.690 127.870 200.070 ;
        RECT 128.130 199.390 128.390 199.710 ;
        RECT 128.190 195.290 128.330 199.390 ;
        RECT 128.590 198.710 128.850 199.030 ;
        RECT 128.650 197.670 128.790 198.710 ;
        RECT 128.590 197.350 128.850 197.670 ;
        RECT 129.970 195.990 130.230 196.310 ;
        RECT 128.130 194.970 128.390 195.290 ;
        RECT 127.730 194.550 128.330 194.690 ;
        RECT 127.670 192.250 127.930 192.570 ;
        RECT 127.210 189.530 127.470 189.850 ;
        RECT 127.270 186.110 127.410 189.530 ;
        RECT 127.730 189.170 127.870 192.250 ;
        RECT 127.670 188.850 127.930 189.170 ;
        RECT 127.670 188.170 127.930 188.490 ;
        RECT 127.730 187.325 127.870 188.170 ;
        RECT 127.660 186.955 127.940 187.325 ;
        RECT 127.670 186.470 127.930 186.790 ;
        RECT 127.210 185.790 127.470 186.110 ;
        RECT 127.270 178.970 127.410 185.790 ;
        RECT 127.730 184.410 127.870 186.470 ;
        RECT 128.190 184.490 128.330 194.550 ;
        RECT 129.050 193.270 129.310 193.590 ;
        RECT 129.110 192.230 129.250 193.270 ;
        RECT 129.050 191.910 129.310 192.230 ;
        RECT 130.030 191.970 130.170 195.990 ;
        RECT 133.250 195.290 133.390 202.110 ;
        RECT 134.170 201.750 134.310 202.595 ;
        RECT 134.570 202.450 134.830 202.770 ;
        RECT 134.630 202.285 134.770 202.450 ;
        RECT 134.560 201.915 134.840 202.285 ;
        RECT 134.110 201.430 134.370 201.750 ;
        RECT 135.090 200.730 135.230 204.490 ;
        RECT 135.550 202.430 135.690 206.870 ;
        RECT 136.010 204.810 136.150 207.550 ;
        RECT 137.790 206.870 138.050 207.190 ;
        RECT 135.950 204.490 136.210 204.810 ;
        RECT 137.330 204.490 137.590 204.810 ;
        RECT 137.390 203.530 137.530 204.490 ;
        RECT 136.930 203.390 137.530 203.530 ;
        RECT 136.930 202.770 137.070 203.390 ;
        RECT 137.850 202.850 137.990 206.870 ;
        RECT 139.450 206.335 140.990 206.705 ;
        RECT 139.160 204.635 139.440 205.005 ;
        RECT 138.250 204.150 138.510 204.470 ;
        RECT 136.870 202.450 137.130 202.770 ;
        RECT 137.390 202.710 137.990 202.850 ;
        RECT 135.490 202.110 135.750 202.430 ;
        RECT 136.410 201.430 136.670 201.750 ;
        RECT 135.030 200.410 135.290 200.730 ;
        RECT 136.470 199.710 136.610 201.430 ;
        RECT 136.410 199.390 136.670 199.710 ;
        RECT 135.490 197.010 135.750 197.330 ;
        RECT 134.110 195.990 134.370 196.310 ;
        RECT 134.570 195.990 134.830 196.310 ;
        RECT 130.890 194.970 131.150 195.290 ;
        RECT 133.190 194.970 133.450 195.290 ;
        RECT 130.950 193.590 131.090 194.970 ;
        RECT 131.810 193.950 132.070 194.270 ;
        RECT 130.890 193.270 131.150 193.590 ;
        RECT 130.030 191.890 131.550 191.970 ;
        RECT 128.590 191.570 128.850 191.890 ;
        RECT 130.030 191.830 131.610 191.890 ;
        RECT 131.350 191.570 131.610 191.830 ;
        RECT 128.650 187.130 128.790 191.570 ;
        RECT 131.350 190.890 131.610 191.210 ;
        RECT 130.890 190.550 131.150 190.870 ;
        RECT 129.510 189.530 129.770 189.850 ;
        RECT 129.570 189.080 129.710 189.530 ;
        RECT 130.950 189.170 131.090 190.550 ;
        RECT 129.110 188.940 129.710 189.080 ;
        RECT 129.110 188.490 129.250 188.940 ;
        RECT 130.890 188.850 131.150 189.170 ;
        RECT 129.050 188.170 129.310 188.490 ;
        RECT 130.430 188.060 130.690 188.150 ;
        RECT 130.030 187.920 130.690 188.060 ;
        RECT 128.590 186.810 128.850 187.130 ;
        RECT 129.040 186.955 129.320 187.325 ;
        RECT 129.110 186.700 129.250 186.955 ;
        RECT 129.510 186.700 129.770 186.790 ;
        RECT 129.110 186.560 129.770 186.700 ;
        RECT 127.670 184.090 127.930 184.410 ;
        RECT 128.190 184.350 128.790 184.490 ;
        RECT 128.130 182.390 128.390 182.710 ;
        RECT 127.210 178.650 127.470 178.970 ;
        RECT 126.810 177.550 127.870 177.690 ;
        RECT 128.190 177.610 128.330 182.390 ;
        RECT 126.290 174.230 126.550 174.550 ;
        RECT 126.350 173.530 126.490 174.230 ;
        RECT 126.290 173.210 126.550 173.530 ;
        RECT 126.750 166.410 127.010 166.730 ;
        RECT 127.210 166.410 127.470 166.730 ;
        RECT 126.810 166.130 126.950 166.410 ;
        RECT 126.350 165.990 126.950 166.130 ;
        RECT 125.430 164.530 126.030 164.670 ;
        RECT 125.370 163.350 125.630 163.670 ;
        RECT 124.510 159.870 125.110 160.010 ;
        RECT 122.150 159.270 122.410 159.590 ;
        RECT 121.230 158.590 121.490 158.910 ;
        RECT 124.510 158.650 124.650 159.870 ;
        RECT 124.910 158.930 125.170 159.250 ;
        RECT 124.050 158.510 124.650 158.650 ;
        RECT 119.850 156.890 120.110 157.210 ;
        RECT 118.930 153.490 119.190 153.810 ;
        RECT 119.910 153.210 120.050 156.890 ;
        RECT 124.050 156.870 124.190 158.510 ;
        RECT 124.450 157.910 124.710 158.230 ;
        RECT 123.990 156.550 124.250 156.870 ;
        RECT 124.510 156.190 124.650 157.910 ;
        RECT 123.990 155.870 124.250 156.190 ;
        RECT 124.450 155.870 124.710 156.190 ;
        RECT 124.050 155.420 124.190 155.870 ;
        RECT 124.050 155.280 124.650 155.420 ;
        RECT 122.660 154.655 124.200 155.025 ;
        RECT 124.510 153.810 124.650 155.280 ;
        RECT 124.970 154.490 125.110 158.930 ;
        RECT 124.910 154.170 125.170 154.490 ;
        RECT 120.310 153.490 120.570 153.810 ;
        RECT 120.770 153.490 121.030 153.810 ;
        RECT 124.450 153.490 124.710 153.810 ;
        RECT 118.990 153.070 120.050 153.210 ;
        RECT 118.470 150.430 118.730 150.750 ;
        RECT 118.530 147.350 118.670 150.430 ;
        RECT 118.470 147.030 118.730 147.350 ;
        RECT 118.470 146.240 118.730 146.330 ;
        RECT 118.070 146.100 118.730 146.240 ;
        RECT 118.470 146.010 118.730 146.100 ;
        RECT 117.090 145.330 117.350 145.650 ;
        RECT 116.170 141.590 116.430 141.910 ;
        RECT 116.230 139.530 116.370 141.590 ;
        RECT 117.150 139.870 117.290 145.330 ;
        RECT 118.010 141.590 118.270 141.910 ;
        RECT 117.090 139.550 117.350 139.870 ;
        RECT 116.170 139.210 116.430 139.530 ;
        RECT 118.070 138.170 118.210 141.590 ;
        RECT 118.010 137.850 118.270 138.170 ;
        RECT 117.090 137.170 117.350 137.490 ;
        RECT 117.150 131.710 117.290 137.170 ;
        RECT 118.530 137.150 118.670 146.010 ;
        RECT 118.470 136.830 118.730 137.150 ;
        RECT 118.470 135.130 118.730 135.450 ;
        RECT 118.010 131.730 118.270 132.050 ;
        RECT 117.090 131.390 117.350 131.710 ;
        RECT 116.630 131.050 116.890 131.370 ;
        RECT 116.170 128.330 116.430 128.650 ;
        RECT 116.230 127.290 116.370 128.330 ;
        RECT 116.170 126.970 116.430 127.290 ;
        RECT 115.710 118.470 115.970 118.790 ;
        RECT 114.330 118.130 114.590 118.450 ;
        RECT 113.870 117.450 114.130 117.770 ;
        RECT 115.250 114.390 115.510 114.710 ;
        RECT 115.710 114.390 115.970 114.710 ;
        RECT 115.310 113.010 115.450 114.390 ;
        RECT 115.770 113.350 115.910 114.390 ;
        RECT 115.710 113.030 115.970 113.350 ;
        RECT 115.250 112.690 115.510 113.010 ;
        RECT 111.110 112.350 111.370 112.670 ;
        RECT 113.410 112.350 113.670 112.670 ;
        RECT 111.170 109.950 111.310 112.350 ;
        RECT 112.030 109.970 112.290 110.290 ;
        RECT 111.110 109.630 111.370 109.950 ;
        RECT 110.650 107.590 110.910 107.910 ;
        RECT 108.350 102.150 109.470 102.210 ;
        RECT 108.410 102.070 109.470 102.150 ;
        RECT 105.590 101.470 105.850 101.790 ;
        RECT 107.890 101.470 108.150 101.790 ;
        RECT 110.190 101.470 110.450 101.790 ;
        RECT 110.650 101.700 110.910 101.790 ;
        RECT 111.170 101.700 111.310 109.630 ;
        RECT 112.090 107.230 112.230 109.970 ;
        RECT 115.310 107.230 115.450 112.690 ;
        RECT 116.170 111.670 116.430 111.990 ;
        RECT 116.230 110.630 116.370 111.670 ;
        RECT 116.170 110.310 116.430 110.630 ;
        RECT 116.230 107.230 116.370 110.310 ;
        RECT 112.030 106.910 112.290 107.230 ;
        RECT 115.250 106.910 115.510 107.230 ;
        RECT 116.170 106.910 116.430 107.230 ;
        RECT 112.950 106.570 113.210 106.890 ;
        RECT 113.010 104.850 113.150 106.570 ;
        RECT 113.870 106.230 114.130 106.550 ;
        RECT 114.330 106.230 114.590 106.550 ;
        RECT 113.930 105.530 114.070 106.230 ;
        RECT 113.870 105.210 114.130 105.530 ;
        RECT 112.950 104.530 113.210 104.850 ;
        RECT 110.650 101.560 111.310 101.700 ;
        RECT 110.650 101.470 110.910 101.560 ;
        RECT 103.750 101.130 104.010 101.450 ;
        RECT 99.150 99.770 99.410 100.090 ;
        RECT 102.830 99.770 103.090 100.090 ;
        RECT 97.310 99.090 97.570 99.410 ;
        RECT 98.230 99.090 98.490 99.410 ;
        RECT 96.850 98.750 97.110 99.070 ;
        RECT 105.130 98.980 105.390 99.070 ;
        RECT 105.650 98.980 105.790 101.470 ;
        RECT 106.970 100.790 107.230 101.110 ;
        RECT 107.030 99.750 107.170 100.790 ;
        RECT 110.250 100.090 110.390 101.470 ;
        RECT 110.190 99.770 110.450 100.090 ;
        RECT 106.970 99.430 107.230 99.750 ;
        RECT 105.130 98.840 105.790 98.980 ;
        RECT 105.130 98.750 105.390 98.840 ;
        RECT 95.470 98.070 95.730 98.390 ;
        RECT 95.010 95.350 95.270 95.670 ;
        RECT 91.850 87.790 92.450 87.930 ;
        RECT 91.790 87.190 92.050 87.510 ;
        RECT 91.850 86.685 91.990 87.190 ;
        RECT 91.780 86.315 92.060 86.685 ;
        RECT 91.790 86.170 92.050 86.315 ;
        RECT 92.310 85.890 92.450 87.790 ;
        RECT 91.850 85.750 92.450 85.890 ;
        RECT 92.770 87.790 93.370 87.930 ;
        RECT 93.690 94.420 94.290 94.560 ;
        RECT 91.330 84.470 91.590 84.790 ;
        RECT 90.870 83.450 91.130 83.770 ;
        RECT 87.650 83.110 87.910 83.430 ;
        RECT 88.570 83.110 88.830 83.430 ;
        RECT 85.350 79.710 85.610 80.030 ;
        RECT 83.970 77.220 84.230 77.310 ;
        RECT 83.970 77.080 84.630 77.220 ;
        RECT 83.970 76.990 84.230 77.080 ;
        RECT 83.970 76.310 84.230 76.630 ;
        RECT 84.030 72.890 84.170 76.310 ;
        RECT 83.970 72.570 84.230 72.890 ;
        RECT 82.590 71.890 82.850 72.210 ;
        RECT 81.670 68.830 81.930 69.150 ;
        RECT 80.810 67.930 81.410 68.070 ;
        RECT 80.810 66.770 80.950 67.930 ;
        RECT 82.650 66.770 82.790 71.890 ;
        RECT 84.030 71.870 84.170 72.570 ;
        RECT 83.970 71.550 84.230 71.870 ;
        RECT 84.490 69.830 84.630 77.080 ;
        RECT 85.410 76.970 85.550 79.710 ;
        RECT 87.190 77.330 87.450 77.650 ;
        RECT 85.350 76.650 85.610 76.970 ;
        RECT 85.410 75.610 85.550 76.650 ;
        RECT 85.810 76.310 86.070 76.630 ;
        RECT 85.350 75.290 85.610 75.610 ;
        RECT 84.890 73.590 85.150 73.910 ;
        RECT 84.950 72.890 85.090 73.590 ;
        RECT 85.410 72.970 85.550 75.290 ;
        RECT 85.870 74.250 86.010 76.310 ;
        RECT 87.250 74.590 87.390 77.330 ;
        RECT 86.730 74.270 86.990 74.590 ;
        RECT 87.190 74.270 87.450 74.590 ;
        RECT 85.810 73.930 86.070 74.250 ;
        RECT 84.890 72.570 85.150 72.890 ;
        RECT 85.410 72.830 86.010 72.970 ;
        RECT 85.870 72.210 86.010 72.830 ;
        RECT 86.270 72.230 86.530 72.550 ;
        RECT 85.810 71.890 86.070 72.210 ;
        RECT 84.430 69.510 84.690 69.830 ;
        RECT 84.490 69.150 84.630 69.510 ;
        RECT 86.330 69.490 86.470 72.230 ;
        RECT 86.790 72.210 86.930 74.270 ;
        RECT 87.710 72.550 87.850 83.110 ;
        RECT 90.870 81.750 91.130 82.070 ;
        RECT 90.930 80.370 91.070 81.750 ;
        RECT 90.870 80.050 91.130 80.370 ;
        RECT 89.080 78.495 90.620 78.865 ;
        RECT 90.870 77.330 91.130 77.650 ;
        RECT 88.110 73.590 88.370 73.910 ;
        RECT 87.650 72.230 87.910 72.550 ;
        RECT 86.730 71.890 86.990 72.210 ;
        RECT 86.270 69.170 86.530 69.490 ;
        RECT 87.710 69.150 87.850 72.230 ;
        RECT 84.430 68.830 84.690 69.150 ;
        RECT 87.650 68.830 87.910 69.150 ;
        RECT 83.510 68.150 83.770 68.470 ;
        RECT 84.430 68.380 84.690 68.470 ;
        RECT 84.030 68.240 84.690 68.380 ;
        RECT 83.570 67.450 83.710 68.150 ;
        RECT 83.510 67.130 83.770 67.450 ;
        RECT 77.070 66.450 77.330 66.770 ;
        RECT 79.370 66.450 79.630 66.770 ;
        RECT 80.750 66.450 81.010 66.770 ;
        RECT 82.590 66.450 82.850 66.770 ;
        RECT 83.510 66.680 83.770 66.770 ;
        RECT 84.030 66.680 84.170 68.240 ;
        RECT 84.430 68.150 84.690 68.240 ;
        RECT 84.430 67.130 84.690 67.450 ;
        RECT 84.490 66.770 84.630 67.130 ;
        RECT 88.170 66.770 88.310 73.590 ;
        RECT 89.080 73.055 90.620 73.425 ;
        RECT 88.570 72.570 88.830 72.890 ;
        RECT 88.630 69.150 88.770 72.570 ;
        RECT 89.490 71.780 89.750 71.870 ;
        RECT 89.090 71.640 89.750 71.780 ;
        RECT 89.090 71.045 89.230 71.640 ;
        RECT 89.490 71.550 89.750 71.640 ;
        RECT 89.020 70.675 89.300 71.045 ;
        RECT 89.090 70.170 89.230 70.675 ;
        RECT 90.930 70.170 91.070 77.330 ;
        RECT 91.330 76.310 91.590 76.630 ;
        RECT 91.390 71.870 91.530 76.310 ;
        RECT 91.850 74.445 91.990 85.750 ;
        RECT 92.250 84.470 92.510 84.790 ;
        RECT 92.310 82.410 92.450 84.470 ;
        RECT 92.250 82.090 92.510 82.410 ;
        RECT 92.250 79.710 92.510 80.030 ;
        RECT 92.310 78.330 92.450 79.710 ;
        RECT 92.250 78.010 92.510 78.330 ;
        RECT 91.780 74.075 92.060 74.445 ;
        RECT 92.770 72.800 92.910 87.790 ;
        RECT 93.170 87.190 93.430 87.510 ;
        RECT 93.230 86.490 93.370 87.190 ;
        RECT 93.170 86.170 93.430 86.490 ;
        RECT 93.690 78.240 93.830 94.420 ;
        RECT 94.550 94.330 94.810 94.650 ;
        RECT 95.530 93.970 95.670 98.070 ;
        RECT 104.210 96.710 104.470 97.030 ;
        RECT 100.990 96.030 101.250 96.350 ;
        RECT 94.090 93.880 94.350 93.970 ;
        RECT 94.090 93.740 94.750 93.880 ;
        RECT 94.090 93.650 94.350 93.740 ;
        RECT 94.610 85.890 94.750 93.740 ;
        RECT 95.470 93.650 95.730 93.970 ;
        RECT 95.930 93.650 96.190 93.970 ;
        RECT 95.010 92.970 95.270 93.290 ;
        RECT 95.070 86.490 95.210 92.970 ;
        RECT 95.990 92.950 96.130 93.650 ;
        RECT 96.850 93.310 97.110 93.630 ;
        RECT 95.930 92.630 96.190 92.950 ;
        RECT 95.470 87.870 95.730 88.190 ;
        RECT 95.010 86.170 95.270 86.490 ;
        RECT 94.610 85.750 95.210 85.890 ;
        RECT 95.070 85.470 95.210 85.750 ;
        RECT 95.010 85.150 95.270 85.470 ;
        RECT 95.530 85.325 95.670 87.870 ;
        RECT 95.990 87.850 96.130 92.630 ;
        RECT 96.910 89.210 97.050 93.310 ;
        RECT 98.690 92.630 98.950 92.950 ;
        RECT 98.750 91.930 98.890 92.630 ;
        RECT 101.050 91.930 101.190 96.030 ;
        RECT 104.270 94.310 104.410 96.710 ;
        RECT 105.190 94.310 105.330 98.750 ;
        RECT 105.870 97.535 107.410 97.905 ;
        RECT 110.250 97.370 110.390 99.770 ;
        RECT 110.710 99.410 110.850 101.470 ;
        RECT 110.650 99.090 110.910 99.410 ;
        RECT 113.010 98.730 113.150 104.530 ;
        RECT 113.410 104.190 113.670 104.510 ;
        RECT 113.470 102.570 113.610 104.190 ;
        RECT 113.470 102.430 114.070 102.570 ;
        RECT 113.930 99.410 114.070 102.430 ;
        RECT 114.390 100.090 114.530 106.230 ;
        RECT 116.690 105.610 116.830 131.050 ;
        RECT 118.070 126.950 118.210 131.730 ;
        RECT 118.010 126.630 118.270 126.950 ;
        RECT 118.530 126.270 118.670 135.130 ;
        RECT 118.470 125.950 118.730 126.270 ;
        RECT 118.990 125.590 119.130 153.070 ;
        RECT 119.390 152.470 119.650 152.790 ;
        RECT 119.450 145.310 119.590 152.470 ;
        RECT 119.850 150.090 120.110 150.410 ;
        RECT 119.390 144.990 119.650 145.310 ;
        RECT 119.390 141.930 119.650 142.250 ;
        RECT 119.450 126.950 119.590 141.930 ;
        RECT 119.910 135.450 120.050 150.090 ;
        RECT 120.370 143.270 120.510 153.490 ;
        RECT 120.830 146.330 120.970 153.490 ;
        RECT 121.230 153.150 121.490 153.470 ;
        RECT 121.290 148.030 121.430 153.150 ;
        RECT 121.690 152.470 121.950 152.790 ;
        RECT 121.750 148.710 121.890 152.470 ;
        RECT 122.150 149.750 122.410 150.070 ;
        RECT 122.210 149.050 122.350 149.750 ;
        RECT 122.660 149.215 124.200 149.585 ;
        RECT 122.150 148.730 122.410 149.050 ;
        RECT 121.690 148.390 121.950 148.710 ;
        RECT 124.510 148.370 124.650 153.490 ;
        RECT 125.430 152.790 125.570 163.350 ;
        RECT 125.890 153.470 126.030 164.530 ;
        RECT 125.830 153.150 126.090 153.470 ;
        RECT 125.370 152.470 125.630 152.790 ;
        RECT 124.910 149.750 125.170 150.070 ;
        RECT 124.970 149.050 125.110 149.750 ;
        RECT 124.910 148.730 125.170 149.050 ;
        RECT 125.430 148.450 125.570 152.470 ;
        RECT 124.450 148.050 124.710 148.370 ;
        RECT 124.970 148.310 125.570 148.450 ;
        RECT 121.230 147.710 121.490 148.030 ;
        RECT 122.150 147.030 122.410 147.350 ;
        RECT 120.770 146.010 121.030 146.330 ;
        RECT 122.210 145.310 122.350 147.030 ;
        RECT 122.150 144.990 122.410 145.310 ;
        RECT 122.660 143.775 124.200 144.145 ;
        RECT 120.310 142.950 120.570 143.270 ;
        RECT 124.510 142.930 124.650 148.050 ;
        RECT 124.970 146.330 125.110 148.310 ;
        RECT 125.370 147.710 125.630 148.030 ;
        RECT 125.430 146.330 125.570 147.710 ;
        RECT 125.830 147.030 126.090 147.350 ;
        RECT 124.910 146.010 125.170 146.330 ;
        RECT 125.370 146.010 125.630 146.330 ;
        RECT 122.150 142.610 122.410 142.930 ;
        RECT 124.450 142.610 124.710 142.930 ;
        RECT 121.230 141.930 121.490 142.250 ;
        RECT 121.290 140.890 121.430 141.930 ;
        RECT 121.230 140.570 121.490 140.890 ;
        RECT 121.690 139.210 121.950 139.530 ;
        RECT 121.750 138.170 121.890 139.210 ;
        RECT 121.690 137.850 121.950 138.170 ;
        RECT 119.850 135.130 120.110 135.450 ;
        RECT 119.390 126.630 119.650 126.950 ;
        RECT 119.390 125.950 119.650 126.270 ;
        RECT 117.550 125.270 117.810 125.590 ;
        RECT 118.470 125.270 118.730 125.590 ;
        RECT 118.930 125.270 119.190 125.590 ;
        RECT 117.610 118.450 117.750 125.270 ;
        RECT 117.550 118.130 117.810 118.450 ;
        RECT 118.530 118.110 118.670 125.270 ;
        RECT 119.450 124.570 119.590 125.950 ;
        RECT 119.390 124.250 119.650 124.570 ;
        RECT 119.910 123.550 120.050 135.130 ;
        RECT 122.210 134.430 122.350 142.610 ;
        RECT 122.660 138.335 124.200 138.705 ;
        RECT 122.150 134.110 122.410 134.430 ;
        RECT 124.450 133.430 124.710 133.750 ;
        RECT 122.660 132.895 124.200 133.265 ;
        RECT 121.230 131.390 121.490 131.710 ;
        RECT 121.290 130.010 121.430 131.390 ;
        RECT 121.230 129.690 121.490 130.010 ;
        RECT 124.510 129.410 124.650 133.430 ;
        RECT 124.970 132.050 125.110 146.010 ;
        RECT 125.890 144.630 126.030 147.030 ;
        RECT 125.830 144.310 126.090 144.630 ;
        RECT 125.370 134.110 125.630 134.430 ;
        RECT 124.910 131.730 125.170 132.050 ;
        RECT 125.430 130.010 125.570 134.110 ;
        RECT 126.350 132.730 126.490 165.990 ;
        RECT 127.270 165.450 127.410 166.410 ;
        RECT 126.810 165.310 127.410 165.450 ;
        RECT 126.810 164.690 126.950 165.310 ;
        RECT 126.750 164.370 127.010 164.690 ;
        RECT 127.210 164.670 127.470 164.690 ;
        RECT 127.730 164.670 127.870 177.550 ;
        RECT 128.130 177.290 128.390 177.610 ;
        RECT 128.190 175.570 128.330 177.290 ;
        RECT 128.130 175.250 128.390 175.570 ;
        RECT 128.650 170.210 128.790 184.350 ;
        RECT 129.110 183.390 129.250 186.560 ;
        RECT 129.510 186.470 129.770 186.560 ;
        RECT 130.030 186.450 130.170 187.920 ;
        RECT 130.430 187.830 130.690 187.920 ;
        RECT 129.970 186.130 130.230 186.450 ;
        RECT 129.510 185.110 129.770 185.430 ;
        RECT 129.050 183.070 129.310 183.390 ;
        RECT 129.110 178.290 129.250 183.070 ;
        RECT 129.050 177.970 129.310 178.290 ;
        RECT 129.570 172.510 129.710 185.110 ;
        RECT 130.030 183.390 130.170 186.130 ;
        RECT 131.410 185.430 131.550 190.890 ;
        RECT 131.870 188.830 132.010 193.950 ;
        RECT 133.190 193.270 133.450 193.590 ;
        RECT 133.250 190.870 133.390 193.270 ;
        RECT 134.170 192.230 134.310 195.990 ;
        RECT 134.630 193.930 134.770 195.990 ;
        RECT 134.570 193.610 134.830 193.930 ;
        RECT 135.550 192.570 135.690 197.010 ;
        RECT 136.410 194.970 136.670 195.290 ;
        RECT 136.470 193.590 136.610 194.970 ;
        RECT 136.410 193.270 136.670 193.590 ;
        RECT 136.870 193.270 137.130 193.590 ;
        RECT 135.490 192.250 135.750 192.570 ;
        RECT 133.650 191.910 133.910 192.230 ;
        RECT 134.110 191.910 134.370 192.230 ;
        RECT 133.190 190.550 133.450 190.870 ;
        RECT 132.270 189.530 132.530 189.850 ;
        RECT 131.810 188.510 132.070 188.830 ;
        RECT 132.330 187.130 132.470 189.530 ;
        RECT 132.270 186.810 132.530 187.130 ;
        RECT 131.350 185.110 131.610 185.430 ;
        RECT 131.410 184.410 131.550 185.110 ;
        RECT 132.330 184.410 132.470 186.810 ;
        RECT 133.250 186.110 133.390 190.550 ;
        RECT 133.710 189.850 133.850 191.910 ;
        RECT 134.170 189.850 134.310 191.910 ;
        RECT 134.570 191.570 134.830 191.890 ;
        RECT 133.650 189.530 133.910 189.850 ;
        RECT 134.110 189.530 134.370 189.850 ;
        RECT 134.630 188.830 134.770 191.570 ;
        RECT 136.930 189.850 137.070 193.270 ;
        RECT 136.870 189.530 137.130 189.850 ;
        RECT 134.570 188.510 134.830 188.830 ;
        RECT 134.110 186.130 134.370 186.450 ;
        RECT 133.190 185.790 133.450 186.110 ;
        RECT 134.170 184.410 134.310 186.130 ;
        RECT 134.630 184.410 134.770 188.510 ;
        RECT 136.930 188.150 137.070 189.530 ;
        RECT 137.390 189.365 137.530 202.710 ;
        RECT 138.310 198.770 138.450 204.150 ;
        RECT 139.230 203.450 139.370 204.635 ;
        RECT 141.930 204.490 142.190 204.810 ;
        RECT 139.630 204.150 139.890 204.470 ;
        RECT 141.010 204.150 141.270 204.470 ;
        RECT 139.170 203.130 139.430 203.450 ;
        RECT 138.710 202.340 138.970 202.430 ;
        RECT 138.710 202.285 139.370 202.340 ;
        RECT 138.710 202.200 139.440 202.285 ;
        RECT 138.710 202.110 138.970 202.200 ;
        RECT 139.160 201.915 139.440 202.200 ;
        RECT 138.710 201.660 138.970 201.750 ;
        RECT 139.690 201.660 139.830 204.150 ;
        RECT 141.070 201.750 141.210 204.150 ;
        RECT 141.990 203.450 142.130 204.490 ;
        RECT 142.390 204.150 142.650 204.470 ;
        RECT 144.230 204.150 144.490 204.470 ;
        RECT 141.930 203.130 142.190 203.450 ;
        RECT 138.710 201.520 139.830 201.660 ;
        RECT 141.010 201.660 141.270 201.750 ;
        RECT 141.010 201.520 141.670 201.660 ;
        RECT 138.710 201.430 138.970 201.520 ;
        RECT 141.010 201.430 141.270 201.520 ;
        RECT 138.770 200.730 138.910 201.430 ;
        RECT 139.450 200.895 140.990 201.265 ;
        RECT 141.530 200.730 141.670 201.520 ;
        RECT 141.990 200.730 142.130 203.130 ;
        RECT 138.710 200.410 138.970 200.730 ;
        RECT 141.470 200.410 141.730 200.730 ;
        RECT 141.930 200.410 142.190 200.730 ;
        RECT 142.450 200.130 142.590 204.150 ;
        RECT 144.290 203.450 144.430 204.150 ;
        RECT 144.230 203.130 144.490 203.450 ;
        RECT 143.310 202.790 143.570 203.110 ;
        RECT 142.850 201.770 143.110 202.090 ;
        RECT 142.910 200.390 143.050 201.770 ;
        RECT 141.530 200.050 142.590 200.130 ;
        RECT 142.850 200.070 143.110 200.390 ;
        RECT 141.470 199.990 142.590 200.050 ;
        RECT 141.470 199.730 141.730 199.990 ;
        RECT 142.450 199.710 142.590 199.990 ;
        RECT 142.390 199.390 142.650 199.710 ;
        RECT 137.850 198.630 138.450 198.770 ;
        RECT 141.930 198.710 142.190 199.030 ;
        RECT 142.390 198.710 142.650 199.030 ;
        RECT 137.850 193.930 137.990 198.630 ;
        RECT 139.450 195.455 140.990 195.825 ;
        RECT 141.990 194.270 142.130 198.710 ;
        RECT 142.450 194.270 142.590 198.710 ;
        RECT 142.850 195.990 143.110 196.310 ;
        RECT 138.250 193.950 138.510 194.270 ;
        RECT 141.010 193.950 141.270 194.270 ;
        RECT 141.930 193.950 142.190 194.270 ;
        RECT 142.390 193.950 142.650 194.270 ;
        RECT 137.790 193.610 138.050 193.930 ;
        RECT 137.320 188.995 137.600 189.365 ;
        RECT 137.390 188.830 137.530 188.995 ;
        RECT 137.330 188.510 137.590 188.830 ;
        RECT 135.030 187.830 135.290 188.150 ;
        RECT 136.870 187.830 137.130 188.150 ;
        RECT 137.330 187.830 137.590 188.150 ;
        RECT 131.350 184.090 131.610 184.410 ;
        RECT 132.270 184.090 132.530 184.410 ;
        RECT 134.110 184.090 134.370 184.410 ;
        RECT 134.570 184.090 134.830 184.410 ;
        RECT 135.090 183.390 135.230 187.830 ;
        RECT 137.390 186.450 137.530 187.830 ;
        RECT 137.330 186.130 137.590 186.450 ;
        RECT 135.490 185.450 135.750 185.770 ;
        RECT 129.970 183.070 130.230 183.390 ;
        RECT 131.350 183.070 131.610 183.390 ;
        RECT 135.030 183.070 135.290 183.390 ;
        RECT 129.970 180.350 130.230 180.670 ;
        RECT 130.030 178.630 130.170 180.350 ;
        RECT 129.970 178.310 130.230 178.630 ;
        RECT 130.030 174.550 130.170 178.310 ;
        RECT 129.970 174.230 130.230 174.550 ;
        RECT 129.050 172.190 129.310 172.510 ;
        RECT 129.510 172.190 129.770 172.510 ;
        RECT 129.110 170.810 129.250 172.190 ;
        RECT 130.030 172.170 130.630 172.250 ;
        RECT 130.030 172.110 130.690 172.170 ;
        RECT 129.050 170.490 129.310 170.810 ;
        RECT 128.650 170.070 129.250 170.210 ;
        RECT 130.030 170.130 130.170 172.110 ;
        RECT 130.430 171.850 130.690 172.110 ;
        RECT 130.890 171.510 131.150 171.830 ;
        RECT 130.950 170.470 131.090 171.510 ;
        RECT 131.410 170.810 131.550 183.070 ;
        RECT 132.730 180.350 132.990 180.670 ;
        RECT 132.790 178.290 132.930 180.350 ;
        RECT 134.570 180.010 134.830 180.330 ;
        RECT 132.730 177.970 132.990 178.290 ;
        RECT 133.190 177.630 133.450 177.950 ;
        RECT 133.250 176.250 133.390 177.630 ;
        RECT 134.110 176.950 134.370 177.270 ;
        RECT 133.190 175.930 133.450 176.250 ;
        RECT 133.250 172.850 133.390 175.930 ;
        RECT 134.170 175.230 134.310 176.950 ;
        RECT 134.630 176.250 134.770 180.010 ;
        RECT 135.030 179.670 135.290 179.990 ;
        RECT 135.090 177.950 135.230 179.670 ;
        RECT 135.550 177.950 135.690 185.450 ;
        RECT 137.390 183.730 137.530 186.130 ;
        RECT 137.790 185.450 138.050 185.770 ;
        RECT 137.850 184.410 137.990 185.450 ;
        RECT 137.790 184.090 138.050 184.410 ;
        RECT 137.330 183.410 137.590 183.730 ;
        RECT 136.410 177.970 136.670 178.290 ;
        RECT 135.030 177.630 135.290 177.950 ;
        RECT 135.490 177.630 135.750 177.950 ;
        RECT 134.570 175.930 134.830 176.250 ;
        RECT 136.470 175.570 136.610 177.970 ;
        RECT 137.330 177.630 137.590 177.950 ;
        RECT 137.390 176.250 137.530 177.630 ;
        RECT 138.310 176.250 138.450 193.950 ;
        RECT 141.070 190.780 141.210 193.950 ;
        RECT 142.910 193.930 143.050 195.990 ;
        RECT 142.850 193.610 143.110 193.930 ;
        RECT 142.390 193.270 142.650 193.590 ;
        RECT 141.070 190.640 141.670 190.780 ;
        RECT 139.450 190.015 140.990 190.385 ;
        RECT 141.530 187.130 141.670 190.640 ;
        RECT 141.470 186.810 141.730 187.130 ;
        RECT 141.930 186.470 142.190 186.790 ;
        RECT 141.470 186.130 141.730 186.450 ;
        RECT 139.450 184.575 140.990 184.945 ;
        RECT 141.530 184.410 141.670 186.130 ;
        RECT 141.470 184.090 141.730 184.410 ;
        RECT 141.470 182.390 141.730 182.710 ;
        RECT 138.710 180.350 138.970 180.670 ;
        RECT 138.770 177.270 138.910 180.350 ;
        RECT 139.450 179.135 140.990 179.505 ;
        RECT 140.550 178.650 140.810 178.970 ;
        RECT 140.610 177.950 140.750 178.650 ;
        RECT 141.530 178.630 141.670 182.390 ;
        RECT 141.470 178.310 141.730 178.630 ;
        RECT 140.550 177.630 140.810 177.950 ;
        RECT 141.470 177.630 141.730 177.950 ;
        RECT 138.710 176.950 138.970 177.270 ;
        RECT 137.330 175.930 137.590 176.250 ;
        RECT 138.250 175.930 138.510 176.250 ;
        RECT 136.410 175.250 136.670 175.570 ;
        RECT 134.110 174.910 134.370 175.230 ;
        RECT 133.190 172.530 133.450 172.850 ;
        RECT 133.250 170.810 133.390 172.530 ;
        RECT 137.330 171.510 137.590 171.830 ;
        RECT 131.350 170.490 131.610 170.810 ;
        RECT 133.190 170.490 133.450 170.810 ;
        RECT 130.890 170.150 131.150 170.470 ;
        RECT 128.130 166.750 128.390 167.070 ;
        RECT 128.190 164.690 128.330 166.750 ;
        RECT 128.590 166.070 128.850 166.390 ;
        RECT 128.650 164.690 128.790 166.070 ;
        RECT 127.210 164.530 127.870 164.670 ;
        RECT 127.210 164.370 127.470 164.530 ;
        RECT 128.130 164.370 128.390 164.690 ;
        RECT 128.590 164.370 128.850 164.690 ;
        RECT 129.110 164.670 129.250 170.070 ;
        RECT 129.970 169.810 130.230 170.130 ;
        RECT 129.510 169.470 129.770 169.790 ;
        RECT 129.570 167.410 129.710 169.470 ;
        RECT 137.390 169.110 137.530 171.510 ;
        RECT 137.330 168.790 137.590 169.110 ;
        RECT 137.790 168.790 138.050 169.110 ;
        RECT 137.850 167.750 137.990 168.790 ;
        RECT 137.790 167.430 138.050 167.750 ;
        RECT 129.510 167.090 129.770 167.410 ;
        RECT 137.850 166.730 137.990 167.430 ;
        RECT 137.790 166.410 138.050 166.730 ;
        RECT 129.110 164.530 130.170 164.670 ;
        RECT 126.810 161.630 126.950 164.370 ;
        RECT 127.670 163.350 127.930 163.670 ;
        RECT 127.730 162.650 127.870 163.350 ;
        RECT 127.670 162.330 127.930 162.650 ;
        RECT 128.190 161.630 128.330 164.370 ;
        RECT 129.050 163.690 129.310 164.010 ;
        RECT 126.750 161.310 127.010 161.630 ;
        RECT 128.130 161.310 128.390 161.630 ;
        RECT 126.810 159.250 126.950 161.310 ;
        RECT 128.190 159.250 128.330 161.310 ;
        RECT 128.590 160.630 128.850 160.950 ;
        RECT 128.650 159.930 128.790 160.630 ;
        RECT 128.590 159.610 128.850 159.930 ;
        RECT 129.110 159.330 129.250 163.690 ;
        RECT 129.510 160.970 129.770 161.290 ;
        RECT 129.570 159.590 129.710 160.970 ;
        RECT 128.650 159.250 129.250 159.330 ;
        RECT 129.510 159.270 129.770 159.590 ;
        RECT 126.750 158.930 127.010 159.250 ;
        RECT 128.130 158.930 128.390 159.250 ;
        RECT 128.590 159.190 129.250 159.250 ;
        RECT 128.590 158.930 128.850 159.190 ;
        RECT 129.050 153.150 129.310 153.470 ;
        RECT 129.110 151.090 129.250 153.150 ;
        RECT 129.050 150.770 129.310 151.090 ;
        RECT 129.510 148.730 129.770 149.050 ;
        RECT 129.570 145.310 129.710 148.730 ;
        RECT 129.510 144.990 129.770 145.310 ;
        RECT 129.050 142.270 129.310 142.590 ;
        RECT 128.130 141.590 128.390 141.910 ;
        RECT 126.750 138.870 127.010 139.190 ;
        RECT 126.810 137.490 126.950 138.870 ;
        RECT 128.190 138.170 128.330 141.590 ;
        RECT 129.110 140.890 129.250 142.270 ;
        RECT 129.050 140.570 129.310 140.890 ;
        RECT 130.030 138.170 130.170 164.530 ;
        RECT 134.570 164.030 134.830 164.350 ;
        RECT 137.790 164.030 138.050 164.350 ;
        RECT 134.630 161.290 134.770 164.030 ;
        RECT 137.850 162.650 137.990 164.030 ;
        RECT 137.790 162.330 138.050 162.650 ;
        RECT 134.570 160.970 134.830 161.290 ;
        RECT 131.350 160.630 131.610 160.950 ;
        RECT 131.410 158.230 131.550 160.630 ;
        RECT 134.630 159.930 134.770 160.970 ;
        RECT 134.570 159.610 134.830 159.930 ;
        RECT 131.350 157.910 131.610 158.230 ;
        RECT 131.410 156.190 131.550 157.910 ;
        RECT 131.350 155.870 131.610 156.190 ;
        RECT 135.030 155.870 135.290 156.190 ;
        RECT 138.250 155.870 138.510 156.190 ;
        RECT 130.430 155.190 130.690 155.510 ;
        RECT 130.890 155.190 131.150 155.510 ;
        RECT 130.490 153.130 130.630 155.190 ;
        RECT 130.950 153.810 131.090 155.190 ;
        RECT 130.890 153.490 131.150 153.810 ;
        RECT 130.430 152.810 130.690 153.130 ;
        RECT 131.810 152.810 132.070 153.130 ;
        RECT 130.430 150.770 130.690 151.090 ;
        RECT 130.490 138.170 130.630 150.770 ;
        RECT 131.350 150.430 131.610 150.750 ;
        RECT 130.890 148.050 131.150 148.370 ;
        RECT 130.950 147.350 131.090 148.050 ;
        RECT 130.890 147.030 131.150 147.350 ;
        RECT 130.950 144.970 131.090 147.030 ;
        RECT 131.410 146.330 131.550 150.430 ;
        RECT 131.350 146.010 131.610 146.330 ;
        RECT 131.870 145.730 132.010 152.810 ;
        RECT 135.090 152.790 135.230 155.870 ;
        RECT 137.330 155.190 137.590 155.510 ;
        RECT 133.190 152.470 133.450 152.790 ;
        RECT 135.030 152.470 135.290 152.790 ;
        RECT 132.270 150.430 132.530 150.750 ;
        RECT 132.730 150.430 132.990 150.750 ;
        RECT 132.330 146.330 132.470 150.430 ;
        RECT 132.790 149.050 132.930 150.430 ;
        RECT 132.730 148.730 132.990 149.050 ;
        RECT 132.270 146.010 132.530 146.330 ;
        RECT 131.410 145.590 132.010 145.730 ;
        RECT 130.890 144.650 131.150 144.970 ;
        RECT 128.130 137.850 128.390 138.170 ;
        RECT 129.970 137.850 130.230 138.170 ;
        RECT 130.430 137.850 130.690 138.170 ;
        RECT 126.750 137.170 127.010 137.490 ;
        RECT 127.210 133.430 127.470 133.750 ;
        RECT 126.290 132.410 126.550 132.730 ;
        RECT 125.370 129.690 125.630 130.010 ;
        RECT 124.050 129.270 124.650 129.410 ;
        RECT 124.050 128.310 124.190 129.270 ;
        RECT 124.450 128.670 124.710 128.990 ;
        RECT 123.990 127.990 124.250 128.310 ;
        RECT 122.660 127.455 124.200 127.825 ;
        RECT 121.690 126.290 121.950 126.610 ;
        RECT 121.230 125.270 121.490 125.590 ;
        RECT 119.850 123.230 120.110 123.550 ;
        RECT 121.290 121.170 121.430 125.270 ;
        RECT 121.750 121.170 121.890 126.290 ;
        RECT 122.150 123.230 122.410 123.550 ;
        RECT 119.390 120.850 119.650 121.170 ;
        RECT 121.230 120.850 121.490 121.170 ;
        RECT 121.690 120.850 121.950 121.170 ;
        RECT 119.450 119.130 119.590 120.850 ;
        RECT 121.230 119.830 121.490 120.150 ;
        RECT 119.390 118.810 119.650 119.130 ;
        RECT 118.010 117.790 118.270 118.110 ;
        RECT 118.470 117.790 118.730 118.110 ;
        RECT 118.070 116.410 118.210 117.790 ;
        RECT 118.010 116.090 118.270 116.410 ;
        RECT 121.290 116.070 121.430 119.830 ;
        RECT 121.690 118.470 121.950 118.790 ;
        RECT 121.230 115.750 121.490 116.070 ;
        RECT 117.550 115.410 117.810 115.730 ;
        RECT 118.930 115.410 119.190 115.730 ;
        RECT 117.610 113.690 117.750 115.410 ;
        RECT 117.550 113.370 117.810 113.690 ;
        RECT 118.990 110.970 119.130 115.410 ;
        RECT 119.850 115.070 120.110 115.390 ;
        RECT 118.930 110.650 119.190 110.970 ;
        RECT 117.090 109.630 117.350 109.950 ;
        RECT 117.150 107.570 117.290 109.630 ;
        RECT 117.090 107.250 117.350 107.570 ;
        RECT 118.470 106.910 118.730 107.230 ;
        RECT 115.770 105.470 116.830 105.610 ;
        RECT 115.770 104.510 115.910 105.470 ;
        RECT 115.710 104.190 115.970 104.510 ;
        RECT 116.630 104.190 116.890 104.510 ;
        RECT 115.250 103.510 115.510 103.830 ;
        RECT 115.310 101.790 115.450 103.510 ;
        RECT 116.690 102.810 116.830 104.190 ;
        RECT 118.530 102.810 118.670 106.910 ;
        RECT 119.390 106.230 119.650 106.550 ;
        RECT 119.450 105.530 119.590 106.230 ;
        RECT 119.390 105.210 119.650 105.530 ;
        RECT 119.910 104.510 120.050 115.070 ;
        RECT 121.750 112.670 121.890 118.470 ;
        RECT 121.690 112.350 121.950 112.670 ;
        RECT 121.680 106.715 121.960 107.085 ;
        RECT 121.690 106.570 121.950 106.715 ;
        RECT 119.850 104.190 120.110 104.510 ;
        RECT 116.630 102.490 116.890 102.810 ;
        RECT 118.470 102.490 118.730 102.810 ;
        RECT 121.230 102.490 121.490 102.810 ;
        RECT 115.250 101.470 115.510 101.790 ;
        RECT 114.790 100.790 115.050 101.110 ;
        RECT 114.330 99.770 114.590 100.090 ;
        RECT 114.850 99.410 114.990 100.790 ;
        RECT 116.630 99.770 116.890 100.090 ;
        RECT 113.870 99.090 114.130 99.410 ;
        RECT 114.790 99.090 115.050 99.410 ;
        RECT 112.950 98.410 113.210 98.730 ;
        RECT 113.930 98.640 114.070 99.090 ;
        RECT 116.170 98.640 116.430 98.730 ;
        RECT 113.930 98.500 116.430 98.640 ;
        RECT 116.170 98.410 116.430 98.500 ;
        RECT 110.190 97.050 110.450 97.370 ;
        RECT 110.650 96.710 110.910 97.030 ;
        RECT 107.890 96.030 108.150 96.350 ;
        RECT 104.210 93.990 104.470 94.310 ;
        RECT 105.130 93.990 105.390 94.310 ;
        RECT 104.210 92.630 104.470 92.950 ;
        RECT 98.690 91.610 98.950 91.930 ;
        RECT 100.990 91.610 101.250 91.930 ;
        RECT 96.850 88.890 97.110 89.210 ;
        RECT 104.270 88.870 104.410 92.630 ;
        RECT 105.870 92.095 107.410 92.465 ;
        RECT 107.950 91.930 108.090 96.030 ;
        RECT 110.190 95.350 110.450 95.670 ;
        RECT 110.250 91.930 110.390 95.350 ;
        RECT 110.710 93.970 110.850 96.710 ;
        RECT 113.010 96.350 113.150 98.410 ;
        RECT 112.950 96.030 113.210 96.350 ;
        RECT 115.710 96.030 115.970 96.350 ;
        RECT 112.030 95.350 112.290 95.670 ;
        RECT 112.090 94.650 112.230 95.350 ;
        RECT 115.770 94.650 115.910 96.030 ;
        RECT 112.030 94.330 112.290 94.650 ;
        RECT 115.710 94.330 115.970 94.650 ;
        RECT 110.650 93.650 110.910 93.970 ;
        RECT 115.250 93.650 115.510 93.970 ;
        RECT 107.890 91.610 108.150 91.930 ;
        RECT 110.190 91.610 110.450 91.930 ;
        RECT 105.130 90.250 105.390 90.570 ;
        RECT 104.210 88.550 104.470 88.870 ;
        RECT 96.850 88.210 97.110 88.530 ;
        RECT 102.830 88.210 103.090 88.530 ;
        RECT 95.930 87.530 96.190 87.850 ;
        RECT 96.390 87.190 96.650 87.510 ;
        RECT 95.920 86.315 96.200 86.685 ;
        RECT 95.990 86.150 96.130 86.315 ;
        RECT 95.930 85.830 96.190 86.150 ;
        RECT 95.070 82.410 95.210 85.150 ;
        RECT 95.460 84.955 95.740 85.325 ;
        RECT 95.530 83.770 95.670 84.955 ;
        RECT 95.930 84.470 96.190 84.790 ;
        RECT 95.470 83.450 95.730 83.770 ;
        RECT 95.010 82.090 95.270 82.410 ;
        RECT 95.990 81.050 96.130 84.470 ;
        RECT 96.450 82.750 96.590 87.190 ;
        RECT 96.910 86.490 97.050 88.210 ;
        RECT 96.850 86.170 97.110 86.490 ;
        RECT 99.150 84.470 99.410 84.790 ;
        RECT 99.210 83.770 99.350 84.470 ;
        RECT 99.150 83.450 99.410 83.770 ;
        RECT 102.890 83.090 103.030 88.210 ;
        RECT 103.290 87.190 103.550 87.510 ;
        RECT 103.350 86.150 103.490 87.190 ;
        RECT 103.290 85.830 103.550 86.150 ;
        RECT 104.270 83.090 104.410 88.550 ;
        RECT 105.190 86.490 105.330 90.250 ;
        RECT 110.250 88.530 110.390 91.610 ;
        RECT 115.310 91.250 115.450 93.650 ;
        RECT 115.250 90.930 115.510 91.250 ;
        RECT 115.770 90.910 115.910 94.330 ;
        RECT 116.230 93.970 116.370 98.410 ;
        RECT 116.690 93.970 116.830 99.770 ;
        RECT 117.550 99.430 117.810 99.750 ;
        RECT 117.090 95.350 117.350 95.670 ;
        RECT 116.170 93.650 116.430 93.970 ;
        RECT 116.630 93.650 116.890 93.970 ;
        RECT 115.710 90.590 115.970 90.910 ;
        RECT 116.230 90.570 116.370 93.650 ;
        RECT 116.690 90.910 116.830 93.650 ;
        RECT 117.150 93.290 117.290 95.350 ;
        RECT 117.090 92.970 117.350 93.290 ;
        RECT 116.630 90.590 116.890 90.910 ;
        RECT 116.170 90.250 116.430 90.570 ;
        RECT 110.190 88.210 110.450 88.530 ;
        RECT 115.250 88.210 115.510 88.530 ;
        RECT 109.730 87.870 109.990 88.190 ;
        RECT 105.870 86.655 107.410 87.025 ;
        RECT 105.130 86.170 105.390 86.490 ;
        RECT 107.890 85.150 108.150 85.470 ;
        RECT 107.950 83.770 108.090 85.150 ;
        RECT 108.350 84.810 108.610 85.130 ;
        RECT 108.410 83.770 108.550 84.810 ;
        RECT 107.890 83.450 108.150 83.770 ;
        RECT 108.350 83.450 108.610 83.770 ;
        RECT 109.790 83.090 109.930 87.870 ;
        RECT 111.570 87.530 111.830 87.850 ;
        RECT 110.190 85.150 110.450 85.470 ;
        RECT 110.250 83.090 110.390 85.150 ;
        RECT 111.630 83.770 111.770 87.530 ;
        RECT 112.030 87.190 112.290 87.510 ;
        RECT 112.090 86.490 112.230 87.190 ;
        RECT 115.310 86.490 115.450 88.210 ;
        RECT 112.030 86.170 112.290 86.490 ;
        RECT 115.250 86.170 115.510 86.490 ;
        RECT 117.150 85.470 117.290 92.970 ;
        RECT 117.610 88.530 117.750 99.430 ;
        RECT 121.290 99.410 121.430 102.490 ;
        RECT 121.230 99.090 121.490 99.410 ;
        RECT 118.010 96.370 118.270 96.690 ;
        RECT 118.070 91.590 118.210 96.370 ;
        RECT 122.210 96.350 122.350 123.230 ;
        RECT 124.510 122.870 124.650 128.670 ;
        RECT 126.350 126.950 126.490 132.410 ;
        RECT 126.290 126.630 126.550 126.950 ;
        RECT 124.910 125.270 125.170 125.590 ;
        RECT 124.450 122.550 124.710 122.870 ;
        RECT 122.660 122.015 124.200 122.385 ;
        RECT 124.510 121.510 124.650 122.550 ;
        RECT 124.450 121.190 124.710 121.510 ;
        RECT 124.970 121.250 125.110 125.270 ;
        RECT 125.370 122.890 125.630 123.210 ;
        RECT 125.430 121.850 125.570 122.890 ;
        RECT 125.370 121.530 125.630 121.850 ;
        RECT 122.610 120.850 122.870 121.170 ;
        RECT 124.970 121.110 125.570 121.250 ;
        RECT 122.670 118.110 122.810 120.850 ;
        RECT 125.430 120.490 125.570 121.110 ;
        RECT 126.290 120.850 126.550 121.170 ;
        RECT 125.370 120.170 125.630 120.490 ;
        RECT 123.070 119.830 123.330 120.150 ;
        RECT 123.130 118.450 123.270 119.830 ;
        RECT 123.070 118.130 123.330 118.450 ;
        RECT 122.610 117.790 122.870 118.110 ;
        RECT 123.530 118.020 123.790 118.110 ;
        RECT 123.530 117.880 124.650 118.020 ;
        RECT 123.530 117.790 123.790 117.880 ;
        RECT 122.660 116.575 124.200 116.945 ;
        RECT 124.510 116.410 124.650 117.880 ;
        RECT 125.430 117.770 125.570 120.170 ;
        RECT 125.370 117.450 125.630 117.770 ;
        RECT 125.830 117.450 126.090 117.770 ;
        RECT 124.910 117.170 125.170 117.430 ;
        RECT 125.890 117.170 126.030 117.450 ;
        RECT 124.910 117.110 126.030 117.170 ;
        RECT 124.970 117.030 126.030 117.110 ;
        RECT 124.450 116.090 124.710 116.410 ;
        RECT 126.350 115.730 126.490 120.850 ;
        RECT 127.270 120.570 127.410 133.430 ;
        RECT 129.510 130.710 129.770 131.030 ;
        RECT 129.570 128.990 129.710 130.710 ;
        RECT 129.510 128.670 129.770 128.990 ;
        RECT 127.670 125.270 127.930 125.590 ;
        RECT 127.730 121.170 127.870 125.270 ;
        RECT 127.670 120.850 127.930 121.170 ;
        RECT 127.270 120.430 127.870 120.570 ;
        RECT 127.210 117.110 127.470 117.430 ;
        RECT 127.270 115.810 127.410 117.110 ;
        RECT 127.730 116.370 127.870 120.430 ;
        RECT 130.030 116.410 130.170 137.850 ;
        RECT 131.410 131.370 131.550 145.590 ;
        RECT 132.270 142.610 132.530 142.930 ;
        RECT 132.330 140.550 132.470 142.610 ;
        RECT 132.730 141.590 132.990 141.910 ;
        RECT 132.270 140.230 132.530 140.550 ;
        RECT 131.810 138.870 132.070 139.190 ;
        RECT 131.870 138.170 132.010 138.870 ;
        RECT 132.790 138.170 132.930 141.590 ;
        RECT 131.810 137.850 132.070 138.170 ;
        RECT 132.730 137.850 132.990 138.170 ;
        RECT 131.810 136.150 132.070 136.470 ;
        RECT 131.350 131.050 131.610 131.370 ;
        RECT 131.350 127.990 131.610 128.310 ;
        RECT 131.410 127.290 131.550 127.990 ;
        RECT 131.870 127.290 132.010 136.150 ;
        RECT 133.250 134.430 133.390 152.470 ;
        RECT 133.650 151.110 133.910 151.430 ;
        RECT 133.710 146.330 133.850 151.110 ;
        RECT 134.110 149.750 134.370 150.070 ;
        RECT 134.170 147.690 134.310 149.750 ;
        RECT 135.090 148.370 135.230 152.470 ;
        RECT 136.870 150.090 137.130 150.410 ;
        RECT 135.490 149.750 135.750 150.070 ;
        RECT 135.550 149.050 135.690 149.750 ;
        RECT 135.490 148.730 135.750 149.050 ;
        RECT 135.030 148.050 135.290 148.370 ;
        RECT 134.110 147.370 134.370 147.690 ;
        RECT 134.170 146.330 134.310 147.370 ;
        RECT 133.650 146.010 133.910 146.330 ;
        RECT 134.110 146.010 134.370 146.330 ;
        RECT 133.710 143.690 133.850 146.010 ;
        RECT 135.550 145.310 135.690 148.730 ;
        RECT 136.930 147.770 137.070 150.090 ;
        RECT 137.390 148.710 137.530 155.190 ;
        RECT 138.310 151.770 138.450 155.870 ;
        RECT 137.790 151.450 138.050 151.770 ;
        RECT 138.250 151.450 138.510 151.770 ;
        RECT 137.330 148.390 137.590 148.710 ;
        RECT 136.930 147.630 137.530 147.770 ;
        RECT 137.390 145.730 137.530 147.630 ;
        RECT 137.850 146.330 137.990 151.450 ;
        RECT 137.790 146.010 138.050 146.330 ;
        RECT 137.390 145.590 137.990 145.730 ;
        RECT 135.490 144.990 135.750 145.310 ;
        RECT 135.950 144.990 136.210 145.310 ;
        RECT 136.410 144.990 136.670 145.310 ;
        RECT 133.710 143.550 134.310 143.690 ;
        RECT 136.010 143.610 136.150 144.990 ;
        RECT 133.650 142.610 133.910 142.930 ;
        RECT 133.710 140.550 133.850 142.610 ;
        RECT 133.650 140.230 133.910 140.550 ;
        RECT 134.170 139.870 134.310 143.550 ;
        RECT 135.950 143.290 136.210 143.610 ;
        RECT 136.010 139.870 136.150 143.290 ;
        RECT 136.470 142.330 136.610 144.990 ;
        RECT 137.850 143.270 137.990 145.590 ;
        RECT 137.790 142.950 138.050 143.270 ;
        RECT 136.470 142.190 137.070 142.330 ;
        RECT 136.410 141.590 136.670 141.910 ;
        RECT 136.470 139.870 136.610 141.590 ;
        RECT 134.110 139.550 134.370 139.870 ;
        RECT 135.950 139.550 136.210 139.870 ;
        RECT 136.410 139.550 136.670 139.870 ;
        RECT 135.030 138.870 135.290 139.190 ;
        RECT 135.490 138.870 135.750 139.190 ;
        RECT 135.090 138.170 135.230 138.870 ;
        RECT 135.030 137.850 135.290 138.170 ;
        RECT 135.030 137.170 135.290 137.490 ;
        RECT 135.090 136.810 135.230 137.170 ;
        RECT 135.030 136.490 135.290 136.810 ;
        RECT 135.550 136.470 135.690 138.870 ;
        RECT 136.930 136.890 137.070 142.190 ;
        RECT 136.010 136.750 137.070 136.890 ;
        RECT 135.490 136.150 135.750 136.470 ;
        RECT 133.190 134.110 133.450 134.430 ;
        RECT 133.250 132.050 133.390 134.110 ;
        RECT 133.190 131.730 133.450 132.050 ;
        RECT 134.570 131.390 134.830 131.710 ;
        RECT 134.630 129.670 134.770 131.390 ;
        RECT 134.570 129.350 134.830 129.670 ;
        RECT 136.010 129.410 136.150 136.750 ;
        RECT 136.410 136.150 136.670 136.470 ;
        RECT 136.870 136.150 137.130 136.470 ;
        RECT 136.470 132.730 136.610 136.150 ;
        RECT 136.410 132.410 136.670 132.730 ;
        RECT 136.410 131.390 136.670 131.710 ;
        RECT 136.470 130.010 136.610 131.390 ;
        RECT 136.410 129.690 136.670 130.010 ;
        RECT 136.010 129.270 136.610 129.410 ;
        RECT 134.110 128.670 134.370 128.990 ;
        RECT 131.350 126.970 131.610 127.290 ;
        RECT 131.810 126.970 132.070 127.290 ;
        RECT 131.350 125.270 131.610 125.590 ;
        RECT 132.270 125.270 132.530 125.590 ;
        RECT 127.730 116.230 128.330 116.370 ;
        RECT 127.670 115.810 127.930 116.070 ;
        RECT 127.270 115.750 127.930 115.810 ;
        RECT 126.290 115.410 126.550 115.730 ;
        RECT 127.270 115.670 127.870 115.750 ;
        RECT 126.350 113.690 126.490 115.410 ;
        RECT 126.290 113.370 126.550 113.690 ;
        RECT 122.660 111.135 124.200 111.505 ;
        RECT 126.290 107.250 126.550 107.570 ;
        RECT 124.450 106.910 124.710 107.230 ;
        RECT 122.660 105.695 124.200 106.065 ;
        RECT 124.510 102.810 124.650 106.910 ;
        RECT 124.910 106.230 125.170 106.550 ;
        RECT 125.370 106.230 125.630 106.550 ;
        RECT 124.970 103.830 125.110 106.230 ;
        RECT 125.430 104.510 125.570 106.230 ;
        RECT 126.350 105.530 126.490 107.250 ;
        RECT 127.670 107.140 127.930 107.230 ;
        RECT 128.190 107.140 128.330 116.230 ;
        RECT 129.970 116.090 130.230 116.410 ;
        RECT 131.410 107.570 131.550 125.270 ;
        RECT 132.330 121.170 132.470 125.270 ;
        RECT 133.650 124.250 133.910 124.570 ;
        RECT 132.270 120.850 132.530 121.170 ;
        RECT 132.270 117.790 132.530 118.110 ;
        RECT 132.330 116.410 132.470 117.790 ;
        RECT 132.730 117.110 132.990 117.430 ;
        RECT 132.270 116.090 132.530 116.410 ;
        RECT 132.790 112.670 132.930 117.110 ;
        RECT 132.730 112.350 132.990 112.670 ;
        RECT 131.350 107.250 131.610 107.570 ;
        RECT 127.670 107.000 128.330 107.140 ;
        RECT 127.670 106.910 127.930 107.000 ;
        RECT 129.510 106.910 129.770 107.230 ;
        RECT 130.890 106.910 131.150 107.230 ;
        RECT 126.290 105.210 126.550 105.530 ;
        RECT 125.830 104.870 126.090 105.190 ;
        RECT 125.370 104.190 125.630 104.510 ;
        RECT 124.910 103.510 125.170 103.830 ;
        RECT 124.450 102.490 124.710 102.810 ;
        RECT 124.970 101.110 125.110 103.510 ;
        RECT 125.430 102.810 125.570 104.190 ;
        RECT 125.370 102.490 125.630 102.810 ;
        RECT 124.910 100.790 125.170 101.110 ;
        RECT 122.660 100.255 124.200 100.625 ;
        RECT 123.070 98.750 123.330 99.070 ;
        RECT 123.130 96.690 123.270 98.750 ;
        RECT 123.070 96.370 123.330 96.690 ;
        RECT 122.150 96.030 122.410 96.350 ;
        RECT 124.450 95.350 124.710 95.670 ;
        RECT 122.660 94.815 124.200 95.185 ;
        RECT 124.510 94.650 124.650 95.350 ;
        RECT 124.450 94.330 124.710 94.650 ;
        RECT 122.150 92.630 122.410 92.950 ;
        RECT 118.010 91.270 118.270 91.590 ;
        RECT 121.690 89.910 121.950 90.230 ;
        RECT 119.390 88.550 119.650 88.870 ;
        RECT 117.550 88.210 117.810 88.530 ;
        RECT 118.930 88.210 119.190 88.530 ;
        RECT 117.550 87.190 117.810 87.510 ;
        RECT 117.090 85.150 117.350 85.470 ;
        RECT 114.330 84.470 114.590 84.790 ;
        RECT 114.390 83.770 114.530 84.470 ;
        RECT 111.570 83.450 111.830 83.770 ;
        RECT 114.330 83.450 114.590 83.770 ;
        RECT 102.830 82.770 103.090 83.090 ;
        RECT 104.210 82.770 104.470 83.090 ;
        RECT 109.730 82.770 109.990 83.090 ;
        RECT 110.190 82.770 110.450 83.090 ;
        RECT 110.650 82.770 110.910 83.090 ;
        RECT 96.390 82.430 96.650 82.750 ;
        RECT 97.770 81.750 98.030 82.070 ;
        RECT 95.930 80.730 96.190 81.050 ;
        RECT 97.830 80.030 97.970 81.750 ;
        RECT 102.890 81.050 103.030 82.770 ;
        RECT 105.870 81.215 107.410 81.585 ;
        RECT 102.830 80.730 103.090 81.050 ;
        RECT 96.390 79.710 96.650 80.030 ;
        RECT 97.770 79.710 98.030 80.030 ;
        RECT 96.450 78.330 96.590 79.710 ;
        RECT 110.250 78.330 110.390 82.770 ;
        RECT 110.710 82.410 110.850 82.770 ;
        RECT 110.650 82.090 110.910 82.410 ;
        RECT 92.310 72.660 92.910 72.800 ;
        RECT 93.230 78.100 93.830 78.240 ;
        RECT 91.790 71.890 92.050 72.210 ;
        RECT 91.330 71.550 91.590 71.870 ;
        RECT 91.850 71.530 91.990 71.890 ;
        RECT 91.790 71.210 92.050 71.530 ;
        RECT 89.030 69.850 89.290 70.170 ;
        RECT 90.870 69.850 91.130 70.170 ;
        RECT 91.850 69.830 91.990 71.210 ;
        RECT 92.310 71.190 92.450 72.660 ;
        RECT 92.710 71.890 92.970 72.210 ;
        RECT 92.250 70.870 92.510 71.190 ;
        RECT 90.410 69.570 90.670 69.830 ;
        RECT 90.410 69.510 91.070 69.570 ;
        RECT 91.790 69.510 92.050 69.830 ;
        RECT 90.470 69.430 91.070 69.510 ;
        RECT 88.570 68.830 88.830 69.150 ;
        RECT 89.030 68.830 89.290 69.150 ;
        RECT 89.090 68.380 89.230 68.830 ;
        RECT 90.930 68.810 91.070 69.430 ;
        RECT 91.330 68.830 91.590 69.150 ;
        RECT 90.870 68.490 91.130 68.810 ;
        RECT 88.630 68.240 89.230 68.380 ;
        RECT 88.630 67.450 88.770 68.240 ;
        RECT 89.080 67.615 90.620 67.985 ;
        RECT 88.570 67.360 88.830 67.450 ;
        RECT 88.570 67.220 89.230 67.360 ;
        RECT 88.570 67.130 88.830 67.220 ;
        RECT 83.510 66.540 84.170 66.680 ;
        RECT 83.510 66.450 83.770 66.540 ;
        RECT 84.430 66.450 84.690 66.770 ;
        RECT 88.110 66.450 88.370 66.770 ;
        RECT 74.770 65.770 75.030 66.090 ;
        RECT 83.050 65.770 83.310 66.090 ;
        RECT 74.830 64.640 74.970 65.770 ;
        RECT 79.370 65.430 79.630 65.750 ;
        RECT 79.830 65.430 80.090 65.750 ;
        RECT 75.230 64.640 75.490 64.730 ;
        RECT 74.830 64.500 75.490 64.640 ;
        RECT 75.230 64.410 75.490 64.500 ;
        RECT 73.850 63.480 74.510 63.620 ;
        RECT 73.850 63.390 74.110 63.480 ;
        RECT 77.990 63.390 78.250 63.710 ;
        RECT 78.450 63.390 78.710 63.710 ;
        RECT 71.550 63.050 71.810 63.370 ;
        RECT 69.250 61.100 70.370 61.240 ;
        RECT 69.250 61.010 69.510 61.100 ;
        RECT 71.610 59.290 71.750 63.050 ;
        RECT 75.690 62.710 75.950 63.030 ;
        RECT 73.390 61.240 73.650 61.330 ;
        RECT 73.390 61.100 74.510 61.240 ;
        RECT 73.390 61.010 73.650 61.100 ;
        RECT 72.290 59.455 73.830 59.825 ;
        RECT 71.550 58.970 71.810 59.290 ;
        RECT 68.330 58.040 68.990 58.180 ;
        RECT 68.330 57.950 68.590 58.040 ;
        RECT 70.170 57.950 70.430 58.270 ;
        RECT 70.230 56.200 70.370 57.950 ;
        RECT 72.990 56.510 73.590 56.650 ;
        RECT 72.990 56.200 73.130 56.510 ;
        RECT 55.050 55.830 56.110 55.970 ;
        RECT 50.840 54.200 51.130 54.830 ;
        RECT 53.600 54.200 53.890 55.000 ;
        RECT 56.360 54.810 56.640 56.200 ;
        RECT 59.120 54.850 59.400 56.200 ;
        RECT 56.360 54.200 56.650 54.810 ;
        RECT 59.120 54.200 59.410 54.850 ;
        RECT 61.880 54.710 62.160 56.200 ;
        RECT 61.880 54.200 62.170 54.710 ;
        RECT 64.640 54.700 64.920 56.200 ;
        RECT 64.640 54.200 64.930 54.700 ;
        RECT 67.400 54.500 67.680 56.200 ;
        RECT 70.160 54.660 70.440 56.200 ;
        RECT 72.920 54.900 73.200 56.200 ;
        RECT 73.450 55.970 73.590 56.510 ;
        RECT 74.370 55.970 74.510 61.100 ;
        RECT 75.230 60.670 75.490 60.990 ;
        RECT 75.290 59.290 75.430 60.670 ;
        RECT 75.230 58.970 75.490 59.290 ;
        RECT 75.750 56.200 75.890 62.710 ;
        RECT 78.050 58.690 78.190 63.390 ;
        RECT 78.510 59.290 78.650 63.390 ;
        RECT 79.430 62.010 79.570 65.430 ;
        RECT 79.890 63.710 80.030 65.430 ;
        RECT 79.830 63.390 80.090 63.710 ;
        RECT 79.370 61.690 79.630 62.010 ;
        RECT 83.110 61.330 83.250 65.770 ;
        RECT 83.510 65.430 83.770 65.750 ;
        RECT 80.750 61.240 81.010 61.330 ;
        RECT 80.750 61.100 81.410 61.240 ;
        RECT 80.750 61.010 81.010 61.100 ;
        RECT 78.450 58.970 78.710 59.290 ;
        RECT 78.050 58.550 78.650 58.690 ;
        RECT 78.510 56.200 78.650 58.550 ;
        RECT 81.270 56.200 81.410 61.100 ;
        RECT 83.050 61.010 83.310 61.330 ;
        RECT 83.570 58.270 83.710 65.430 ;
        RECT 83.970 63.390 84.230 63.710 ;
        RECT 84.430 63.390 84.690 63.710 ;
        RECT 85.810 63.390 86.070 63.710 ;
        RECT 89.090 63.450 89.230 67.220 ;
        RECT 90.930 66.770 91.070 68.490 ;
        RECT 91.390 66.770 91.530 68.830 ;
        RECT 92.770 68.070 92.910 71.890 ;
        RECT 93.230 71.725 93.370 78.100 ;
        RECT 96.390 78.010 96.650 78.330 ;
        RECT 110.190 78.010 110.450 78.330 ;
        RECT 93.630 77.330 93.890 77.650 ;
        RECT 94.550 77.330 94.810 77.650 ;
        RECT 102.830 77.330 103.090 77.650 ;
        RECT 107.890 77.330 108.150 77.650 ;
        RECT 108.350 77.330 108.610 77.650 ;
        RECT 93.160 71.355 93.440 71.725 ;
        RECT 92.770 67.930 93.370 68.070 ;
        RECT 90.870 66.450 91.130 66.770 ;
        RECT 91.330 66.450 91.590 66.770 ;
        RECT 93.230 66.090 93.370 67.930 ;
        RECT 93.170 65.770 93.430 66.090 ;
        RECT 93.690 65.750 93.830 77.330 ;
        RECT 94.610 72.890 94.750 77.330 ;
        RECT 95.010 74.950 95.270 75.270 ;
        RECT 94.550 72.570 94.810 72.890 ;
        RECT 94.090 71.890 94.350 72.210 ;
        RECT 93.630 65.430 93.890 65.750 ;
        RECT 83.510 57.950 83.770 58.270 ;
        RECT 84.030 56.200 84.170 63.390 ;
        RECT 84.490 61.330 84.630 63.390 ;
        RECT 84.430 61.010 84.690 61.330 ;
        RECT 85.870 59.290 86.010 63.390 ;
        RECT 88.630 63.310 89.230 63.450 ;
        RECT 90.870 63.390 91.130 63.710 ;
        RECT 93.170 63.390 93.430 63.710 ;
        RECT 88.630 61.330 88.770 63.310 ;
        RECT 89.080 62.175 90.620 62.545 ;
        RECT 88.110 61.010 88.370 61.330 ;
        RECT 88.570 61.010 88.830 61.330 ;
        RECT 87.190 60.670 87.450 60.990 ;
        RECT 87.250 59.290 87.390 60.670 ;
        RECT 85.810 58.970 86.070 59.290 ;
        RECT 87.190 58.970 87.450 59.290 ;
        RECT 86.730 57.950 86.990 58.270 ;
        RECT 86.790 56.200 86.930 57.950 ;
        RECT 88.170 56.480 88.310 61.010 ;
        RECT 90.930 59.290 91.070 63.390 ;
        RECT 93.230 61.330 93.370 63.390 ;
        RECT 92.710 61.240 92.970 61.330 ;
        RECT 92.310 61.100 92.970 61.240 ;
        RECT 90.870 58.970 91.130 59.290 ;
        RECT 89.080 56.735 90.620 57.105 ;
        RECT 88.170 56.340 89.690 56.480 ;
        RECT 89.550 56.200 89.690 56.340 ;
        RECT 92.310 56.200 92.450 61.100 ;
        RECT 92.710 61.010 92.970 61.100 ;
        RECT 93.170 61.010 93.430 61.330 ;
        RECT 94.150 58.270 94.290 71.890 ;
        RECT 94.550 71.550 94.810 71.870 ;
        RECT 94.610 71.045 94.750 71.550 ;
        RECT 94.540 70.675 94.820 71.045 ;
        RECT 95.070 69.150 95.210 74.950 ;
        RECT 102.890 74.590 103.030 77.330 ;
        RECT 105.870 75.775 107.410 76.145 ;
        RECT 96.390 74.270 96.650 74.590 ;
        RECT 97.770 74.270 98.030 74.590 ;
        RECT 102.830 74.270 103.090 74.590 ;
        RECT 96.450 72.890 96.590 74.270 ;
        RECT 96.850 73.590 97.110 73.910 ;
        RECT 96.390 72.570 96.650 72.890 ;
        RECT 96.910 72.210 97.050 73.590 ;
        RECT 96.850 71.890 97.110 72.210 ;
        RECT 95.470 70.870 95.730 71.190 ;
        RECT 97.310 70.870 97.570 71.190 ;
        RECT 95.530 70.170 95.670 70.870 ;
        RECT 97.370 70.170 97.510 70.870 ;
        RECT 97.830 70.170 97.970 74.270 ;
        RECT 107.950 74.250 108.090 77.330 ;
        RECT 108.410 75.610 108.550 77.330 ;
        RECT 109.270 76.990 109.530 77.310 ;
        RECT 108.350 75.290 108.610 75.610 ;
        RECT 107.890 73.930 108.150 74.250 ;
        RECT 98.230 71.890 98.490 72.210 ;
        RECT 98.680 72.035 98.960 72.405 ;
        RECT 98.690 71.890 98.950 72.035 ;
        RECT 98.290 71.100 98.430 71.890 ;
        RECT 107.950 71.870 108.090 73.930 ;
        RECT 108.410 72.890 108.550 75.290 ;
        RECT 109.330 74.590 109.470 76.990 ;
        RECT 110.710 76.970 110.850 82.090 ;
        RECT 113.410 80.390 113.670 80.710 ;
        RECT 110.650 76.650 110.910 76.970 ;
        RECT 111.110 76.310 111.370 76.630 ;
        RECT 111.170 75.270 111.310 76.310 ;
        RECT 111.110 74.950 111.370 75.270 ;
        RECT 109.270 74.270 109.530 74.590 ;
        RECT 109.330 73.910 109.470 74.270 ;
        RECT 113.470 74.250 113.610 80.390 ;
        RECT 116.630 77.330 116.890 77.650 ;
        RECT 116.690 75.610 116.830 77.330 ;
        RECT 117.150 76.630 117.290 85.150 ;
        RECT 117.610 85.130 117.750 87.190 ;
        RECT 117.550 84.810 117.810 85.130 ;
        RECT 118.990 80.030 119.130 88.210 ;
        RECT 118.930 79.710 119.190 80.030 ;
        RECT 118.470 77.330 118.730 77.650 ;
        RECT 117.090 76.310 117.350 76.630 ;
        RECT 116.630 75.290 116.890 75.610 ;
        RECT 113.410 73.930 113.670 74.250 ;
        RECT 109.270 73.590 109.530 73.910 ;
        RECT 110.190 73.590 110.450 73.910 ;
        RECT 108.350 72.570 108.610 72.890 ;
        RECT 109.330 72.210 109.470 73.590 ;
        RECT 110.250 72.890 110.390 73.590 ;
        RECT 110.190 72.570 110.450 72.890 ;
        RECT 109.270 71.890 109.530 72.210 ;
        RECT 107.890 71.550 108.150 71.870 ;
        RECT 98.290 70.960 99.810 71.100 ;
        RECT 95.470 69.850 95.730 70.170 ;
        RECT 97.310 69.850 97.570 70.170 ;
        RECT 97.770 69.850 98.030 70.170 ;
        RECT 95.010 68.830 95.270 69.150 ;
        RECT 97.370 67.450 97.510 69.850 ;
        RECT 99.150 68.490 99.410 68.810 ;
        RECT 97.310 67.130 97.570 67.450 ;
        RECT 96.850 66.790 97.110 67.110 ;
        RECT 95.010 66.450 95.270 66.770 ;
        RECT 94.550 65.430 94.810 65.750 ;
        RECT 94.610 61.330 94.750 65.430 ;
        RECT 95.070 64.730 95.210 66.450 ;
        RECT 95.010 64.410 95.270 64.730 ;
        RECT 96.910 63.710 97.050 66.790 ;
        RECT 96.850 63.390 97.110 63.710 ;
        RECT 99.210 61.330 99.350 68.490 ;
        RECT 94.550 61.010 94.810 61.330 ;
        RECT 98.690 61.240 98.950 61.330 ;
        RECT 97.830 61.100 98.950 61.240 ;
        RECT 94.090 57.950 94.350 58.270 ;
        RECT 95.010 57.950 95.270 58.270 ;
        RECT 95.070 56.200 95.210 57.950 ;
        RECT 97.830 56.200 97.970 61.100 ;
        RECT 98.690 61.010 98.950 61.100 ;
        RECT 99.150 61.010 99.410 61.330 ;
        RECT 99.670 57.930 99.810 70.960 ;
        RECT 102.370 70.870 102.630 71.190 ;
        RECT 105.130 70.870 105.390 71.190 ;
        RECT 102.430 70.170 102.570 70.870 ;
        RECT 102.370 69.850 102.630 70.170 ;
        RECT 100.990 68.830 101.250 69.150 ;
        RECT 101.050 66.770 101.190 68.830 ;
        RECT 100.990 66.450 101.250 66.770 ;
        RECT 104.670 66.450 104.930 66.770 ;
        RECT 104.730 64.730 104.870 66.450 ;
        RECT 104.670 64.410 104.930 64.730 ;
        RECT 101.450 63.620 101.710 63.710 ;
        RECT 101.050 63.480 101.710 63.620 ;
        RECT 100.530 60.670 100.790 60.990 ;
        RECT 100.590 59.290 100.730 60.670 ;
        RECT 100.530 58.970 100.790 59.290 ;
        RECT 101.050 58.690 101.190 63.480 ;
        RECT 101.450 63.390 101.710 63.480 ;
        RECT 101.910 63.390 102.170 63.710 ;
        RECT 100.590 58.550 101.190 58.690 ;
        RECT 99.610 57.610 99.870 57.930 ;
        RECT 100.590 56.200 100.730 58.550 ;
        RECT 101.970 58.270 102.110 63.390 ;
        RECT 105.190 61.670 105.330 70.870 ;
        RECT 105.870 70.335 107.410 70.705 ;
        RECT 107.950 70.170 108.090 71.550 ;
        RECT 108.350 70.870 108.610 71.190 ;
        RECT 107.890 69.850 108.150 70.170 ;
        RECT 108.410 69.570 108.550 70.870 ;
        RECT 113.470 70.170 113.610 73.930 ;
        RECT 116.630 72.570 116.890 72.890 ;
        RECT 116.690 70.250 116.830 72.570 ;
        RECT 117.150 71.190 117.290 76.310 ;
        RECT 118.530 72.890 118.670 77.330 ;
        RECT 118.930 73.590 119.190 73.910 ;
        RECT 118.990 72.890 119.130 73.590 ;
        RECT 118.470 72.570 118.730 72.890 ;
        RECT 118.930 72.570 119.190 72.890 ;
        RECT 117.550 71.210 117.810 71.530 ;
        RECT 117.090 70.870 117.350 71.190 ;
        RECT 113.410 69.850 113.670 70.170 ;
        RECT 116.230 70.110 116.830 70.250 ;
        RECT 107.950 69.430 108.550 69.570 ;
        RECT 107.950 67.110 108.090 69.430 ;
        RECT 110.650 69.060 110.910 69.150 ;
        RECT 110.650 68.920 111.310 69.060 ;
        RECT 110.650 68.830 110.910 68.920 ;
        RECT 108.350 68.150 108.610 68.470 ;
        RECT 110.650 68.150 110.910 68.470 ;
        RECT 107.890 66.790 108.150 67.110 ;
        RECT 105.870 64.895 107.410 65.265 ;
        RECT 108.410 63.710 108.550 68.150 ;
        RECT 110.710 66.430 110.850 68.150 ;
        RECT 111.170 66.770 111.310 68.920 ;
        RECT 111.570 68.830 111.830 69.150 ;
        RECT 111.630 67.110 111.770 68.830 ;
        RECT 113.470 68.810 113.610 69.850 ;
        RECT 116.230 69.830 116.370 70.110 ;
        RECT 116.170 69.510 116.430 69.830 ;
        RECT 116.630 69.510 116.890 69.830 ;
        RECT 116.690 68.890 116.830 69.510 ;
        RECT 117.610 68.890 117.750 71.210 ;
        RECT 118.470 70.870 118.730 71.190 ;
        RECT 118.530 69.150 118.670 70.870 ;
        RECT 119.450 69.830 119.590 88.550 ;
        RECT 119.850 87.190 120.110 87.510 ;
        RECT 119.910 86.490 120.050 87.190 ;
        RECT 119.850 86.170 120.110 86.490 ;
        RECT 119.850 80.730 120.110 81.050 ;
        RECT 119.910 74.590 120.050 80.730 ;
        RECT 121.750 80.030 121.890 89.910 ;
        RECT 122.210 88.870 122.350 92.630 ;
        RECT 122.660 89.375 124.200 89.745 ;
        RECT 122.150 88.550 122.410 88.870 ;
        RECT 124.970 86.490 125.110 100.790 ;
        RECT 125.370 98.070 125.630 98.390 ;
        RECT 125.430 87.850 125.570 98.070 ;
        RECT 125.890 88.190 126.030 104.870 ;
        RECT 126.350 101.450 126.490 105.210 ;
        RECT 129.570 101.450 129.710 106.910 ;
        RECT 130.430 104.530 130.690 104.850 ;
        RECT 130.490 102.470 130.630 104.530 ;
        RECT 130.430 102.150 130.690 102.470 ;
        RECT 130.950 101.790 131.090 106.910 ;
        RECT 130.890 101.470 131.150 101.790 ;
        RECT 126.290 101.130 126.550 101.450 ;
        RECT 129.510 101.130 129.770 101.450 ;
        RECT 129.050 97.050 129.310 97.370 ;
        RECT 128.130 96.030 128.390 96.350 ;
        RECT 128.190 95.670 128.330 96.030 ;
        RECT 128.130 95.350 128.390 95.670 ;
        RECT 128.190 93.970 128.330 95.350 ;
        RECT 129.110 94.650 129.250 97.050 ;
        RECT 129.570 95.670 129.710 101.130 ;
        RECT 131.410 99.070 131.550 107.250 ;
        RECT 133.190 99.090 133.450 99.410 ;
        RECT 131.350 98.750 131.610 99.070 ;
        RECT 129.970 98.070 130.230 98.390 ;
        RECT 130.030 97.030 130.170 98.070 ;
        RECT 129.970 96.710 130.230 97.030 ;
        RECT 130.030 96.350 130.170 96.710 ;
        RECT 130.430 96.370 130.690 96.690 ;
        RECT 129.970 96.030 130.230 96.350 ;
        RECT 129.510 95.350 129.770 95.670 ;
        RECT 129.050 94.330 129.310 94.650 ;
        RECT 128.130 93.650 128.390 93.970 ;
        RECT 129.510 93.880 129.770 93.970 ;
        RECT 130.030 93.880 130.170 96.030 ;
        RECT 130.490 94.650 130.630 96.370 ;
        RECT 133.250 94.650 133.390 99.090 ;
        RECT 130.430 94.330 130.690 94.650 ;
        RECT 133.190 94.330 133.450 94.650 ;
        RECT 133.710 93.970 133.850 124.250 ;
        RECT 134.170 123.550 134.310 128.670 ;
        RECT 135.030 127.990 135.290 128.310 ;
        RECT 135.090 127.290 135.230 127.990 ;
        RECT 135.030 126.970 135.290 127.290 ;
        RECT 135.030 126.290 135.290 126.610 ;
        RECT 135.950 126.290 136.210 126.610 ;
        RECT 134.110 123.230 134.370 123.550 ;
        RECT 134.170 121.850 134.310 123.230 ;
        RECT 134.570 122.550 134.830 122.870 ;
        RECT 134.110 121.530 134.370 121.850 ;
        RECT 134.170 120.490 134.310 121.530 ;
        RECT 134.630 121.510 134.770 122.550 ;
        RECT 135.090 121.850 135.230 126.290 ;
        RECT 136.010 124.230 136.150 126.290 ;
        RECT 135.950 123.910 136.210 124.230 ;
        RECT 135.030 121.530 135.290 121.850 ;
        RECT 134.570 121.190 134.830 121.510 ;
        RECT 136.470 121.170 136.610 129.270 ;
        RECT 136.930 126.950 137.070 136.150 ;
        RECT 137.850 133.750 137.990 142.950 ;
        RECT 138.770 142.500 138.910 176.950 ;
        RECT 140.610 174.460 140.750 177.630 ;
        RECT 141.530 176.250 141.670 177.630 ;
        RECT 141.470 175.930 141.730 176.250 ;
        RECT 141.990 175.230 142.130 186.470 ;
        RECT 142.450 184.070 142.590 193.270 ;
        RECT 142.910 192.570 143.050 193.610 ;
        RECT 142.850 192.250 143.110 192.570 ;
        RECT 143.370 192.230 143.510 202.790 ;
        RECT 143.770 199.390 144.030 199.710 ;
        RECT 143.830 193.930 143.970 199.390 ;
        RECT 143.770 193.610 144.030 193.930 ;
        RECT 143.310 191.910 143.570 192.230 ;
        RECT 143.830 191.970 143.970 193.610 ;
        RECT 144.750 192.765 144.890 212.200 ;
        RECT 152.110 208.890 152.250 212.200 ;
        RECT 156.240 209.055 157.780 209.425 ;
        RECT 152.050 208.570 152.310 208.890 ;
        RECT 152.510 206.870 152.770 207.190 ;
        RECT 152.570 206.170 152.710 206.870 ;
        RECT 152.510 205.850 152.770 206.170 ;
        RECT 146.070 204.150 146.330 204.470 ;
        RECT 146.130 202.965 146.270 204.150 ;
        RECT 156.240 203.615 157.780 203.985 ;
        RECT 146.060 202.595 146.340 202.965 ;
        RECT 146.130 201.750 146.270 202.595 ;
        RECT 149.750 202.450 150.010 202.770 ;
        RECT 148.360 201.915 148.640 202.285 ;
        RECT 146.070 201.430 146.330 201.750 ;
        RECT 146.530 199.390 146.790 199.710 ;
        RECT 146.590 198.010 146.730 199.390 ;
        RECT 148.430 198.010 148.570 201.915 ;
        RECT 146.530 197.690 146.790 198.010 ;
        RECT 148.370 197.690 148.630 198.010 ;
        RECT 145.150 197.410 145.410 197.670 ;
        RECT 145.150 197.350 145.810 197.410 ;
        RECT 146.070 197.350 146.330 197.670 ;
        RECT 145.210 197.270 145.810 197.350 ;
        RECT 145.670 196.310 145.810 197.270 ;
        RECT 145.150 195.990 145.410 196.310 ;
        RECT 145.610 195.990 145.870 196.310 ;
        RECT 145.210 195.290 145.350 195.990 ;
        RECT 145.150 194.970 145.410 195.290 ;
        RECT 146.130 194.950 146.270 197.350 ;
        RECT 147.910 197.010 148.170 197.330 ;
        RECT 146.070 194.630 146.330 194.950 ;
        RECT 146.070 193.950 146.330 194.270 ;
        RECT 144.680 192.395 144.960 192.765 ;
        RECT 143.830 191.890 144.430 191.970 ;
        RECT 142.850 191.570 143.110 191.890 ;
        RECT 143.830 191.830 144.490 191.890 ;
        RECT 144.230 191.570 144.490 191.830 ;
        RECT 142.910 185.430 143.050 191.570 ;
        RECT 146.130 190.870 146.270 193.950 ;
        RECT 146.530 193.610 146.790 193.930 ;
        RECT 145.610 190.550 145.870 190.870 ;
        RECT 146.070 190.550 146.330 190.870 ;
        RECT 143.310 188.510 143.570 188.830 ;
        RECT 142.850 185.110 143.110 185.430 ;
        RECT 142.390 183.750 142.650 184.070 ;
        RECT 142.910 183.390 143.050 185.110 ;
        RECT 142.850 183.070 143.110 183.390 ;
        RECT 142.390 182.390 142.650 182.710 ;
        RECT 142.450 181.690 142.590 182.390 ;
        RECT 142.910 181.690 143.050 183.070 ;
        RECT 142.390 181.370 142.650 181.690 ;
        RECT 142.850 181.370 143.110 181.690 ;
        RECT 143.370 180.330 143.510 188.510 ;
        RECT 144.690 186.470 144.950 186.790 ;
        RECT 144.230 185.790 144.490 186.110 ;
        RECT 143.770 183.750 144.030 184.070 ;
        RECT 143.310 180.010 143.570 180.330 ;
        RECT 141.930 174.910 142.190 175.230 ;
        RECT 140.610 174.320 141.670 174.460 ;
        RECT 139.450 173.695 140.990 174.065 ;
        RECT 139.450 168.255 140.990 168.625 ;
        RECT 139.450 162.815 140.990 163.185 ;
        RECT 140.090 161.650 140.350 161.970 ;
        RECT 139.170 161.310 139.430 161.630 ;
        RECT 139.230 159.930 139.370 161.310 ;
        RECT 140.150 159.930 140.290 161.650 ;
        RECT 139.170 159.610 139.430 159.930 ;
        RECT 140.090 159.610 140.350 159.930 ;
        RECT 139.450 157.375 140.990 157.745 ;
        RECT 139.450 151.935 140.990 152.305 ;
        RECT 140.090 150.430 140.350 150.750 ;
        RECT 140.150 149.050 140.290 150.430 ;
        RECT 140.090 148.730 140.350 149.050 ;
        RECT 141.530 148.370 141.670 174.320 ;
        RECT 142.850 174.230 143.110 174.550 ;
        RECT 142.390 172.190 142.650 172.510 ;
        RECT 141.930 171.850 142.190 172.170 ;
        RECT 141.990 170.810 142.130 171.850 ;
        RECT 142.450 170.810 142.590 172.190 ;
        RECT 141.930 170.490 142.190 170.810 ;
        RECT 142.390 170.490 142.650 170.810 ;
        RECT 142.910 170.470 143.050 174.230 ;
        RECT 143.370 172.930 143.510 180.010 ;
        RECT 143.830 178.970 143.970 183.750 ;
        RECT 143.770 178.650 144.030 178.970 ;
        RECT 143.770 177.290 144.030 177.610 ;
        RECT 143.830 175.910 143.970 177.290 ;
        RECT 144.290 176.250 144.430 185.790 ;
        RECT 144.750 184.410 144.890 186.470 ;
        RECT 145.670 186.450 145.810 190.550 ;
        RECT 146.130 186.450 146.270 190.550 ;
        RECT 146.590 188.490 146.730 193.610 ;
        RECT 147.970 193.590 148.110 197.010 ;
        RECT 147.450 193.270 147.710 193.590 ;
        RECT 147.910 193.270 148.170 193.590 ;
        RECT 147.510 192.570 147.650 193.270 ;
        RECT 147.450 192.250 147.710 192.570 ;
        RECT 147.970 192.230 148.110 193.270 ;
        RECT 147.910 191.910 148.170 192.230 ;
        RECT 148.430 191.890 148.570 197.690 ;
        RECT 149.290 197.010 149.550 197.330 ;
        RECT 148.830 195.990 149.090 196.310 ;
        RECT 148.890 191.890 149.030 195.990 ;
        RECT 149.350 195.290 149.490 197.010 ;
        RECT 149.290 194.970 149.550 195.290 ;
        RECT 148.370 191.570 148.630 191.890 ;
        RECT 148.830 191.570 149.090 191.890 ;
        RECT 146.530 188.170 146.790 188.490 ;
        RECT 145.610 186.130 145.870 186.450 ;
        RECT 146.070 186.130 146.330 186.450 ;
        RECT 144.690 184.090 144.950 184.410 ;
        RECT 146.130 183.390 146.270 186.130 ;
        RECT 146.070 183.070 146.330 183.390 ;
        RECT 144.230 175.930 144.490 176.250 ;
        RECT 143.770 175.590 144.030 175.910 ;
        RECT 143.830 173.530 143.970 175.590 ;
        RECT 145.150 174.910 145.410 175.230 ;
        RECT 143.770 173.210 144.030 173.530 ;
        RECT 143.370 172.790 143.970 172.930 ;
        RECT 142.850 170.150 143.110 170.470 ;
        RECT 141.930 169.810 142.190 170.130 ;
        RECT 141.990 167.750 142.130 169.810 ;
        RECT 142.390 169.470 142.650 169.790 ;
        RECT 143.310 169.470 143.570 169.790 ;
        RECT 141.930 167.430 142.190 167.750 ;
        RECT 141.990 164.690 142.130 167.430 ;
        RECT 142.450 166.390 142.590 169.470 ;
        RECT 142.850 166.750 143.110 167.070 ;
        RECT 142.390 166.070 142.650 166.390 ;
        RECT 142.390 165.050 142.650 165.370 ;
        RECT 141.930 164.370 142.190 164.690 ;
        RECT 141.930 163.690 142.190 164.010 ;
        RECT 141.990 161.630 142.130 163.690 ;
        RECT 141.930 161.310 142.190 161.630 ;
        RECT 142.450 150.750 142.590 165.050 ;
        RECT 142.910 158.570 143.050 166.750 ;
        RECT 143.370 166.730 143.510 169.470 ;
        RECT 143.310 166.410 143.570 166.730 ;
        RECT 143.370 162.650 143.510 166.410 ;
        RECT 143.310 162.330 143.570 162.650 ;
        RECT 142.850 158.250 143.110 158.570 ;
        RECT 143.830 150.870 143.970 172.790 ;
        RECT 144.690 172.190 144.950 172.510 ;
        RECT 144.750 170.470 144.890 172.190 ;
        RECT 144.690 170.150 144.950 170.470 ;
        RECT 144.750 168.090 144.890 170.150 ;
        RECT 145.210 169.110 145.350 174.910 ;
        RECT 145.610 169.810 145.870 170.130 ;
        RECT 145.150 168.790 145.410 169.110 ;
        RECT 144.690 167.770 144.950 168.090 ;
        RECT 144.230 167.430 144.490 167.750 ;
        RECT 144.290 167.070 144.430 167.430 ;
        RECT 144.230 166.750 144.490 167.070 ;
        RECT 145.670 162.650 145.810 169.810 ;
        RECT 145.610 162.330 145.870 162.650 ;
        RECT 145.670 159.590 145.810 162.330 ;
        RECT 146.590 161.630 146.730 188.170 ;
        RECT 149.810 186.790 149.950 202.450 ;
        RECT 152.050 199.050 152.310 199.370 ;
        RECT 151.130 198.710 151.390 199.030 ;
        RECT 150.210 195.990 150.470 196.310 ;
        RECT 150.270 195.290 150.410 195.990 ;
        RECT 150.210 194.970 150.470 195.290 ;
        RECT 151.190 194.270 151.330 198.710 ;
        RECT 152.110 197.330 152.250 199.050 ;
        RECT 156.240 198.175 157.780 198.545 ;
        RECT 152.050 197.010 152.310 197.330 ;
        RECT 151.130 193.950 151.390 194.270 ;
        RECT 151.190 188.150 151.330 193.950 ;
        RECT 156.240 192.735 157.780 193.105 ;
        RECT 151.130 187.830 151.390 188.150 ;
        RECT 149.750 186.470 150.010 186.790 ;
        RECT 146.990 185.110 147.250 185.430 ;
        RECT 147.450 185.110 147.710 185.430 ;
        RECT 147.050 184.410 147.190 185.110 ;
        RECT 146.990 184.090 147.250 184.410 ;
        RECT 146.990 183.130 147.250 183.390 ;
        RECT 147.510 183.130 147.650 185.110 ;
        RECT 149.810 184.410 149.950 186.470 ;
        RECT 150.670 185.790 150.930 186.110 ;
        RECT 150.210 185.110 150.470 185.430 ;
        RECT 149.750 184.090 150.010 184.410 ;
        RECT 146.990 183.070 147.650 183.130 ;
        RECT 147.050 182.990 147.650 183.070 ;
        RECT 147.050 178.630 147.190 182.990 ;
        RECT 147.450 182.390 147.710 182.710 ;
        RECT 147.910 182.390 148.170 182.710 ;
        RECT 147.510 179.990 147.650 182.390 ;
        RECT 147.970 181.690 148.110 182.390 ;
        RECT 147.910 181.370 148.170 181.690 ;
        RECT 149.810 180.580 149.950 184.090 ;
        RECT 150.270 181.350 150.410 185.110 ;
        RECT 150.730 181.350 150.870 185.790 ;
        RECT 151.190 183.390 151.330 187.830 ;
        RECT 156.240 187.295 157.780 187.665 ;
        RECT 151.130 183.070 151.390 183.390 ;
        RECT 150.210 181.030 150.470 181.350 ;
        RECT 150.670 181.030 150.930 181.350 ;
        RECT 151.190 181.010 151.330 183.070 ;
        RECT 153.890 182.730 154.150 183.050 ;
        RECT 153.950 181.690 154.090 182.730 ;
        RECT 156.240 181.855 157.780 182.225 ;
        RECT 153.890 181.370 154.150 181.690 ;
        RECT 151.130 180.690 151.390 181.010 ;
        RECT 151.590 180.690 151.850 181.010 ;
        RECT 149.810 180.440 150.410 180.580 ;
        RECT 147.450 179.670 147.710 179.990 ;
        RECT 149.290 178.650 149.550 178.970 ;
        RECT 146.990 178.310 147.250 178.630 ;
        RECT 147.450 177.630 147.710 177.950 ;
        RECT 146.990 177.290 147.250 177.610 ;
        RECT 147.050 176.250 147.190 177.290 ;
        RECT 146.990 175.930 147.250 176.250 ;
        RECT 147.510 172.510 147.650 177.630 ;
        RECT 147.450 172.190 147.710 172.510 ;
        RECT 148.830 172.420 149.090 172.510 ;
        RECT 149.350 172.420 149.490 178.650 ;
        RECT 149.810 174.550 149.950 180.440 ;
        RECT 150.270 180.410 150.410 180.440 ;
        RECT 151.650 180.410 151.790 180.690 ;
        RECT 150.270 180.270 151.790 180.410 ;
        RECT 152.050 176.950 152.310 177.270 ;
        RECT 154.810 176.950 155.070 177.270 ;
        RECT 152.110 176.250 152.250 176.950 ;
        RECT 154.870 176.250 155.010 176.950 ;
        RECT 156.240 176.415 157.780 176.785 ;
        RECT 152.050 175.930 152.310 176.250 ;
        RECT 154.810 175.930 155.070 176.250 ;
        RECT 151.130 175.250 151.390 175.570 ;
        RECT 149.750 174.230 150.010 174.550 ;
        RECT 150.210 174.230 150.470 174.550 ;
        RECT 148.830 172.280 149.490 172.420 ;
        RECT 148.830 172.190 149.090 172.280 ;
        RECT 146.990 168.790 147.250 169.110 ;
        RECT 147.050 167.070 147.190 168.790 ;
        RECT 147.510 167.410 147.650 172.190 ;
        RECT 147.910 171.850 148.170 172.170 ;
        RECT 147.970 168.090 148.110 171.850 ;
        RECT 149.350 170.470 149.490 172.280 ;
        RECT 150.270 170.810 150.410 174.230 ;
        RECT 151.190 171.830 151.330 175.250 ;
        RECT 152.050 174.230 152.310 174.550 ;
        RECT 151.130 171.510 151.390 171.830 ;
        RECT 151.190 170.810 151.330 171.510 ;
        RECT 150.210 170.490 150.470 170.810 ;
        RECT 151.130 170.490 151.390 170.810 ;
        RECT 149.290 170.150 149.550 170.470 ;
        RECT 148.370 169.470 148.630 169.790 ;
        RECT 148.430 168.090 148.570 169.470 ;
        RECT 147.910 167.770 148.170 168.090 ;
        RECT 148.370 167.770 148.630 168.090 ;
        RECT 147.450 167.090 147.710 167.410 ;
        RECT 146.990 166.750 147.250 167.070 ;
        RECT 147.450 164.030 147.710 164.350 ;
        RECT 147.510 162.650 147.650 164.030 ;
        RECT 148.430 162.650 148.570 167.770 ;
        RECT 149.350 165.030 149.490 170.150 ;
        RECT 149.290 164.710 149.550 165.030 ;
        RECT 150.270 164.670 150.410 170.490 ;
        RECT 152.110 170.130 152.250 174.230 ;
        RECT 156.240 170.975 157.780 171.345 ;
        RECT 152.050 169.810 152.310 170.130 ;
        RECT 150.670 168.790 150.930 169.110 ;
        RECT 154.810 168.790 155.070 169.110 ;
        RECT 150.730 166.730 150.870 168.790 ;
        RECT 152.510 166.750 152.770 167.070 ;
        RECT 154.870 166.810 155.010 168.790 ;
        RECT 150.670 166.410 150.930 166.730 ;
        RECT 150.270 164.530 150.870 164.670 ;
        RECT 149.290 163.350 149.550 163.670 ;
        RECT 147.450 162.330 147.710 162.650 ;
        RECT 148.370 162.330 148.630 162.650 ;
        RECT 146.530 161.310 146.790 161.630 ;
        RECT 145.610 159.270 145.870 159.590 ;
        RECT 146.590 154.150 146.730 161.310 ;
        RECT 147.510 159.930 147.650 162.330 ;
        RECT 149.350 159.930 149.490 163.350 ;
        RECT 147.450 159.610 147.710 159.930 ;
        RECT 149.290 159.610 149.550 159.930 ;
        RECT 150.730 159.590 150.870 164.530 ;
        RECT 152.050 163.350 152.310 163.670 ;
        RECT 152.110 159.930 152.250 163.350 ;
        RECT 152.570 162.650 152.710 166.750 ;
        RECT 153.890 166.410 154.150 166.730 ;
        RECT 154.410 166.670 155.010 166.810 ;
        RECT 153.950 165.370 154.090 166.410 ;
        RECT 153.890 165.050 154.150 165.370 ;
        RECT 152.510 162.330 152.770 162.650 ;
        RECT 152.050 159.610 152.310 159.930 ;
        RECT 150.670 159.270 150.930 159.590 ;
        RECT 152.570 159.250 152.710 162.330 ;
        RECT 152.510 158.930 152.770 159.250 ;
        RECT 153.430 159.160 153.690 159.250 ;
        RECT 154.410 159.160 154.550 166.670 ;
        RECT 156.240 165.535 157.780 165.905 ;
        RECT 154.810 164.710 155.070 165.030 ;
        RECT 154.870 159.930 155.010 164.710 ;
        RECT 156.240 160.095 157.780 160.465 ;
        RECT 154.810 159.610 155.070 159.930 ;
        RECT 154.810 159.160 155.070 159.250 ;
        RECT 153.430 159.020 155.070 159.160 ;
        RECT 153.430 158.930 153.690 159.020 ;
        RECT 154.810 158.930 155.070 159.020 ;
        RECT 152.570 156.190 152.710 158.930 ;
        RECT 151.130 155.870 151.390 156.190 ;
        RECT 152.510 155.870 152.770 156.190 ;
        RECT 147.910 155.530 148.170 155.850 ;
        RECT 146.530 153.830 146.790 154.150 ;
        RECT 147.450 152.470 147.710 152.790 ;
        RECT 142.390 150.430 142.650 150.750 ;
        RECT 143.370 150.730 143.970 150.870 ;
        RECT 143.370 150.490 143.510 150.730 ;
        RECT 142.910 150.350 143.510 150.490 ;
        RECT 146.070 150.430 146.330 150.750 ;
        RECT 141.470 148.050 141.730 148.370 ;
        RECT 139.450 146.495 140.990 146.865 ;
        RECT 140.550 146.010 140.810 146.330 ;
        RECT 140.610 145.310 140.750 146.010 ;
        RECT 141.530 145.990 141.670 148.050 ;
        RECT 142.390 147.710 142.650 148.030 ;
        RECT 142.450 145.990 142.590 147.710 ;
        RECT 141.470 145.670 141.730 145.990 ;
        RECT 142.390 145.670 142.650 145.990 ;
        RECT 140.550 144.990 140.810 145.310 ;
        RECT 141.470 142.950 141.730 143.270 ;
        RECT 138.310 142.360 138.910 142.500 ;
        RECT 137.790 133.430 138.050 133.750 ;
        RECT 137.330 131.730 137.590 132.050 ;
        RECT 137.390 128.990 137.530 131.730 ;
        RECT 137.790 130.710 138.050 131.030 ;
        RECT 137.330 128.670 137.590 128.990 ;
        RECT 136.870 126.630 137.130 126.950 ;
        RECT 137.330 122.550 137.590 122.870 ;
        RECT 137.390 121.170 137.530 122.550 ;
        RECT 136.410 120.850 136.670 121.170 ;
        RECT 137.330 120.850 137.590 121.170 ;
        RECT 135.490 120.510 135.750 120.830 ;
        RECT 134.110 120.170 134.370 120.490 ;
        RECT 135.550 119.130 135.690 120.510 ;
        RECT 137.850 120.150 137.990 130.710 ;
        RECT 138.310 129.330 138.450 142.360 ;
        RECT 138.710 141.590 138.970 141.910 ;
        RECT 138.770 137.830 138.910 141.590 ;
        RECT 139.450 141.055 140.990 141.425 ;
        RECT 139.630 140.405 139.890 140.550 ;
        RECT 139.620 140.035 139.900 140.405 ;
        RECT 140.550 138.870 140.810 139.190 ;
        RECT 141.010 139.045 141.270 139.190 ;
        RECT 138.710 137.510 138.970 137.830 ;
        RECT 140.610 137.490 140.750 138.870 ;
        RECT 141.000 138.675 141.280 139.045 ;
        RECT 141.530 138.170 141.670 142.950 ;
        RECT 142.390 142.270 142.650 142.590 ;
        RECT 141.930 141.590 142.190 141.910 ;
        RECT 141.990 140.890 142.130 141.590 ;
        RECT 141.930 140.570 142.190 140.890 ;
        RECT 142.450 139.610 142.590 142.270 ;
        RECT 141.990 139.470 142.590 139.610 ;
        RECT 141.990 139.190 142.130 139.470 ;
        RECT 141.930 138.870 142.190 139.190 ;
        RECT 141.470 137.850 141.730 138.170 ;
        RECT 140.550 137.170 140.810 137.490 ;
        RECT 142.910 137.150 143.050 150.350 ;
        RECT 143.310 149.750 143.570 150.070 ;
        RECT 144.230 149.750 144.490 150.070 ;
        RECT 143.370 149.050 143.510 149.750 ;
        RECT 143.310 148.730 143.570 149.050 ;
        RECT 144.290 148.710 144.430 149.750 ;
        RECT 144.230 148.390 144.490 148.710 ;
        RECT 144.230 147.370 144.490 147.690 ;
        RECT 143.770 147.030 144.030 147.350 ;
        RECT 143.310 142.610 143.570 142.930 ;
        RECT 143.370 139.045 143.510 142.610 ;
        RECT 143.300 138.675 143.580 139.045 ;
        RECT 143.830 138.170 143.970 147.030 ;
        RECT 144.290 143.270 144.430 147.370 ;
        RECT 145.150 144.310 145.410 144.630 ;
        RECT 145.210 143.270 145.350 144.310 ;
        RECT 146.130 143.270 146.270 150.430 ;
        RECT 146.990 147.030 147.250 147.350 ;
        RECT 147.050 146.330 147.190 147.030 ;
        RECT 146.990 146.010 147.250 146.330 ;
        RECT 144.230 142.950 144.490 143.270 ;
        RECT 145.150 142.950 145.410 143.270 ;
        RECT 146.070 142.950 146.330 143.270 ;
        RECT 144.230 141.930 144.490 142.250 ;
        RECT 144.290 140.210 144.430 141.930 ;
        RECT 145.610 141.590 145.870 141.910 ;
        RECT 144.680 140.290 144.960 140.405 ;
        RECT 144.230 139.890 144.490 140.210 ;
        RECT 144.680 140.150 145.350 140.290 ;
        RECT 144.680 140.035 144.960 140.150 ;
        RECT 145.210 139.870 145.350 140.150 ;
        RECT 145.150 139.550 145.410 139.870 ;
        RECT 144.690 139.210 144.950 139.530 ;
        RECT 144.750 138.170 144.890 139.210 ;
        RECT 145.150 138.870 145.410 139.190 ;
        RECT 143.770 137.850 144.030 138.170 ;
        RECT 144.690 137.850 144.950 138.170 ;
        RECT 141.470 136.830 141.730 137.150 ;
        RECT 142.850 136.830 143.110 137.150 ;
        RECT 139.450 135.615 140.990 135.985 ;
        RECT 138.710 134.110 138.970 134.430 ;
        RECT 140.550 134.110 140.810 134.430 ;
        RECT 138.770 132.050 138.910 134.110 ;
        RECT 140.610 132.390 140.750 134.110 ;
        RECT 141.530 132.390 141.670 136.830 ;
        RECT 142.910 132.810 143.050 136.830 ;
        RECT 143.830 134.430 143.970 137.850 ;
        RECT 144.750 137.490 144.890 137.850 ;
        RECT 145.210 137.490 145.350 138.870 ;
        RECT 145.670 138.170 145.810 141.590 ;
        RECT 147.510 140.210 147.650 152.470 ;
        RECT 147.970 151.770 148.110 155.530 ;
        RECT 147.910 151.450 148.170 151.770 ;
        RECT 151.190 150.750 151.330 155.870 ;
        RECT 155.270 155.190 155.530 155.510 ;
        RECT 155.330 153.810 155.470 155.190 ;
        RECT 156.240 154.655 157.780 155.025 ;
        RECT 155.270 153.490 155.530 153.810 ;
        RECT 152.050 152.470 152.310 152.790 ;
        RECT 148.830 150.430 149.090 150.750 ;
        RECT 151.130 150.430 151.390 150.750 ;
        RECT 148.890 145.310 149.030 150.430 ;
        RECT 149.290 150.090 149.550 150.410 ;
        RECT 149.350 149.050 149.490 150.090 ;
        RECT 152.110 150.070 152.250 152.470 ;
        RECT 152.050 149.750 152.310 150.070 ;
        RECT 149.290 148.730 149.550 149.050 ;
        RECT 155.330 148.030 155.470 153.490 ;
        RECT 156.240 149.215 157.780 149.585 ;
        RECT 155.270 147.710 155.530 148.030 ;
        RECT 148.830 144.990 149.090 145.310 ;
        RECT 149.750 144.650 150.010 144.970 ;
        RECT 149.810 143.610 149.950 144.650 ;
        RECT 156.240 143.775 157.780 144.145 ;
        RECT 149.750 143.290 150.010 143.610 ;
        RECT 147.450 139.890 147.710 140.210 ;
        RECT 146.530 139.550 146.790 139.870 ;
        RECT 146.070 138.870 146.330 139.190 ;
        RECT 145.610 137.850 145.870 138.170 ;
        RECT 144.690 137.170 144.950 137.490 ;
        RECT 145.150 137.170 145.410 137.490 ;
        RECT 146.130 136.470 146.270 138.870 ;
        RECT 146.070 136.150 146.330 136.470 ;
        RECT 146.590 135.450 146.730 139.550 ;
        RECT 148.830 139.210 149.090 139.530 ;
        RECT 148.890 138.170 149.030 139.210 ;
        RECT 156.240 138.335 157.780 138.705 ;
        RECT 148.830 137.850 149.090 138.170 ;
        RECT 151.130 137.510 151.390 137.830 ;
        RECT 146.530 135.130 146.790 135.450 ;
        RECT 151.190 134.430 151.330 137.510 ;
        RECT 143.770 134.110 144.030 134.430 ;
        RECT 151.130 134.110 151.390 134.430 ;
        RECT 154.350 134.110 154.610 134.430 ;
        RECT 143.310 133.430 143.570 133.750 ;
        RECT 142.450 132.670 143.050 132.810 ;
        RECT 140.550 132.070 140.810 132.390 ;
        RECT 141.470 132.070 141.730 132.390 ;
        RECT 138.710 131.730 138.970 132.050 ;
        RECT 139.450 130.175 140.990 130.545 ;
        RECT 138.250 129.010 138.510 129.330 ;
        RECT 141.530 128.900 141.670 132.070 ;
        RECT 142.450 132.050 142.590 132.670 ;
        RECT 142.850 132.070 143.110 132.390 ;
        RECT 142.390 131.730 142.650 132.050 ;
        RECT 142.910 128.990 143.050 132.070 ;
        RECT 141.930 128.900 142.190 128.990 ;
        RECT 141.530 128.760 142.190 128.900 ;
        RECT 140.550 127.990 140.810 128.310 ;
        RECT 140.610 127.290 140.750 127.990 ;
        RECT 141.530 127.290 141.670 128.760 ;
        RECT 141.930 128.670 142.190 128.760 ;
        RECT 142.850 128.670 143.110 128.990 ;
        RECT 141.930 127.990 142.190 128.310 ;
        RECT 140.550 126.970 140.810 127.290 ;
        RECT 141.470 126.970 141.730 127.290 ;
        RECT 141.990 126.950 142.130 127.990 ;
        RECT 142.910 127.290 143.050 128.670 ;
        RECT 143.370 128.650 143.510 133.430 ;
        RECT 146.990 131.730 147.250 132.050 ;
        RECT 143.770 130.710 144.030 131.030 ;
        RECT 143.830 130.010 143.970 130.710 ;
        RECT 147.050 130.010 147.190 131.730 ;
        RECT 151.130 130.710 151.390 131.030 ;
        RECT 143.770 129.690 144.030 130.010 ;
        RECT 146.990 129.690 147.250 130.010 ;
        RECT 151.190 128.990 151.330 130.710 ;
        RECT 154.410 128.990 154.550 134.110 ;
        RECT 156.240 132.895 157.780 133.265 ;
        RECT 151.130 128.670 151.390 128.990 ;
        RECT 154.350 128.670 154.610 128.990 ;
        RECT 143.310 128.330 143.570 128.650 ;
        RECT 143.370 127.290 143.510 128.330 ;
        RECT 146.070 127.990 146.330 128.310 ;
        RECT 146.130 127.290 146.270 127.990 ;
        RECT 142.850 126.970 143.110 127.290 ;
        RECT 143.310 126.970 143.570 127.290 ;
        RECT 146.070 126.970 146.330 127.290 ;
        RECT 141.930 126.630 142.190 126.950 ;
        RECT 145.150 126.290 145.410 126.610 ;
        RECT 143.770 125.610 144.030 125.930 ;
        RECT 144.230 125.610 144.490 125.930 ;
        RECT 138.710 125.270 138.970 125.590 ;
        RECT 138.770 123.890 138.910 125.270 ;
        RECT 139.450 124.735 140.990 125.105 ;
        RECT 141.010 124.250 141.270 124.570 ;
        RECT 139.170 123.910 139.430 124.230 ;
        RECT 138.710 123.570 138.970 123.890 ;
        RECT 138.250 122.890 138.510 123.210 ;
        RECT 138.310 121.170 138.450 122.890 ;
        RECT 138.770 121.170 138.910 123.570 ;
        RECT 139.230 121.170 139.370 123.910 ;
        RECT 141.070 123.550 141.210 124.250 ;
        RECT 143.830 123.890 143.970 125.610 ;
        RECT 143.770 123.800 144.030 123.890 ;
        RECT 142.910 123.660 144.030 123.800 ;
        RECT 141.010 123.230 141.270 123.550 ;
        RECT 141.930 122.890 142.190 123.210 ;
        RECT 138.250 120.850 138.510 121.170 ;
        RECT 138.710 120.850 138.970 121.170 ;
        RECT 139.170 120.850 139.430 121.170 ;
        RECT 137.790 119.830 138.050 120.150 ;
        RECT 135.490 118.810 135.750 119.130 ;
        RECT 138.310 118.110 138.450 120.850 ;
        RECT 141.990 120.490 142.130 122.890 ;
        RECT 141.930 120.170 142.190 120.490 ;
        RECT 141.470 119.830 141.730 120.150 ;
        RECT 139.450 119.295 140.990 119.665 ;
        RECT 139.170 118.810 139.430 119.130 ;
        RECT 135.490 117.790 135.750 118.110 ;
        RECT 138.250 117.790 138.510 118.110 ;
        RECT 135.550 116.410 135.690 117.790 ;
        RECT 136.870 117.450 137.130 117.770 ;
        RECT 137.790 117.450 138.050 117.770 ;
        RECT 134.570 116.090 134.830 116.410 ;
        RECT 135.490 116.090 135.750 116.410 ;
        RECT 136.930 116.370 137.070 117.450 ;
        RECT 137.850 116.370 137.990 117.450 ;
        RECT 136.470 116.230 137.070 116.370 ;
        RECT 137.390 116.230 137.990 116.370 ;
        RECT 134.110 115.070 134.370 115.390 ;
        RECT 134.170 113.690 134.310 115.070 ;
        RECT 134.630 113.690 134.770 116.090 ;
        RECT 134.110 113.370 134.370 113.690 ;
        RECT 134.570 113.370 134.830 113.690 ;
        RECT 134.170 110.970 134.310 113.370 ;
        RECT 135.030 112.010 135.290 112.330 ;
        RECT 134.110 110.650 134.370 110.970 ;
        RECT 135.090 110.290 135.230 112.010 ;
        RECT 136.470 111.990 136.610 116.230 ;
        RECT 136.870 114.390 137.130 114.710 ;
        RECT 136.930 113.010 137.070 114.390 ;
        RECT 137.390 113.690 137.530 116.230 ;
        RECT 138.250 115.750 138.510 116.070 ;
        RECT 137.790 115.070 138.050 115.390 ;
        RECT 137.330 113.370 137.590 113.690 ;
        RECT 136.870 112.690 137.130 113.010 ;
        RECT 136.870 112.010 137.130 112.330 ;
        RECT 136.410 111.670 136.670 111.990 ;
        RECT 135.030 109.970 135.290 110.290 ;
        RECT 136.930 109.610 137.070 112.010 ;
        RECT 137.390 110.630 137.530 113.370 ;
        RECT 137.850 113.350 137.990 115.070 ;
        RECT 137.790 113.030 138.050 113.350 ;
        RECT 137.790 112.350 138.050 112.670 ;
        RECT 137.850 110.970 137.990 112.350 ;
        RECT 137.790 110.650 138.050 110.970 ;
        RECT 137.330 110.310 137.590 110.630 ;
        RECT 138.310 109.950 138.450 115.750 ;
        RECT 139.230 115.730 139.370 118.810 ;
        RECT 141.530 118.790 141.670 119.830 ;
        RECT 141.470 118.470 141.730 118.790 ;
        RECT 139.170 115.410 139.430 115.730 ;
        RECT 138.710 114.390 138.970 114.710 ;
        RECT 138.770 110.630 138.910 114.390 ;
        RECT 139.450 113.855 140.990 114.225 ;
        RECT 141.530 112.410 141.670 118.470 ;
        RECT 142.910 113.690 143.050 123.660 ;
        RECT 143.770 123.570 144.030 123.660 ;
        RECT 144.290 122.870 144.430 125.610 ;
        RECT 145.210 124.570 145.350 126.290 ;
        RECT 145.610 125.610 145.870 125.930 ;
        RECT 144.690 124.250 144.950 124.570 ;
        RECT 145.150 124.250 145.410 124.570 ;
        RECT 144.230 122.550 144.490 122.870 ;
        RECT 144.290 121.850 144.430 122.550 ;
        RECT 144.750 121.850 144.890 124.250 ;
        RECT 144.230 121.530 144.490 121.850 ;
        RECT 144.690 121.530 144.950 121.850 ;
        RECT 145.670 120.830 145.810 125.610 ;
        RECT 145.150 120.510 145.410 120.830 ;
        RECT 145.610 120.510 145.870 120.830 ;
        RECT 143.310 118.810 143.570 119.130 ;
        RECT 143.370 117.430 143.510 118.810 ;
        RECT 144.690 117.450 144.950 117.770 ;
        RECT 143.310 117.110 143.570 117.430 ;
        RECT 143.770 117.110 144.030 117.430 ;
        RECT 143.830 116.370 143.970 117.110 ;
        RECT 143.370 116.230 143.970 116.370 ;
        RECT 142.850 113.370 143.110 113.690 ;
        RECT 141.530 112.270 142.590 112.410 ;
        RECT 142.450 111.990 142.590 112.270 ;
        RECT 143.370 111.990 143.510 116.230 ;
        RECT 143.770 115.070 144.030 115.390 ;
        RECT 143.830 113.690 143.970 115.070 ;
        RECT 144.230 114.390 144.490 114.710 ;
        RECT 143.770 113.370 144.030 113.690 ;
        RECT 144.290 113.090 144.430 114.390 ;
        RECT 144.750 113.690 144.890 117.450 ;
        RECT 145.210 117.430 145.350 120.510 ;
        RECT 145.150 117.110 145.410 117.430 ;
        RECT 144.690 113.370 144.950 113.690 ;
        RECT 144.290 113.010 144.890 113.090 ;
        RECT 144.290 112.950 144.950 113.010 ;
        RECT 144.690 112.690 144.950 112.950 ;
        RECT 142.390 111.670 142.650 111.990 ;
        RECT 143.310 111.670 143.570 111.990 ;
        RECT 143.770 111.670 144.030 111.990 ;
        RECT 138.710 110.310 138.970 110.630 ;
        RECT 138.250 109.630 138.510 109.950 ;
        RECT 136.870 109.290 137.130 109.610 ;
        RECT 138.310 104.850 138.450 109.630 ;
        RECT 139.450 108.415 140.990 108.785 ;
        RECT 142.450 107.570 142.590 111.670 ;
        RECT 142.390 107.250 142.650 107.570 ;
        RECT 143.370 107.230 143.510 111.670 ;
        RECT 143.310 106.910 143.570 107.230 ;
        RECT 138.250 104.530 138.510 104.850 ;
        RECT 143.310 104.530 143.570 104.850 ;
        RECT 139.450 102.975 140.990 103.345 ;
        RECT 137.330 102.150 137.590 102.470 ;
        RECT 135.030 101.470 135.290 101.790 ;
        RECT 135.090 99.490 135.230 101.470 ;
        RECT 135.490 100.790 135.750 101.110 ;
        RECT 135.550 100.090 135.690 100.790 ;
        RECT 137.390 100.090 137.530 102.150 ;
        RECT 141.470 101.810 141.730 102.130 ;
        RECT 135.490 99.770 135.750 100.090 ;
        RECT 137.330 99.770 137.590 100.090 ;
        RECT 137.390 99.490 137.530 99.770 ;
        RECT 135.090 99.410 135.690 99.490 ;
        RECT 135.090 99.350 135.750 99.410 ;
        RECT 135.490 99.090 135.750 99.350 ;
        RECT 136.930 99.350 137.530 99.490 ;
        RECT 134.110 98.410 134.370 98.730 ;
        RECT 134.170 96.690 134.310 98.410 ;
        RECT 134.570 98.070 134.830 98.390 ;
        RECT 135.030 98.070 135.290 98.390 ;
        RECT 134.630 97.370 134.770 98.070 ;
        RECT 134.570 97.050 134.830 97.370 ;
        RECT 134.110 96.370 134.370 96.690 ;
        RECT 134.170 93.970 134.310 96.370 ;
        RECT 135.090 96.090 135.230 98.070 ;
        RECT 135.550 96.350 135.690 99.090 ;
        RECT 136.930 96.690 137.070 99.350 ;
        RECT 137.790 99.090 138.050 99.410 ;
        RECT 137.330 98.410 137.590 98.730 ;
        RECT 136.870 96.370 137.130 96.690 ;
        RECT 137.390 96.350 137.530 98.410 ;
        RECT 137.850 96.350 137.990 99.090 ;
        RECT 139.450 97.535 140.990 97.905 ;
        RECT 141.010 97.280 141.270 97.370 ;
        RECT 141.530 97.280 141.670 101.810 ;
        RECT 141.930 100.790 142.190 101.110 ;
        RECT 141.990 100.090 142.130 100.790 ;
        RECT 143.370 100.090 143.510 104.530 ;
        RECT 141.930 99.770 142.190 100.090 ;
        RECT 143.310 99.770 143.570 100.090 ;
        RECT 141.930 98.750 142.190 99.070 ;
        RECT 141.990 97.370 142.130 98.750 ;
        RECT 141.010 97.140 141.670 97.280 ;
        RECT 141.010 97.050 141.270 97.140 ;
        RECT 141.930 97.050 142.190 97.370 ;
        RECT 134.630 96.010 135.230 96.090 ;
        RECT 135.490 96.030 135.750 96.350 ;
        RECT 137.330 96.030 137.590 96.350 ;
        RECT 137.790 96.030 138.050 96.350 ;
        RECT 138.710 96.030 138.970 96.350 ;
        RECT 141.010 96.030 141.270 96.350 ;
        RECT 134.570 95.950 135.230 96.010 ;
        RECT 134.570 95.690 134.830 95.950 ;
        RECT 129.510 93.740 130.170 93.880 ;
        RECT 129.510 93.650 129.770 93.740 ;
        RECT 132.270 93.650 132.530 93.970 ;
        RECT 133.650 93.650 133.910 93.970 ;
        RECT 134.110 93.650 134.370 93.970 ;
        RECT 128.130 90.590 128.390 90.910 ;
        RECT 128.190 88.530 128.330 90.590 ;
        RECT 128.130 88.210 128.390 88.530 ;
        RECT 125.830 87.870 126.090 88.190 ;
        RECT 127.670 87.870 127.930 88.190 ;
        RECT 125.370 87.530 125.630 87.850 ;
        RECT 124.910 86.170 125.170 86.490 ;
        RECT 122.150 84.470 122.410 84.790 ;
        RECT 121.690 79.710 121.950 80.030 ;
        RECT 120.310 79.030 120.570 79.350 ;
        RECT 120.770 79.030 121.030 79.350 ;
        RECT 120.370 77.990 120.510 79.030 ;
        RECT 120.310 77.670 120.570 77.990 ;
        RECT 119.850 74.270 120.110 74.590 ;
        RECT 120.830 72.210 120.970 79.030 ;
        RECT 121.230 74.270 121.490 74.590 ;
        RECT 120.770 71.890 121.030 72.210 ;
        RECT 119.390 69.510 119.650 69.830 ;
        RECT 113.410 68.490 113.670 68.810 ;
        RECT 116.690 68.750 117.750 68.890 ;
        RECT 118.470 68.830 118.730 69.150 ;
        RECT 120.830 68.810 120.970 71.890 ;
        RECT 115.710 68.150 115.970 68.470 ;
        RECT 111.570 66.790 111.830 67.110 ;
        RECT 111.110 66.450 111.370 66.770 ;
        RECT 110.650 66.110 110.910 66.430 ;
        RECT 106.510 63.390 106.770 63.710 ;
        RECT 108.350 63.390 108.610 63.710 ;
        RECT 105.130 61.350 105.390 61.670 ;
        RECT 106.570 61.330 106.710 63.390 ;
        RECT 103.750 61.240 104.010 61.330 ;
        RECT 103.350 61.100 104.010 61.240 ;
        RECT 101.910 57.950 102.170 58.270 ;
        RECT 103.350 56.200 103.490 61.100 ;
        RECT 103.750 61.010 104.010 61.100 ;
        RECT 106.510 61.010 106.770 61.330 ;
        RECT 108.810 61.010 109.070 61.330 ;
        RECT 112.490 61.240 112.750 61.330 ;
        RECT 111.630 61.100 112.750 61.240 ;
        RECT 105.870 59.455 107.410 59.825 ;
        RECT 106.510 58.180 106.770 58.270 ;
        RECT 106.110 58.040 106.770 58.180 ;
        RECT 106.110 56.200 106.250 58.040 ;
        RECT 106.510 57.950 106.770 58.040 ;
        RECT 108.870 56.200 109.010 61.010 ;
        RECT 109.270 59.990 109.530 60.310 ;
        RECT 109.330 59.290 109.470 59.990 ;
        RECT 109.270 58.970 109.530 59.290 ;
        RECT 111.630 56.200 111.770 61.100 ;
        RECT 112.490 61.010 112.750 61.100 ;
        RECT 114.790 58.180 115.050 58.270 ;
        RECT 115.770 58.180 115.910 68.150 ;
        RECT 116.630 61.240 116.890 61.330 ;
        RECT 117.610 61.240 117.750 68.750 ;
        RECT 120.770 68.490 121.030 68.810 ;
        RECT 118.470 68.150 118.730 68.470 ;
        RECT 119.850 68.380 120.110 68.470 ;
        RECT 118.990 68.240 120.110 68.380 ;
        RECT 118.530 66.090 118.670 68.150 ;
        RECT 118.470 65.770 118.730 66.090 ;
        RECT 118.530 62.010 118.670 65.770 ;
        RECT 118.990 63.710 119.130 68.240 ;
        RECT 119.850 68.150 120.110 68.240 ;
        RECT 121.290 66.770 121.430 74.270 ;
        RECT 121.750 69.150 121.890 79.710 ;
        RECT 122.210 76.970 122.350 84.470 ;
        RECT 122.660 83.935 124.200 84.305 ;
        RECT 123.530 81.750 123.790 82.070 ;
        RECT 123.590 81.050 123.730 81.750 ;
        RECT 123.530 80.730 123.790 81.050 ;
        RECT 123.530 79.710 123.790 80.030 ;
        RECT 123.590 79.350 123.730 79.710 ;
        RECT 125.430 79.690 125.570 87.530 ;
        RECT 127.210 85.150 127.470 85.470 ;
        RECT 127.270 83.770 127.410 85.150 ;
        RECT 127.210 83.450 127.470 83.770 ;
        RECT 127.730 82.070 127.870 87.870 ;
        RECT 132.330 86.490 132.470 93.650 ;
        RECT 132.730 92.630 132.990 92.950 ;
        RECT 132.790 90.570 132.930 92.630 ;
        RECT 132.730 90.250 132.990 90.570 ;
        RECT 133.710 89.210 133.850 93.650 ;
        RECT 133.650 88.890 133.910 89.210 ;
        RECT 135.550 87.850 135.690 96.030 ;
        RECT 137.390 94.310 137.530 96.030 ;
        RECT 137.330 93.990 137.590 94.310 ;
        RECT 137.390 91.930 137.530 93.990 ;
        RECT 137.850 93.970 137.990 96.030 ;
        RECT 138.770 94.650 138.910 96.030 ;
        RECT 141.070 94.650 141.210 96.030 ;
        RECT 138.710 94.330 138.970 94.650 ;
        RECT 141.010 94.330 141.270 94.650 ;
        RECT 137.790 93.650 138.050 93.970 ;
        RECT 137.330 91.610 137.590 91.930 ;
        RECT 135.490 87.530 135.750 87.850 ;
        RECT 137.850 86.490 137.990 93.650 ;
        RECT 141.470 93.310 141.730 93.630 ;
        RECT 139.450 92.095 140.990 92.465 ;
        RECT 141.530 91.250 141.670 93.310 ;
        RECT 141.990 91.590 142.130 97.050 ;
        RECT 143.830 96.690 143.970 111.670 ;
        RECT 144.750 108.250 144.890 112.690 ;
        RECT 145.210 112.330 145.350 117.110 ;
        RECT 145.670 112.670 145.810 120.510 ;
        RECT 146.130 118.110 146.270 126.970 ;
        RECT 147.450 126.630 147.710 126.950 ;
        RECT 146.990 126.290 147.250 126.610 ;
        RECT 147.050 126.010 147.190 126.290 ;
        RECT 146.590 125.870 147.190 126.010 ;
        RECT 146.590 125.590 146.730 125.870 ;
        RECT 146.530 125.270 146.790 125.590 ;
        RECT 146.590 118.790 146.730 125.270 ;
        RECT 146.530 118.470 146.790 118.790 ;
        RECT 147.510 118.450 147.650 126.630 ;
        RECT 150.670 125.610 150.930 125.930 ;
        RECT 150.730 121.510 150.870 125.610 ;
        RECT 151.130 125.270 151.390 125.590 ;
        RECT 151.190 123.550 151.330 125.270 ;
        RECT 154.410 123.550 154.550 128.670 ;
        RECT 156.240 127.455 157.780 127.825 ;
        RECT 151.130 123.230 151.390 123.550 ;
        RECT 154.350 123.230 154.610 123.550 ;
        RECT 150.670 121.190 150.930 121.510 ;
        RECT 154.410 121.170 154.550 123.230 ;
        RECT 156.240 122.015 157.780 122.385 ;
        RECT 154.350 120.850 154.610 121.170 ;
        RECT 151.130 118.810 151.390 119.130 ;
        RECT 147.450 118.130 147.710 118.450 ;
        RECT 146.070 117.790 146.330 118.110 ;
        RECT 146.530 117.790 146.790 118.110 ;
        RECT 146.590 116.410 146.730 117.790 ;
        RECT 146.530 116.090 146.790 116.410 ;
        RECT 151.190 116.370 151.330 118.810 ;
        RECT 154.410 118.450 154.550 120.850 ;
        RECT 154.350 118.130 154.610 118.450 ;
        RECT 152.970 117.450 153.230 117.770 ;
        RECT 153.030 116.410 153.170 117.450 ;
        RECT 151.190 116.230 152.250 116.370 ;
        RECT 145.610 112.350 145.870 112.670 ;
        RECT 145.150 112.010 145.410 112.330 ;
        RECT 146.590 110.290 146.730 116.090 ;
        RECT 149.750 115.750 150.010 116.070 ;
        RECT 146.530 109.970 146.790 110.290 ;
        RECT 144.690 107.930 144.950 108.250 ;
        RECT 144.230 103.510 144.490 103.830 ;
        RECT 144.290 101.790 144.430 103.510 ;
        RECT 149.810 102.130 149.950 115.750 ;
        RECT 152.110 115.730 152.250 116.230 ;
        RECT 152.970 116.090 153.230 116.410 ;
        RECT 154.410 116.070 154.550 118.130 ;
        RECT 156.240 116.575 157.780 116.945 ;
        RECT 154.350 115.750 154.610 116.070 ;
        RECT 152.050 115.410 152.310 115.730 ;
        RECT 154.410 113.690 154.550 115.750 ;
        RECT 154.350 113.370 154.610 113.690 ;
        RECT 156.240 111.135 157.780 111.505 ;
        RECT 156.240 105.695 157.780 106.065 ;
        RECT 149.750 101.810 150.010 102.130 ;
        RECT 144.230 101.470 144.490 101.790 ;
        RECT 145.610 96.710 145.870 97.030 ;
        RECT 143.770 96.370 144.030 96.690 ;
        RECT 142.850 95.690 143.110 96.010 ;
        RECT 143.770 95.690 144.030 96.010 ;
        RECT 141.930 91.270 142.190 91.590 ;
        RECT 141.470 90.930 141.730 91.250 ;
        RECT 138.710 90.590 138.970 90.910 ;
        RECT 132.270 86.170 132.530 86.490 ;
        RECT 137.790 86.170 138.050 86.490 ;
        RECT 138.770 85.810 138.910 90.590 ;
        RECT 139.450 86.655 140.990 87.025 ;
        RECT 138.710 85.490 138.970 85.810 ;
        RECT 132.730 85.150 132.990 85.470 ;
        RECT 134.110 85.150 134.370 85.470 ;
        RECT 137.330 85.150 137.590 85.470 ;
        RECT 128.590 84.470 128.850 84.790 ;
        RECT 127.670 81.750 127.930 82.070 ;
        RECT 127.730 80.710 127.870 81.750 ;
        RECT 128.650 81.050 128.790 84.470 ;
        RECT 132.790 83.770 132.930 85.150 ;
        RECT 134.170 83.770 134.310 85.150 ;
        RECT 132.730 83.450 132.990 83.770 ;
        RECT 134.110 83.450 134.370 83.770 ;
        RECT 135.030 82.770 135.290 83.090 ;
        RECT 135.950 82.770 136.210 83.090 ;
        RECT 128.590 80.730 128.850 81.050 ;
        RECT 127.670 80.450 127.930 80.710 ;
        RECT 126.810 80.390 127.930 80.450 ;
        RECT 125.830 80.050 126.090 80.370 ;
        RECT 126.810 80.310 127.870 80.390 ;
        RECT 124.450 79.370 124.710 79.690 ;
        RECT 125.370 79.370 125.630 79.690 ;
        RECT 123.530 79.030 123.790 79.350 ;
        RECT 122.660 78.495 124.200 78.865 ;
        RECT 122.150 76.650 122.410 76.970 ;
        RECT 124.510 74.590 124.650 79.370 ;
        RECT 125.890 77.990 126.030 80.050 ;
        RECT 125.830 77.670 126.090 77.990 ;
        RECT 125.890 75.270 126.030 77.670 ;
        RECT 126.810 76.630 126.950 80.310 ;
        RECT 127.210 79.710 127.470 80.030 ;
        RECT 133.650 79.710 133.910 80.030 ;
        RECT 134.570 79.710 134.830 80.030 ;
        RECT 127.270 78.330 127.410 79.710 ;
        RECT 130.430 79.030 130.690 79.350 ;
        RECT 130.890 79.030 131.150 79.350 ;
        RECT 130.490 78.330 130.630 79.030 ;
        RECT 127.210 78.010 127.470 78.330 ;
        RECT 130.430 78.010 130.690 78.330 ;
        RECT 126.750 76.310 127.010 76.630 ;
        RECT 126.810 75.270 126.950 76.310 ;
        RECT 125.830 74.950 126.090 75.270 ;
        RECT 126.750 74.950 127.010 75.270 ;
        RECT 125.890 74.590 126.030 74.950 ;
        RECT 124.450 74.270 124.710 74.590 ;
        RECT 125.830 74.500 126.090 74.590 ;
        RECT 125.830 74.360 126.490 74.500 ;
        RECT 125.830 74.270 126.090 74.360 ;
        RECT 125.830 73.590 126.090 73.910 ;
        RECT 122.660 73.055 124.200 73.425 ;
        RECT 125.370 71.550 125.630 71.870 ;
        RECT 125.430 69.830 125.570 71.550 ;
        RECT 125.370 69.510 125.630 69.830 ;
        RECT 124.910 69.170 125.170 69.490 ;
        RECT 121.690 68.830 121.950 69.150 ;
        RECT 123.530 68.380 123.790 68.470 ;
        RECT 123.530 68.240 124.650 68.380 ;
        RECT 123.530 68.150 123.790 68.240 ;
        RECT 122.660 67.615 124.200 67.985 ;
        RECT 124.510 67.110 124.650 68.240 ;
        RECT 124.450 66.790 124.710 67.110 ;
        RECT 124.970 66.770 125.110 69.170 ;
        RECT 125.890 66.770 126.030 73.590 ;
        RECT 126.350 72.210 126.490 74.360 ;
        RECT 126.810 72.290 126.950 74.950 ;
        RECT 127.270 73.910 127.410 78.010 ;
        RECT 129.050 74.500 129.310 74.590 ;
        RECT 128.650 74.360 129.310 74.500 ;
        RECT 127.210 73.590 127.470 73.910 ;
        RECT 126.810 72.210 127.410 72.290 ;
        RECT 126.290 71.890 126.550 72.210 ;
        RECT 126.810 72.150 127.470 72.210 ;
        RECT 127.210 71.890 127.470 72.150 ;
        RECT 128.650 71.870 128.790 74.360 ;
        RECT 129.050 74.270 129.310 74.360 ;
        RECT 129.970 73.930 130.230 74.250 ;
        RECT 129.050 73.590 129.310 73.910 ;
        RECT 129.110 72.890 129.250 73.590 ;
        RECT 129.050 72.570 129.310 72.890 ;
        RECT 129.510 72.570 129.770 72.890 ;
        RECT 128.590 71.550 128.850 71.870 ;
        RECT 127.210 70.870 127.470 71.190 ;
        RECT 127.270 69.830 127.410 70.870 ;
        RECT 127.210 69.510 127.470 69.830 ;
        RECT 128.650 68.810 128.790 71.550 ;
        RECT 129.050 71.100 129.310 71.190 ;
        RECT 129.570 71.100 129.710 72.570 ;
        RECT 130.030 71.190 130.170 73.930 ;
        RECT 130.430 71.890 130.690 72.210 ;
        RECT 129.050 70.960 129.710 71.100 ;
        RECT 129.050 70.870 129.310 70.960 ;
        RECT 129.970 70.870 130.230 71.190 ;
        RECT 128.590 68.490 128.850 68.810 ;
        RECT 129.110 66.770 129.250 70.870 ;
        RECT 130.490 69.490 130.630 71.890 ;
        RECT 130.430 69.170 130.690 69.490 ;
        RECT 121.230 66.450 121.490 66.770 ;
        RECT 124.910 66.450 125.170 66.770 ;
        RECT 125.830 66.450 126.090 66.770 ;
        RECT 129.050 66.450 129.310 66.770 ;
        RECT 121.690 65.770 121.950 66.090 ;
        RECT 118.930 63.390 119.190 63.710 ;
        RECT 120.310 63.620 120.570 63.710 ;
        RECT 119.910 63.480 120.570 63.620 ;
        RECT 118.470 61.690 118.730 62.010 ;
        RECT 119.390 61.350 119.650 61.670 ;
        RECT 116.630 61.100 117.750 61.240 ;
        RECT 116.630 61.010 116.890 61.100 ;
        RECT 118.470 60.670 118.730 60.990 ;
        RECT 118.530 59.290 118.670 60.670 ;
        RECT 118.470 58.970 118.730 59.290 ;
        RECT 114.790 58.040 115.910 58.180 ;
        RECT 114.790 57.950 115.050 58.040 ;
        RECT 116.630 57.950 116.890 58.270 ;
        RECT 114.390 56.510 114.990 56.650 ;
        RECT 114.390 56.200 114.530 56.510 ;
        RECT 73.450 55.830 74.510 55.970 ;
        RECT 67.400 54.200 67.690 54.500 ;
        RECT 70.160 54.200 70.450 54.660 ;
        RECT 72.920 54.200 73.210 54.900 ;
        RECT 75.680 54.730 75.960 56.200 ;
        RECT 78.440 54.900 78.720 56.200 ;
        RECT 75.680 54.200 75.970 54.730 ;
        RECT 78.440 54.200 78.730 54.900 ;
        RECT 81.200 54.700 81.480 56.200 ;
        RECT 83.960 54.950 84.240 56.200 ;
        RECT 81.200 54.200 81.490 54.700 ;
        RECT 83.960 54.200 84.250 54.950 ;
        RECT 86.720 54.810 87.000 56.200 ;
        RECT 89.480 54.830 89.760 56.200 ;
        RECT 92.240 54.860 92.520 56.200 ;
        RECT 86.720 54.200 87.010 54.810 ;
        RECT 89.480 54.200 89.770 54.830 ;
        RECT 92.240 54.200 92.530 54.860 ;
        RECT 95.000 54.780 95.280 56.200 ;
        RECT 97.760 54.780 98.040 56.200 ;
        RECT 100.520 54.830 100.800 56.200 ;
        RECT 95.000 54.200 95.290 54.780 ;
        RECT 97.760 54.200 98.050 54.780 ;
        RECT 100.520 54.200 100.810 54.830 ;
        RECT 103.280 54.730 103.560 56.200 ;
        RECT 103.280 54.200 103.570 54.730 ;
        RECT 106.040 54.660 106.320 56.200 ;
        RECT 106.040 54.200 106.330 54.660 ;
        RECT 108.800 54.560 109.080 56.200 ;
        RECT 108.800 54.200 109.090 54.560 ;
        RECT 111.560 54.500 111.840 56.200 ;
        RECT 114.320 54.500 114.600 56.200 ;
        RECT 114.850 55.970 114.990 56.510 ;
        RECT 116.690 55.970 116.830 57.950 ;
        RECT 117.150 56.510 117.750 56.650 ;
        RECT 117.150 56.200 117.290 56.510 ;
        RECT 114.850 55.830 116.830 55.970 ;
        RECT 117.080 54.500 117.360 56.200 ;
        RECT 117.610 55.970 117.750 56.510 ;
        RECT 119.450 55.970 119.590 61.350 ;
        RECT 119.910 56.200 120.050 63.480 ;
        RECT 120.310 63.390 120.570 63.480 ;
        RECT 121.750 58.270 121.890 65.770 ;
        RECT 122.150 65.430 122.410 65.750 ;
        RECT 124.910 65.430 125.170 65.750 ;
        RECT 127.670 65.430 127.930 65.750 ;
        RECT 122.210 63.710 122.350 65.430 ;
        RECT 122.150 63.390 122.410 63.710 ;
        RECT 122.660 62.175 124.200 62.545 ;
        RECT 124.970 62.010 125.110 65.430 ;
        RECT 126.290 63.620 126.550 63.710 ;
        RECT 125.890 63.480 126.550 63.620 ;
        RECT 124.910 61.690 125.170 62.010 ;
        RECT 125.370 59.990 125.630 60.310 ;
        RECT 125.430 59.290 125.570 59.990 ;
        RECT 125.370 58.970 125.630 59.290 ;
        RECT 125.890 58.690 126.030 63.480 ;
        RECT 126.290 63.390 126.550 63.480 ;
        RECT 127.210 63.390 127.470 63.710 ;
        RECT 127.270 61.330 127.410 63.390 ;
        RECT 127.210 61.010 127.470 61.330 ;
        RECT 125.430 58.550 126.030 58.690 ;
        RECT 121.230 57.950 121.490 58.270 ;
        RECT 121.690 57.950 121.950 58.270 ;
        RECT 117.610 55.830 119.590 55.970 ;
        RECT 119.840 54.500 120.120 56.200 ;
        RECT 121.290 55.970 121.430 57.950 ;
        RECT 122.660 56.735 124.200 57.105 ;
        RECT 122.210 56.340 122.810 56.480 ;
        RECT 122.210 55.970 122.350 56.340 ;
        RECT 122.670 56.200 122.810 56.340 ;
        RECT 125.430 56.200 125.570 58.550 ;
        RECT 127.730 58.270 127.870 65.430 ;
        RECT 129.510 63.390 129.770 63.710 ;
        RECT 129.570 59.290 129.710 63.390 ;
        RECT 130.490 61.670 130.630 69.170 ;
        RECT 130.950 69.150 131.090 79.030 ;
        RECT 132.730 76.990 132.990 77.310 ;
        RECT 131.350 76.310 131.610 76.630 ;
        RECT 132.270 76.310 132.530 76.630 ;
        RECT 131.410 75.270 131.550 76.310 ;
        RECT 131.350 74.950 131.610 75.270 ;
        RECT 132.330 72.210 132.470 76.310 ;
        RECT 132.790 75.610 132.930 76.990 ;
        RECT 132.730 75.290 132.990 75.610 ;
        RECT 132.790 74.590 132.930 75.290 ;
        RECT 133.190 74.950 133.450 75.270 ;
        RECT 133.250 74.590 133.390 74.950 ;
        RECT 132.730 74.270 132.990 74.590 ;
        RECT 133.190 74.270 133.450 74.590 ;
        RECT 132.730 73.590 132.990 73.910 ;
        RECT 132.790 72.890 132.930 73.590 ;
        RECT 132.730 72.570 132.990 72.890 ;
        RECT 132.270 71.890 132.530 72.210 ;
        RECT 132.730 69.510 132.990 69.830 ;
        RECT 130.890 68.830 131.150 69.150 ;
        RECT 130.950 66.770 131.090 68.830 ;
        RECT 132.790 66.770 132.930 69.510 ;
        RECT 130.890 66.450 131.150 66.770 ;
        RECT 132.730 66.450 132.990 66.770 ;
        RECT 133.250 63.710 133.390 74.270 ;
        RECT 133.710 73.820 133.850 79.710 ;
        RECT 134.630 75.610 134.770 79.710 ;
        RECT 134.570 75.290 134.830 75.610 ;
        RECT 133.710 73.680 134.310 73.820 ;
        RECT 133.650 71.890 133.910 72.210 ;
        RECT 133.710 69.830 133.850 71.890 ;
        RECT 133.650 69.510 133.910 69.830 ;
        RECT 134.170 67.450 134.310 73.680 ;
        RECT 134.630 72.890 134.770 75.290 ;
        RECT 134.570 72.570 134.830 72.890 ;
        RECT 135.090 71.870 135.230 82.770 ;
        RECT 136.010 81.050 136.150 82.770 ;
        RECT 137.390 82.750 137.530 85.150 ;
        RECT 137.330 82.430 137.590 82.750 ;
        RECT 138.770 81.050 138.910 85.490 ;
        RECT 141.530 83.770 141.670 90.930 ;
        RECT 142.390 87.190 142.650 87.510 ;
        RECT 142.450 85.470 142.590 87.190 ;
        RECT 142.390 85.150 142.650 85.470 ;
        RECT 141.470 83.450 141.730 83.770 ;
        RECT 141.470 82.090 141.730 82.410 ;
        RECT 139.450 81.215 140.990 81.585 ;
        RECT 135.950 80.730 136.210 81.050 ;
        RECT 138.710 80.730 138.970 81.050 ;
        RECT 138.710 79.710 138.970 80.030 ;
        RECT 136.870 77.330 137.130 77.650 ;
        RECT 135.490 76.310 135.750 76.630 ;
        RECT 135.030 71.550 135.290 71.870 ;
        RECT 135.550 71.190 135.690 76.310 ;
        RECT 135.950 75.290 136.210 75.610 ;
        RECT 135.490 70.870 135.750 71.190 ;
        RECT 135.550 67.450 135.690 70.870 ;
        RECT 136.010 68.470 136.150 75.290 ;
        RECT 136.930 74.840 137.070 77.330 ;
        RECT 138.770 74.930 138.910 79.710 ;
        RECT 141.530 76.630 141.670 82.090 ;
        RECT 142.390 80.730 142.650 81.050 ;
        RECT 141.470 76.310 141.730 76.630 ;
        RECT 139.450 75.775 140.990 76.145 ;
        RECT 136.930 74.700 137.990 74.840 ;
        RECT 136.410 74.270 136.670 74.590 ;
        RECT 136.470 72.890 136.610 74.270 ;
        RECT 137.330 73.590 137.590 73.910 ;
        RECT 137.390 72.890 137.530 73.590 ;
        RECT 136.410 72.570 136.670 72.890 ;
        RECT 137.330 72.570 137.590 72.890 ;
        RECT 136.870 68.830 137.130 69.150 ;
        RECT 135.950 68.150 136.210 68.470 ;
        RECT 136.930 68.070 137.070 68.830 ;
        RECT 137.850 68.810 137.990 74.700 ;
        RECT 138.710 74.610 138.970 74.930 ;
        RECT 141.010 74.270 141.270 74.590 ;
        RECT 141.070 72.890 141.210 74.270 ;
        RECT 141.010 72.570 141.270 72.890 ;
        RECT 141.470 71.210 141.730 71.530 ;
        RECT 138.710 70.870 138.970 71.190 ;
        RECT 138.770 70.170 138.910 70.870 ;
        RECT 139.450 70.335 140.990 70.705 ;
        RECT 138.710 69.850 138.970 70.170 ;
        RECT 141.530 69.150 141.670 71.210 ;
        RECT 141.470 68.830 141.730 69.150 ;
        RECT 137.790 68.490 138.050 68.810 ;
        RECT 136.470 67.930 137.070 68.070 ;
        RECT 134.110 67.130 134.370 67.450 ;
        RECT 135.490 67.130 135.750 67.450 ;
        RECT 132.730 63.390 132.990 63.710 ;
        RECT 133.190 63.390 133.450 63.710 ;
        RECT 130.430 61.350 130.690 61.670 ;
        RECT 129.970 61.010 130.230 61.330 ;
        RECT 129.510 58.970 129.770 59.290 ;
        RECT 127.670 57.950 127.930 58.270 ;
        RECT 128.190 56.510 128.790 56.650 ;
        RECT 128.190 56.200 128.330 56.510 ;
        RECT 121.290 55.830 122.350 55.970 ;
        RECT 122.600 54.500 122.880 56.200 ;
        RECT 125.360 54.690 125.640 56.200 ;
        RECT 111.560 54.200 111.850 54.500 ;
        RECT 114.320 54.200 114.610 54.500 ;
        RECT 117.080 54.200 117.370 54.500 ;
        RECT 119.840 54.200 120.130 54.500 ;
        RECT 122.600 54.200 122.890 54.500 ;
        RECT 125.360 54.200 125.650 54.690 ;
        RECT 128.120 54.640 128.400 56.200 ;
        RECT 128.650 55.970 128.790 56.510 ;
        RECT 130.030 55.970 130.170 61.010 ;
        RECT 132.270 60.670 132.530 60.990 ;
        RECT 132.330 59.290 132.470 60.670 ;
        RECT 132.790 59.290 132.930 63.390 ;
        RECT 134.170 62.010 134.310 67.130 ;
        RECT 136.470 66.430 136.610 67.930 ;
        RECT 136.410 66.110 136.670 66.430 ;
        RECT 136.410 63.390 136.670 63.710 ;
        RECT 134.110 61.690 134.370 62.010 ;
        RECT 134.110 61.010 134.370 61.330 ;
        RECT 132.270 58.970 132.530 59.290 ;
        RECT 132.730 58.970 132.990 59.290 ;
        RECT 131.810 58.180 132.070 58.270 ;
        RECT 130.950 58.040 132.070 58.180 ;
        RECT 130.950 56.200 131.090 58.040 ;
        RECT 131.810 57.950 132.070 58.040 ;
        RECT 134.170 58.010 134.310 61.010 ;
        RECT 133.710 57.870 134.310 58.010 ;
        RECT 133.710 56.200 133.850 57.870 ;
        RECT 136.470 56.200 136.610 63.390 ;
        RECT 137.850 58.270 137.990 68.490 ;
        RECT 142.450 66.770 142.590 80.730 ;
        RECT 142.910 80.030 143.050 95.690 ;
        RECT 143.830 94.310 143.970 95.690 ;
        RECT 143.770 93.990 144.030 94.310 ;
        RECT 143.830 92.950 143.970 93.990 ;
        RECT 145.670 93.970 145.810 96.710 ;
        RECT 147.910 96.030 148.170 96.350 ;
        RECT 146.070 95.350 146.330 95.670 ;
        RECT 145.610 93.650 145.870 93.970 ;
        RECT 145.150 93.310 145.410 93.630 ;
        RECT 143.770 92.630 144.030 92.950 ;
        RECT 145.210 90.910 145.350 93.310 ;
        RECT 146.130 91.250 146.270 95.350 ;
        RECT 147.450 93.650 147.710 93.970 ;
        RECT 146.530 92.630 146.790 92.950 ;
        RECT 146.590 91.250 146.730 92.630 ;
        RECT 146.070 90.930 146.330 91.250 ;
        RECT 146.530 90.930 146.790 91.250 ;
        RECT 145.150 90.590 145.410 90.910 ;
        RECT 146.990 90.590 147.250 90.910 ;
        RECT 145.150 88.210 145.410 88.530 ;
        RECT 144.690 87.870 144.950 88.190 ;
        RECT 144.750 86.490 144.890 87.870 ;
        RECT 144.690 86.170 144.950 86.490 ;
        RECT 142.850 79.710 143.110 80.030 ;
        RECT 145.210 78.330 145.350 88.210 ;
        RECT 147.050 83.770 147.190 90.590 ;
        RECT 147.510 90.230 147.650 93.650 ;
        RECT 147.970 91.930 148.110 96.030 ;
        RECT 149.810 94.650 149.950 101.810 ;
        RECT 156.240 100.255 157.780 100.625 ;
        RECT 151.130 95.690 151.390 96.010 ;
        RECT 151.190 94.650 151.330 95.690 ;
        RECT 156.240 94.815 157.780 95.185 ;
        RECT 149.750 94.330 150.010 94.650 ;
        RECT 151.130 94.330 151.390 94.650 ;
        RECT 147.910 91.610 148.170 91.930 ;
        RECT 147.450 89.910 147.710 90.230 ;
        RECT 156.240 89.375 157.780 89.745 ;
        RECT 147.910 87.190 148.170 87.510 ;
        RECT 148.370 87.190 148.630 87.510 ;
        RECT 148.830 87.190 149.090 87.510 ;
        RECT 147.970 86.490 148.110 87.190 ;
        RECT 147.910 86.170 148.170 86.490 ;
        RECT 148.430 85.130 148.570 87.190 ;
        RECT 148.890 86.150 149.030 87.190 ;
        RECT 148.830 85.830 149.090 86.150 ;
        RECT 148.370 84.810 148.630 85.130 ;
        RECT 146.990 83.450 147.250 83.770 ;
        RECT 148.430 82.750 148.570 84.810 ;
        RECT 148.890 83.090 149.030 85.830 ;
        RECT 150.670 85.150 150.930 85.470 ;
        RECT 148.830 82.770 149.090 83.090 ;
        RECT 150.730 82.750 150.870 85.150 ;
        RECT 156.240 83.935 157.780 84.305 ;
        RECT 148.370 82.430 148.630 82.750 ;
        RECT 150.670 82.430 150.930 82.750 ;
        RECT 148.830 80.390 149.090 80.710 ;
        RECT 147.910 79.710 148.170 80.030 ;
        RECT 145.150 78.010 145.410 78.330 ;
        RECT 147.970 77.650 148.110 79.710 ;
        RECT 148.890 78.330 149.030 80.390 ;
        RECT 150.210 79.710 150.470 80.030 ;
        RECT 148.830 78.010 149.090 78.330 ;
        RECT 148.890 77.650 149.030 78.010 ;
        RECT 150.270 77.650 150.410 79.710 ;
        RECT 150.730 78.330 150.870 82.430 ;
        RECT 151.590 80.730 151.850 81.050 ;
        RECT 150.670 78.010 150.930 78.330 ;
        RECT 147.910 77.330 148.170 77.650 ;
        RECT 148.830 77.330 149.090 77.650 ;
        RECT 150.210 77.330 150.470 77.650 ;
        RECT 147.450 76.650 147.710 76.970 ;
        RECT 147.510 75.610 147.650 76.650 ;
        RECT 147.450 75.290 147.710 75.610 ;
        RECT 144.690 73.590 144.950 73.910 ;
        RECT 144.750 72.890 144.890 73.590 ;
        RECT 144.690 72.570 144.950 72.890 ;
        RECT 142.850 70.870 143.110 71.190 ;
        RECT 142.910 70.170 143.050 70.870 ;
        RECT 147.970 70.170 148.110 77.330 ;
        RECT 148.370 73.590 148.630 73.910 ;
        RECT 148.430 72.890 148.570 73.590 ;
        RECT 148.370 72.570 148.630 72.890 ;
        RECT 148.890 71.870 149.030 77.330 ;
        RECT 151.650 75.610 151.790 80.730 ;
        RECT 153.890 79.030 154.150 79.350 ;
        RECT 152.050 77.670 152.310 77.990 ;
        RECT 151.590 75.290 151.850 75.610 ;
        RECT 148.830 71.550 149.090 71.870 ;
        RECT 152.110 71.530 152.250 77.670 ;
        RECT 153.950 77.310 154.090 79.030 ;
        RECT 156.240 78.495 157.780 78.865 ;
        RECT 153.890 76.990 154.150 77.310 ;
        RECT 154.350 76.310 154.610 76.630 ;
        RECT 154.410 74.250 154.550 76.310 ;
        RECT 154.350 73.930 154.610 74.250 ;
        RECT 156.240 73.055 157.780 73.425 ;
        RECT 148.370 71.210 148.630 71.530 ;
        RECT 152.050 71.210 152.310 71.530 ;
        RECT 142.850 69.850 143.110 70.170 ;
        RECT 147.910 69.850 148.170 70.170 ;
        RECT 145.610 68.830 145.870 69.150 ;
        RECT 144.230 68.150 144.490 68.470 ;
        RECT 145.150 68.150 145.410 68.470 ;
        RECT 141.930 66.450 142.190 66.770 ;
        RECT 142.390 66.450 142.650 66.770 ;
        RECT 139.450 64.895 140.990 65.265 ;
        RECT 138.710 63.390 138.970 63.710 ;
        RECT 138.250 60.670 138.510 60.990 ;
        RECT 138.310 59.290 138.450 60.670 ;
        RECT 138.250 58.970 138.510 59.290 ;
        RECT 138.770 58.610 138.910 63.390 ;
        RECT 141.470 61.010 141.730 61.330 ;
        RECT 139.450 59.455 140.990 59.825 ;
        RECT 138.710 58.290 138.970 58.610 ;
        RECT 137.790 57.950 138.050 58.270 ;
        RECT 139.230 56.510 139.830 56.650 ;
        RECT 139.230 56.200 139.370 56.510 ;
        RECT 128.650 55.830 130.170 55.970 ;
        RECT 130.880 54.640 131.160 56.200 ;
        RECT 128.120 54.200 128.410 54.640 ;
        RECT 130.880 54.200 131.170 54.640 ;
        RECT 133.640 54.540 133.920 56.200 ;
        RECT 136.400 54.690 136.680 56.200 ;
        RECT 133.640 54.200 133.930 54.540 ;
        RECT 136.400 54.200 136.690 54.690 ;
        RECT 139.160 54.590 139.440 56.200 ;
        RECT 139.690 55.970 139.830 56.510 ;
        RECT 141.530 55.970 141.670 61.010 ;
        RECT 141.990 56.200 142.130 66.450 ;
        RECT 144.290 63.710 144.430 68.150 ;
        RECT 145.210 67.110 145.350 68.150 ;
        RECT 145.150 66.790 145.410 67.110 ;
        RECT 144.230 63.390 144.490 63.710 ;
        RECT 145.670 61.330 145.810 68.830 ;
        RECT 148.430 68.810 148.570 71.210 ;
        RECT 148.370 68.490 148.630 68.810 ;
        RECT 150.210 68.490 150.470 68.810 ;
        RECT 150.270 67.450 150.410 68.490 ;
        RECT 156.240 67.615 157.780 67.985 ;
        RECT 150.210 67.130 150.470 67.450 ;
        RECT 150.210 63.390 150.470 63.710 ;
        RECT 146.530 63.050 146.790 63.370 ;
        RECT 145.610 61.010 145.870 61.330 ;
        RECT 144.230 60.670 144.490 60.990 ;
        RECT 144.290 59.290 144.430 60.670 ;
        RECT 146.590 59.290 146.730 63.050 ;
        RECT 147.450 61.010 147.710 61.330 ;
        RECT 144.230 58.970 144.490 59.290 ;
        RECT 146.530 58.970 146.790 59.290 ;
        RECT 144.690 57.950 144.950 58.270 ;
        RECT 144.750 56.200 144.890 57.950 ;
        RECT 147.510 56.200 147.650 61.010 ;
        RECT 150.270 56.200 150.410 63.390 ;
        RECT 156.240 62.175 157.780 62.545 ;
        RECT 156.240 56.735 157.780 57.105 ;
        RECT 139.690 55.830 141.670 55.970 ;
        RECT 139.160 54.200 139.450 54.590 ;
        RECT 141.920 54.540 142.200 56.200 ;
        RECT 144.680 54.690 144.960 56.200 ;
        RECT 141.920 54.200 142.210 54.540 ;
        RECT 144.680 54.200 144.970 54.690 ;
        RECT 147.440 54.500 147.720 56.200 ;
        RECT 150.200 54.640 150.480 56.200 ;
        RECT 147.440 54.200 147.730 54.500 ;
        RECT 150.200 54.200 150.490 54.640 ;
        RECT 28.770 49.740 29.050 54.200 ;
        RECT 31.530 51.790 31.810 54.200 ;
        RECT 34.290 52.390 34.570 54.200 ;
        RECT 37.050 52.890 37.330 54.200 ;
        RECT 39.810 53.440 40.090 54.200 ;
        RECT 42.570 53.990 42.850 54.200 ;
        RECT 42.570 53.710 43.840 53.990 ;
        RECT 39.810 53.160 41.240 53.440 ;
        RECT 37.050 52.610 39.240 52.890 ;
        RECT 34.290 52.110 37.640 52.390 ;
        RECT 31.530 51.510 36.140 51.790 ;
        RECT 35.860 49.790 36.140 51.510 ;
        RECT 33.850 49.740 34.760 49.745 ;
        RECT 28.770 49.460 34.760 49.740 ;
        RECT 33.850 48.895 34.760 49.460 ;
        RECT 35.860 48.910 36.720 49.790 ;
        RECT 37.360 49.770 37.640 52.110 ;
        RECT 38.960 49.785 39.240 52.610 ;
        RECT 37.360 48.910 38.210 49.770 ;
        RECT 38.935 48.975 39.805 49.785 ;
        RECT 40.960 49.735 41.240 53.160 ;
        RECT 43.560 49.815 43.840 53.710 ;
        RECT 40.900 48.985 41.710 49.735 ;
        RECT 43.560 49.060 44.355 49.815 ;
        RECT 38.960 48.960 39.775 48.975 ;
        RECT 30.280 32.060 32.280 46.760 ;
        RECT 33.880 33.205 34.730 48.895 ;
        RECT 30.280 30.060 35.310 32.060 ;
        RECT 30.280 21.060 32.280 30.060 ;
        RECT 35.880 22.725 36.720 48.910 ;
        RECT 30.280 19.060 36.810 21.060 ;
        RECT 30.280 12.860 32.280 19.060 ;
        RECT 37.390 14.080 38.210 48.910 ;
        RECT 38.965 32.585 39.775 48.960 ;
        RECT 40.930 33.705 41.680 48.985 ;
        RECT 43.605 47.785 44.355 49.060 ;
        RECT 45.330 49.240 45.610 54.200 ;
        RECT 48.090 49.760 48.370 54.200 ;
        RECT 45.830 49.240 46.580 49.760 ;
        RECT 45.330 48.960 46.580 49.240 ;
        RECT 43.605 47.035 45.380 47.785 ;
        RECT 42.430 33.860 43.830 38.040 ;
        RECT 44.630 34.585 45.380 47.035 ;
        RECT 45.830 33.980 46.580 48.960 ;
        RECT 47.980 38.135 48.730 49.760 ;
        RECT 49.830 49.240 50.580 49.765 ;
        RECT 50.850 49.240 51.130 54.200 ;
        RECT 53.610 50.340 53.890 54.200 ;
        RECT 56.370 51.990 56.650 54.200 ;
        RECT 52.160 50.060 53.890 50.340 ;
        RECT 54.210 51.710 56.650 51.990 ;
        RECT 52.160 49.760 52.440 50.060 ;
        RECT 54.210 49.765 54.490 51.710 ;
        RECT 59.130 51.490 59.410 54.200 ;
        RECT 56.160 51.210 59.410 51.490 ;
        RECT 56.160 49.785 56.440 51.210 ;
        RECT 61.890 50.940 62.170 54.200 ;
        RECT 58.010 50.660 62.170 50.940 ;
        RECT 58.010 49.815 58.290 50.660 ;
        RECT 64.650 50.390 64.930 54.200 ;
        RECT 60.200 50.110 64.930 50.390 ;
        RECT 51.630 49.735 52.955 49.760 ;
        RECT 49.810 48.960 51.130 49.240 ;
        RECT 51.625 48.985 52.955 49.735 ;
        RECT 49.830 39.635 50.580 48.960 ;
        RECT 52.205 41.185 52.955 48.985 ;
        RECT 53.705 49.010 54.490 49.765 ;
        RECT 55.625 49.035 57.040 49.785 ;
        RECT 53.705 42.885 54.455 49.010 ;
        RECT 53.705 42.135 55.780 42.885 ;
        RECT 52.205 40.435 54.805 41.185 ;
        RECT 49.830 38.885 53.755 39.635 ;
        RECT 47.980 37.385 50.880 38.135 ;
        RECT 42.430 32.760 45.610 33.860 ;
        RECT 45.830 33.340 49.580 33.980 ;
        RECT 50.105 33.935 50.855 37.385 ;
        RECT 45.830 33.335 46.580 33.340 ;
        RECT 50.105 33.280 52.735 33.935 ;
        RECT 50.105 33.235 50.855 33.280 ;
        RECT 38.965 31.775 40.210 32.585 ;
        RECT 30.280 10.860 38.810 12.860 ;
        RECT 30.280 7.050 32.280 10.860 ;
        RECT 39.400 7.335 40.210 31.775 ;
        RECT 42.430 30.460 43.830 32.760 ;
        RECT 53.005 31.035 53.755 38.885 ;
        RECT 42.430 29.360 50.260 30.460 ;
        RECT 50.905 29.785 53.755 31.035 ;
        RECT 42.430 7.060 43.830 29.360 ;
        RECT 47.600 25.460 49.000 29.360 ;
        RECT 52.005 28.285 52.655 28.315 ;
        RECT 54.055 28.285 54.805 40.435 ;
        RECT 50.955 27.535 54.805 28.285 ;
        RECT 50.955 26.685 52.780 27.535 ;
        RECT 50.955 25.950 52.730 26.685 ;
        RECT 47.600 24.710 51.705 25.460 ;
        RECT 47.600 21.880 49.000 24.710 ;
        RECT 55.030 24.260 55.780 42.135 ;
        RECT 51.035 23.510 55.780 24.260 ;
        RECT 51.035 23.495 53.815 23.510 ;
        RECT 51.035 23.125 51.925 23.495 ;
        RECT 53.065 23.125 53.815 23.495 ;
        RECT 55.030 23.485 55.780 23.510 ;
        RECT 51.035 22.375 53.815 23.125 ;
        RECT 51.175 22.365 51.925 22.375 ;
        RECT 47.600 21.130 51.705 21.880 ;
        RECT 47.600 18.300 49.000 21.130 ;
        RECT 56.290 20.640 57.040 49.035 ;
        RECT 51.035 19.890 57.040 20.640 ;
        RECT 51.115 19.535 51.865 19.890 ;
        RECT 52.715 19.885 55.045 19.890 ;
        RECT 54.295 19.535 55.045 19.885 ;
        RECT 51.115 18.785 55.075 19.535 ;
        RECT 51.115 18.755 51.865 18.785 ;
        RECT 47.600 17.550 51.705 18.300 ;
        RECT 47.600 14.720 49.000 17.550 ;
        RECT 55.855 17.080 56.605 17.105 ;
        RECT 57.550 17.080 58.300 49.815 ;
        RECT 60.200 49.685 60.480 50.110 ;
        RECT 61.425 49.780 63.905 49.785 ;
        RECT 67.410 49.780 67.690 54.200 ;
        RECT 70.170 52.190 70.450 54.200 ;
        RECT 72.930 52.790 73.210 54.200 ;
        RECT 75.690 53.440 75.970 54.200 ;
        RECT 78.450 53.940 78.730 54.200 ;
        RECT 78.450 53.660 80.490 53.940 ;
        RECT 75.690 53.160 78.840 53.440 ;
        RECT 72.930 52.510 77.340 52.790 ;
        RECT 70.170 51.910 75.390 52.190 ;
        RECT 75.110 50.585 75.390 51.910 ;
        RECT 77.060 50.630 77.340 52.510 ;
        RECT 59.675 48.935 60.880 49.685 ;
        RECT 61.425 49.500 67.690 49.780 ;
        RECT 75.070 49.735 75.980 50.585 ;
        RECT 77.060 49.760 77.940 50.630 ;
        RECT 78.560 50.610 78.840 53.160 ;
        RECT 80.210 50.625 80.490 53.660 ;
        RECT 81.210 52.740 81.490 54.200 ;
        RECT 81.210 52.460 82.440 52.740 ;
        RECT 78.560 49.760 79.430 50.610 ;
        RECT 80.155 49.815 81.025 50.625 ;
        RECT 82.160 50.575 82.440 52.460 ;
        RECT 82.120 49.825 82.930 50.575 ;
        RECT 83.970 50.140 84.250 54.200 ;
        RECT 86.730 51.940 87.010 54.200 ;
        RECT 86.730 51.660 87.340 51.940 ;
        RECT 84.825 50.140 85.575 50.655 ;
        RECT 87.060 50.600 87.340 51.660 ;
        RECT 89.490 50.600 89.770 54.200 ;
        RECT 92.250 52.490 92.530 54.200 ;
        RECT 95.010 53.140 95.290 54.200 ;
        RECT 91.560 52.210 92.530 52.490 ;
        RECT 93.360 52.860 95.290 53.140 ;
        RECT 91.560 50.605 91.840 52.210 ;
        RECT 83.970 49.860 85.590 50.140 ;
        RECT 61.425 49.035 63.905 49.500 ;
        RECT 50.955 16.330 58.300 17.080 ;
        RECT 50.985 15.955 51.735 16.330 ;
        RECT 55.855 15.955 56.605 16.330 ;
        RECT 50.985 15.205 56.635 15.955 ;
        RECT 50.985 15.175 51.735 15.205 ;
        RECT 47.600 13.970 51.705 14.720 ;
        RECT 47.600 11.140 49.000 13.970 ;
        RECT 58.385 13.520 59.135 13.535 ;
        RECT 60.130 13.520 60.880 48.935 ;
        RECT 50.935 12.770 60.880 13.520 ;
        RECT 50.965 12.385 51.715 12.770 ;
        RECT 58.385 12.385 59.135 12.770 ;
        RECT 50.965 11.635 59.165 12.385 ;
        RECT 50.965 11.605 51.715 11.635 ;
        RECT 47.600 10.390 51.705 11.140 ;
        RECT 47.600 7.060 49.000 10.390 ;
        RECT 61.905 9.920 62.655 9.945 ;
        RECT 63.155 9.920 63.905 49.035 ;
        RECT 64.450 43.250 65.950 45.780 ;
        RECT 64.420 41.750 65.980 43.250 ;
        RECT 64.450 26.300 65.950 41.750 ;
        RECT 71.500 32.900 73.500 47.600 ;
        RECT 75.100 34.045 75.950 49.735 ;
        RECT 71.500 30.900 76.530 32.900 ;
        RECT 64.420 24.800 65.980 26.300 ;
        RECT 64.450 13.450 65.950 24.800 ;
        RECT 71.500 21.900 73.500 30.900 ;
        RECT 77.100 23.565 77.940 49.760 ;
        RECT 71.500 19.900 78.030 21.900 ;
        RECT 71.500 13.700 73.500 19.900 ;
        RECT 78.610 14.920 79.430 49.760 ;
        RECT 80.185 33.425 80.995 49.815 ;
        RECT 82.150 34.545 82.900 49.825 ;
        RECT 84.825 48.625 85.575 49.860 ;
        RECT 84.825 47.875 86.600 48.625 ;
        RECT 83.650 34.700 85.050 38.880 ;
        RECT 85.850 35.425 86.600 47.875 ;
        RECT 87.050 34.820 87.800 50.600 ;
        RECT 89.200 38.975 89.950 50.600 ;
        RECT 91.050 49.810 91.840 50.605 ;
        RECT 93.360 50.600 93.640 52.860 ;
        RECT 97.770 52.590 98.050 54.200 ;
        RECT 95.410 52.310 98.050 52.590 ;
        RECT 95.410 50.605 95.690 52.310 ;
        RECT 100.530 52.090 100.810 54.200 ;
        RECT 97.360 51.810 100.810 52.090 ;
        RECT 97.360 50.625 97.640 51.810 ;
        RECT 103.290 51.570 103.570 54.200 ;
        RECT 99.260 51.290 103.570 51.570 ;
        RECT 99.260 50.655 99.540 51.290 ;
        RECT 106.050 51.110 106.330 54.200 ;
        RECT 92.850 50.575 94.175 50.600 ;
        RECT 92.845 49.825 94.175 50.575 ;
        RECT 93.360 49.810 94.175 49.825 ;
        RECT 91.050 40.475 91.800 49.810 ;
        RECT 93.425 42.025 94.175 49.810 ;
        RECT 94.925 49.810 95.690 50.605 ;
        RECT 96.845 49.875 98.260 50.625 ;
        RECT 97.360 49.860 98.260 49.875 ;
        RECT 94.925 43.725 95.675 49.810 ;
        RECT 94.925 42.975 97.000 43.725 ;
        RECT 93.425 41.275 96.025 42.025 ;
        RECT 91.050 39.725 94.975 40.475 ;
        RECT 89.200 38.225 92.100 38.975 ;
        RECT 83.650 33.600 86.830 34.700 ;
        RECT 87.050 34.180 90.800 34.820 ;
        RECT 91.325 34.775 92.075 38.225 ;
        RECT 87.050 34.175 87.800 34.180 ;
        RECT 91.325 34.120 93.955 34.775 ;
        RECT 91.325 34.075 92.075 34.120 ;
        RECT 80.185 32.615 81.430 33.425 ;
        RECT 64.420 11.950 65.980 13.450 ;
        RECT 64.450 11.000 65.950 11.950 ;
        RECT 71.500 11.700 80.030 13.700 ;
        RECT 50.965 9.170 63.990 9.920 ;
        RECT 50.995 8.785 51.745 9.170 ;
        RECT 61.905 8.785 62.655 9.170 ;
        RECT 50.995 8.035 62.685 8.785 ;
        RECT 50.995 8.005 51.745 8.035 ;
        RECT 71.500 7.890 73.500 11.700 ;
        RECT 80.620 8.175 81.430 32.615 ;
        RECT 83.650 31.300 85.050 33.600 ;
        RECT 94.225 31.875 94.975 39.725 ;
        RECT 83.650 30.200 91.480 31.300 ;
        RECT 92.125 30.625 94.975 31.875 ;
        RECT 83.650 7.900 85.050 30.200 ;
        RECT 88.820 26.300 90.220 30.200 ;
        RECT 93.225 29.125 93.875 29.155 ;
        RECT 95.275 29.125 96.025 41.275 ;
        RECT 92.175 28.375 96.025 29.125 ;
        RECT 92.175 27.525 94.000 28.375 ;
        RECT 92.175 26.790 93.950 27.525 ;
        RECT 88.820 25.550 92.925 26.300 ;
        RECT 88.820 22.720 90.220 25.550 ;
        RECT 96.250 25.100 97.000 42.975 ;
        RECT 92.255 24.350 97.000 25.100 ;
        RECT 92.255 24.335 95.035 24.350 ;
        RECT 92.255 23.965 93.145 24.335 ;
        RECT 94.285 23.965 95.035 24.335 ;
        RECT 96.250 24.325 97.000 24.350 ;
        RECT 92.255 23.215 95.035 23.965 ;
        RECT 92.395 23.205 93.145 23.215 ;
        RECT 88.820 21.970 92.925 22.720 ;
        RECT 88.820 19.140 90.220 21.970 ;
        RECT 97.510 21.480 98.260 49.860 ;
        RECT 92.255 20.730 98.260 21.480 ;
        RECT 98.770 49.860 99.540 50.655 ;
        RECT 101.400 50.830 106.330 51.110 ;
        RECT 101.400 50.525 101.680 50.830 ;
        RECT 92.335 20.375 93.085 20.730 ;
        RECT 93.935 20.725 96.265 20.730 ;
        RECT 95.515 20.375 96.265 20.725 ;
        RECT 92.335 19.625 96.295 20.375 ;
        RECT 92.335 19.595 93.085 19.625 ;
        RECT 88.820 18.390 92.925 19.140 ;
        RECT 88.820 15.560 90.220 18.390 ;
        RECT 97.075 17.920 97.825 17.945 ;
        RECT 98.770 17.920 99.520 49.860 ;
        RECT 100.895 49.775 102.100 50.525 ;
        RECT 102.645 50.460 105.125 50.625 ;
        RECT 108.810 50.460 109.090 54.200 ;
        RECT 111.570 52.890 111.850 54.200 ;
        RECT 114.330 53.340 114.610 54.200 ;
        RECT 117.090 53.340 117.370 54.200 ;
        RECT 119.850 53.390 120.130 54.200 ;
        RECT 114.330 53.060 116.740 53.340 ;
        RECT 117.090 53.060 119.290 53.340 ;
        RECT 119.850 53.110 120.840 53.390 ;
        RECT 111.570 52.610 115.240 52.890 ;
        RECT 114.960 51.985 115.240 52.610 ;
        RECT 114.950 51.135 115.860 51.985 ;
        RECT 116.460 51.440 116.740 53.060 ;
        RECT 116.980 51.440 117.820 52.030 ;
        RECT 119.010 52.010 119.290 53.060 ;
        RECT 120.560 52.025 120.840 53.110 ;
        RECT 116.460 51.160 117.840 51.440 ;
        RECT 102.645 50.180 109.090 50.460 ;
        RECT 102.645 49.875 105.125 50.180 ;
        RECT 92.175 17.170 99.520 17.920 ;
        RECT 92.205 16.795 92.955 17.170 ;
        RECT 97.075 16.795 97.825 17.170 ;
        RECT 92.205 16.045 97.855 16.795 ;
        RECT 92.205 16.015 92.955 16.045 ;
        RECT 88.820 14.810 92.925 15.560 ;
        RECT 88.820 11.980 90.220 14.810 ;
        RECT 99.605 14.360 100.355 14.375 ;
        RECT 101.350 14.360 102.100 49.775 ;
        RECT 92.155 13.610 102.100 14.360 ;
        RECT 92.185 13.225 92.935 13.610 ;
        RECT 99.605 13.225 100.355 13.610 ;
        RECT 92.185 12.475 100.385 13.225 ;
        RECT 92.185 12.445 92.935 12.475 ;
        RECT 88.820 11.230 92.925 11.980 ;
        RECT 88.820 7.900 90.220 11.230 ;
        RECT 103.125 10.760 103.875 10.785 ;
        RECT 104.375 10.760 105.125 49.875 ;
        RECT 105.700 43.300 107.200 45.830 ;
        RECT 105.670 41.800 107.230 43.300 ;
        RECT 105.700 26.350 107.200 41.800 ;
        RECT 111.380 34.300 113.380 49.000 ;
        RECT 114.980 35.445 115.830 51.135 ;
        RECT 111.380 32.300 116.410 34.300 ;
        RECT 105.670 24.850 107.230 26.350 ;
        RECT 105.700 13.500 107.200 24.850 ;
        RECT 111.380 23.300 113.380 32.300 ;
        RECT 116.980 24.965 117.820 51.160 ;
        RECT 111.380 21.300 117.910 23.300 ;
        RECT 111.380 15.100 113.380 21.300 ;
        RECT 118.490 16.320 119.310 52.010 ;
        RECT 120.035 51.215 120.905 52.025 ;
        RECT 122.610 51.975 122.890 54.200 ;
        RECT 125.370 52.055 125.650 54.200 ;
        RECT 128.130 52.590 128.410 54.200 ;
        RECT 130.890 52.590 131.170 54.200 ;
        RECT 133.650 53.040 133.930 54.200 ;
        RECT 136.410 53.440 136.690 54.200 ;
        RECT 139.170 53.990 139.450 54.200 ;
        RECT 122.000 51.225 122.890 51.975 ;
        RECT 120.065 34.825 120.875 51.215 ;
        RECT 122.030 51.210 122.890 51.225 ;
        RECT 124.705 51.260 125.650 52.055 ;
        RECT 127.410 52.310 128.410 52.590 ;
        RECT 129.560 52.310 131.170 52.590 ;
        RECT 131.410 52.760 133.930 53.040 ;
        RECT 134.610 53.160 136.690 53.440 ;
        RECT 138.110 53.710 139.450 53.990 ;
        RECT 127.410 52.000 127.690 52.310 ;
        RECT 129.560 52.000 129.840 52.310 ;
        RECT 131.410 52.005 131.690 52.760 ;
        RECT 134.610 52.590 134.890 53.160 ;
        RECT 138.110 52.990 138.390 53.710 ;
        RECT 141.930 53.490 142.210 54.200 ;
        RECT 122.030 35.945 122.780 51.210 ;
        RECT 124.705 50.025 125.455 51.260 ;
        RECT 126.930 51.210 127.690 52.000 ;
        RECT 124.705 49.275 126.480 50.025 ;
        RECT 123.530 36.100 124.930 40.280 ;
        RECT 125.730 36.825 126.480 49.275 ;
        RECT 126.930 36.220 127.680 51.210 ;
        RECT 129.080 51.160 129.840 52.000 ;
        RECT 130.930 51.260 131.690 52.005 ;
        RECT 133.160 52.310 134.890 52.590 ;
        RECT 135.210 52.710 138.390 52.990 ;
        RECT 138.910 53.210 142.210 53.490 ;
        RECT 133.160 52.000 133.440 52.310 ;
        RECT 135.210 52.005 135.490 52.710 ;
        RECT 138.910 52.490 139.190 53.210 ;
        RECT 144.690 52.990 144.970 54.200 ;
        RECT 137.210 52.210 139.190 52.490 ;
        RECT 139.710 52.710 144.970 52.990 ;
        RECT 137.210 52.025 137.490 52.210 ;
        RECT 132.730 51.975 134.055 52.000 ;
        RECT 129.080 40.375 129.830 51.160 ;
        RECT 130.930 41.875 131.680 51.260 ;
        RECT 132.725 51.225 134.055 51.975 ;
        RECT 133.305 43.425 134.055 51.225 ;
        RECT 134.805 45.125 135.555 52.005 ;
        RECT 136.725 51.275 138.140 52.025 ;
        RECT 134.805 44.375 136.880 45.125 ;
        RECT 133.305 42.675 135.905 43.425 ;
        RECT 130.930 41.125 134.855 41.875 ;
        RECT 129.080 39.625 131.980 40.375 ;
        RECT 123.530 35.000 126.710 36.100 ;
        RECT 126.930 35.580 130.680 36.220 ;
        RECT 131.205 36.175 131.955 39.625 ;
        RECT 126.930 35.575 127.680 35.580 ;
        RECT 131.205 35.520 133.835 36.175 ;
        RECT 131.205 35.475 131.955 35.520 ;
        RECT 120.065 34.015 121.310 34.825 ;
        RECT 105.670 12.000 107.230 13.500 ;
        RECT 111.380 13.100 119.910 15.100 ;
        RECT 105.700 11.050 107.200 12.000 ;
        RECT 92.185 10.010 105.210 10.760 ;
        RECT 92.215 9.625 92.965 10.010 ;
        RECT 103.125 9.625 103.875 10.010 ;
        RECT 92.215 8.875 103.905 9.625 ;
        RECT 111.380 9.290 113.380 13.100 ;
        RECT 120.500 9.575 121.310 34.015 ;
        RECT 123.530 32.700 124.930 35.000 ;
        RECT 134.105 33.275 134.855 41.125 ;
        RECT 123.530 31.600 131.360 32.700 ;
        RECT 132.005 32.025 134.855 33.275 ;
        RECT 123.530 9.300 124.930 31.600 ;
        RECT 128.700 27.700 130.100 31.600 ;
        RECT 133.105 30.525 133.755 30.555 ;
        RECT 135.155 30.525 135.905 42.675 ;
        RECT 132.055 29.775 135.905 30.525 ;
        RECT 132.055 28.925 133.880 29.775 ;
        RECT 132.055 28.190 133.830 28.925 ;
        RECT 128.700 26.950 132.805 27.700 ;
        RECT 128.700 24.120 130.100 26.950 ;
        RECT 136.130 26.500 136.880 44.375 ;
        RECT 132.135 25.750 136.880 26.500 ;
        RECT 132.135 25.735 134.915 25.750 ;
        RECT 132.135 25.365 133.025 25.735 ;
        RECT 134.165 25.365 134.915 25.735 ;
        RECT 136.130 25.725 136.880 25.750 ;
        RECT 132.135 24.615 134.915 25.365 ;
        RECT 132.275 24.605 133.025 24.615 ;
        RECT 128.700 23.370 132.805 24.120 ;
        RECT 128.700 20.540 130.100 23.370 ;
        RECT 137.390 22.880 138.140 51.275 ;
        RECT 132.135 22.130 138.140 22.880 ;
        RECT 138.650 51.940 139.400 52.055 ;
        RECT 139.710 51.940 139.990 52.710 ;
        RECT 147.450 52.490 147.730 54.200 ;
        RECT 138.650 51.660 139.990 51.940 ;
        RECT 141.310 52.210 147.730 52.490 ;
        RECT 141.310 51.925 141.590 52.210 ;
        RECT 132.215 21.775 132.965 22.130 ;
        RECT 133.815 22.125 136.145 22.130 ;
        RECT 135.395 21.775 136.145 22.125 ;
        RECT 132.215 21.025 136.175 21.775 ;
        RECT 132.215 20.995 132.965 21.025 ;
        RECT 128.700 19.790 132.805 20.540 ;
        RECT 128.700 16.960 130.100 19.790 ;
        RECT 136.955 19.320 137.705 19.345 ;
        RECT 138.650 19.320 139.400 51.660 ;
        RECT 140.775 51.175 141.980 51.925 ;
        RECT 142.525 51.490 145.005 52.025 ;
        RECT 150.210 51.490 150.490 54.200 ;
        RECT 142.525 51.275 150.490 51.490 ;
        RECT 142.610 51.210 150.490 51.275 ;
        RECT 132.055 18.570 139.400 19.320 ;
        RECT 132.085 18.195 132.835 18.570 ;
        RECT 136.955 18.195 137.705 18.570 ;
        RECT 132.085 17.445 137.735 18.195 ;
        RECT 132.085 17.415 132.835 17.445 ;
        RECT 128.700 16.210 132.805 16.960 ;
        RECT 128.700 13.380 130.100 16.210 ;
        RECT 139.485 15.760 140.235 15.775 ;
        RECT 141.230 15.760 141.980 51.175 ;
        RECT 132.035 15.010 141.980 15.760 ;
        RECT 132.065 14.625 132.815 15.010 ;
        RECT 139.485 14.625 140.235 15.010 ;
        RECT 132.065 13.875 140.265 14.625 ;
        RECT 132.065 13.845 132.815 13.875 ;
        RECT 128.700 12.630 132.805 13.380 ;
        RECT 128.700 9.300 130.100 12.630 ;
        RECT 143.005 12.160 143.755 12.185 ;
        RECT 144.255 12.160 145.005 51.210 ;
        RECT 145.650 43.250 147.150 45.780 ;
        RECT 145.620 41.750 147.180 43.250 ;
        RECT 145.650 26.300 147.150 41.750 ;
        RECT 145.620 24.800 147.180 26.300 ;
        RECT 145.650 13.450 147.150 24.800 ;
        RECT 132.065 11.410 145.090 12.160 ;
        RECT 145.620 11.950 147.180 13.450 ;
        RECT 132.095 11.025 132.845 11.410 ;
        RECT 143.005 11.025 143.755 11.410 ;
        RECT 132.095 10.275 143.785 11.025 ;
        RECT 145.650 11.000 147.150 11.950 ;
        RECT 132.095 10.245 132.845 10.275 ;
        RECT 123.530 9.290 130.100 9.300 ;
        RECT 142.830 9.290 144.230 9.880 ;
        RECT 92.215 8.845 92.965 8.875 ;
        RECT 83.650 7.890 90.220 7.900 ;
        RECT 102.950 7.890 104.350 8.480 ;
        RECT 42.430 7.050 49.000 7.060 ;
        RECT 61.730 7.050 63.130 7.640 ;
        RECT 30.280 5.050 63.180 7.050 ;
        RECT 71.500 5.890 104.400 7.890 ;
        RECT 111.380 7.290 144.280 9.290 ;
        RECT 127.830 6.595 129.870 6.615 ;
        RECT 87.465 5.515 89.740 5.535 ;
        RECT 44.415 4.505 46.585 4.525 ;
        RECT 41.610 2.285 46.610 4.505 ;
        RECT 84.360 3.190 89.765 5.515 ;
        RECT 124.125 4.505 129.895 6.595 ;
        RECT 127.830 4.485 129.870 4.505 ;
        RECT 87.465 3.170 89.740 3.190 ;
        RECT 44.415 2.265 46.585 2.285 ;
      LAYER met3 ;
        RECT 81.230 223.890 81.610 224.210 ;
        RECT 84.910 223.890 85.290 224.210 ;
        RECT 88.590 223.890 88.970 224.210 ;
        RECT 78.435 220.900 78.765 220.915 ;
        RECT 79.190 220.900 79.510 220.940 ;
        RECT 78.435 220.600 79.510 220.900 ;
        RECT 78.435 220.585 78.765 220.600 ;
        RECT 79.190 220.560 79.510 220.600 ;
        RECT 26.935 217.950 27.265 217.965 ;
        RECT 81.270 217.950 81.570 223.890 ;
        RECT 26.935 217.650 81.570 217.950 ;
        RECT 26.935 217.635 27.265 217.650 ;
        RECT 34.285 217.250 34.615 217.265 ;
        RECT 84.950 217.250 85.250 223.890 ;
        RECT 85.785 220.200 86.115 220.215 ;
        RECT 86.590 220.200 86.910 220.240 ;
        RECT 85.785 219.900 86.910 220.200 ;
        RECT 85.785 219.885 86.115 219.900 ;
        RECT 86.590 219.860 86.910 219.900 ;
        RECT 34.285 216.950 85.250 217.250 ;
        RECT 34.285 216.935 34.615 216.950 ;
        RECT 41.635 216.550 41.965 216.565 ;
        RECT 88.630 216.550 88.930 223.890 ;
        RECT 93.135 219.550 93.465 219.565 ;
        RECT 94.040 219.550 94.360 219.590 ;
        RECT 93.135 219.250 94.360 219.550 ;
        RECT 93.135 219.235 93.465 219.250 ;
        RECT 94.040 219.210 94.360 219.250 ;
        RECT 100.535 218.850 100.865 218.865 ;
        RECT 101.490 218.850 101.810 218.890 ;
        RECT 100.535 218.550 101.810 218.850 ;
        RECT 100.535 218.535 100.865 218.550 ;
        RECT 101.490 218.510 101.810 218.550 ;
        RECT 107.885 218.150 108.215 218.165 ;
        RECT 108.690 218.150 109.010 218.190 ;
        RECT 107.885 217.850 109.010 218.150 ;
        RECT 107.885 217.835 108.215 217.850 ;
        RECT 108.690 217.810 109.010 217.850 ;
        RECT 115.235 217.400 115.565 217.415 ;
        RECT 116.040 217.400 116.360 217.440 ;
        RECT 115.235 217.100 116.360 217.400 ;
        RECT 115.235 217.085 115.565 217.100 ;
        RECT 116.040 217.060 116.360 217.100 ;
        RECT 41.635 216.250 88.930 216.550 ;
        RECT 122.585 216.750 122.915 216.765 ;
        RECT 123.390 216.750 123.710 216.790 ;
        RECT 122.585 216.450 123.710 216.750 ;
        RECT 122.585 216.435 122.915 216.450 ;
        RECT 123.390 216.410 123.710 216.450 ;
        RECT 41.635 216.235 41.965 216.250 ;
        RECT 129.935 216.100 130.265 216.115 ;
        RECT 130.840 216.100 131.160 216.140 ;
        RECT 48.960 215.540 49.340 215.860 ;
        RECT 49.000 214.915 49.300 215.540 ;
        RECT 56.340 215.510 56.660 215.890 ;
        RECT 63.690 215.510 64.010 215.890 ;
        RECT 129.935 215.800 131.160 216.100 ;
        RECT 129.935 215.785 130.265 215.800 ;
        RECT 130.840 215.760 131.160 215.800 ;
        RECT 56.350 214.915 56.650 215.510 ;
        RECT 63.700 214.965 64.000 215.510 ;
        RECT 137.275 215.460 137.605 215.475 ;
        RECT 138.560 215.460 138.880 215.500 ;
        RECT 137.275 215.160 138.880 215.460 ;
        RECT 137.275 215.145 137.605 215.160 ;
        RECT 138.560 215.120 138.880 215.160 ;
        RECT 48.985 214.585 49.315 214.915 ;
        RECT 56.335 214.585 56.665 214.915 ;
        RECT 63.685 214.635 64.015 214.965 ;
        RECT 71.050 214.915 71.350 214.950 ;
        RECT 71.035 214.900 71.365 214.915 ;
        RECT 71.940 214.900 72.260 214.940 ;
        RECT 71.035 214.600 72.260 214.900 ;
        RECT 71.035 214.585 71.365 214.600 ;
        RECT 71.940 214.560 72.260 214.600 ;
        RECT 144.665 214.790 144.995 214.805 ;
        RECT 145.870 214.790 146.190 214.830 ;
        RECT 144.665 214.490 146.190 214.790 ;
        RECT 144.665 214.475 144.995 214.490 ;
        RECT 145.870 214.450 146.190 214.490 ;
        RECT 152.545 214.140 152.875 214.155 ;
        RECT 153.500 214.140 153.820 214.180 ;
        RECT 152.545 213.840 153.820 214.140 ;
        RECT 152.545 213.825 152.875 213.840 ;
        RECT 153.500 213.800 153.820 213.840 ;
        RECT 55.480 209.075 57.060 209.405 ;
        RECT 89.060 209.075 90.640 209.405 ;
        RECT 122.640 209.075 124.220 209.405 ;
        RECT 156.220 209.075 157.800 209.405 ;
        RECT 38.690 206.355 40.270 206.685 ;
        RECT 72.270 206.355 73.850 206.685 ;
        RECT 105.850 206.355 107.430 206.685 ;
        RECT 139.430 206.355 141.010 206.685 ;
        RECT 30.115 206.340 30.445 206.345 ;
        RECT 30.115 206.330 30.700 206.340 ;
        RECT 30.115 206.030 30.900 206.330 ;
        RECT 30.115 206.020 30.700 206.030 ;
        RECT 30.115 206.015 30.445 206.020 ;
        RECT 123.955 204.970 124.285 204.985 ;
        RECT 139.135 204.970 139.465 204.985 ;
        RECT 123.955 204.670 139.465 204.970 ;
        RECT 123.955 204.655 124.285 204.670 ;
        RECT 139.135 204.655 139.465 204.670 ;
        RECT 55.480 203.635 57.060 203.965 ;
        RECT 89.060 203.635 90.640 203.965 ;
        RECT 122.640 203.635 124.220 203.965 ;
        RECT 156.220 203.635 157.800 203.965 ;
        RECT 29.195 202.940 29.525 202.945 ;
        RECT 29.195 202.930 29.780 202.940 ;
        RECT 134.075 202.930 134.405 202.945 ;
        RECT 146.035 202.930 146.365 202.945 ;
        RECT 29.195 202.630 29.980 202.930 ;
        RECT 134.075 202.630 146.365 202.930 ;
        RECT 29.195 202.620 29.780 202.630 ;
        RECT 29.195 202.615 29.525 202.620 ;
        RECT 134.075 202.615 134.405 202.630 ;
        RECT 146.035 202.615 146.365 202.630 ;
        RECT 79.795 202.250 80.125 202.265 ;
        RECT 102.795 202.250 103.125 202.265 ;
        RECT 114.755 202.250 115.085 202.265 ;
        RECT 79.795 201.950 115.085 202.250 ;
        RECT 79.795 201.935 80.125 201.950 ;
        RECT 102.795 201.935 103.125 201.950 ;
        RECT 114.755 201.935 115.085 201.950 ;
        RECT 134.535 202.250 134.865 202.265 ;
        RECT 139.135 202.250 139.465 202.265 ;
        RECT 148.335 202.250 148.665 202.265 ;
        RECT 134.535 201.950 148.665 202.250 ;
        RECT 134.535 201.935 134.865 201.950 ;
        RECT 139.135 201.935 139.465 201.950 ;
        RECT 148.335 201.935 148.665 201.950 ;
        RECT 52.195 201.570 52.525 201.585 ;
        RECT 58.635 201.570 58.965 201.585 ;
        RECT 52.195 201.270 58.965 201.570 ;
        RECT 52.195 201.255 52.525 201.270 ;
        RECT 58.635 201.255 58.965 201.270 ;
        RECT 38.690 200.915 40.270 201.245 ;
        RECT 72.270 200.915 73.850 201.245 ;
        RECT 105.850 200.915 107.430 201.245 ;
        RECT 139.430 200.915 141.010 201.245 ;
        RECT 40.695 199.530 41.025 199.545 ;
        RECT 42.995 199.530 43.325 199.545 ;
        RECT 40.695 199.230 43.325 199.530 ;
        RECT 40.695 199.215 41.025 199.230 ;
        RECT 42.995 199.215 43.325 199.230 ;
        RECT 55.480 198.195 57.060 198.525 ;
        RECT 89.060 198.195 90.640 198.525 ;
        RECT 122.640 198.195 124.220 198.525 ;
        RECT 156.220 198.195 157.800 198.525 ;
        RECT 38.690 195.475 40.270 195.805 ;
        RECT 72.270 195.475 73.850 195.805 ;
        RECT 105.850 195.475 107.430 195.805 ;
        RECT 139.430 195.475 141.010 195.805 ;
        RECT 103.255 193.410 103.585 193.425 ;
        RECT 106.015 193.410 106.345 193.425 ;
        RECT 103.255 193.110 106.345 193.410 ;
        RECT 103.255 193.095 103.585 193.110 ;
        RECT 106.015 193.095 106.345 193.110 ;
        RECT 55.480 192.755 57.060 193.085 ;
        RECT 89.060 192.755 90.640 193.085 ;
        RECT 122.640 192.755 124.220 193.085 ;
        RECT 156.220 192.755 157.800 193.085 ;
        RECT 106.015 192.730 106.345 192.745 ;
        RECT 107.855 192.730 108.185 192.745 ;
        RECT 144.655 192.740 144.985 192.745 ;
        RECT 144.400 192.730 144.985 192.740 ;
        RECT 106.015 192.430 108.185 192.730 ;
        RECT 144.200 192.430 144.985 192.730 ;
        RECT 106.015 192.415 106.345 192.430 ;
        RECT 107.855 192.415 108.185 192.430 ;
        RECT 144.400 192.420 144.985 192.430 ;
        RECT 144.655 192.415 144.985 192.420 ;
        RECT 38.690 190.035 40.270 190.365 ;
        RECT 72.270 190.035 73.850 190.365 ;
        RECT 105.850 190.035 107.430 190.365 ;
        RECT 139.430 190.035 141.010 190.365 ;
        RECT 126.255 189.330 126.585 189.345 ;
        RECT 137.295 189.330 137.625 189.345 ;
        RECT 126.255 189.030 137.625 189.330 ;
        RECT 126.255 189.015 126.585 189.030 ;
        RECT 137.295 189.015 137.625 189.030 ;
        RECT 55.480 187.315 57.060 187.645 ;
        RECT 89.060 187.315 90.640 187.645 ;
        RECT 122.640 187.315 124.220 187.645 ;
        RECT 156.220 187.315 157.800 187.645 ;
        RECT 127.635 187.290 127.965 187.305 ;
        RECT 129.015 187.290 129.345 187.305 ;
        RECT 127.635 186.990 129.345 187.290 ;
        RECT 127.635 186.975 127.965 186.990 ;
        RECT 129.015 186.975 129.345 186.990 ;
        RECT 38.690 184.595 40.270 184.925 ;
        RECT 72.270 184.595 73.850 184.925 ;
        RECT 105.850 184.595 107.430 184.925 ;
        RECT 139.430 184.595 141.010 184.925 ;
        RECT 55.480 181.875 57.060 182.205 ;
        RECT 89.060 181.875 90.640 182.205 ;
        RECT 122.640 181.875 124.220 182.205 ;
        RECT 156.220 181.875 157.800 182.205 ;
        RECT 38.690 179.155 40.270 179.485 ;
        RECT 72.270 179.155 73.850 179.485 ;
        RECT 105.850 179.155 107.430 179.485 ;
        RECT 139.430 179.155 141.010 179.485 ;
        RECT 51.735 178.450 52.065 178.465 ;
        RECT 60.475 178.450 60.805 178.465 ;
        RECT 97.735 178.450 98.065 178.465 ;
        RECT 51.735 178.150 98.065 178.450 ;
        RECT 51.735 178.135 52.065 178.150 ;
        RECT 60.475 178.135 60.805 178.150 ;
        RECT 97.735 178.135 98.065 178.150 ;
        RECT 51.735 177.770 52.065 177.785 ;
        RECT 58.175 177.770 58.505 177.785 ;
        RECT 51.735 177.470 58.505 177.770 ;
        RECT 51.735 177.455 52.065 177.470 ;
        RECT 58.175 177.455 58.505 177.470 ;
        RECT 55.480 176.435 57.060 176.765 ;
        RECT 89.060 176.435 90.640 176.765 ;
        RECT 122.640 176.435 124.220 176.765 ;
        RECT 156.220 176.435 157.800 176.765 ;
        RECT 51.735 175.730 52.065 175.745 ;
        RECT 59.555 175.730 59.885 175.745 ;
        RECT 51.735 175.430 59.885 175.730 ;
        RECT 51.735 175.415 52.065 175.430 ;
        RECT 59.555 175.415 59.885 175.430 ;
        RECT 54.495 174.370 54.825 174.385 ;
        RECT 59.095 174.370 59.425 174.385 ;
        RECT 54.495 174.070 59.425 174.370 ;
        RECT 54.495 174.055 54.825 174.070 ;
        RECT 59.095 174.055 59.425 174.070 ;
        RECT 38.690 173.715 40.270 174.045 ;
        RECT 72.270 173.715 73.850 174.045 ;
        RECT 105.850 173.715 107.430 174.045 ;
        RECT 139.430 173.715 141.010 174.045 ;
        RECT 55.480 170.995 57.060 171.325 ;
        RECT 89.060 170.995 90.640 171.325 ;
        RECT 122.640 170.995 124.220 171.325 ;
        RECT 156.220 170.995 157.800 171.325 ;
        RECT 38.690 168.275 40.270 168.605 ;
        RECT 72.270 168.275 73.850 168.605 ;
        RECT 105.850 168.275 107.430 168.605 ;
        RECT 139.430 168.275 141.010 168.605 ;
        RECT 55.480 165.555 57.060 165.885 ;
        RECT 89.060 165.555 90.640 165.885 ;
        RECT 122.640 165.555 124.220 165.885 ;
        RECT 156.220 165.555 157.800 165.885 ;
        RECT 74.735 164.170 75.065 164.185 ;
        RECT 110.155 164.170 110.485 164.185 ;
        RECT 74.735 163.870 110.485 164.170 ;
        RECT 74.735 163.855 75.065 163.870 ;
        RECT 110.155 163.855 110.485 163.870 ;
        RECT 38.690 162.835 40.270 163.165 ;
        RECT 72.270 162.835 73.850 163.165 ;
        RECT 105.850 162.835 107.430 163.165 ;
        RECT 139.430 162.835 141.010 163.165 ;
        RECT 55.480 160.115 57.060 160.445 ;
        RECT 89.060 160.115 90.640 160.445 ;
        RECT 122.640 160.115 124.220 160.445 ;
        RECT 156.220 160.115 157.800 160.445 ;
        RECT 38.690 157.395 40.270 157.725 ;
        RECT 72.270 157.395 73.850 157.725 ;
        RECT 105.850 157.395 107.430 157.725 ;
        RECT 139.430 157.395 141.010 157.725 ;
        RECT 55.480 154.675 57.060 155.005 ;
        RECT 89.060 154.675 90.640 155.005 ;
        RECT 122.640 154.675 124.220 155.005 ;
        RECT 156.220 154.675 157.800 155.005 ;
        RECT 84.855 153.290 85.185 153.305 ;
        RECT 112.455 153.290 112.785 153.305 ;
        RECT 84.855 152.990 112.785 153.290 ;
        RECT 84.855 152.975 85.185 152.990 ;
        RECT 112.455 152.975 112.785 152.990 ;
        RECT 38.690 151.955 40.270 152.285 ;
        RECT 72.270 151.955 73.850 152.285 ;
        RECT 105.850 151.955 107.430 152.285 ;
        RECT 139.430 151.955 141.010 152.285 ;
        RECT 94.515 151.250 94.845 151.265 ;
        RECT 111.535 151.250 111.865 151.265 ;
        RECT 94.515 150.950 111.865 151.250 ;
        RECT 94.515 150.935 94.845 150.950 ;
        RECT 111.535 150.935 111.865 150.950 ;
        RECT 55.480 149.235 57.060 149.565 ;
        RECT 89.060 149.235 90.640 149.565 ;
        RECT 122.640 149.235 124.220 149.565 ;
        RECT 156.220 149.235 157.800 149.565 ;
        RECT 38.690 146.515 40.270 146.845 ;
        RECT 72.270 146.515 73.850 146.845 ;
        RECT 105.850 146.515 107.430 146.845 ;
        RECT 139.430 146.515 141.010 146.845 ;
        RECT 55.480 143.795 57.060 144.125 ;
        RECT 89.060 143.795 90.640 144.125 ;
        RECT 122.640 143.795 124.220 144.125 ;
        RECT 156.220 143.795 157.800 144.125 ;
        RECT 38.690 141.075 40.270 141.405 ;
        RECT 72.270 141.075 73.850 141.405 ;
        RECT 105.850 141.075 107.430 141.405 ;
        RECT 139.430 141.075 141.010 141.405 ;
        RECT 62.315 140.370 62.645 140.385 ;
        RECT 72.435 140.370 72.765 140.385 ;
        RECT 62.315 140.070 72.765 140.370 ;
        RECT 62.315 140.055 62.645 140.070 ;
        RECT 72.435 140.055 72.765 140.070 ;
        RECT 139.595 140.370 139.925 140.385 ;
        RECT 144.655 140.370 144.985 140.385 ;
        RECT 139.595 140.070 144.985 140.370 ;
        RECT 139.595 140.055 139.925 140.070 ;
        RECT 144.655 140.055 144.985 140.070 ;
        RECT 100.495 139.690 100.825 139.705 ;
        RECT 144.400 139.690 144.780 139.700 ;
        RECT 100.495 139.390 144.780 139.690 ;
        RECT 100.495 139.375 100.825 139.390 ;
        RECT 144.400 139.380 144.780 139.390 ;
        RECT 140.975 139.010 141.305 139.025 ;
        RECT 143.275 139.010 143.605 139.025 ;
        RECT 140.975 138.710 143.605 139.010 ;
        RECT 140.975 138.695 141.305 138.710 ;
        RECT 143.275 138.695 143.605 138.710 ;
        RECT 55.480 138.355 57.060 138.685 ;
        RECT 89.060 138.355 90.640 138.685 ;
        RECT 122.640 138.355 124.220 138.685 ;
        RECT 156.220 138.355 157.800 138.685 ;
        RECT 38.690 135.635 40.270 135.965 ;
        RECT 72.270 135.635 73.850 135.965 ;
        RECT 105.850 135.635 107.430 135.965 ;
        RECT 139.430 135.635 141.010 135.965 ;
        RECT 73.355 134.250 73.685 134.265 ;
        RECT 93.135 134.250 93.465 134.265 ;
        RECT 97.275 134.250 97.605 134.265 ;
        RECT 73.355 133.950 97.605 134.250 ;
        RECT 73.355 133.935 73.685 133.950 ;
        RECT 93.135 133.935 93.465 133.950 ;
        RECT 97.275 133.935 97.605 133.950 ;
        RECT 55.480 132.915 57.060 133.245 ;
        RECT 89.060 132.915 90.640 133.245 ;
        RECT 122.640 132.915 124.220 133.245 ;
        RECT 156.220 132.915 157.800 133.245 ;
        RECT 38.690 130.195 40.270 130.525 ;
        RECT 72.270 130.195 73.850 130.525 ;
        RECT 105.850 130.195 107.430 130.525 ;
        RECT 139.430 130.195 141.010 130.525 ;
        RECT 55.480 127.475 57.060 127.805 ;
        RECT 89.060 127.475 90.640 127.805 ;
        RECT 122.640 127.475 124.220 127.805 ;
        RECT 156.220 127.475 157.800 127.805 ;
        RECT 69.215 126.090 69.545 126.105 ;
        RECT 71.055 126.090 71.385 126.105 ;
        RECT 83.475 126.090 83.805 126.105 ;
        RECT 111.535 126.090 111.865 126.105 ;
        RECT 69.215 125.790 111.865 126.090 ;
        RECT 69.215 125.775 69.545 125.790 ;
        RECT 71.055 125.775 71.385 125.790 ;
        RECT 83.475 125.775 83.805 125.790 ;
        RECT 111.535 125.775 111.865 125.790 ;
        RECT 38.690 124.755 40.270 125.085 ;
        RECT 72.270 124.755 73.850 125.085 ;
        RECT 105.850 124.755 107.430 125.085 ;
        RECT 139.430 124.755 141.010 125.085 ;
        RECT 55.480 122.035 57.060 122.365 ;
        RECT 89.060 122.035 90.640 122.365 ;
        RECT 122.640 122.035 124.220 122.365 ;
        RECT 156.220 122.035 157.800 122.365 ;
        RECT 38.690 119.315 40.270 119.645 ;
        RECT 72.270 119.315 73.850 119.645 ;
        RECT 105.850 119.315 107.430 119.645 ;
        RECT 139.430 119.315 141.010 119.645 ;
        RECT 55.480 116.595 57.060 116.925 ;
        RECT 89.060 116.595 90.640 116.925 ;
        RECT 122.640 116.595 124.220 116.925 ;
        RECT 156.220 116.595 157.800 116.925 ;
        RECT 38.690 113.875 40.270 114.205 ;
        RECT 72.270 113.875 73.850 114.205 ;
        RECT 105.850 113.875 107.430 114.205 ;
        RECT 139.430 113.875 141.010 114.205 ;
        RECT 55.480 111.155 57.060 111.485 ;
        RECT 89.060 111.155 90.640 111.485 ;
        RECT 122.640 111.155 124.220 111.485 ;
        RECT 156.220 111.155 157.800 111.485 ;
        RECT 38.690 108.435 40.270 108.765 ;
        RECT 72.270 108.435 73.850 108.765 ;
        RECT 105.850 108.435 107.430 108.765 ;
        RECT 139.430 108.435 141.010 108.765 ;
        RECT 30.320 107.050 30.700 107.060 ;
        RECT 121.655 107.050 121.985 107.065 ;
        RECT 30.320 106.750 121.985 107.050 ;
        RECT 30.320 106.740 30.700 106.750 ;
        RECT 121.655 106.735 121.985 106.750 ;
        RECT 55.480 105.715 57.060 106.045 ;
        RECT 89.060 105.715 90.640 106.045 ;
        RECT 122.640 105.715 124.220 106.045 ;
        RECT 156.220 105.715 157.800 106.045 ;
        RECT 38.690 102.995 40.270 103.325 ;
        RECT 72.270 102.995 73.850 103.325 ;
        RECT 105.850 102.995 107.430 103.325 ;
        RECT 139.430 102.995 141.010 103.325 ;
        RECT 55.480 100.275 57.060 100.605 ;
        RECT 89.060 100.275 90.640 100.605 ;
        RECT 122.640 100.275 124.220 100.605 ;
        RECT 156.220 100.275 157.800 100.605 ;
        RECT 38.690 97.555 40.270 97.885 ;
        RECT 72.270 97.555 73.850 97.885 ;
        RECT 105.850 97.555 107.430 97.885 ;
        RECT 139.430 97.555 141.010 97.885 ;
        RECT 55.480 94.835 57.060 95.165 ;
        RECT 89.060 94.835 90.640 95.165 ;
        RECT 122.640 94.835 124.220 95.165 ;
        RECT 156.220 94.835 157.800 95.165 ;
        RECT 38.690 92.115 40.270 92.445 ;
        RECT 72.270 92.115 73.850 92.445 ;
        RECT 105.850 92.115 107.430 92.445 ;
        RECT 139.430 92.115 141.010 92.445 ;
        RECT 29.400 90.730 29.780 90.740 ;
        RECT 69.215 90.730 69.545 90.745 ;
        RECT 29.400 90.430 69.545 90.730 ;
        RECT 29.400 90.420 29.780 90.430 ;
        RECT 69.215 90.415 69.545 90.430 ;
        RECT 79.335 90.050 79.665 90.065 ;
        RECT 84.855 90.050 85.185 90.065 ;
        RECT 79.335 89.750 85.185 90.050 ;
        RECT 79.335 89.735 79.665 89.750 ;
        RECT 84.855 89.735 85.185 89.750 ;
        RECT 55.480 89.395 57.060 89.725 ;
        RECT 89.060 89.395 90.640 89.725 ;
        RECT 122.640 89.395 124.220 89.725 ;
        RECT 156.220 89.395 157.800 89.725 ;
        RECT 38.690 86.675 40.270 87.005 ;
        RECT 72.270 86.675 73.850 87.005 ;
        RECT 105.850 86.675 107.430 87.005 ;
        RECT 139.430 86.675 141.010 87.005 ;
        RECT 91.755 86.650 92.085 86.665 ;
        RECT 95.895 86.650 96.225 86.665 ;
        RECT 91.755 86.350 96.225 86.650 ;
        RECT 91.755 86.335 92.085 86.350 ;
        RECT 95.895 86.335 96.225 86.350 ;
        RECT 90.375 85.290 90.705 85.305 ;
        RECT 95.435 85.290 95.765 85.305 ;
        RECT 90.375 84.990 95.765 85.290 ;
        RECT 90.375 84.975 90.705 84.990 ;
        RECT 95.435 84.975 95.765 84.990 ;
        RECT 55.480 83.955 57.060 84.285 ;
        RECT 89.060 83.955 90.640 84.285 ;
        RECT 122.640 83.955 124.220 84.285 ;
        RECT 156.220 83.955 157.800 84.285 ;
        RECT 38.690 81.235 40.270 81.565 ;
        RECT 72.270 81.235 73.850 81.565 ;
        RECT 105.850 81.235 107.430 81.565 ;
        RECT 139.430 81.235 141.010 81.565 ;
        RECT 55.480 78.515 57.060 78.845 ;
        RECT 89.060 78.515 90.640 78.845 ;
        RECT 122.640 78.515 124.220 78.845 ;
        RECT 156.220 78.515 157.800 78.845 ;
        RECT 38.690 75.795 40.270 76.125 ;
        RECT 72.270 75.795 73.850 76.125 ;
        RECT 105.850 75.795 107.430 76.125 ;
        RECT 139.430 75.795 141.010 76.125 ;
        RECT 34.715 74.410 35.045 74.425 ;
        RECT 37.935 74.410 38.265 74.425 ;
        RECT 58.175 74.410 58.505 74.425 ;
        RECT 91.755 74.410 92.085 74.425 ;
        RECT 34.715 74.110 92.085 74.410 ;
        RECT 34.715 74.095 35.045 74.110 ;
        RECT 37.935 74.095 38.265 74.110 ;
        RECT 58.175 74.095 58.505 74.110 ;
        RECT 91.755 74.095 92.085 74.110 ;
        RECT 55.480 73.075 57.060 73.405 ;
        RECT 89.060 73.075 90.640 73.405 ;
        RECT 122.640 73.075 124.220 73.405 ;
        RECT 156.220 73.075 157.800 73.405 ;
        RECT 73.815 72.370 74.145 72.385 ;
        RECT 98.655 72.370 98.985 72.385 ;
        RECT 73.815 72.070 98.985 72.370 ;
        RECT 73.815 72.055 74.145 72.070 ;
        RECT 98.655 72.055 98.985 72.070 ;
        RECT 44.835 71.690 45.165 71.705 ;
        RECT 55.875 71.690 56.205 71.705 ;
        RECT 93.135 71.690 93.465 71.705 ;
        RECT 44.835 71.390 93.465 71.690 ;
        RECT 44.835 71.375 45.165 71.390 ;
        RECT 55.875 71.375 56.205 71.390 ;
        RECT 93.135 71.375 93.465 71.390 ;
        RECT 88.995 71.010 89.325 71.025 ;
        RECT 94.515 71.010 94.845 71.025 ;
        RECT 88.995 70.710 94.845 71.010 ;
        RECT 88.995 70.695 89.325 70.710 ;
        RECT 94.515 70.695 94.845 70.710 ;
        RECT 38.690 70.355 40.270 70.685 ;
        RECT 72.270 70.355 73.850 70.685 ;
        RECT 105.850 70.355 107.430 70.685 ;
        RECT 139.430 70.355 141.010 70.685 ;
        RECT 55.480 67.635 57.060 67.965 ;
        RECT 89.060 67.635 90.640 67.965 ;
        RECT 122.640 67.635 124.220 67.965 ;
        RECT 156.220 67.635 157.800 67.965 ;
        RECT 42.075 66.930 42.405 66.945 ;
        RECT 47.135 66.930 47.465 66.945 ;
        RECT 52.195 66.930 52.525 66.945 ;
        RECT 42.075 66.630 52.525 66.930 ;
        RECT 42.075 66.615 42.405 66.630 ;
        RECT 47.135 66.615 47.465 66.630 ;
        RECT 52.195 66.615 52.525 66.630 ;
        RECT 38.690 64.915 40.270 65.245 ;
        RECT 72.270 64.915 73.850 65.245 ;
        RECT 105.850 64.915 107.430 65.245 ;
        RECT 139.430 64.915 141.010 65.245 ;
        RECT 55.480 62.195 57.060 62.525 ;
        RECT 89.060 62.195 90.640 62.525 ;
        RECT 122.640 62.195 124.220 62.525 ;
        RECT 156.220 62.195 157.800 62.525 ;
        RECT 38.690 59.475 40.270 59.805 ;
        RECT 72.270 59.475 73.850 59.805 ;
        RECT 105.850 59.475 107.430 59.805 ;
        RECT 139.430 59.475 141.010 59.805 ;
        RECT 55.480 56.755 57.060 57.085 ;
        RECT 89.060 56.755 90.640 57.085 ;
        RECT 122.640 56.755 124.220 57.085 ;
        RECT 156.220 56.755 157.800 57.085 ;
        RECT 26.955 46.400 28.445 46.425 ;
        RECT 26.950 44.900 32.100 46.400 ;
        RECT 26.955 44.875 28.445 44.900 ;
        RECT 5.005 40.400 6.495 40.425 ;
        RECT 38.750 40.400 40.250 54.010 ;
        RECT 72.280 52.410 77.970 53.910 ;
        RECT 68.300 47.095 73.350 47.100 ;
        RECT 68.275 45.605 73.350 47.095 ;
        RECT 68.300 45.600 73.350 45.605 ;
        RECT 76.470 40.400 77.970 52.410 ;
        RECT 105.980 40.450 107.480 53.940 ;
        RECT 109.155 48.650 110.645 48.675 ;
        RECT 109.150 47.150 113.100 48.650 ;
        RECT 109.155 47.125 110.645 47.150 ;
        RECT 105.550 40.400 107.550 40.450 ;
        RECT 139.480 40.400 140.980 53.940 ;
        RECT 5.000 38.900 147.400 40.400 ;
        RECT 5.005 38.875 6.495 38.900 ;
        RECT 127.805 6.305 133.445 6.595 ;
        RECT 149.450 6.305 150.950 6.330 ;
        RECT 87.440 5.095 93.665 5.515 ;
        RECT 102.710 5.095 104.190 5.120 ;
        RECT 44.390 4.170 51.510 4.505 ;
        RECT 52.235 4.170 53.770 4.195 ;
        RECT 44.390 2.625 53.775 4.170 ;
        RECT 87.440 3.605 104.195 5.095 ;
        RECT 127.805 4.795 150.955 6.305 ;
        RECT 127.805 4.505 133.445 4.795 ;
        RECT 149.450 4.770 150.950 4.795 ;
        RECT 87.440 3.190 93.665 3.605 ;
        RECT 102.710 3.580 104.190 3.605 ;
        RECT 44.390 2.285 51.510 2.625 ;
        RECT 52.235 2.600 53.770 2.625 ;
      LAYER met4 ;
        RECT 3.990 224.500 4.290 224.760 ;
        RECT 3.950 224.000 4.350 224.500 ;
        RECT 7.670 224.000 7.970 224.760 ;
        RECT 11.350 224.000 11.650 224.760 ;
        RECT 15.030 224.000 15.330 224.760 ;
        RECT 18.710 224.000 19.010 224.760 ;
        RECT 22.390 224.000 22.690 224.760 ;
        RECT 26.070 224.000 26.370 224.760 ;
        RECT 29.750 224.000 30.050 224.760 ;
        RECT 33.430 224.000 33.730 224.760 ;
        RECT 37.110 224.000 37.410 224.760 ;
        RECT 40.790 224.000 41.090 224.760 ;
        RECT 44.470 224.000 44.770 224.760 ;
        RECT 48.150 224.000 48.450 224.760 ;
        RECT 51.830 224.000 52.130 224.760 ;
        RECT 55.510 224.000 55.810 224.760 ;
        RECT 59.190 224.000 59.490 224.760 ;
        RECT 62.870 224.000 63.170 224.760 ;
        RECT 66.550 224.000 66.850 224.760 ;
        RECT 70.230 224.000 70.530 224.760 ;
        RECT 73.910 224.000 74.210 224.760 ;
        RECT 77.590 224.000 77.890 224.760 ;
        RECT 81.270 224.215 81.570 224.760 ;
        RECT 84.950 224.215 85.250 224.760 ;
        RECT 88.630 224.215 88.930 224.760 ;
        RECT 92.310 224.300 92.610 224.760 ;
        RECT 95.990 224.300 96.290 224.760 ;
        RECT 99.670 224.300 99.970 224.760 ;
        RECT 103.350 224.300 103.650 224.760 ;
        RECT 3.950 223.700 77.890 224.000 ;
        RECT 81.255 223.885 81.585 224.215 ;
        RECT 84.935 223.885 85.265 224.215 ;
        RECT 88.615 223.885 88.945 224.215 ;
        RECT 3.950 223.600 74.200 223.700 ;
        RECT 7.650 222.500 74.200 223.600 ;
        RECT 107.030 223.400 107.330 224.760 ;
        RECT 75.150 223.100 107.330 223.400 ;
        RECT 9.000 220.760 10.500 222.500 ;
        RECT 75.150 219.200 75.450 223.100 ;
        RECT 110.710 222.800 111.010 224.760 ;
        RECT 49.000 218.900 75.450 219.200 ;
        RECT 75.950 222.500 111.010 222.800 ;
        RECT 49.000 215.865 49.300 218.900 ;
        RECT 75.950 218.550 76.250 222.500 ;
        RECT 114.390 222.200 114.690 224.760 ;
        RECT 56.350 218.250 76.250 218.550 ;
        RECT 76.750 221.900 114.690 222.200 ;
        RECT 56.350 215.865 56.650 218.250 ;
        RECT 63.700 215.865 64.000 215.900 ;
        RECT 48.985 215.535 49.315 215.865 ;
        RECT 56.335 215.535 56.665 215.865 ;
        RECT 63.685 215.850 64.015 215.865 ;
        RECT 70.250 215.850 70.550 215.900 ;
        RECT 76.750 215.850 77.050 221.900 ;
        RECT 118.070 221.550 118.370 224.760 ;
        RECT 77.600 221.250 118.370 221.550 ;
        RECT 77.600 215.850 77.900 221.250 ;
        RECT 79.185 220.900 79.515 220.915 ;
        RECT 121.750 220.900 122.050 224.760 ;
        RECT 79.185 220.600 122.050 220.900 ;
        RECT 79.185 220.585 79.515 220.600 ;
        RECT 86.585 220.200 86.915 220.215 ;
        RECT 125.430 220.200 125.730 224.760 ;
        RECT 86.585 219.900 125.730 220.200 ;
        RECT 86.585 219.885 86.915 219.900 ;
        RECT 94.035 219.550 94.365 219.565 ;
        RECT 129.110 219.550 129.410 224.760 ;
        RECT 94.035 219.250 129.410 219.550 ;
        RECT 94.035 219.235 94.365 219.250 ;
        RECT 101.485 218.850 101.815 218.865 ;
        RECT 132.790 218.850 133.090 224.760 ;
        RECT 101.485 218.550 133.090 218.850 ;
        RECT 101.485 218.535 101.815 218.550 ;
        RECT 108.685 218.150 109.015 218.165 ;
        RECT 136.470 218.150 136.770 224.760 ;
        RECT 108.685 217.850 136.770 218.150 ;
        RECT 108.685 217.835 109.015 217.850 ;
        RECT 116.035 217.400 116.365 217.415 ;
        RECT 140.150 217.400 140.450 224.760 ;
        RECT 116.035 217.100 140.450 217.400 ;
        RECT 116.035 217.085 116.365 217.100 ;
        RECT 123.385 216.750 123.715 216.765 ;
        RECT 143.830 216.750 144.130 224.760 ;
        RECT 123.385 216.450 144.130 216.750 ;
        RECT 123.385 216.435 123.715 216.450 ;
        RECT 63.685 215.550 77.050 215.850 ;
        RECT 77.550 215.550 77.900 215.850 ;
        RECT 130.835 216.100 131.165 216.115 ;
        RECT 147.510 216.100 147.810 224.760 ;
        RECT 130.835 215.800 147.810 216.100 ;
        RECT 130.835 215.785 131.165 215.800 ;
        RECT 63.685 215.535 64.015 215.550 ;
        RECT 71.935 214.900 72.265 214.915 ;
        RECT 77.600 214.900 77.900 215.550 ;
        RECT 138.555 215.460 138.885 215.475 ;
        RECT 151.190 215.460 151.490 224.760 ;
        RECT 138.555 215.160 151.490 215.460 ;
        RECT 138.555 215.145 138.885 215.160 ;
        RECT 71.935 214.600 77.900 214.900 ;
        RECT 145.865 214.790 146.195 214.805 ;
        RECT 154.870 214.790 155.170 224.760 ;
        RECT 71.935 214.585 72.265 214.600 ;
        RECT 145.865 214.490 155.170 214.790 ;
        RECT 145.865 214.475 146.195 214.490 ;
        RECT 153.495 214.140 153.825 214.155 ;
        RECT 158.550 214.140 158.850 224.760 ;
        RECT 153.495 213.840 158.850 214.140 ;
        RECT 153.495 213.825 153.825 213.840 ;
        RECT 38.750 209.480 40.250 209.500 ;
        RECT 89.130 209.480 90.630 209.500 ;
        RECT 139.480 209.480 140.980 209.530 ;
        RECT 30.345 206.015 30.675 206.345 ;
        RECT 29.425 202.615 29.755 202.945 ;
        RECT 29.440 90.745 29.740 202.615 ;
        RECT 30.360 107.065 30.660 206.015 ;
        RECT 30.345 106.735 30.675 107.065 ;
        RECT 29.425 90.415 29.755 90.745 ;
        RECT 38.680 56.680 40.280 209.480 ;
        RECT 55.470 56.680 57.070 209.480 ;
        RECT 72.260 56.680 73.860 209.480 ;
        RECT 89.050 56.680 90.650 209.480 ;
        RECT 105.840 209.250 107.440 209.480 ;
        RECT 122.630 209.470 124.230 209.480 ;
        RECT 105.840 56.680 107.480 209.250 ;
        RECT 122.630 56.680 124.270 209.470 ;
        RECT 139.420 56.680 141.020 209.480 ;
        RECT 144.425 192.415 144.755 192.745 ;
        RECT 144.440 139.705 144.740 192.415 ;
        RECT 144.425 139.375 144.755 139.705 ;
        RECT 156.210 56.680 157.810 209.480 ;
        RECT 38.750 53.985 40.250 56.680 ;
        RECT 38.745 52.475 40.255 53.985 ;
        RECT 55.490 48.650 56.990 56.680 ;
        RECT 72.310 53.915 73.810 56.680 ;
        RECT 72.305 52.405 73.815 53.915 ;
        RECT 89.130 48.650 90.630 56.680 ;
        RECT 105.980 53.915 107.480 56.680 ;
        RECT 105.975 52.405 107.485 53.915 ;
        RECT 122.770 48.650 124.270 56.680 ;
        RECT 139.480 53.915 140.980 56.680 ;
        RECT 139.475 52.405 140.985 53.915 ;
        RECT 156.250 48.650 157.750 56.680 ;
        RECT 10.500 47.150 157.750 48.650 ;
        RECT 26.950 44.900 28.450 47.150 ;
        RECT 68.300 45.600 69.800 47.150 ;
        RECT 2.500 38.900 6.500 40.400 ;
        RECT 149.445 6.300 157.300 6.305 ;
        RECT 108.150 5.095 109.850 5.100 ;
        RECT 60.880 4.170 64.470 4.175 ;
        RECT 52.230 2.625 64.470 4.170 ;
        RECT 102.705 3.900 109.850 5.095 ;
        RECT 149.445 4.795 157.310 6.300 ;
        RECT 102.705 3.605 135.230 3.900 ;
        RECT 108.100 3.000 135.230 3.605 ;
        RECT 62.925 2.280 64.470 2.625 ;
        RECT 62.925 1.430 113.150 2.280 ;
        RECT 63.200 1.380 113.150 1.430 ;
        RECT 112.250 1.000 113.150 1.380 ;
        RECT 134.330 1.000 135.230 3.000 ;
        RECT 156.410 1.000 157.310 4.795 ;
  END
END tt_um_rejunity_ay8913
END LIBRARY

