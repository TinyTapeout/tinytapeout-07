module tt_ctrl (ctrl_ena,
    ctrl_sel_inc,
    ctrl_sel_rst_n,
    k_one,
    k_zero,
    pad_ui_in,
    pad_uio_in,
    pad_uio_oe_n,
    pad_uio_out,
    pad_uo_out,
    spine_bot_iw,
    spine_bot_ow,
    spine_top_iw,
    spine_top_ow);
 input ctrl_ena;
 input ctrl_sel_inc;
 input ctrl_sel_rst_n;
 output k_one;
 output k_zero;
 input [9:0] pad_ui_in;
 input [7:0] pad_uio_in;
 output [7:0] pad_uio_oe_n;
 output [7:0] pad_uio_out;
 output [7:0] pad_uo_out;
 output [29:0] spine_bot_iw;
 input [25:0] spine_bot_ow;
 output [29:0] spine_top_iw;
 input [25:0] spine_top_ow;

 wire \ctrl_ibuf_I[0].z ;
 wire \ctrl_ibuf_I[1].z ;
 wire \ctrl_ibuf_I[2].z ;
 wire \genblk1[0].tbuf_pol_spine_ow_I.t ;
 wire \genblk1[0].tbuf_pol_spine_ow_I.tx ;
 wire \genblk1[0].tbuf_spine_ow_I[0].a ;
 wire \genblk1[0].tie_I.hi ;
 wire \genblk1[1].tbuf_pol_spine_ow_I.t ;
 wire \genblk1[1].tbuf_pol_spine_ow_I.tx ;
 wire \genblk1[1].tbuf_spine_ow_I[0].a ;
 wire \genblk1[1].tie_I.hi ;
 wire \genblk2[0].ctrl_ena_buf_I.e ;
 wire \genblk2[0].ctrl_ena_buf_I.genblk1.l ;
 wire \genblk2[0].ctrl_ena_buf_I.z ;
 wire \genblk2[0].pad_ui_in_buf_I[0].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[0].z ;
 wire \genblk2[0].pad_ui_in_buf_I[1].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[1].z ;
 wire \genblk2[0].pad_ui_in_buf_I[2].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[2].z ;
 wire \genblk2[0].pad_ui_in_buf_I[3].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[3].z ;
 wire \genblk2[0].pad_ui_in_buf_I[4].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[4].z ;
 wire \genblk2[0].pad_ui_in_buf_I[5].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[5].z ;
 wire \genblk2[0].pad_ui_in_buf_I[6].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[6].z ;
 wire \genblk2[0].pad_ui_in_buf_I[7].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[7].z ;
 wire \genblk2[0].pad_ui_in_buf_I[8].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[8].z ;
 wire \genblk2[0].pad_ui_in_buf_I[9].genblk1.l ;
 wire \genblk2[0].pad_ui_in_buf_I[9].z ;
 wire \genblk2[0].pad_uio_in_buf_I[0].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[0].z ;
 wire \genblk2[0].pad_uio_in_buf_I[1].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[1].z ;
 wire \genblk2[0].pad_uio_in_buf_I[2].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[2].z ;
 wire \genblk2[0].pad_uio_in_buf_I[3].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[3].z ;
 wire \genblk2[0].pad_uio_in_buf_I[4].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[4].z ;
 wire \genblk2[0].pad_uio_in_buf_I[5].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[5].z ;
 wire \genblk2[0].pad_uio_in_buf_I[6].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[6].z ;
 wire \genblk2[0].pad_uio_in_buf_I[7].genblk1.l ;
 wire \genblk2[0].pad_uio_in_buf_I[7].z ;
 wire \genblk2[0].sel_cnt_buf_I[0].a ;
 wire \genblk2[0].sel_cnt_buf_I[0].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[0].z ;
 wire \genblk2[0].sel_cnt_buf_I[1].a ;
 wire \genblk2[0].sel_cnt_buf_I[1].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[1].z ;
 wire \genblk2[0].sel_cnt_buf_I[2].a ;
 wire \genblk2[0].sel_cnt_buf_I[2].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[2].z ;
 wire \genblk2[0].sel_cnt_buf_I[3].a ;
 wire \genblk2[0].sel_cnt_buf_I[3].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[3].z ;
 wire \genblk2[0].sel_cnt_buf_I[4].a ;
 wire \genblk2[0].sel_cnt_buf_I[4].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[4].z ;
 wire \genblk2[0].sel_cnt_buf_I[5].a ;
 wire \genblk2[0].sel_cnt_buf_I[5].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[5].z ;
 wire \genblk2[0].sel_cnt_buf_I[6].a ;
 wire \genblk2[0].sel_cnt_buf_I[6].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[6].z ;
 wire \genblk2[0].sel_cnt_buf_I[7].a ;
 wire \genblk2[0].sel_cnt_buf_I[7].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[7].z ;
 wire \genblk2[0].sel_cnt_buf_I[8].a ;
 wire \genblk2[0].sel_cnt_buf_I[8].genblk1.l ;
 wire \genblk2[0].sel_cnt_buf_I[8].z ;
 wire \genblk2[0].tie_guard_I[0].hi ;
 wire \genblk2[0].tie_guard_I[0].lo ;
 wire \genblk2[0].tie_guard_I[1].hi ;
 wire \genblk2[0].tie_guard_I[1].lo ;
 wire \genblk2[1].ctrl_ena_buf_I.e ;
 wire \genblk2[1].ctrl_ena_buf_I.genblk1.l ;
 wire \genblk2[1].ctrl_ena_buf_I.z ;
 wire \genblk2[1].pad_ui_in_buf_I[0].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[0].z ;
 wire \genblk2[1].pad_ui_in_buf_I[1].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[1].z ;
 wire \genblk2[1].pad_ui_in_buf_I[2].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[2].z ;
 wire \genblk2[1].pad_ui_in_buf_I[3].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[3].z ;
 wire \genblk2[1].pad_ui_in_buf_I[4].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[4].z ;
 wire \genblk2[1].pad_ui_in_buf_I[5].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[5].z ;
 wire \genblk2[1].pad_ui_in_buf_I[6].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[6].z ;
 wire \genblk2[1].pad_ui_in_buf_I[7].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[7].z ;
 wire \genblk2[1].pad_ui_in_buf_I[8].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[8].z ;
 wire \genblk2[1].pad_ui_in_buf_I[9].genblk1.l ;
 wire \genblk2[1].pad_ui_in_buf_I[9].z ;
 wire \genblk2[1].pad_uio_in_buf_I[0].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[0].z ;
 wire \genblk2[1].pad_uio_in_buf_I[1].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[1].z ;
 wire \genblk2[1].pad_uio_in_buf_I[2].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[2].z ;
 wire \genblk2[1].pad_uio_in_buf_I[3].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[3].z ;
 wire \genblk2[1].pad_uio_in_buf_I[4].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[4].z ;
 wire \genblk2[1].pad_uio_in_buf_I[5].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[5].z ;
 wire \genblk2[1].pad_uio_in_buf_I[6].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[6].z ;
 wire \genblk2[1].pad_uio_in_buf_I[7].genblk1.l ;
 wire \genblk2[1].pad_uio_in_buf_I[7].z ;
 wire \genblk2[1].sel_cnt_buf_I[0].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[0].z ;
 wire \genblk2[1].sel_cnt_buf_I[1].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[1].z ;
 wire \genblk2[1].sel_cnt_buf_I[2].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[2].z ;
 wire \genblk2[1].sel_cnt_buf_I[3].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[3].z ;
 wire \genblk2[1].sel_cnt_buf_I[4].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[4].z ;
 wire \genblk2[1].sel_cnt_buf_I[5].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[5].z ;
 wire \genblk2[1].sel_cnt_buf_I[6].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[6].z ;
 wire \genblk2[1].sel_cnt_buf_I[7].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[7].z ;
 wire \genblk2[1].sel_cnt_buf_I[8].genblk1.l ;
 wire \genblk2[1].sel_cnt_buf_I[8].z ;
 wire \genblk2[1].tie_guard_I[0].hi ;
 wire \genblk2[1].tie_guard_I[0].lo ;
 wire \genblk2[1].tie_guard_I[1].hi ;
 wire \genblk2[1].tie_guard_I[1].lo ;
 wire \sel_cnt_gen[0].cnt_bit_I.d ;
 wire \sel_cnt_gen[1].cnt_bit_I.d ;
 wire \sel_cnt_gen[2].cnt_bit_I.d ;
 wire \sel_cnt_gen[3].cnt_bit_I.d ;
 wire \sel_cnt_gen[4].cnt_bit_I.d ;
 wire \sel_cnt_gen[5].cnt_bit_I.d ;
 wire \sel_cnt_gen[5].cnt_bit_I.q ;
 wire \sel_cnt_gen[6].cnt_bit_I.d ;
 wire \sel_cnt_gen[7].cnt_bit_I.d ;
 wire \sel_cnt_gen[8].cnt_bit_I.d ;
 wire \sel_cnt_gen[9].cnt_bit_I.d ;
 wire \side_sel_buf_I.z ;
 wire \uio_oe_ibuf_I[0].z ;
 wire \uio_oe_ibuf_I[10].z ;
 wire \uio_oe_ibuf_I[11].z ;
 wire \uio_oe_ibuf_I[12].z ;
 wire \uio_oe_ibuf_I[13].z ;
 wire \uio_oe_ibuf_I[14].z ;
 wire \uio_oe_ibuf_I[15].z ;
 wire \uio_oe_ibuf_I[1].z ;
 wire \uio_oe_ibuf_I[2].z ;
 wire \uio_oe_ibuf_I[3].z ;
 wire \uio_oe_ibuf_I[4].z ;
 wire \uio_oe_ibuf_I[5].z ;
 wire \uio_oe_ibuf_I[6].z ;
 wire \uio_oe_ibuf_I[7].z ;
 wire \uio_oe_ibuf_I[8].z ;
 wire \uio_oe_ibuf_I[9].z ;
 wire \uio_oe_mux_I[0].x ;
 wire \uio_oe_mux_I[1].x ;
 wire \uio_oe_mux_I[2].x ;
 wire \uio_oe_mux_I[3].x ;
 wire \uio_oe_mux_I[4].x ;
 wire \uio_oe_mux_I[5].x ;
 wire \uio_oe_mux_I[6].x ;
 wire \uio_oe_mux_I[7].x ;
 wire \uio_oe_obuf_I[0].z ;
 wire \uio_oe_obuf_I[1].z ;
 wire \uio_oe_obuf_I[2].z ;
 wire \uio_oe_obuf_I[3].z ;
 wire \uio_oe_obuf_I[4].z ;
 wire \uio_oe_obuf_I[5].z ;
 wire \uio_oe_obuf_I[6].z ;
 wire \uio_oe_obuf_I[7].z ;
 wire \uio_out_ibuf_I[0].z ;
 wire \uio_out_ibuf_I[10].z ;
 wire \uio_out_ibuf_I[11].z ;
 wire \uio_out_ibuf_I[12].z ;
 wire \uio_out_ibuf_I[13].z ;
 wire \uio_out_ibuf_I[14].z ;
 wire \uio_out_ibuf_I[15].z ;
 wire \uio_out_ibuf_I[1].z ;
 wire \uio_out_ibuf_I[2].z ;
 wire \uio_out_ibuf_I[3].z ;
 wire \uio_out_ibuf_I[4].z ;
 wire \uio_out_ibuf_I[5].z ;
 wire \uio_out_ibuf_I[6].z ;
 wire \uio_out_ibuf_I[7].z ;
 wire \uio_out_ibuf_I[8].z ;
 wire \uio_out_ibuf_I[9].z ;
 wire \uio_out_mux_I[0].x ;
 wire \uio_out_mux_I[1].x ;
 wire \uio_out_mux_I[2].x ;
 wire \uio_out_mux_I[3].x ;
 wire \uio_out_mux_I[4].x ;
 wire \uio_out_mux_I[5].x ;
 wire \uio_out_mux_I[6].x ;
 wire \uio_out_mux_I[7].x ;
 wire \uio_out_obuf_I[0].z ;
 wire \uio_out_obuf_I[1].z ;
 wire \uio_out_obuf_I[2].z ;
 wire \uio_out_obuf_I[3].z ;
 wire \uio_out_obuf_I[4].z ;
 wire \uio_out_obuf_I[5].z ;
 wire \uio_out_obuf_I[6].z ;
 wire \uio_out_obuf_I[7].z ;
 wire \uo_out_ibuf_I[0].z ;
 wire \uo_out_ibuf_I[10].z ;
 wire \uo_out_ibuf_I[11].z ;
 wire \uo_out_ibuf_I[12].z ;
 wire \uo_out_ibuf_I[13].z ;
 wire \uo_out_ibuf_I[14].z ;
 wire \uo_out_ibuf_I[15].z ;
 wire \uo_out_ibuf_I[1].z ;
 wire \uo_out_ibuf_I[2].z ;
 wire \uo_out_ibuf_I[3].z ;
 wire \uo_out_ibuf_I[4].z ;
 wire \uo_out_ibuf_I[5].z ;
 wire \uo_out_ibuf_I[6].z ;
 wire \uo_out_ibuf_I[7].z ;
 wire \uo_out_ibuf_I[8].z ;
 wire \uo_out_ibuf_I[9].z ;
 wire \uo_out_mux_I[0].x ;
 wire \uo_out_mux_I[1].x ;
 wire \uo_out_mux_I[2].x ;
 wire \uo_out_mux_I[3].x ;
 wire \uo_out_mux_I[4].x ;
 wire \uo_out_mux_I[5].x ;
 wire \uo_out_mux_I[6].x ;
 wire \uo_out_mux_I[7].x ;
 wire \uo_out_obuf_I[0].z ;
 wire \uo_out_obuf_I[1].z ;
 wire \uo_out_obuf_I[2].z ;
 wire \uo_out_obuf_I[3].z ;
 wire \uo_out_obuf_I[4].z ;
 wire \uo_out_obuf_I[5].z ;
 wire \uo_out_obuf_I[6].z ;
 wire \uo_out_obuf_I[7].z ;

 sky130_fd_sc_hd__nand2_1 _0_ (.A(\ctrl_ibuf_I[0].z ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .Y(\genblk1[0].tbuf_pol_spine_ow_I.t ));
 sky130_fd_sc_hd__nand2_1 _1_ (.A(\ctrl_ibuf_I[0].z ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .Y(\genblk1[1].tbuf_pol_spine_ow_I.t ));
 sky130_fd_sc_hd__diode_2 \ctrl_diode_I[0].cell0_I  (.DIODE(ctrl_ena));
 sky130_fd_sc_hd__diode_2 \ctrl_diode_I[1].cell0_I  (.DIODE(ctrl_sel_inc));
 sky130_fd_sc_hd__diode_2 \ctrl_diode_I[2].cell0_I  (.DIODE(ctrl_sel_rst_n));
 sky130_fd_sc_hd__buf_2 \ctrl_ibuf_I[0].genblk1.cell0_I  (.A(ctrl_ena),
    .X(\ctrl_ibuf_I[0].z ));
 sky130_fd_sc_hd__buf_2 \ctrl_ibuf_I[1].genblk1.cell0_I  (.A(ctrl_sel_inc),
    .X(\ctrl_ibuf_I[1].z ));
 sky130_fd_sc_hd__buf_2 \ctrl_ibuf_I[2].genblk1.cell0_I  (.A(ctrl_sel_rst_n),
    .X(\ctrl_ibuf_I[2].z ));
 sky130_fd_sc_hd__bufinv_8 \genblk1[0].tbuf_pol_spine_ow_I.cell0_I  (.A(\genblk1[0].tbuf_pol_spine_ow_I.t ),
    .Y(\genblk1[0].tbuf_pol_spine_ow_I.tx ));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[1]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[11]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[12]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[13]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[14]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[15]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[16]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[17]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[18]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[19]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[20]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[2]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[21]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[22]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[23]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[24]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[3]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[4]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[5]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[6]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[7]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[8]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[9]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[0].tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\genblk1[0].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[0].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_bot_ow[10]));
 sky130_fd_sc_hd__conb_1 \genblk1[0].tie_I.cell_I  (.HI(\genblk1[0].tie_I.hi ),
    .LO(\genblk1[0].tbuf_spine_ow_I[0].a ));
 sky130_fd_sc_hd__bufinv_8 \genblk1[1].tbuf_pol_spine_ow_I.cell0_I  (.A(\genblk1[1].tbuf_pol_spine_ow_I.t ),
    .Y(\genblk1[1].tbuf_pol_spine_ow_I.tx ));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[0].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[1]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[10].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[11]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[11].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[12]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[12].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[13]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[13].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[14]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[14].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[15]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[15].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[16]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[16].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[17]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[17].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[18]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[18].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[19]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[19].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[20]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[1].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[2]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[20].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[21]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[21].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[22]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[22].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[23]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[23].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[24]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[2].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[3]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[3].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[4]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[4].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[5]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[5].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[6]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[6].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[7]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[7].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[8]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[8].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[9]));
 sky130_fd_sc_hd__ebufn_1 \genblk1[1].tbuf_spine_ow_I[9].genblk1.cell0_I  (.A(\genblk1[1].tbuf_spine_ow_I[0].a ),
    .TE_B(\genblk1[1].tbuf_pol_spine_ow_I.tx ),
    .Z(spine_top_ow[10]));
 sky130_fd_sc_hd__conb_1 \genblk1[1].tie_I.cell_I  (.HI(\genblk1[1].tie_I.hi ),
    .LO(\genblk1[1].tbuf_spine_ow_I[0].a ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].ctrl_ena_buf_I.genblk1.cell0_I  (.A(\ctrl_ibuf_I[0].z ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].ctrl_ena_buf_I.genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].ctrl_ena_buf_I.genblk1.cell1_I  (.A(\genblk2[0].ctrl_ena_buf_I.genblk1.l ),
    .X(\genblk2[0].ctrl_ena_buf_I.z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[0].genblk1.cell0_I  (.A(pad_ui_in[0]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[0].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[0].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[1].genblk1.cell0_I  (.A(pad_ui_in[1]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[1].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[1].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[2].genblk1.cell0_I  (.A(pad_ui_in[2]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[2].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[2].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[3].genblk1.cell0_I  (.A(pad_ui_in[3]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[3].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[3].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[4].genblk1.cell0_I  (.A(pad_ui_in[4]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[4].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[4].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[5].genblk1.cell0_I  (.A(pad_ui_in[5]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[5].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[5].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[6].genblk1.cell0_I  (.A(pad_ui_in[6]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[6].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[6].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[7].genblk1.cell0_I  (.A(pad_ui_in[7]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[7].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[7].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[8].genblk1.cell0_I  (.A(pad_ui_in[8]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[8].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[8].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[8].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[8].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_ui_in_buf_I[9].genblk1.cell0_I  (.A(pad_ui_in[9]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_ui_in_buf_I[9].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_ui_in_buf_I[9].genblk1.cell1_I  (.A(\genblk2[0].pad_ui_in_buf_I[9].genblk1.l ),
    .X(\genblk2[0].pad_ui_in_buf_I[9].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[0].genblk1.cell0_I  (.A(pad_uio_in[0]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[0].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[0].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[1].genblk1.cell0_I  (.A(pad_uio_in[1]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[1].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[1].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[2].genblk1.cell0_I  (.A(pad_uio_in[2]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[2].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[2].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[3].genblk1.cell0_I  (.A(pad_uio_in[3]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[3].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[3].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[4].genblk1.cell0_I  (.A(pad_uio_in[4]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[4].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[4].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[5].genblk1.cell0_I  (.A(pad_uio_in[5]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[5].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[5].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[6].genblk1.cell0_I  (.A(pad_uio_in[6]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[6].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[6].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].pad_uio_in_buf_I[7].genblk1.cell0_I  (.A(pad_uio_in[7]),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].pad_uio_in_buf_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].pad_uio_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[0].pad_uio_in_buf_I[7].genblk1.l ),
    .X(\genblk2[0].pad_uio_in_buf_I[7].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[0].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[0].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[0].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[0].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[0].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[1].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[1].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[1].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[1].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[1].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[2].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[2].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[2].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[2].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[2].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[3].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[3].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[3].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[3].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[3].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[4].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[4].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[4].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[4].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[4].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[5].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[5].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[5].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[5].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[5].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[6].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[6].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[6].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[6].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[6].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[7].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[7].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[7].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[7].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[7].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[0].sel_cnt_buf_I[8].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[8].a ),
    .B(\genblk2[0].ctrl_ena_buf_I.e ),
    .X(\genblk2[0].sel_cnt_buf_I[8].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[0].sel_cnt_buf_I[8].genblk1.cell1_I  (.A(\genblk2[0].sel_cnt_buf_I[8].genblk1.l ),
    .X(\genblk2[0].sel_cnt_buf_I[8].z ));
 sky130_fd_sc_hd__conb_1 \genblk2[0].tie_guard_I[0].cell_I  (.HI(\genblk2[0].tie_guard_I[0].hi ),
    .LO(\genblk2[0].tie_guard_I[0].lo ));
 sky130_fd_sc_hd__conb_1 \genblk2[0].tie_guard_I[1].cell_I  (.HI(\genblk2[0].tie_guard_I[1].hi ),
    .LO(\genblk2[0].tie_guard_I[1].lo ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].ctrl_ena_buf_I.genblk1.cell0_I  (.A(\ctrl_ibuf_I[0].z ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].ctrl_ena_buf_I.genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].ctrl_ena_buf_I.genblk1.cell1_I  (.A(\genblk2[1].ctrl_ena_buf_I.genblk1.l ),
    .X(\genblk2[1].ctrl_ena_buf_I.z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[0].genblk1.cell0_I  (.A(pad_ui_in[0]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[0].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[0].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[1].genblk1.cell0_I  (.A(pad_ui_in[1]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[1].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[1].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[2].genblk1.cell0_I  (.A(pad_ui_in[2]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[2].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[2].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[3].genblk1.cell0_I  (.A(pad_ui_in[3]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[3].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[3].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[4].genblk1.cell0_I  (.A(pad_ui_in[4]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[4].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[4].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[5].genblk1.cell0_I  (.A(pad_ui_in[5]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[5].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[5].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[6].genblk1.cell0_I  (.A(pad_ui_in[6]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[6].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[6].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[7].genblk1.cell0_I  (.A(pad_ui_in[7]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[7].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[7].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[8].genblk1.cell0_I  (.A(pad_ui_in[8]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[8].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[8].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[8].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[8].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_ui_in_buf_I[9].genblk1.cell0_I  (.A(pad_ui_in[9]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_ui_in_buf_I[9].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_ui_in_buf_I[9].genblk1.cell1_I  (.A(\genblk2[1].pad_ui_in_buf_I[9].genblk1.l ),
    .X(\genblk2[1].pad_ui_in_buf_I[9].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[0].genblk1.cell0_I  (.A(pad_uio_in[0]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[0].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[0].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[0].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[1].genblk1.cell0_I  (.A(pad_uio_in[1]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[1].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[1].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[1].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[2].genblk1.cell0_I  (.A(pad_uio_in[2]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[2].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[2].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[2].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[3].genblk1.cell0_I  (.A(pad_uio_in[3]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[3].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[3].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[3].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[4].genblk1.cell0_I  (.A(pad_uio_in[4]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[4].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[4].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[4].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[5].genblk1.cell0_I  (.A(pad_uio_in[5]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[5].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[5].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[5].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[6].genblk1.cell0_I  (.A(pad_uio_in[6]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[6].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[6].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[6].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].pad_uio_in_buf_I[7].genblk1.cell0_I  (.A(pad_uio_in[7]),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].pad_uio_in_buf_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].pad_uio_in_buf_I[7].genblk1.cell1_I  (.A(\genblk2[1].pad_uio_in_buf_I[7].genblk1.l ),
    .X(\genblk2[1].pad_uio_in_buf_I[7].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[0].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[0].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[0].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[0].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[0].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[0].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[1].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[1].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[1].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[1].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[1].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[1].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[2].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[2].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[2].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[2].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[2].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[2].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[3].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[3].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[3].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[3].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[3].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[3].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[4].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[4].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[4].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[4].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[4].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[4].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[5].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[5].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[5].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[5].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[5].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[5].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[6].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[6].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[6].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[6].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[6].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[6].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[7].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[7].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[7].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[7].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[7].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[7].z ));
 sky130_fd_sc_hd__and2_2 \genblk2[1].sel_cnt_buf_I[8].genblk1.cell0_I  (.A(\genblk2[0].sel_cnt_buf_I[8].a ),
    .B(\genblk2[1].ctrl_ena_buf_I.e ),
    .X(\genblk2[1].sel_cnt_buf_I[8].genblk1.l ));
 sky130_fd_sc_hd__buf_8 \genblk2[1].sel_cnt_buf_I[8].genblk1.cell1_I  (.A(\genblk2[1].sel_cnt_buf_I[8].genblk1.l ),
    .X(\genblk2[1].sel_cnt_buf_I[8].z ));
 sky130_fd_sc_hd__conb_1 \genblk2[1].tie_guard_I[0].cell_I  (.HI(\genblk2[1].tie_guard_I[0].hi ),
    .LO(\genblk2[1].tie_guard_I[0].lo ));
 sky130_fd_sc_hd__conb_1 \genblk2[1].tie_guard_I[1].cell_I  (.HI(\genblk2[1].tie_guard_I[1].hi ),
    .LO(\genblk2[1].tie_guard_I[1].lo ));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[0].cell0_I  (.DIODE(pad_ui_in[0]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[1].cell0_I  (.DIODE(pad_ui_in[1]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[2].cell0_I  (.DIODE(pad_ui_in[2]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[3].cell0_I  (.DIODE(pad_ui_in[3]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[4].cell0_I  (.DIODE(pad_ui_in[4]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[5].cell0_I  (.DIODE(pad_ui_in[5]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[6].cell0_I  (.DIODE(pad_ui_in[6]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[7].cell0_I  (.DIODE(pad_ui_in[7]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[8].cell0_I  (.DIODE(pad_ui_in[8]));
 sky130_fd_sc_hd__diode_2 \pad_ui_in_diode_I[9].cell0_I  (.DIODE(pad_ui_in[9]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[0].cell0_I  (.DIODE(pad_uio_in[0]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[1].cell0_I  (.DIODE(pad_uio_in[1]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[2].cell0_I  (.DIODE(pad_uio_in[2]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[3].cell0_I  (.DIODE(pad_uio_in[3]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[4].cell0_I  (.DIODE(pad_uio_in[4]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[5].cell0_I  (.DIODE(pad_uio_in[5]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[6].cell0_I  (.DIODE(pad_uio_in[6]));
 sky130_fd_sc_hd__diode_2 \pad_uio_in_diode_I[7].cell0_I  (.DIODE(pad_uio_in[7]));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[0].cnt_bit_I.cell0_I  (.CLK(\ctrl_ibuf_I[1].z ),
    .D(\sel_cnt_gen[0].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[0].a ),
    .Q_N(\sel_cnt_gen[0].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[1].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[0].cnt_bit_I.d ),
    .D(\sel_cnt_gen[1].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[1].a ),
    .Q_N(\sel_cnt_gen[1].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[2].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[1].cnt_bit_I.d ),
    .D(\sel_cnt_gen[2].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[2].a ),
    .Q_N(\sel_cnt_gen[2].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[3].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[2].cnt_bit_I.d ),
    .D(\sel_cnt_gen[3].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[3].a ),
    .Q_N(\sel_cnt_gen[3].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[4].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[3].cnt_bit_I.d ),
    .D(\sel_cnt_gen[4].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[4].a ),
    .Q_N(\sel_cnt_gen[4].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[5].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[4].cnt_bit_I.d ),
    .D(\sel_cnt_gen[5].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\sel_cnt_gen[5].cnt_bit_I.q ),
    .Q_N(\sel_cnt_gen[5].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[6].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[5].cnt_bit_I.d ),
    .D(\sel_cnt_gen[6].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[5].a ),
    .Q_N(\sel_cnt_gen[6].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[7].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[6].cnt_bit_I.d ),
    .D(\sel_cnt_gen[7].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[6].a ),
    .Q_N(\sel_cnt_gen[7].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[8].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[7].cnt_bit_I.d ),
    .D(\sel_cnt_gen[8].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[7].a ),
    .Q_N(\sel_cnt_gen[8].cnt_bit_I.d ));
 sky130_fd_sc_hd__dfrbp_2 \sel_cnt_gen[9].cnt_bit_I.cell0_I  (.CLK(\sel_cnt_gen[8].cnt_bit_I.d ),
    .D(\sel_cnt_gen[9].cnt_bit_I.d ),
    .RESET_B(\ctrl_ibuf_I[2].z ),
    .Q(\genblk2[0].sel_cnt_buf_I[8].a ),
    .Q_N(\sel_cnt_gen[9].cnt_bit_I.d ));
 sky130_fd_sc_hd__bufinv_8 \side_ena0_buf_I.genblk1.cell0_I  (.A(\sel_cnt_gen[5].cnt_bit_I.q ),
    .Y(\genblk2[0].ctrl_ena_buf_I.e ));
 sky130_fd_sc_hd__buf_8 \side_ena1_buf_I.genblk1.cell0_I  (.A(\sel_cnt_gen[5].cnt_bit_I.q ),
    .X(\genblk2[1].ctrl_ena_buf_I.e ));
 sky130_fd_sc_hd__buf_8 \side_sel_buf_I.genblk1.cell0_I  (.A(\sel_cnt_gen[5].cnt_bit_I.q ),
    .X(\side_sel_buf_I.z ));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[0].cell0_I  (.DIODE(spine_bot_ow[0]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[10].cell0_I  (.DIODE(spine_bot_ow[10]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[11].cell0_I  (.DIODE(spine_bot_ow[11]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[12].cell0_I  (.DIODE(spine_bot_ow[12]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[13].cell0_I  (.DIODE(spine_bot_ow[13]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[14].cell0_I  (.DIODE(spine_bot_ow[14]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[15].cell0_I  (.DIODE(spine_bot_ow[15]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[16].cell0_I  (.DIODE(spine_bot_ow[16]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[17].cell0_I  (.DIODE(spine_bot_ow[17]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[18].cell0_I  (.DIODE(spine_bot_ow[18]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[19].cell0_I  (.DIODE(spine_bot_ow[19]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[1].cell0_I  (.DIODE(spine_bot_ow[1]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[20].cell0_I  (.DIODE(spine_bot_ow[20]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[21].cell0_I  (.DIODE(spine_bot_ow[21]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[22].cell0_I  (.DIODE(spine_bot_ow[22]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[23].cell0_I  (.DIODE(spine_bot_ow[23]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[24].cell0_I  (.DIODE(spine_bot_ow[24]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[25].cell0_I  (.DIODE(spine_bot_ow[25]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[26].cell0_I  (.DIODE(spine_top_ow[0]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[27].cell0_I  (.DIODE(spine_top_ow[1]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[28].cell0_I  (.DIODE(spine_top_ow[2]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[29].cell0_I  (.DIODE(spine_top_ow[3]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[2].cell0_I  (.DIODE(spine_bot_ow[2]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[30].cell0_I  (.DIODE(spine_top_ow[4]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[31].cell0_I  (.DIODE(spine_top_ow[5]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[32].cell0_I  (.DIODE(spine_top_ow[6]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[33].cell0_I  (.DIODE(spine_top_ow[7]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[34].cell0_I  (.DIODE(spine_top_ow[8]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[35].cell0_I  (.DIODE(spine_top_ow[9]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[36].cell0_I  (.DIODE(spine_top_ow[10]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[37].cell0_I  (.DIODE(spine_top_ow[11]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[38].cell0_I  (.DIODE(spine_top_ow[12]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[39].cell0_I  (.DIODE(spine_top_ow[13]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[3].cell0_I  (.DIODE(spine_bot_ow[3]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[40].cell0_I  (.DIODE(spine_top_ow[14]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[41].cell0_I  (.DIODE(spine_top_ow[15]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[42].cell0_I  (.DIODE(spine_top_ow[16]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[43].cell0_I  (.DIODE(spine_top_ow[17]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[44].cell0_I  (.DIODE(spine_top_ow[18]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[45].cell0_I  (.DIODE(spine_top_ow[19]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[46].cell0_I  (.DIODE(spine_top_ow[20]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[47].cell0_I  (.DIODE(spine_top_ow[21]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[48].cell0_I  (.DIODE(spine_top_ow[22]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[49].cell0_I  (.DIODE(spine_top_ow[23]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[4].cell0_I  (.DIODE(spine_bot_ow[4]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[50].cell0_I  (.DIODE(spine_top_ow[24]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[51].cell0_I  (.DIODE(spine_top_ow[25]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[5].cell0_I  (.DIODE(spine_bot_ow[5]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[6].cell0_I  (.DIODE(spine_bot_ow[6]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[7].cell0_I  (.DIODE(spine_bot_ow[7]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[8].cell0_I  (.DIODE(spine_bot_ow[8]));
 sky130_fd_sc_hd__diode_2 \spine_diode_I[9].cell0_I  (.DIODE(spine_bot_ow[9]));
 sky130_fd_sc_hd__conb_1 \tie_I.cell_I  (.HI(k_one),
    .LO(k_zero));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[0].genblk1.cell0_I  (.A(spine_bot_ow[17]),
    .X(\uio_oe_ibuf_I[0].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[10].genblk1.cell0_I  (.A(spine_top_ow[19]),
    .X(\uio_oe_ibuf_I[10].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[11].genblk1.cell0_I  (.A(spine_top_ow[20]),
    .X(\uio_oe_ibuf_I[11].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[12].genblk1.cell0_I  (.A(spine_top_ow[21]),
    .X(\uio_oe_ibuf_I[12].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[13].genblk1.cell0_I  (.A(spine_top_ow[22]),
    .X(\uio_oe_ibuf_I[13].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[14].genblk1.cell0_I  (.A(spine_top_ow[23]),
    .X(\uio_oe_ibuf_I[14].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[15].genblk1.cell0_I  (.A(spine_top_ow[24]),
    .X(\uio_oe_ibuf_I[15].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[1].genblk1.cell0_I  (.A(spine_bot_ow[18]),
    .X(\uio_oe_ibuf_I[1].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[2].genblk1.cell0_I  (.A(spine_bot_ow[19]),
    .X(\uio_oe_ibuf_I[2].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[3].genblk1.cell0_I  (.A(spine_bot_ow[20]),
    .X(\uio_oe_ibuf_I[3].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[4].genblk1.cell0_I  (.A(spine_bot_ow[21]),
    .X(\uio_oe_ibuf_I[4].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[5].genblk1.cell0_I  (.A(spine_bot_ow[22]),
    .X(\uio_oe_ibuf_I[5].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[6].genblk1.cell0_I  (.A(spine_bot_ow[23]),
    .X(\uio_oe_ibuf_I[6].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[7].genblk1.cell0_I  (.A(spine_bot_ow[24]),
    .X(\uio_oe_ibuf_I[7].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[8].genblk1.cell0_I  (.A(spine_top_ow[17]),
    .X(\uio_oe_ibuf_I[8].z ));
 sky130_fd_sc_hd__buf_2 \uio_oe_ibuf_I[9].genblk1.cell0_I  (.A(spine_top_ow[18]),
    .X(\uio_oe_ibuf_I[9].z ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[0].cell0_I  (.A0(\uio_oe_ibuf_I[0].z ),
    .A1(\uio_oe_ibuf_I[8].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[0].x ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[1].cell0_I  (.A0(\uio_oe_ibuf_I[1].z ),
    .A1(\uio_oe_ibuf_I[9].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[1].x ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[2].cell0_I  (.A0(\uio_oe_ibuf_I[2].z ),
    .A1(\uio_oe_ibuf_I[10].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[2].x ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[3].cell0_I  (.A0(\uio_oe_ibuf_I[3].z ),
    .A1(\uio_oe_ibuf_I[11].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[3].x ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[4].cell0_I  (.A0(\uio_oe_ibuf_I[4].z ),
    .A1(\uio_oe_ibuf_I[12].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[4].x ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[5].cell0_I  (.A0(\uio_oe_ibuf_I[5].z ),
    .A1(\uio_oe_ibuf_I[13].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[5].x ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[6].cell0_I  (.A0(\uio_oe_ibuf_I[6].z ),
    .A1(\uio_oe_ibuf_I[14].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[6].x ));
 sky130_fd_sc_hd__mux2_2 \uio_oe_mux_I[7].cell0_I  (.A0(\uio_oe_ibuf_I[7].z ),
    .A1(\uio_oe_ibuf_I[15].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_oe_mux_I[7].x ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[0].genblk1.cell0_I  (.A(\uio_oe_mux_I[0].x ),
    .Y(\uio_oe_obuf_I[0].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[1].genblk1.cell0_I  (.A(\uio_oe_mux_I[1].x ),
    .Y(\uio_oe_obuf_I[1].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[2].genblk1.cell0_I  (.A(\uio_oe_mux_I[2].x ),
    .Y(\uio_oe_obuf_I[2].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[3].genblk1.cell0_I  (.A(\uio_oe_mux_I[3].x ),
    .Y(\uio_oe_obuf_I[3].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[4].genblk1.cell0_I  (.A(\uio_oe_mux_I[4].x ),
    .Y(\uio_oe_obuf_I[4].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[5].genblk1.cell0_I  (.A(\uio_oe_mux_I[5].x ),
    .Y(\uio_oe_obuf_I[5].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[6].genblk1.cell0_I  (.A(\uio_oe_mux_I[6].x ),
    .Y(\uio_oe_obuf_I[6].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_oe_obuf_I[7].genblk1.cell0_I  (.A(\uio_oe_mux_I[7].x ),
    .Y(\uio_oe_obuf_I[7].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[0].genblk1.cell0_I  (.A(spine_bot_ow[9]),
    .Y(\uio_out_ibuf_I[0].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[10].genblk1.cell0_I  (.A(spine_top_ow[11]),
    .Y(\uio_out_ibuf_I[10].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[11].genblk1.cell0_I  (.A(spine_top_ow[12]),
    .Y(\uio_out_ibuf_I[11].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[12].genblk1.cell0_I  (.A(spine_top_ow[13]),
    .Y(\uio_out_ibuf_I[12].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[13].genblk1.cell0_I  (.A(spine_top_ow[14]),
    .Y(\uio_out_ibuf_I[13].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[14].genblk1.cell0_I  (.A(spine_top_ow[15]),
    .Y(\uio_out_ibuf_I[14].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[15].genblk1.cell0_I  (.A(spine_top_ow[16]),
    .Y(\uio_out_ibuf_I[15].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[1].genblk1.cell0_I  (.A(spine_bot_ow[10]),
    .Y(\uio_out_ibuf_I[1].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[2].genblk1.cell0_I  (.A(spine_bot_ow[11]),
    .Y(\uio_out_ibuf_I[2].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[3].genblk1.cell0_I  (.A(spine_bot_ow[12]),
    .Y(\uio_out_ibuf_I[3].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[4].genblk1.cell0_I  (.A(spine_bot_ow[13]),
    .Y(\uio_out_ibuf_I[4].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[5].genblk1.cell0_I  (.A(spine_bot_ow[14]),
    .Y(\uio_out_ibuf_I[5].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[6].genblk1.cell0_I  (.A(spine_bot_ow[15]),
    .Y(\uio_out_ibuf_I[6].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[7].genblk1.cell0_I  (.A(spine_bot_ow[16]),
    .Y(\uio_out_ibuf_I[7].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[8].genblk1.cell0_I  (.A(spine_top_ow[9]),
    .Y(\uio_out_ibuf_I[8].z ));
 sky130_fd_sc_hd__inv_2 \uio_out_ibuf_I[9].genblk1.cell0_I  (.A(spine_top_ow[10]),
    .Y(\uio_out_ibuf_I[9].z ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[0].cell0_I  (.A0(\uio_out_ibuf_I[0].z ),
    .A1(\uio_out_ibuf_I[8].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[0].x ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[1].cell0_I  (.A0(\uio_out_ibuf_I[1].z ),
    .A1(\uio_out_ibuf_I[9].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[1].x ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[2].cell0_I  (.A0(\uio_out_ibuf_I[2].z ),
    .A1(\uio_out_ibuf_I[10].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[2].x ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[3].cell0_I  (.A0(\uio_out_ibuf_I[3].z ),
    .A1(\uio_out_ibuf_I[11].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[3].x ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[4].cell0_I  (.A0(\uio_out_ibuf_I[4].z ),
    .A1(\uio_out_ibuf_I[12].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[4].x ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[5].cell0_I  (.A0(\uio_out_ibuf_I[5].z ),
    .A1(\uio_out_ibuf_I[13].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[5].x ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[6].cell0_I  (.A0(\uio_out_ibuf_I[6].z ),
    .A1(\uio_out_ibuf_I[14].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[6].x ));
 sky130_fd_sc_hd__mux2_2 \uio_out_mux_I[7].cell0_I  (.A0(\uio_out_ibuf_I[7].z ),
    .A1(\uio_out_ibuf_I[15].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uio_out_mux_I[7].x ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[0].genblk1.cell0_I  (.A(\uio_out_mux_I[0].x ),
    .Y(\uio_out_obuf_I[0].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[1].genblk1.cell0_I  (.A(\uio_out_mux_I[1].x ),
    .Y(\uio_out_obuf_I[1].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[2].genblk1.cell0_I  (.A(\uio_out_mux_I[2].x ),
    .Y(\uio_out_obuf_I[2].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[3].genblk1.cell0_I  (.A(\uio_out_mux_I[3].x ),
    .Y(\uio_out_obuf_I[3].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[4].genblk1.cell0_I  (.A(\uio_out_mux_I[4].x ),
    .Y(\uio_out_obuf_I[4].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[5].genblk1.cell0_I  (.A(\uio_out_mux_I[5].x ),
    .Y(\uio_out_obuf_I[5].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[6].genblk1.cell0_I  (.A(\uio_out_mux_I[6].x ),
    .Y(\uio_out_obuf_I[6].z ));
 sky130_fd_sc_hd__bufinv_8 \uio_out_obuf_I[7].genblk1.cell0_I  (.A(\uio_out_mux_I[7].x ),
    .Y(\uio_out_obuf_I[7].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[0].genblk1.cell0_I  (.A(spine_bot_ow[1]),
    .Y(\uo_out_ibuf_I[0].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[10].genblk1.cell0_I  (.A(spine_top_ow[3]),
    .Y(\uo_out_ibuf_I[10].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[11].genblk1.cell0_I  (.A(spine_top_ow[4]),
    .Y(\uo_out_ibuf_I[11].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[12].genblk1.cell0_I  (.A(spine_top_ow[5]),
    .Y(\uo_out_ibuf_I[12].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[13].genblk1.cell0_I  (.A(spine_top_ow[6]),
    .Y(\uo_out_ibuf_I[13].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[14].genblk1.cell0_I  (.A(spine_top_ow[7]),
    .Y(\uo_out_ibuf_I[14].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[15].genblk1.cell0_I  (.A(spine_top_ow[8]),
    .Y(\uo_out_ibuf_I[15].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[1].genblk1.cell0_I  (.A(spine_bot_ow[2]),
    .Y(\uo_out_ibuf_I[1].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[2].genblk1.cell0_I  (.A(spine_bot_ow[3]),
    .Y(\uo_out_ibuf_I[2].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[3].genblk1.cell0_I  (.A(spine_bot_ow[4]),
    .Y(\uo_out_ibuf_I[3].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[4].genblk1.cell0_I  (.A(spine_bot_ow[5]),
    .Y(\uo_out_ibuf_I[4].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[5].genblk1.cell0_I  (.A(spine_bot_ow[6]),
    .Y(\uo_out_ibuf_I[5].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[6].genblk1.cell0_I  (.A(spine_bot_ow[7]),
    .Y(\uo_out_ibuf_I[6].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[7].genblk1.cell0_I  (.A(spine_bot_ow[8]),
    .Y(\uo_out_ibuf_I[7].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[8].genblk1.cell0_I  (.A(spine_top_ow[1]),
    .Y(\uo_out_ibuf_I[8].z ));
 sky130_fd_sc_hd__inv_2 \uo_out_ibuf_I[9].genblk1.cell0_I  (.A(spine_top_ow[2]),
    .Y(\uo_out_ibuf_I[9].z ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[0].cell0_I  (.A0(\uo_out_ibuf_I[0].z ),
    .A1(\uo_out_ibuf_I[8].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[0].x ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[1].cell0_I  (.A0(\uo_out_ibuf_I[1].z ),
    .A1(\uo_out_ibuf_I[9].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[1].x ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[2].cell0_I  (.A0(\uo_out_ibuf_I[2].z ),
    .A1(\uo_out_ibuf_I[10].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[2].x ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[3].cell0_I  (.A0(\uo_out_ibuf_I[3].z ),
    .A1(\uo_out_ibuf_I[11].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[3].x ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[4].cell0_I  (.A0(\uo_out_ibuf_I[4].z ),
    .A1(\uo_out_ibuf_I[12].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[4].x ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[5].cell0_I  (.A0(\uo_out_ibuf_I[5].z ),
    .A1(\uo_out_ibuf_I[13].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[5].x ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[6].cell0_I  (.A0(\uo_out_ibuf_I[6].z ),
    .A1(\uo_out_ibuf_I[14].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[6].x ));
 sky130_fd_sc_hd__mux2_2 \uo_out_mux_I[7].cell0_I  (.A0(\uo_out_ibuf_I[7].z ),
    .A1(\uo_out_ibuf_I[15].z ),
    .S(\side_sel_buf_I.z ),
    .X(\uo_out_mux_I[7].x ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[0].genblk1.cell0_I  (.A(\uo_out_mux_I[0].x ),
    .Y(\uo_out_obuf_I[0].z ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[1].genblk1.cell0_I  (.A(\uo_out_mux_I[1].x ),
    .Y(\uo_out_obuf_I[1].z ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[2].genblk1.cell0_I  (.A(\uo_out_mux_I[2].x ),
    .Y(\uo_out_obuf_I[2].z ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[3].genblk1.cell0_I  (.A(\uo_out_mux_I[3].x ),
    .Y(\uo_out_obuf_I[3].z ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[4].genblk1.cell0_I  (.A(\uo_out_mux_I[4].x ),
    .Y(\uo_out_obuf_I[4].z ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[5].genblk1.cell0_I  (.A(\uo_out_mux_I[5].x ),
    .Y(\uo_out_obuf_I[5].z ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[6].genblk1.cell0_I  (.A(\uo_out_mux_I[6].x ),
    .Y(\uo_out_obuf_I[6].z ));
 sky130_fd_sc_hd__bufinv_8 \uo_out_obuf_I[7].genblk1.cell0_I  (.A(\uo_out_mux_I[7].x ),
    .Y(\uo_out_obuf_I[7].z ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_343 ();
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(spine_bot_ow[21]));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_112 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_381 ();
 assign spine_bot_iw[1] = \genblk2[0].ctrl_ena_buf_I.z ;
 assign spine_bot_iw[11] = \genblk2[0].pad_ui_in_buf_I[0].z ;
 assign spine_bot_iw[12] = \genblk2[0].pad_ui_in_buf_I[1].z ;
 assign spine_bot_iw[13] = \genblk2[0].pad_ui_in_buf_I[2].z ;
 assign spine_bot_iw[14] = \genblk2[0].pad_ui_in_buf_I[3].z ;
 assign spine_bot_iw[15] = \genblk2[0].pad_ui_in_buf_I[4].z ;
 assign spine_bot_iw[16] = \genblk2[0].pad_ui_in_buf_I[5].z ;
 assign spine_bot_iw[17] = \genblk2[0].pad_ui_in_buf_I[6].z ;
 assign spine_bot_iw[18] = \genblk2[0].pad_ui_in_buf_I[7].z ;
 assign spine_bot_iw[19] = \genblk2[0].pad_ui_in_buf_I[8].z ;
 assign spine_bot_iw[20] = \genblk2[0].pad_ui_in_buf_I[9].z ;
 assign spine_bot_iw[21] = \genblk2[0].pad_uio_in_buf_I[0].z ;
 assign spine_bot_iw[22] = \genblk2[0].pad_uio_in_buf_I[1].z ;
 assign spine_bot_iw[23] = \genblk2[0].pad_uio_in_buf_I[2].z ;
 assign spine_bot_iw[24] = \genblk2[0].pad_uio_in_buf_I[3].z ;
 assign spine_bot_iw[25] = \genblk2[0].pad_uio_in_buf_I[4].z ;
 assign spine_bot_iw[26] = \genblk2[0].pad_uio_in_buf_I[5].z ;
 assign spine_bot_iw[27] = \genblk2[0].pad_uio_in_buf_I[6].z ;
 assign spine_bot_iw[28] = \genblk2[0].pad_uio_in_buf_I[7].z ;
 assign spine_bot_iw[2] = \genblk2[0].sel_cnt_buf_I[0].z ;
 assign spine_bot_iw[3] = \genblk2[0].sel_cnt_buf_I[1].z ;
 assign spine_bot_iw[4] = \genblk2[0].sel_cnt_buf_I[2].z ;
 assign spine_bot_iw[5] = \genblk2[0].sel_cnt_buf_I[3].z ;
 assign spine_bot_iw[6] = \genblk2[0].sel_cnt_buf_I[4].z ;
 assign spine_bot_iw[7] = \genblk2[0].sel_cnt_buf_I[5].z ;
 assign spine_bot_iw[8] = \genblk2[0].sel_cnt_buf_I[6].z ;
 assign spine_bot_iw[9] = \genblk2[0].sel_cnt_buf_I[7].z ;
 assign spine_bot_iw[10] = \genblk2[0].sel_cnt_buf_I[8].z ;
 assign spine_bot_iw[0] = \genblk2[0].tie_guard_I[0].lo ;
 assign spine_bot_iw[29] = \genblk2[0].tie_guard_I[1].lo ;
 assign spine_top_iw[1] = \genblk2[1].ctrl_ena_buf_I.z ;
 assign spine_top_iw[11] = \genblk2[1].pad_ui_in_buf_I[0].z ;
 assign spine_top_iw[12] = \genblk2[1].pad_ui_in_buf_I[1].z ;
 assign spine_top_iw[13] = \genblk2[1].pad_ui_in_buf_I[2].z ;
 assign spine_top_iw[14] = \genblk2[1].pad_ui_in_buf_I[3].z ;
 assign spine_top_iw[15] = \genblk2[1].pad_ui_in_buf_I[4].z ;
 assign spine_top_iw[16] = \genblk2[1].pad_ui_in_buf_I[5].z ;
 assign spine_top_iw[17] = \genblk2[1].pad_ui_in_buf_I[6].z ;
 assign spine_top_iw[18] = \genblk2[1].pad_ui_in_buf_I[7].z ;
 assign spine_top_iw[19] = \genblk2[1].pad_ui_in_buf_I[8].z ;
 assign spine_top_iw[20] = \genblk2[1].pad_ui_in_buf_I[9].z ;
 assign spine_top_iw[21] = \genblk2[1].pad_uio_in_buf_I[0].z ;
 assign spine_top_iw[22] = \genblk2[1].pad_uio_in_buf_I[1].z ;
 assign spine_top_iw[23] = \genblk2[1].pad_uio_in_buf_I[2].z ;
 assign spine_top_iw[24] = \genblk2[1].pad_uio_in_buf_I[3].z ;
 assign spine_top_iw[25] = \genblk2[1].pad_uio_in_buf_I[4].z ;
 assign spine_top_iw[26] = \genblk2[1].pad_uio_in_buf_I[5].z ;
 assign spine_top_iw[27] = \genblk2[1].pad_uio_in_buf_I[6].z ;
 assign spine_top_iw[28] = \genblk2[1].pad_uio_in_buf_I[7].z ;
 assign spine_top_iw[2] = \genblk2[1].sel_cnt_buf_I[0].z ;
 assign spine_top_iw[3] = \genblk2[1].sel_cnt_buf_I[1].z ;
 assign spine_top_iw[4] = \genblk2[1].sel_cnt_buf_I[2].z ;
 assign spine_top_iw[5] = \genblk2[1].sel_cnt_buf_I[3].z ;
 assign spine_top_iw[6] = \genblk2[1].sel_cnt_buf_I[4].z ;
 assign spine_top_iw[7] = \genblk2[1].sel_cnt_buf_I[5].z ;
 assign spine_top_iw[8] = \genblk2[1].sel_cnt_buf_I[6].z ;
 assign spine_top_iw[9] = \genblk2[1].sel_cnt_buf_I[7].z ;
 assign spine_top_iw[10] = \genblk2[1].sel_cnt_buf_I[8].z ;
 assign spine_top_iw[0] = \genblk2[1].tie_guard_I[0].lo ;
 assign spine_top_iw[29] = \genblk2[1].tie_guard_I[1].lo ;
 assign pad_uio_oe_n[0] = \uio_oe_obuf_I[0].z ;
 assign pad_uio_oe_n[1] = \uio_oe_obuf_I[1].z ;
 assign pad_uio_oe_n[2] = \uio_oe_obuf_I[2].z ;
 assign pad_uio_oe_n[3] = \uio_oe_obuf_I[3].z ;
 assign pad_uio_oe_n[4] = \uio_oe_obuf_I[4].z ;
 assign pad_uio_oe_n[5] = \uio_oe_obuf_I[5].z ;
 assign pad_uio_oe_n[6] = \uio_oe_obuf_I[6].z ;
 assign pad_uio_oe_n[7] = \uio_oe_obuf_I[7].z ;
 assign pad_uio_out[0] = \uio_out_obuf_I[0].z ;
 assign pad_uio_out[1] = \uio_out_obuf_I[1].z ;
 assign pad_uio_out[2] = \uio_out_obuf_I[2].z ;
 assign pad_uio_out[3] = \uio_out_obuf_I[3].z ;
 assign pad_uio_out[4] = \uio_out_obuf_I[4].z ;
 assign pad_uio_out[5] = \uio_out_obuf_I[5].z ;
 assign pad_uio_out[6] = \uio_out_obuf_I[6].z ;
 assign pad_uio_out[7] = \uio_out_obuf_I[7].z ;
 assign pad_uo_out[0] = \uo_out_obuf_I[0].z ;
 assign pad_uo_out[1] = \uo_out_obuf_I[1].z ;
 assign pad_uo_out[2] = \uo_out_obuf_I[2].z ;
 assign pad_uo_out[3] = \uo_out_obuf_I[3].z ;
 assign pad_uo_out[4] = \uo_out_obuf_I[4].z ;
 assign pad_uo_out[5] = \uo_out_obuf_I[5].z ;
 assign pad_uo_out[6] = \uo_out_obuf_I[6].z ;
 assign pad_uo_out[7] = \uo_out_obuf_I[7].z ;
endmodule
