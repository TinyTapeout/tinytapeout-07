VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mos_bandgap
  CLASS BLOCK ;
  FOREIGN tt_um_mos_bandgap ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.250000 ;
    ANTENNADIFFAREA 4.060000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 115.000000 ;
    ANTENNADIFFAREA 69.352196 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 86.170 73.370 99.050 98.210 ;
      LAYER nwell ;
        RECT 101.170 86.370 113.130 98.210 ;
        RECT 115.170 86.370 127.130 98.210 ;
        RECT 129.170 86.370 141.130 98.210 ;
      LAYER pwell ;
        RECT 105.170 72.370 112.130 84.160 ;
        RECT 118.170 72.370 125.130 84.160 ;
        RECT 143.170 73.370 156.050 98.210 ;
      LAYER nwell ;
        RECT 105.170 58.370 112.130 70.210 ;
        RECT 118.070 59.070 125.030 63.910 ;
        RECT 129.170 58.370 136.130 70.210 ;
      LAYER pwell ;
        RECT 128.420 23.920 130.430 32.620 ;
        RECT 127.870 12.270 130.970 23.100 ;
      LAYER nwell ;
        RECT 132.470 18.320 135.660 33.730 ;
        RECT 138.820 18.320 142.010 33.730 ;
      LAYER pwell ;
        RECT 132.620 15.470 141.820 17.930 ;
      LAYER nwell ;
        RECT 143.420 16.520 146.610 33.990 ;
      LAYER pwell ;
        RECT 139.420 15.420 139.970 15.470 ;
        RECT 131.920 12.320 142.750 15.420 ;
        RECT 147.420 12.320 150.520 30.020 ;
      LAYER li1 ;
        RECT 86.350 97.860 98.870 98.030 ;
        RECT 86.350 73.720 86.520 97.860 ;
        RECT 86.960 74.150 87.740 76.420 ;
        RECT 97.530 74.200 98.220 76.360 ;
        RECT 90.770 73.720 93.770 73.770 ;
        RECT 98.700 73.720 98.870 97.860 ;
        RECT 101.350 97.860 112.950 98.030 ;
        RECT 101.350 96.670 101.520 97.860 ;
        RECT 102.150 97.345 112.150 97.515 ;
        RECT 101.170 87.370 101.570 96.670 ;
        RECT 101.350 86.720 101.520 87.370 ;
        RECT 101.920 87.090 102.090 97.130 ;
        RECT 112.210 87.090 112.380 97.130 ;
        RECT 112.780 86.720 112.950 97.860 ;
        RECT 115.350 97.860 126.950 98.030 ;
        RECT 115.350 96.370 115.520 97.860 ;
        RECT 116.150 97.345 126.150 97.515 ;
        RECT 115.170 87.470 115.670 96.370 ;
        RECT 101.350 86.550 112.950 86.720 ;
        RECT 115.350 86.720 115.520 87.470 ;
        RECT 115.920 87.090 116.090 97.130 ;
        RECT 126.210 87.090 126.380 97.130 ;
        RECT 126.780 86.720 126.950 97.860 ;
        RECT 129.350 97.860 140.950 98.030 ;
        RECT 129.350 96.670 129.520 97.860 ;
        RECT 130.150 97.345 140.150 97.515 ;
        RECT 129.270 87.470 129.670 96.670 ;
        RECT 115.350 86.550 126.950 86.720 ;
        RECT 129.350 86.720 129.520 87.470 ;
        RECT 129.920 87.090 130.090 97.130 ;
        RECT 140.210 87.090 140.380 97.130 ;
        RECT 140.780 86.720 140.950 97.860 ;
        RECT 129.350 86.550 140.950 86.720 ;
        RECT 143.350 97.860 155.870 98.030 ;
        RECT 86.350 73.550 98.870 73.720 ;
        RECT 105.350 83.810 111.950 83.980 ;
        RECT 90.770 73.470 93.770 73.550 ;
        RECT 105.350 72.720 105.520 83.810 ;
        RECT 106.150 83.300 111.150 83.470 ;
        RECT 105.920 73.090 106.090 83.130 ;
        RECT 111.210 73.090 111.380 83.130 ;
        RECT 106.170 72.720 111.270 72.770 ;
        RECT 111.780 72.720 111.950 83.810 ;
        RECT 105.350 72.550 111.950 72.720 ;
        RECT 118.350 83.810 124.950 83.980 ;
        RECT 118.350 72.720 118.520 83.810 ;
        RECT 119.150 83.300 124.150 83.470 ;
        RECT 118.920 73.090 119.090 83.130 ;
        RECT 124.210 73.090 124.380 83.130 ;
        RECT 124.780 72.770 124.950 83.810 ;
        RECT 143.350 73.720 143.520 97.860 ;
        RECT 144.000 74.200 144.690 76.360 ;
        RECT 154.530 74.200 155.220 76.360 ;
        RECT 148.270 73.720 150.970 73.870 ;
        RECT 155.700 73.720 155.870 97.860 ;
        RECT 143.350 73.550 155.870 73.720 ;
        RECT 148.270 73.370 150.970 73.550 ;
        RECT 120.170 72.720 124.950 72.770 ;
        RECT 118.350 72.550 124.950 72.720 ;
        RECT 106.170 72.470 111.270 72.550 ;
        RECT 120.170 72.370 124.870 72.550 ;
        RECT 106.970 70.030 110.870 70.370 ;
        RECT 130.570 70.030 133.570 70.070 ;
        RECT 105.350 69.860 111.950 70.030 ;
        RECT 105.350 58.720 105.520 69.860 ;
        RECT 106.970 69.770 110.870 69.860 ;
        RECT 105.920 59.450 106.090 69.490 ;
        RECT 111.210 59.450 111.380 69.490 ;
        RECT 106.150 59.065 111.150 59.235 ;
        RECT 111.780 58.720 111.950 69.860 ;
        RECT 129.350 69.860 135.950 70.030 ;
        RECT 120.170 63.730 122.770 63.870 ;
        RECT 118.250 63.560 124.850 63.730 ;
        RECT 118.250 59.420 118.420 63.560 ;
        RECT 120.170 63.470 122.770 63.560 ;
        RECT 118.820 60.150 118.990 63.190 ;
        RECT 124.110 60.150 124.280 63.190 ;
        RECT 119.050 59.765 124.050 59.935 ;
        RECT 124.680 59.420 124.850 63.560 ;
        RECT 118.250 59.250 124.850 59.420 ;
        RECT 105.350 58.550 111.950 58.720 ;
        RECT 129.350 58.720 129.520 69.860 ;
        RECT 130.570 69.770 133.570 69.860 ;
        RECT 129.920 59.450 130.090 69.490 ;
        RECT 135.210 59.450 135.380 69.490 ;
        RECT 130.150 59.065 135.150 59.235 ;
        RECT 135.780 58.720 135.950 69.860 ;
        RECT 129.350 58.550 135.950 58.720 ;
        RECT 143.600 33.640 146.430 33.810 ;
        RECT 132.650 33.380 135.480 33.550 ;
        RECT 132.650 33.020 132.820 33.380 ;
        RECT 128.600 32.320 130.250 32.440 ;
        RECT 126.770 32.270 130.250 32.320 ;
        RECT 126.770 24.270 128.770 32.270 ;
        RECT 129.250 29.630 129.600 31.790 ;
        RECT 129.250 24.750 129.600 26.910 ;
        RECT 130.080 24.270 130.250 32.270 ;
        RECT 126.770 24.100 130.250 24.270 ;
        RECT 126.770 22.920 129.920 24.100 ;
        RECT 126.770 22.750 130.790 22.920 ;
        RECT 126.770 12.620 128.220 22.750 ;
        RECT 128.900 22.180 129.940 22.350 ;
        RECT 128.560 20.120 128.730 22.120 ;
        RECT 130.110 20.120 130.280 22.120 ;
        RECT 128.900 19.890 129.940 20.060 ;
        RECT 128.560 17.830 128.730 19.830 ;
        RECT 130.110 17.830 130.280 19.830 ;
        RECT 128.900 17.600 129.940 17.770 ;
        RECT 128.560 15.540 128.730 17.540 ;
        RECT 130.110 15.540 130.280 17.540 ;
        RECT 128.900 15.310 129.940 15.480 ;
        RECT 128.560 13.250 128.730 15.250 ;
        RECT 130.110 13.250 130.280 15.250 ;
        RECT 130.620 14.920 130.790 22.750 ;
        RECT 132.520 21.120 132.820 33.020 ;
        RECT 133.545 32.810 134.585 32.980 ;
        RECT 133.160 30.750 133.330 32.750 ;
        RECT 134.800 30.750 134.970 32.750 ;
        RECT 133.545 30.520 134.585 30.690 ;
        RECT 133.160 28.460 133.330 30.460 ;
        RECT 134.800 28.460 134.970 30.460 ;
        RECT 133.545 28.230 134.585 28.400 ;
        RECT 133.160 26.170 133.330 28.170 ;
        RECT 134.800 26.170 134.970 28.170 ;
        RECT 133.545 25.940 134.585 26.110 ;
        RECT 133.160 23.880 133.330 25.880 ;
        RECT 134.800 23.880 134.970 25.880 ;
        RECT 133.545 23.650 134.585 23.820 ;
        RECT 133.160 21.590 133.330 23.590 ;
        RECT 134.800 21.590 134.970 23.590 ;
        RECT 133.545 21.360 134.585 21.530 ;
        RECT 132.650 18.670 132.820 21.120 ;
        RECT 133.160 19.300 133.330 21.300 ;
        RECT 134.800 19.300 134.970 21.300 ;
        RECT 133.545 19.070 134.585 19.240 ;
        RECT 135.310 18.670 135.480 33.380 ;
        RECT 132.650 18.500 135.480 18.670 ;
        RECT 139.000 33.380 141.830 33.550 ;
        RECT 139.000 18.670 139.170 33.380 ;
        RECT 141.660 33.020 141.830 33.380 ;
        RECT 143.600 33.270 143.770 33.640 ;
        RECT 139.895 32.810 140.935 32.980 ;
        RECT 139.510 30.750 139.680 32.750 ;
        RECT 141.150 30.750 141.320 32.750 ;
        RECT 139.895 30.520 140.935 30.690 ;
        RECT 139.510 28.460 139.680 30.460 ;
        RECT 141.150 28.460 141.320 30.460 ;
        RECT 139.895 28.230 140.935 28.400 ;
        RECT 139.510 26.170 139.680 28.170 ;
        RECT 141.150 26.170 141.320 28.170 ;
        RECT 139.895 25.940 140.935 26.110 ;
        RECT 139.510 23.880 139.680 25.880 ;
        RECT 141.150 23.880 141.320 25.880 ;
        RECT 139.895 23.650 140.935 23.820 ;
        RECT 139.510 21.590 139.680 23.590 ;
        RECT 141.150 21.590 141.320 23.590 ;
        RECT 139.895 21.360 140.935 21.530 ;
        RECT 139.510 19.300 139.680 21.300 ;
        RECT 141.150 19.300 141.320 21.300 ;
        RECT 141.660 21.120 141.970 33.020 ;
        RECT 139.895 19.070 140.935 19.240 ;
        RECT 141.660 18.670 141.830 21.120 ;
        RECT 139.000 18.500 141.830 18.670 ;
        RECT 132.800 17.580 137.040 17.750 ;
        RECT 132.800 15.820 132.970 17.580 ;
        RECT 133.650 17.010 136.190 17.180 ;
        RECT 133.310 16.450 133.480 16.950 ;
        RECT 136.360 16.450 136.530 16.950 ;
        RECT 133.650 16.220 136.190 16.390 ;
        RECT 136.870 15.820 137.040 17.580 ;
        RECT 132.800 15.650 137.040 15.820 ;
        RECT 137.400 17.580 141.640 17.750 ;
        RECT 143.570 17.720 143.770 33.270 ;
        RECT 144.495 33.070 145.535 33.240 ;
        RECT 144.110 32.510 144.280 33.010 ;
        RECT 145.750 32.510 145.920 33.010 ;
        RECT 144.495 32.280 145.535 32.450 ;
        RECT 144.110 31.720 144.280 32.220 ;
        RECT 145.750 31.720 145.920 32.220 ;
        RECT 144.495 31.490 145.535 31.660 ;
        RECT 144.110 30.930 144.280 31.430 ;
        RECT 145.750 30.930 145.920 31.430 ;
        RECT 144.495 30.700 145.535 30.870 ;
        RECT 144.110 30.140 144.280 30.640 ;
        RECT 145.750 30.140 145.920 30.640 ;
        RECT 144.495 29.910 145.535 30.080 ;
        RECT 144.110 29.350 144.280 29.850 ;
        RECT 145.750 29.350 145.920 29.850 ;
        RECT 144.495 29.120 145.535 29.290 ;
        RECT 144.110 28.560 144.280 29.060 ;
        RECT 145.750 28.560 145.920 29.060 ;
        RECT 144.495 28.330 145.535 28.500 ;
        RECT 144.110 27.770 144.280 28.270 ;
        RECT 145.750 27.770 145.920 28.270 ;
        RECT 144.495 27.540 145.535 27.710 ;
        RECT 144.110 26.980 144.280 27.480 ;
        RECT 145.750 26.980 145.920 27.480 ;
        RECT 144.495 26.750 145.535 26.920 ;
        RECT 144.110 26.190 144.280 26.690 ;
        RECT 145.750 26.190 145.920 26.690 ;
        RECT 144.495 25.960 145.535 26.130 ;
        RECT 144.110 25.400 144.280 25.900 ;
        RECT 145.750 25.400 145.920 25.900 ;
        RECT 144.495 25.170 145.535 25.340 ;
        RECT 144.110 24.610 144.280 25.110 ;
        RECT 145.750 24.610 145.920 25.110 ;
        RECT 144.495 24.380 145.535 24.550 ;
        RECT 144.110 23.820 144.280 24.320 ;
        RECT 145.750 23.820 145.920 24.320 ;
        RECT 144.495 23.590 145.535 23.760 ;
        RECT 144.110 23.030 144.280 23.530 ;
        RECT 145.750 23.030 145.920 23.530 ;
        RECT 144.495 22.800 145.535 22.970 ;
        RECT 144.110 22.240 144.280 22.740 ;
        RECT 145.750 22.240 145.920 22.740 ;
        RECT 144.495 22.010 145.535 22.180 ;
        RECT 144.110 21.450 144.280 21.950 ;
        RECT 145.750 21.450 145.920 21.950 ;
        RECT 144.495 21.220 145.535 21.390 ;
        RECT 144.110 20.660 144.280 21.160 ;
        RECT 145.750 20.660 145.920 21.160 ;
        RECT 144.495 20.430 145.535 20.600 ;
        RECT 144.110 19.870 144.280 20.370 ;
        RECT 145.750 19.870 145.920 20.370 ;
        RECT 144.495 19.640 145.535 19.810 ;
        RECT 144.110 19.080 144.280 19.580 ;
        RECT 145.750 19.080 145.920 19.580 ;
        RECT 144.495 18.850 145.535 19.020 ;
        RECT 144.110 18.290 144.280 18.790 ;
        RECT 145.750 18.290 145.920 18.790 ;
        RECT 144.495 18.060 145.535 18.230 ;
        RECT 137.400 15.820 137.570 17.580 ;
        RECT 138.250 17.010 140.790 17.180 ;
        RECT 137.910 16.450 138.080 16.950 ;
        RECT 140.960 16.450 141.130 16.950 ;
        RECT 138.250 16.220 140.790 16.390 ;
        RECT 141.470 15.820 141.640 17.580 ;
        RECT 143.600 16.870 143.770 17.720 ;
        RECT 144.110 17.500 144.280 18.000 ;
        RECT 145.750 17.500 145.920 18.000 ;
        RECT 144.495 17.270 145.535 17.440 ;
        RECT 146.260 16.870 146.430 33.640 ;
        RECT 143.600 16.700 146.430 16.870 ;
        RECT 147.600 29.670 150.340 29.840 ;
        RECT 137.400 15.650 141.770 15.820 ;
        RECT 132.820 15.620 133.620 15.650 ;
        RECT 140.970 15.620 141.770 15.650 ;
        RECT 132.100 15.170 142.570 15.240 ;
        RECT 147.600 15.170 147.770 29.670 ;
        RECT 148.450 29.100 149.490 29.270 ;
        RECT 148.110 27.040 148.280 29.040 ;
        RECT 149.660 27.040 149.830 29.040 ;
        RECT 148.450 26.810 149.490 26.980 ;
        RECT 150.170 26.970 150.340 29.670 ;
        RECT 148.110 24.750 148.280 26.750 ;
        RECT 149.660 24.750 149.830 26.750 ;
        RECT 148.450 24.520 149.490 24.690 ;
        RECT 148.110 22.460 148.280 24.460 ;
        RECT 149.660 22.460 149.830 24.460 ;
        RECT 148.450 22.230 149.490 22.400 ;
        RECT 148.110 20.170 148.280 22.170 ;
        RECT 149.660 20.170 149.830 22.170 ;
        RECT 148.450 19.940 149.490 20.110 ;
        RECT 148.110 17.880 148.280 19.880 ;
        RECT 149.660 17.880 149.830 19.880 ;
        RECT 148.450 17.650 149.490 17.820 ;
        RECT 148.110 15.590 148.280 17.590 ;
        RECT 149.660 15.590 149.830 17.590 ;
        RECT 148.450 15.360 149.490 15.530 ;
        RECT 132.100 15.070 147.770 15.170 ;
        RECT 132.100 14.920 132.270 15.070 ;
        RECT 128.900 13.020 129.940 13.190 ;
        RECT 130.620 12.670 132.270 14.920 ;
        RECT 132.900 14.560 134.900 14.730 ;
        RECT 135.190 14.560 137.190 14.730 ;
        RECT 137.480 14.560 139.480 14.730 ;
        RECT 139.770 14.560 141.770 14.730 ;
        RECT 142.400 14.570 147.770 15.070 ;
        RECT 132.670 13.350 132.840 14.390 ;
        RECT 134.960 13.350 135.130 14.390 ;
        RECT 137.250 13.350 137.420 14.390 ;
        RECT 139.540 13.350 139.710 14.390 ;
        RECT 141.830 13.350 142.000 14.390 ;
        RECT 132.900 13.010 134.900 13.180 ;
        RECT 135.190 13.010 137.190 13.180 ;
        RECT 137.480 13.010 139.480 13.180 ;
        RECT 139.770 13.010 141.770 13.180 ;
        RECT 142.370 12.970 147.770 14.570 ;
        RECT 148.110 13.300 148.280 15.300 ;
        RECT 149.660 13.300 149.830 15.300 ;
        RECT 148.450 13.070 149.490 13.240 ;
        RECT 142.400 12.670 147.770 12.970 ;
        RECT 150.170 12.670 150.920 26.970 ;
        RECT 128.470 12.620 130.370 12.670 ;
        RECT 130.620 12.620 150.920 12.670 ;
        RECT 126.770 10.420 150.920 12.620 ;
      LAYER mcon ;
        RECT 97.570 74.270 98.170 76.270 ;
        RECT 102.230 97.345 112.070 97.515 ;
        RECT 101.170 87.370 101.570 96.670 ;
        RECT 101.920 87.170 102.090 97.050 ;
        RECT 112.210 87.170 112.380 97.050 ;
        RECT 116.230 97.345 126.070 97.515 ;
        RECT 115.170 87.470 115.670 96.370 ;
        RECT 115.920 87.170 116.090 97.050 ;
        RECT 126.210 87.170 126.380 97.050 ;
        RECT 130.230 97.345 140.070 97.515 ;
        RECT 129.270 87.470 129.670 96.670 ;
        RECT 129.920 87.170 130.090 97.050 ;
        RECT 140.210 87.170 140.380 97.050 ;
        RECT 106.230 83.300 111.070 83.470 ;
        RECT 105.920 73.170 106.090 83.050 ;
        RECT 111.210 73.170 111.380 83.050 ;
        RECT 119.230 83.300 124.070 83.470 ;
        RECT 118.920 73.170 119.090 83.050 ;
        RECT 124.210 73.170 124.380 83.050 ;
        RECT 144.070 74.270 144.570 76.270 ;
        RECT 154.570 74.270 155.170 76.270 ;
        RECT 105.920 59.530 106.090 69.410 ;
        RECT 111.210 59.530 111.380 69.410 ;
        RECT 106.230 59.065 111.070 59.235 ;
        RECT 118.820 60.230 118.990 63.110 ;
        RECT 124.110 60.230 124.280 63.110 ;
        RECT 119.130 59.765 123.970 59.935 ;
        RECT 129.920 59.530 130.090 69.410 ;
        RECT 135.210 59.530 135.380 69.410 ;
        RECT 130.230 59.065 135.070 59.235 ;
        RECT 127.270 28.020 128.120 31.720 ;
        RECT 128.520 24.720 128.770 31.870 ;
        RECT 129.330 29.715 129.520 31.700 ;
        RECT 129.330 24.840 129.520 26.825 ;
        RECT 127.970 13.470 128.220 22.820 ;
        RECT 128.980 22.180 129.860 22.350 ;
        RECT 128.560 20.200 128.730 22.040 ;
        RECT 130.110 20.200 130.280 22.040 ;
        RECT 128.980 19.890 129.860 20.060 ;
        RECT 128.560 17.910 128.730 19.750 ;
        RECT 130.110 17.910 130.280 19.750 ;
        RECT 128.980 17.600 129.860 17.770 ;
        RECT 128.560 15.620 128.730 17.460 ;
        RECT 130.110 15.620 130.280 17.460 ;
        RECT 128.980 15.310 129.860 15.480 ;
        RECT 128.560 13.330 128.730 15.170 ;
        RECT 130.110 13.330 130.280 15.170 ;
        RECT 132.520 21.120 132.820 33.020 ;
        RECT 133.625 32.810 134.505 32.980 ;
        RECT 133.160 30.830 133.330 32.670 ;
        RECT 134.800 30.830 134.970 32.670 ;
        RECT 133.625 30.520 134.505 30.690 ;
        RECT 133.160 28.540 133.330 30.380 ;
        RECT 134.800 28.540 134.970 30.380 ;
        RECT 133.625 28.230 134.505 28.400 ;
        RECT 133.160 26.250 133.330 28.090 ;
        RECT 134.800 26.250 134.970 28.090 ;
        RECT 133.625 25.940 134.505 26.110 ;
        RECT 133.160 23.960 133.330 25.800 ;
        RECT 134.800 23.960 134.970 25.800 ;
        RECT 133.625 23.650 134.505 23.820 ;
        RECT 133.160 21.670 133.330 23.510 ;
        RECT 134.800 21.670 134.970 23.510 ;
        RECT 133.625 21.360 134.505 21.530 ;
        RECT 133.160 19.380 133.330 21.220 ;
        RECT 134.800 19.380 134.970 21.220 ;
        RECT 133.625 19.070 134.505 19.240 ;
        RECT 139.975 32.810 140.855 32.980 ;
        RECT 139.510 30.830 139.680 32.670 ;
        RECT 141.150 30.830 141.320 32.670 ;
        RECT 139.975 30.520 140.855 30.690 ;
        RECT 139.510 28.540 139.680 30.380 ;
        RECT 141.150 28.540 141.320 30.380 ;
        RECT 139.975 28.230 140.855 28.400 ;
        RECT 139.510 26.250 139.680 28.090 ;
        RECT 141.150 26.250 141.320 28.090 ;
        RECT 139.975 25.940 140.855 26.110 ;
        RECT 139.510 23.960 139.680 25.800 ;
        RECT 141.150 23.960 141.320 25.800 ;
        RECT 139.975 23.650 140.855 23.820 ;
        RECT 139.510 21.670 139.680 23.510 ;
        RECT 141.150 21.670 141.320 23.510 ;
        RECT 139.975 21.360 140.855 21.530 ;
        RECT 139.510 19.380 139.680 21.220 ;
        RECT 141.150 19.380 141.320 21.220 ;
        RECT 141.670 21.120 141.970 33.020 ;
        RECT 139.975 19.070 140.855 19.240 ;
        RECT 133.730 17.010 136.110 17.180 ;
        RECT 133.310 16.530 133.480 16.870 ;
        RECT 136.360 16.530 136.530 16.870 ;
        RECT 133.730 16.220 136.110 16.390 ;
        RECT 143.570 17.720 143.770 33.270 ;
        RECT 144.575 33.070 145.455 33.240 ;
        RECT 144.110 32.590 144.280 32.930 ;
        RECT 145.750 32.590 145.920 32.930 ;
        RECT 144.575 32.280 145.455 32.450 ;
        RECT 144.110 31.800 144.280 32.140 ;
        RECT 145.750 31.800 145.920 32.140 ;
        RECT 144.575 31.490 145.455 31.660 ;
        RECT 144.110 31.010 144.280 31.350 ;
        RECT 145.750 31.010 145.920 31.350 ;
        RECT 144.575 30.700 145.455 30.870 ;
        RECT 144.110 30.220 144.280 30.560 ;
        RECT 145.750 30.220 145.920 30.560 ;
        RECT 144.575 29.910 145.455 30.080 ;
        RECT 144.110 29.430 144.280 29.770 ;
        RECT 145.750 29.430 145.920 29.770 ;
        RECT 144.575 29.120 145.455 29.290 ;
        RECT 144.110 28.640 144.280 28.980 ;
        RECT 145.750 28.640 145.920 28.980 ;
        RECT 144.575 28.330 145.455 28.500 ;
        RECT 144.110 27.850 144.280 28.190 ;
        RECT 145.750 27.850 145.920 28.190 ;
        RECT 144.575 27.540 145.455 27.710 ;
        RECT 144.110 27.060 144.280 27.400 ;
        RECT 145.750 27.060 145.920 27.400 ;
        RECT 144.575 26.750 145.455 26.920 ;
        RECT 144.110 26.270 144.280 26.610 ;
        RECT 145.750 26.270 145.920 26.610 ;
        RECT 144.575 25.960 145.455 26.130 ;
        RECT 144.110 25.480 144.280 25.820 ;
        RECT 145.750 25.480 145.920 25.820 ;
        RECT 144.575 25.170 145.455 25.340 ;
        RECT 144.110 24.690 144.280 25.030 ;
        RECT 145.750 24.690 145.920 25.030 ;
        RECT 144.575 24.380 145.455 24.550 ;
        RECT 144.110 23.900 144.280 24.240 ;
        RECT 145.750 23.900 145.920 24.240 ;
        RECT 144.575 23.590 145.455 23.760 ;
        RECT 144.110 23.110 144.280 23.450 ;
        RECT 145.750 23.110 145.920 23.450 ;
        RECT 144.575 22.800 145.455 22.970 ;
        RECT 144.110 22.320 144.280 22.660 ;
        RECT 145.750 22.320 145.920 22.660 ;
        RECT 144.575 22.010 145.455 22.180 ;
        RECT 144.110 21.530 144.280 21.870 ;
        RECT 145.750 21.530 145.920 21.870 ;
        RECT 144.575 21.220 145.455 21.390 ;
        RECT 144.110 20.740 144.280 21.080 ;
        RECT 145.750 20.740 145.920 21.080 ;
        RECT 144.575 20.430 145.455 20.600 ;
        RECT 144.110 19.950 144.280 20.290 ;
        RECT 145.750 19.950 145.920 20.290 ;
        RECT 144.575 19.640 145.455 19.810 ;
        RECT 144.110 19.160 144.280 19.500 ;
        RECT 145.750 19.160 145.920 19.500 ;
        RECT 144.575 18.850 145.455 19.020 ;
        RECT 144.110 18.370 144.280 18.710 ;
        RECT 145.750 18.370 145.920 18.710 ;
        RECT 144.575 18.060 145.455 18.230 ;
        RECT 138.330 17.010 140.710 17.180 ;
        RECT 137.910 16.530 138.080 16.870 ;
        RECT 140.960 16.530 141.130 16.870 ;
        RECT 138.330 16.220 140.710 16.390 ;
        RECT 144.110 17.580 144.280 17.920 ;
        RECT 145.750 17.580 145.920 17.920 ;
        RECT 144.575 17.270 145.455 17.440 ;
        RECT 148.530 29.100 149.410 29.270 ;
        RECT 148.110 27.120 148.280 28.960 ;
        RECT 149.660 27.120 149.830 28.960 ;
        RECT 148.530 26.810 149.410 26.980 ;
        RECT 148.110 24.830 148.280 26.670 ;
        RECT 149.660 24.830 149.830 26.670 ;
        RECT 148.530 24.520 149.410 24.690 ;
        RECT 148.110 22.540 148.280 24.380 ;
        RECT 149.660 22.540 149.830 24.380 ;
        RECT 148.530 22.230 149.410 22.400 ;
        RECT 148.110 20.250 148.280 22.090 ;
        RECT 149.660 20.250 149.830 22.090 ;
        RECT 148.530 19.940 149.410 20.110 ;
        RECT 148.110 17.960 148.280 19.800 ;
        RECT 149.660 17.960 149.830 19.800 ;
        RECT 148.530 17.650 149.410 17.820 ;
        RECT 148.110 15.670 148.280 17.510 ;
        RECT 149.660 15.670 149.830 17.510 ;
        RECT 148.530 15.360 149.410 15.530 ;
        RECT 128.980 13.020 129.860 13.190 ;
        RECT 132.980 14.560 134.820 14.730 ;
        RECT 135.270 14.560 137.110 14.730 ;
        RECT 137.560 14.560 139.400 14.730 ;
        RECT 139.850 14.560 141.690 14.730 ;
        RECT 132.670 13.430 132.840 14.310 ;
        RECT 134.960 13.430 135.130 14.310 ;
        RECT 137.250 13.430 137.420 14.310 ;
        RECT 139.540 13.430 139.710 14.310 ;
        RECT 141.830 13.430 142.000 14.310 ;
        RECT 132.980 13.010 134.820 13.180 ;
        RECT 135.270 13.010 137.110 13.180 ;
        RECT 137.560 13.010 139.400 13.180 ;
        RECT 139.850 13.010 141.690 13.180 ;
        RECT 147.520 12.970 147.770 14.120 ;
        RECT 148.110 13.380 148.280 15.220 ;
        RECT 149.660 13.380 149.830 15.220 ;
        RECT 148.530 13.070 149.410 13.240 ;
        RECT 150.170 12.970 150.420 14.120 ;
        RECT 128.470 12.370 130.370 12.670 ;
        RECT 132.570 12.420 142.120 12.670 ;
        RECT 147.870 12.470 150.070 12.670 ;
        RECT 130.070 10.720 149.020 11.270 ;
      LAYER met1 ;
        RECT 79.330 105.150 80.830 105.180 ;
        RECT 86.170 105.150 155.170 106.370 ;
        RECT 79.330 103.650 155.170 105.150 ;
        RECT 79.330 103.620 80.830 103.650 ;
        RECT 86.170 101.370 155.170 103.650 ;
        RECT 100.470 96.870 101.170 101.370 ;
        RECT 102.270 97.545 113.770 98.870 ;
        RECT 102.170 97.315 113.770 97.545 ;
        RECT 102.270 97.270 113.770 97.315 ;
        RECT 101.890 96.870 102.120 97.110 ;
        RECT 100.470 87.270 102.170 96.870 ;
        RECT 101.890 87.110 102.120 87.270 ;
        RECT 112.170 87.170 113.770 97.270 ;
        RECT 114.470 96.870 115.170 101.370 ;
        RECT 116.270 97.545 126.170 98.870 ;
        RECT 116.170 97.315 126.170 97.545 ;
        RECT 116.270 97.270 126.170 97.315 ;
        RECT 115.890 96.870 116.120 97.110 ;
        RECT 126.180 97.070 126.410 97.110 ;
        RECT 114.470 87.270 116.170 96.870 ;
        RECT 112.180 87.110 112.410 87.170 ;
        RECT 106.270 83.500 111.070 85.070 ;
        RECT 106.170 83.270 111.130 83.500 ;
        RECT 105.890 83.070 106.120 83.110 ;
        RECT 111.180 83.070 111.410 83.110 ;
        RECT 113.070 83.070 113.770 87.170 ;
        RECT 115.890 87.110 116.120 87.270 ;
        RECT 126.170 87.170 127.570 97.070 ;
        RECT 128.470 96.870 129.170 101.370 ;
        RECT 130.270 97.545 140.170 98.870 ;
        RECT 130.170 97.315 140.170 97.545 ;
        RECT 130.270 97.270 140.170 97.315 ;
        RECT 129.890 96.870 130.120 97.110 ;
        RECT 140.180 96.970 140.410 97.110 ;
        RECT 128.470 87.270 130.170 96.870 ;
        RECT 126.180 87.110 126.410 87.170 ;
        RECT 126.870 85.070 127.570 87.170 ;
        RECT 129.890 87.110 130.120 87.270 ;
        RECT 140.170 87.170 142.570 96.970 ;
        RECT 140.180 87.110 140.410 87.170 ;
        RECT 119.270 83.500 127.570 85.070 ;
        RECT 119.170 83.470 127.570 83.500 ;
        RECT 119.170 83.270 125.470 83.470 ;
        RECT 86.870 69.070 87.870 76.570 ;
        RECT 103.770 76.370 106.120 83.070 ;
        RECT 97.470 74.170 106.120 76.370 ;
        RECT 90.620 73.370 93.920 73.870 ;
        RECT 103.770 73.170 106.120 74.170 ;
        RECT 111.170 82.370 113.770 83.070 ;
        RECT 111.170 73.170 112.470 82.370 ;
        RECT 118.890 82.170 119.120 83.110 ;
        RECT 105.890 73.110 106.120 73.170 ;
        RECT 111.180 73.110 111.410 73.170 ;
        RECT 106.070 72.170 111.570 72.870 ;
        RECT 106.070 71.570 112.570 72.170 ;
        RECT 106.820 69.670 111.020 70.470 ;
        RECT 111.970 69.470 112.570 71.570 ;
        RECT 105.890 69.070 106.120 69.470 ;
        RECT 86.870 65.870 106.170 69.070 ;
        RECT 104.770 59.770 106.170 65.870 ;
        RECT 105.890 59.470 106.120 59.770 ;
        RECT 111.170 59.270 112.570 69.470 ;
        RECT 118.570 63.870 119.175 82.170 ;
        RECT 124.170 73.170 125.470 83.270 ;
        RECT 141.370 82.670 142.570 87.170 ;
        RECT 136.170 76.370 142.570 82.670 ;
        RECT 136.170 74.270 144.670 76.370 ;
        RECT 141.370 74.170 144.670 74.270 ;
        RECT 141.370 74.070 142.570 74.170 ;
        RECT 148.120 73.170 151.120 74.070 ;
        RECT 124.180 73.110 124.410 73.170 ;
        RECT 120.070 71.770 125.070 72.870 ;
        RECT 118.570 60.170 119.170 63.870 ;
        RECT 120.020 63.370 122.920 63.970 ;
        RECT 124.470 63.170 125.070 71.770 ;
        RECT 130.420 70.100 133.620 70.270 ;
        RECT 130.420 69.740 133.630 70.100 ;
        RECT 130.420 69.570 133.620 69.740 ;
        RECT 123.970 59.970 125.070 63.170 ;
        RECT 119.770 59.965 125.070 59.970 ;
        RECT 119.070 59.735 125.070 59.965 ;
        RECT 119.770 59.270 125.070 59.735 ;
        RECT 128.970 59.270 130.170 69.470 ;
        RECT 135.180 69.170 135.410 69.470 ;
        RECT 154.370 69.170 155.570 76.470 ;
        RECT 135.170 67.270 155.570 69.170 ;
        RECT 135.170 59.470 136.070 67.270 ;
        RECT 106.470 59.265 130.170 59.270 ;
        RECT 130.570 59.265 134.770 59.270 ;
        RECT 106.170 59.035 135.130 59.265 ;
        RECT 106.470 58.170 134.770 59.035 ;
        RECT 106.170 57.470 134.770 58.170 ;
        RECT 106.170 55.370 135.170 57.470 ;
        RECT 86.170 50.370 155.170 55.370 ;
        RECT 110.970 46.050 112.470 46.080 ;
        RECT 112.910 46.050 114.410 50.370 ;
        RECT 110.970 44.550 114.410 46.050 ;
        RECT 110.970 44.520 112.470 44.550 ;
        RECT 104.580 35.350 106.080 35.380 ;
        RECT 104.580 35.250 112.700 35.350 ;
        RECT 126.670 35.250 150.920 35.820 ;
        RECT 104.580 33.850 150.920 35.250 ;
        RECT 104.580 33.820 106.080 33.850 ;
        RECT 111.110 33.750 150.920 33.850 ;
        RECT 126.670 33.470 150.920 33.750 ;
        RECT 126.670 24.570 128.870 32.320 ;
        RECT 129.020 29.570 129.970 33.470 ;
        RECT 129.300 26.870 129.550 26.885 ;
        RECT 126.670 12.720 128.320 24.570 ;
        RECT 129.170 24.370 131.020 26.870 ;
        RECT 128.920 22.120 129.920 22.470 ;
        RECT 128.530 21.670 128.760 22.100 ;
        RECT 130.070 21.670 131.020 24.370 ;
        RECT 128.520 20.520 131.020 21.670 ;
        RECT 131.170 20.970 132.920 33.470 ;
        RECT 133.520 32.770 138.870 33.120 ;
        RECT 139.870 32.770 140.970 33.070 ;
        RECT 133.130 32.370 133.360 32.730 ;
        RECT 134.720 32.720 138.870 32.770 ;
        RECT 134.720 32.370 139.220 32.720 ;
        RECT 139.480 32.370 139.710 32.730 ;
        RECT 141.120 32.370 141.350 32.730 ;
        RECT 133.120 31.570 141.350 32.370 ;
        RECT 133.120 31.170 136.720 31.570 ;
        RECT 133.130 30.770 133.360 31.170 ;
        RECT 134.720 31.120 136.720 31.170 ;
        RECT 134.770 30.770 136.720 31.120 ;
        RECT 133.570 30.720 134.570 30.770 ;
        RECT 133.565 30.490 134.570 30.720 ;
        RECT 133.570 30.470 134.570 30.490 ;
        RECT 134.820 30.440 136.720 30.770 ;
        RECT 133.130 30.020 133.360 30.440 ;
        RECT 134.770 30.020 136.720 30.440 ;
        RECT 133.120 28.770 136.720 30.020 ;
        RECT 133.130 28.480 133.360 28.770 ;
        RECT 134.720 28.470 136.720 28.770 ;
        RECT 133.520 28.170 136.720 28.470 ;
        RECT 133.130 27.870 133.360 28.150 ;
        RECT 134.720 27.870 136.720 28.170 ;
        RECT 133.120 26.670 136.720 27.870 ;
        RECT 133.130 26.190 133.360 26.670 ;
        RECT 133.570 26.140 134.570 26.170 ;
        RECT 133.565 25.910 134.570 26.140 ;
        RECT 133.570 25.870 134.570 25.910 ;
        RECT 133.130 25.570 133.360 25.860 ;
        RECT 134.720 25.570 136.720 26.670 ;
        RECT 133.120 24.370 136.720 25.570 ;
        RECT 133.130 23.900 133.360 24.370 ;
        RECT 134.720 23.870 136.720 24.370 ;
        RECT 133.520 23.620 136.720 23.870 ;
        RECT 133.130 23.170 133.360 23.570 ;
        RECT 134.720 23.170 136.720 23.620 ;
        RECT 133.120 21.970 136.720 23.170 ;
        RECT 133.130 21.610 133.360 21.970 ;
        RECT 133.570 21.560 134.570 21.620 ;
        RECT 133.565 21.330 134.570 21.560 ;
        RECT 133.570 21.320 134.570 21.330 ;
        RECT 133.130 20.920 133.360 21.280 ;
        RECT 134.720 20.920 136.720 21.970 ;
        RECT 128.530 20.140 128.760 20.520 ;
        RECT 130.070 20.120 131.020 20.520 ;
        RECT 128.920 19.820 131.020 20.120 ;
        RECT 128.530 19.420 128.760 19.810 ;
        RECT 130.070 19.420 131.020 19.820 ;
        RECT 133.120 19.720 136.720 20.920 ;
        RECT 128.520 18.270 131.020 19.420 ;
        RECT 133.130 19.320 133.360 19.720 ;
        RECT 134.720 19.270 136.720 19.720 ;
        RECT 133.520 19.070 136.720 19.270 ;
        RECT 137.720 31.170 141.350 31.570 ;
        RECT 137.720 29.970 139.220 31.170 ;
        RECT 139.480 30.770 139.710 31.170 ;
        RECT 141.120 30.770 141.350 31.170 ;
        RECT 139.920 30.720 140.970 30.770 ;
        RECT 139.915 30.490 140.970 30.720 ;
        RECT 139.920 30.470 140.970 30.490 ;
        RECT 139.480 29.970 139.710 30.440 ;
        RECT 141.120 29.970 141.350 30.440 ;
        RECT 137.720 28.770 141.350 29.970 ;
        RECT 137.720 27.870 139.220 28.770 ;
        RECT 139.480 28.480 139.710 28.770 ;
        RECT 141.120 28.480 141.350 28.770 ;
        RECT 139.870 28.170 140.970 28.470 ;
        RECT 139.480 27.870 139.710 28.150 ;
        RECT 141.120 27.870 141.350 28.150 ;
        RECT 137.720 26.670 141.350 27.870 ;
        RECT 137.720 25.570 139.220 26.670 ;
        RECT 139.480 26.190 139.710 26.670 ;
        RECT 141.120 26.190 141.350 26.670 ;
        RECT 139.920 26.140 140.970 26.170 ;
        RECT 139.915 25.910 140.970 26.140 ;
        RECT 139.920 25.870 140.970 25.910 ;
        RECT 139.480 25.570 139.710 25.860 ;
        RECT 141.120 25.570 141.350 25.860 ;
        RECT 137.720 24.370 141.350 25.570 ;
        RECT 137.720 23.170 139.220 24.370 ;
        RECT 139.480 23.900 139.710 24.370 ;
        RECT 141.120 23.900 141.350 24.370 ;
        RECT 139.870 23.570 140.970 23.870 ;
        RECT 139.480 23.170 139.710 23.570 ;
        RECT 141.120 23.170 141.350 23.570 ;
        RECT 137.720 21.970 141.350 23.170 ;
        RECT 137.720 20.920 139.220 21.970 ;
        RECT 139.480 21.610 139.710 21.970 ;
        RECT 139.920 21.560 140.970 21.620 ;
        RECT 141.120 21.610 141.350 21.970 ;
        RECT 139.915 21.330 140.970 21.560 ;
        RECT 139.920 21.320 140.970 21.330 ;
        RECT 139.480 20.920 139.710 21.280 ;
        RECT 141.120 20.920 141.350 21.280 ;
        RECT 141.520 20.970 143.820 33.470 ;
        RECT 144.470 33.020 145.520 33.320 ;
        RECT 137.720 19.720 141.350 20.920 ;
        RECT 137.720 19.070 139.220 19.720 ;
        RECT 139.480 19.320 139.710 19.720 ;
        RECT 141.120 19.320 141.350 19.720 ;
        RECT 140.195 19.270 140.745 19.300 ;
        RECT 133.520 19.020 139.220 19.070 ;
        RECT 128.530 17.850 128.760 18.270 ;
        RECT 128.920 17.520 129.920 17.870 ;
        RECT 128.530 17.120 128.760 17.520 ;
        RECT 130.070 17.120 131.020 18.270 ;
        RECT 134.720 18.120 139.220 19.020 ;
        RECT 139.870 18.970 140.970 19.270 ;
        RECT 139.970 18.720 140.920 18.970 ;
        RECT 140.195 18.690 140.745 18.720 ;
        RECT 134.720 17.320 137.070 18.120 ;
        RECT 139.920 17.620 140.920 18.020 ;
        RECT 133.820 17.210 137.070 17.320 ;
        RECT 138.370 17.370 140.920 17.620 ;
        RECT 138.370 17.210 140.770 17.370 ;
        RECT 141.970 17.320 143.820 20.970 ;
        RECT 143.970 20.220 144.320 33.020 ;
        RECT 145.720 32.530 145.950 32.990 ;
        RECT 144.520 32.480 145.570 32.520 ;
        RECT 144.515 32.250 145.570 32.480 ;
        RECT 144.520 32.220 145.570 32.250 ;
        RECT 145.720 31.740 145.950 32.200 ;
        RECT 144.470 31.420 145.520 31.720 ;
        RECT 145.720 30.950 145.950 31.410 ;
        RECT 144.520 30.900 145.570 30.920 ;
        RECT 144.515 30.670 145.570 30.900 ;
        RECT 144.520 30.620 145.570 30.670 ;
        RECT 144.470 29.870 145.520 30.170 ;
        RECT 145.720 30.160 145.950 30.620 ;
        RECT 145.720 29.370 145.950 29.830 ;
        RECT 146.320 29.370 150.920 32.570 ;
        RECT 144.520 29.320 145.570 29.370 ;
        RECT 144.515 29.090 145.570 29.320 ;
        RECT 144.520 29.070 145.570 29.090 ;
        RECT 146.320 29.320 149.670 29.370 ;
        RECT 145.720 28.580 145.950 29.040 ;
        RECT 144.470 28.270 145.520 28.570 ;
        RECT 145.720 27.790 145.950 28.250 ;
        RECT 144.520 27.740 145.570 27.770 ;
        RECT 144.515 27.510 145.570 27.740 ;
        RECT 144.520 27.470 145.570 27.510 ;
        RECT 145.720 27.000 145.950 27.460 ;
        RECT 144.470 26.670 145.520 26.970 ;
        RECT 145.720 26.210 145.950 26.670 ;
        RECT 144.520 26.160 145.570 26.170 ;
        RECT 144.515 25.930 145.570 26.160 ;
        RECT 144.520 25.870 145.570 25.930 ;
        RECT 145.720 25.420 145.950 25.880 ;
        RECT 144.470 25.120 145.520 25.420 ;
        RECT 145.720 24.630 145.950 25.090 ;
        RECT 144.520 24.580 145.570 24.620 ;
        RECT 144.515 24.350 145.570 24.580 ;
        RECT 144.520 24.320 145.570 24.350 ;
        RECT 145.720 23.840 145.950 24.300 ;
        RECT 144.470 23.520 145.520 23.820 ;
        RECT 144.520 23.000 145.570 23.070 ;
        RECT 145.720 23.050 145.950 23.510 ;
        RECT 144.515 22.770 145.570 23.000 ;
        RECT 144.470 21.970 145.520 22.270 ;
        RECT 145.720 22.260 145.950 22.720 ;
        RECT 145.720 21.470 145.950 21.930 ;
        RECT 144.520 21.420 145.570 21.470 ;
        RECT 144.515 21.190 145.570 21.420 ;
        RECT 144.520 21.170 145.570 21.190 ;
        RECT 145.720 20.680 145.950 21.140 ;
        RECT 144.470 20.370 145.520 20.670 ;
        RECT 143.970 19.320 144.370 20.220 ;
        RECT 145.720 19.890 145.950 20.350 ;
        RECT 144.520 19.840 145.570 19.870 ;
        RECT 144.515 19.610 145.570 19.840 ;
        RECT 144.520 19.570 145.570 19.610 ;
        RECT 143.970 17.470 144.320 19.320 ;
        RECT 145.720 19.100 145.950 19.560 ;
        RECT 144.470 18.770 145.520 19.070 ;
        RECT 144.520 18.260 145.570 18.320 ;
        RECT 145.720 18.310 145.950 18.770 ;
        RECT 144.515 18.030 145.570 18.260 ;
        RECT 144.520 18.020 145.570 18.030 ;
        RECT 145.720 17.520 145.950 17.980 ;
        RECT 144.470 17.220 145.520 17.520 ;
        RECT 128.520 15.970 131.020 17.120 ;
        RECT 131.820 16.780 132.820 17.170 ;
        RECT 133.670 17.070 137.070 17.210 ;
        RECT 133.670 16.980 136.170 17.070 ;
        RECT 138.270 16.980 140.770 17.210 ;
        RECT 133.820 16.970 136.120 16.980 ;
        RECT 133.280 16.870 133.510 16.930 ;
        RECT 136.330 16.870 136.560 16.930 ;
        RECT 137.880 16.870 138.110 16.930 ;
        RECT 140.930 16.870 141.160 16.930 ;
        RECT 133.170 16.780 133.570 16.870 ;
        RECT 136.270 16.780 136.670 16.870 ;
        RECT 131.820 16.565 136.670 16.780 ;
        RECT 131.820 16.170 132.820 16.565 ;
        RECT 133.170 16.520 133.570 16.565 ;
        RECT 136.270 16.520 136.670 16.565 ;
        RECT 137.770 16.795 138.170 16.870 ;
        RECT 140.870 16.795 141.270 16.870 ;
        RECT 141.670 16.795 142.670 17.170 ;
        RECT 137.770 16.570 142.670 16.795 ;
        RECT 137.770 16.520 138.170 16.570 ;
        RECT 140.870 16.550 142.670 16.570 ;
        RECT 140.870 16.520 141.270 16.550 ;
        RECT 133.280 16.470 133.510 16.520 ;
        RECT 136.330 16.470 136.560 16.520 ;
        RECT 137.880 16.470 138.110 16.520 ;
        RECT 140.930 16.470 141.160 16.520 ;
        RECT 133.670 16.320 136.170 16.420 ;
        RECT 138.270 16.320 140.770 16.420 ;
        RECT 133.670 16.190 140.770 16.320 ;
        RECT 133.870 15.970 140.520 16.190 ;
        RECT 141.670 16.170 142.670 16.550 ;
        RECT 146.320 16.520 147.620 29.320 ;
        RECT 148.420 29.170 149.470 29.320 ;
        RECT 148.470 29.070 149.470 29.170 ;
        RECT 148.080 28.670 148.310 29.020 ;
        RECT 147.970 28.470 148.320 28.670 ;
        RECT 149.630 28.470 149.860 29.020 ;
        RECT 147.970 27.520 149.860 28.470 ;
        RECT 147.970 26.220 148.320 27.520 ;
        RECT 148.470 26.770 149.470 27.070 ;
        RECT 149.630 27.060 149.860 27.520 ;
        RECT 149.630 26.220 149.860 26.730 ;
        RECT 147.970 25.270 149.860 26.220 ;
        RECT 147.970 23.870 148.320 25.270 ;
        RECT 149.630 24.770 149.860 25.270 ;
        RECT 148.470 24.470 149.470 24.770 ;
        RECT 149.630 23.870 149.860 24.440 ;
        RECT 147.970 22.920 149.860 23.870 ;
        RECT 147.970 21.720 148.320 22.920 ;
        RECT 149.630 22.480 149.860 22.920 ;
        RECT 148.470 22.170 149.470 22.470 ;
        RECT 149.630 21.720 149.860 22.150 ;
        RECT 147.970 20.770 149.860 21.720 ;
        RECT 147.970 19.420 148.320 20.770 ;
        RECT 148.470 19.870 149.470 20.220 ;
        RECT 149.630 20.190 149.860 20.770 ;
        RECT 149.630 19.420 149.860 19.860 ;
        RECT 147.970 18.470 149.860 19.420 ;
        RECT 147.970 17.170 148.320 18.470 ;
        RECT 148.470 17.570 149.470 17.920 ;
        RECT 149.630 17.900 149.860 18.470 ;
        RECT 149.630 17.170 149.860 17.570 ;
        RECT 147.970 16.220 149.860 17.170 ;
        RECT 128.530 15.560 128.760 15.970 ;
        RECT 130.070 15.720 131.020 15.970 ;
        RECT 130.070 15.570 131.400 15.720 ;
        RECT 132.720 15.570 133.720 15.870 ;
        RECT 128.920 15.270 131.400 15.570 ;
        RECT 128.530 14.870 128.760 15.230 ;
        RECT 130.070 15.070 131.400 15.270 ;
        RECT 130.070 14.870 131.020 15.070 ;
        RECT 134.720 15.020 139.970 15.970 ;
        RECT 140.870 15.570 141.870 15.870 ;
        RECT 145.825 15.840 146.715 15.870 ;
        RECT 147.970 15.840 148.320 16.220 ;
        RECT 145.825 14.950 148.320 15.840 ;
        RECT 149.630 15.610 149.860 16.220 ;
        RECT 148.570 15.560 149.470 15.570 ;
        RECT 148.470 15.330 149.470 15.560 ;
        RECT 148.570 15.270 149.470 15.330 ;
        RECT 145.825 14.920 146.715 14.950 ;
        RECT 128.520 13.720 131.020 14.870 ;
        RECT 147.970 14.820 148.320 14.950 ;
        RECT 149.630 14.820 149.860 15.280 ;
        RECT 132.920 14.530 134.880 14.760 ;
        RECT 135.210 14.530 137.170 14.760 ;
        RECT 137.500 14.530 139.460 14.760 ;
        RECT 139.790 14.530 141.750 14.760 ;
        RECT 132.640 14.320 132.870 14.370 ;
        RECT 128.530 13.270 128.760 13.720 ;
        RECT 130.070 13.270 131.020 13.720 ;
        RECT 132.520 13.420 132.920 14.320 ;
        RECT 132.640 13.370 132.870 13.420 ;
        RECT 130.120 13.220 131.020 13.270 ;
        RECT 133.370 13.220 134.270 14.530 ;
        RECT 134.930 14.220 135.160 14.370 ;
        RECT 134.820 13.520 135.270 14.220 ;
        RECT 134.930 13.370 135.160 13.520 ;
        RECT 135.770 13.220 136.670 14.530 ;
        RECT 137.220 14.220 137.450 14.370 ;
        RECT 137.120 13.520 137.570 14.220 ;
        RECT 137.220 13.370 137.450 13.520 ;
        RECT 138.070 13.220 138.970 14.530 ;
        RECT 139.510 14.220 139.740 14.370 ;
        RECT 139.420 13.520 139.870 14.220 ;
        RECT 139.510 13.370 139.740 13.520 ;
        RECT 140.320 13.220 141.220 14.530 ;
        RECT 141.800 14.320 142.030 14.370 ;
        RECT 141.720 13.420 142.120 14.320 ;
        RECT 141.800 13.370 142.030 13.420 ;
        RECT 128.920 12.870 129.920 13.220 ;
        RECT 130.120 13.210 141.720 13.220 ;
        RECT 130.120 12.980 141.750 13.210 ;
        RECT 130.120 12.920 141.720 12.980 ;
        RECT 142.320 12.720 143.670 14.770 ;
        RECT 146.120 12.720 147.820 14.220 ;
        RECT 147.970 13.870 149.920 14.820 ;
        RECT 150.170 14.220 150.920 27.170 ;
        RECT 147.970 13.370 148.320 13.870 ;
        RECT 148.080 13.320 148.310 13.370 ;
        RECT 149.630 13.320 149.860 13.870 ;
        RECT 148.470 12.970 149.470 13.320 ;
        RECT 150.070 12.720 150.920 14.220 ;
        RECT 117.950 12.050 119.450 12.080 ;
        RECT 126.720 12.050 150.920 12.720 ;
        RECT 117.950 10.550 150.920 12.050 ;
        RECT 117.950 10.520 119.450 10.550 ;
        RECT 126.720 10.370 150.920 10.550 ;
      LAYER via ;
        RECT 137.370 102.570 139.870 105.070 ;
        RECT 106.270 97.570 107.970 98.770 ;
        RECT 120.270 97.570 121.970 98.770 ;
        RECT 107.770 83.670 109.470 84.770 ;
        RECT 134.370 97.570 136.070 98.770 ;
        RECT 120.870 83.670 122.570 84.770 ;
        RECT 90.670 73.370 93.870 73.870 ;
        RECT 106.870 69.670 110.970 70.470 ;
        RECT 139.230 74.640 140.330 75.740 ;
        RECT 148.170 73.170 151.070 74.070 ;
        RECT 120.070 63.370 122.870 63.970 ;
        RECT 130.470 69.570 133.570 70.270 ;
        RECT 90.670 51.970 93.870 54.170 ;
        RECT 148.270 51.970 150.970 53.870 ;
        RECT 139.920 32.770 140.920 33.070 ;
        RECT 131.470 30.770 132.320 31.120 ;
        RECT 131.370 30.470 132.320 30.770 ;
        RECT 126.870 12.820 127.670 22.620 ;
        RECT 128.970 22.120 129.870 22.470 ;
        RECT 131.470 26.170 132.320 30.470 ;
        RECT 131.370 25.870 132.320 26.170 ;
        RECT 131.470 21.620 132.320 25.870 ;
        RECT 131.370 21.320 132.320 21.620 ;
        RECT 131.470 21.170 132.320 21.320 ;
        RECT 133.620 30.470 134.520 30.770 ;
        RECT 133.620 25.870 134.520 26.170 ;
        RECT 133.620 21.320 134.520 21.620 ;
        RECT 140.020 30.470 140.920 30.770 ;
        RECT 139.920 28.170 140.920 28.470 ;
        RECT 140.020 25.870 140.920 26.170 ;
        RECT 139.920 23.570 140.920 23.870 ;
        RECT 140.020 21.320 140.920 21.620 ;
        RECT 142.220 23.870 143.070 33.520 ;
        RECT 144.520 33.020 145.470 33.320 ;
        RECT 142.220 23.470 143.120 23.870 ;
        RECT 142.220 22.320 143.070 23.470 ;
        RECT 142.220 21.920 143.120 22.320 ;
        RECT 128.970 17.520 129.870 17.870 ;
        RECT 139.920 18.970 140.920 19.270 ;
        RECT 140.195 18.720 140.745 18.970 ;
        RECT 139.970 17.370 140.820 18.020 ;
        RECT 142.220 20.720 143.070 21.920 ;
        RECT 142.220 17.720 143.120 20.720 ;
        RECT 142.220 17.370 143.470 17.720 ;
        RECT 142.320 17.320 143.470 17.370 ;
        RECT 144.570 32.220 145.520 32.520 ;
        RECT 144.520 31.420 145.470 31.720 ;
        RECT 144.570 30.620 145.520 30.920 ;
        RECT 144.520 29.870 145.470 30.170 ;
        RECT 144.570 29.070 145.520 29.370 ;
        RECT 144.520 28.270 145.470 28.570 ;
        RECT 144.570 27.470 145.520 27.770 ;
        RECT 144.520 26.670 145.470 26.970 ;
        RECT 144.570 25.870 145.520 26.170 ;
        RECT 144.520 25.120 145.470 25.420 ;
        RECT 144.570 24.320 145.520 24.620 ;
        RECT 144.520 23.520 145.470 23.820 ;
        RECT 144.570 22.770 145.520 23.070 ;
        RECT 144.520 21.970 145.470 22.270 ;
        RECT 144.570 21.170 145.520 21.470 ;
        RECT 144.520 20.370 145.470 20.670 ;
        RECT 144.020 19.520 144.320 19.920 ;
        RECT 144.570 19.570 145.520 19.870 ;
        RECT 144.520 18.770 145.470 19.070 ;
        RECT 144.570 18.020 145.520 18.320 ;
        RECT 144.520 17.220 145.470 17.520 ;
        RECT 131.920 16.950 132.620 16.970 ;
        RECT 131.895 16.395 132.620 16.950 ;
        RECT 131.920 16.370 132.620 16.395 ;
        RECT 133.220 16.520 133.520 16.870 ;
        RECT 136.320 16.520 136.620 16.870 ;
        RECT 137.820 16.520 138.120 16.870 ;
        RECT 140.920 16.520 141.220 16.870 ;
        RECT 141.945 16.400 142.495 16.950 ;
        RECT 146.670 16.520 147.270 32.370 ;
        RECT 150.370 29.670 150.770 32.370 ;
        RECT 148.470 29.170 149.420 29.470 ;
        RECT 148.620 29.070 149.370 29.170 ;
        RECT 148.520 26.770 149.420 27.070 ;
        RECT 148.520 24.470 149.420 24.770 ;
        RECT 148.520 22.170 149.420 22.470 ;
        RECT 148.520 19.870 149.420 20.220 ;
        RECT 148.520 17.570 149.420 17.920 ;
        RECT 130.720 15.070 131.370 15.720 ;
        RECT 132.770 15.570 133.670 15.870 ;
        RECT 134.870 15.320 135.270 16.020 ;
        RECT 139.420 15.320 139.820 16.020 ;
        RECT 140.920 15.570 141.820 15.870 ;
        RECT 148.620 15.270 149.420 15.570 ;
        RECT 132.570 13.420 132.870 14.320 ;
        RECT 134.870 13.520 135.220 14.220 ;
        RECT 137.170 13.520 137.520 14.220 ;
        RECT 139.470 13.520 139.820 14.220 ;
        RECT 141.770 13.420 142.070 14.320 ;
        RECT 128.970 12.870 129.870 13.220 ;
        RECT 150.320 14.520 150.720 27.020 ;
        RECT 148.520 12.970 149.420 13.320 ;
        RECT 132.420 12.170 132.920 12.270 ;
        RECT 137.170 12.170 137.520 12.270 ;
        RECT 141.570 12.170 142.070 12.270 ;
        RECT 132.420 11.820 142.070 12.170 ;
        RECT 132.420 11.520 142.020 11.820 ;
      LAYER met2 ;
        RECT 75.005 105.150 76.455 105.170 ;
        RECT 74.980 103.650 80.860 105.150 ;
        RECT 75.005 103.630 76.455 103.650 ;
        RECT 106.170 97.470 136.170 98.970 ;
        RECT 137.070 89.970 140.070 105.570 ;
        RECT 130.670 86.970 140.070 89.970 ;
        RECT 107.670 83.570 122.670 84.870 ;
        RECT 90.470 51.670 94.070 74.070 ;
        RECT 130.670 71.470 133.670 86.970 ;
        RECT 106.470 68.470 133.670 71.470 ;
        RECT 119.970 62.870 122.970 68.470 ;
        RECT 107.915 46.050 109.365 46.070 ;
        RECT 107.890 44.550 112.500 46.050 ;
        RECT 139.230 45.270 140.330 75.770 ;
        RECT 148.070 51.770 151.170 74.470 ;
        RECT 107.915 44.530 109.365 44.550 ;
        RECT 139.230 44.170 153.750 45.270 ;
        RECT 102.555 35.350 104.005 35.370 ;
        RECT 102.530 33.850 106.110 35.350 ;
        RECT 102.555 33.830 104.005 33.850 ;
        RECT 142.220 33.370 143.070 33.570 ;
        RECT 136.330 33.320 138.110 33.360 ;
        RECT 136.320 33.070 140.970 33.320 ;
        RECT 136.330 32.770 140.970 33.070 ;
        RECT 142.220 32.970 145.520 33.370 ;
        RECT 136.330 32.730 140.920 32.770 ;
        RECT 131.470 30.820 132.320 31.170 ;
        RECT 131.370 30.770 132.320 30.820 ;
        RECT 133.620 30.770 134.520 30.820 ;
        RECT 131.320 30.470 134.770 30.770 ;
        RECT 131.370 30.420 132.320 30.470 ;
        RECT 133.620 30.420 134.520 30.470 ;
        RECT 131.470 26.220 132.320 30.420 ;
        RECT 136.330 28.510 138.110 32.730 ;
        RECT 139.920 32.720 140.920 32.730 ;
        RECT 142.220 31.770 143.070 32.970 ;
        RECT 144.520 32.170 150.920 32.570 ;
        RECT 142.220 31.370 145.520 31.770 ;
        RECT 142.220 30.820 143.070 31.370 ;
        RECT 146.320 30.920 150.920 32.170 ;
        RECT 140.020 30.470 143.070 30.820 ;
        RECT 144.520 30.620 150.920 30.920 ;
        RECT 140.020 30.420 140.920 30.470 ;
        RECT 142.220 30.220 143.070 30.470 ;
        RECT 142.220 29.820 145.520 30.220 ;
        RECT 142.220 28.620 143.070 29.820 ;
        RECT 146.370 29.370 150.920 30.620 ;
        RECT 144.520 29.070 149.620 29.370 ;
        RECT 146.320 28.920 149.620 29.070 ;
        RECT 139.920 28.510 140.920 28.520 ;
        RECT 136.330 28.130 140.970 28.510 ;
        RECT 142.220 28.220 145.520 28.620 ;
        RECT 131.370 26.170 132.320 26.220 ;
        RECT 133.620 26.170 134.520 26.220 ;
        RECT 131.320 25.870 134.770 26.170 ;
        RECT 131.370 25.820 132.320 25.870 ;
        RECT 133.620 25.820 134.520 25.870 ;
        RECT 126.870 22.620 127.670 22.670 ;
        RECT 126.870 21.970 130.020 22.620 ;
        RECT 126.870 18.070 127.670 21.970 ;
        RECT 131.470 21.670 132.320 25.820 ;
        RECT 136.330 23.910 138.110 28.130 ;
        RECT 139.920 28.120 140.920 28.130 ;
        RECT 142.220 27.020 143.070 28.220 ;
        RECT 146.320 27.770 147.620 28.920 ;
        RECT 144.520 27.470 147.620 27.770 ;
        RECT 142.220 26.620 145.470 27.020 ;
        RECT 142.220 26.270 143.070 26.620 ;
        RECT 140.020 25.870 143.070 26.270 ;
        RECT 146.320 26.220 147.620 27.470 ;
        RECT 148.470 26.620 150.920 27.170 ;
        RECT 152.650 26.725 153.750 44.170 ;
        RECT 144.520 25.870 147.620 26.220 ;
        RECT 140.020 25.820 140.920 25.870 ;
        RECT 142.220 25.470 143.070 25.870 ;
        RECT 142.220 25.070 145.470 25.470 ;
        RECT 139.920 23.910 140.920 23.920 ;
        RECT 136.330 23.530 140.920 23.910 ;
        RECT 131.370 21.620 132.320 21.670 ;
        RECT 133.620 21.620 134.520 21.670 ;
        RECT 131.320 21.320 134.770 21.620 ;
        RECT 131.370 21.270 132.320 21.320 ;
        RECT 133.620 21.270 134.520 21.320 ;
        RECT 131.470 21.120 132.320 21.270 ;
        RECT 136.330 20.030 138.110 23.530 ;
        RECT 139.920 23.520 140.920 23.530 ;
        RECT 142.220 23.870 143.070 25.070 ;
        RECT 146.320 24.870 147.620 25.870 ;
        RECT 146.320 24.620 149.620 24.870 ;
        RECT 144.520 24.320 149.620 24.620 ;
        RECT 144.520 24.270 147.620 24.320 ;
        RECT 142.220 23.470 145.520 23.870 ;
        RECT 142.220 22.320 143.070 23.470 ;
        RECT 146.320 23.070 147.620 24.270 ;
        RECT 144.520 22.720 147.620 23.070 ;
        RECT 142.220 21.920 145.520 22.320 ;
        RECT 142.220 21.670 143.070 21.920 ;
        RECT 140.020 21.320 143.070 21.670 ;
        RECT 146.320 21.470 147.620 22.720 ;
        RECT 150.170 22.620 150.920 26.620 ;
        RECT 152.630 25.675 153.770 26.725 ;
        RECT 152.650 25.650 153.750 25.675 ;
        RECT 148.470 22.070 150.920 22.620 ;
        RECT 140.020 21.270 140.920 21.320 ;
        RECT 142.220 20.720 143.070 21.320 ;
        RECT 144.520 21.120 147.620 21.470 ;
        RECT 142.220 20.320 145.520 20.720 ;
        RECT 136.340 18.790 138.100 20.030 ;
        RECT 140.195 19.320 140.745 19.890 ;
        RECT 126.870 17.420 130.020 18.070 ;
        RECT 139.920 17.770 140.920 19.320 ;
        RECT 142.220 19.120 143.120 20.320 ;
        RECT 146.320 20.270 147.620 21.120 ;
        RECT 143.320 19.470 144.320 19.970 ;
        RECT 146.320 19.920 149.620 20.270 ;
        RECT 144.520 19.720 149.620 19.920 ;
        RECT 144.520 19.520 147.620 19.720 ;
        RECT 143.320 19.420 144.020 19.470 ;
        RECT 142.220 18.720 145.470 19.120 ;
        RECT 142.220 17.770 143.120 18.720 ;
        RECT 146.320 18.370 147.620 19.520 ;
        RECT 144.520 17.970 147.620 18.370 ;
        RECT 150.170 18.020 150.920 22.070 ;
        RECT 126.870 13.470 127.670 17.420 ;
        RECT 139.970 17.320 140.820 17.770 ;
        RECT 142.220 17.620 143.470 17.770 ;
        RECT 142.220 17.320 145.470 17.620 ;
        RECT 131.900 16.980 132.700 17.250 ;
        RECT 143.370 17.170 145.470 17.320 ;
        RECT 142.000 16.980 142.700 17.150 ;
        RECT 131.895 16.950 132.700 16.980 ;
        RECT 141.945 16.950 142.700 16.980 ;
        RECT 131.895 16.920 136.595 16.950 ;
        RECT 137.845 16.920 142.700 16.950 ;
        RECT 131.895 16.470 136.620 16.920 ;
        RECT 137.820 16.470 142.700 16.920 ;
        RECT 146.320 17.120 147.620 17.970 ;
        RECT 148.470 17.470 150.920 18.020 ;
        RECT 146.320 16.520 149.420 17.120 ;
        RECT 131.895 16.395 136.595 16.470 ;
        RECT 137.845 16.450 142.700 16.470 ;
        RECT 137.845 16.400 142.495 16.450 ;
        RECT 131.895 16.365 132.700 16.395 ;
        RECT 141.945 16.370 142.495 16.400 ;
        RECT 131.900 16.350 132.700 16.365 ;
        RECT 131.920 16.320 132.620 16.350 ;
        RECT 130.720 15.720 131.370 15.750 ;
        RECT 130.720 15.070 132.090 15.720 ;
        RECT 132.370 15.470 133.720 15.920 ;
        RECT 130.720 15.040 131.370 15.070 ;
        RECT 126.870 12.820 130.020 13.470 ;
        RECT 126.870 12.770 127.670 12.820 ;
        RECT 132.370 12.270 133.020 15.470 ;
        RECT 134.770 13.370 135.370 16.120 ;
        RECT 137.070 12.270 137.620 14.370 ;
        RECT 139.320 13.370 139.920 16.120 ;
        RECT 140.820 15.470 142.170 15.920 ;
        RECT 144.805 15.840 145.645 16.015 ;
        RECT 141.520 12.270 142.170 15.470 ;
        RECT 144.780 14.950 146.745 15.840 ;
        RECT 148.620 15.220 149.420 16.520 ;
        RECT 144.805 14.775 145.645 14.950 ;
        RECT 150.170 13.470 150.920 17.470 ;
        RECT 148.470 12.920 150.920 13.470 ;
        RECT 109.275 12.050 110.725 12.070 ;
        RECT 109.250 10.550 119.480 12.050 ;
        RECT 132.370 11.370 142.170 12.270 ;
        RECT 109.275 10.530 110.725 10.550 ;
      LAYER via2 ;
        RECT 75.005 103.675 76.455 105.125 ;
        RECT 107.915 44.575 109.365 46.025 ;
        RECT 102.555 33.875 104.005 35.325 ;
        RECT 147.800 30.300 149.800 32.100 ;
        RECT 152.675 25.675 153.725 26.725 ;
        RECT 136.570 19.270 138.020 20.070 ;
        RECT 140.195 19.295 140.745 19.845 ;
        RECT 131.900 16.400 132.700 17.200 ;
        RECT 142.000 16.500 142.700 17.100 ;
        RECT 131.395 15.070 132.045 15.720 ;
        RECT 144.805 14.820 145.645 15.970 ;
        RECT 109.275 10.575 110.725 12.025 ;
      LAYER met3 ;
        RECT 64.990 103.650 76.480 105.150 ;
        RECT 32.155 64.950 33.645 64.975 ;
        RECT 64.990 64.950 66.490 103.650 ;
        RECT 32.150 63.450 66.490 64.950 ;
        RECT 32.155 63.425 33.645 63.450 ;
        RECT 64.990 35.350 66.490 63.450 ;
        RECT 104.475 46.050 105.965 46.075 ;
        RECT 104.470 44.550 109.390 46.050 ;
        RECT 104.475 44.525 105.965 44.550 ;
        RECT 64.990 33.850 104.030 35.350 ;
        RECT 147.400 31.750 154.900 32.200 ;
        RECT 156.415 31.750 157.305 31.775 ;
        RECT 147.400 30.850 157.310 31.750 ;
        RECT 147.400 30.600 154.900 30.850 ;
        RECT 156.415 30.825 157.305 30.850 ;
        RECT 147.750 30.275 149.850 30.600 ;
        RECT 136.470 20.085 143.420 20.120 ;
        RECT 136.470 19.895 143.985 20.085 ;
        RECT 136.470 19.445 144.020 19.895 ;
        RECT 136.470 19.260 143.985 19.445 ;
        RECT 136.470 19.170 143.420 19.260 ;
        RECT 138.770 18.670 141.620 19.170 ;
        RECT 123.700 16.400 133.000 17.600 ;
        RECT 152.650 17.400 153.750 26.750 ;
        RECT 99.955 12.050 101.445 12.075 ;
        RECT 99.950 10.550 110.750 12.050 ;
        RECT 99.955 10.525 101.445 10.550 ;
        RECT 123.800 8.700 125.000 16.400 ;
        RECT 131.850 16.375 132.750 16.400 ;
        RECT 141.800 16.300 153.750 17.400 ;
        RECT 131.120 14.795 145.670 15.995 ;
        RECT 123.800 7.500 153.730 8.700 ;
      LAYER via3 ;
        RECT 32.155 63.455 33.645 64.945 ;
        RECT 104.475 44.555 105.965 46.045 ;
        RECT 156.415 30.855 157.305 31.745 ;
        RECT 99.955 10.555 101.445 12.045 ;
        RECT 152.500 7.500 153.700 8.700 ;
      LAYER met4 ;
        RECT 3.990 223.850 4.290 224.760 ;
        RECT 7.670 223.850 7.970 224.760 ;
        RECT 11.350 223.850 11.650 224.760 ;
        RECT 15.030 223.850 15.330 224.760 ;
        RECT 18.710 223.850 19.010 224.760 ;
        RECT 22.390 223.850 22.690 224.760 ;
        RECT 26.070 223.850 26.370 224.760 ;
        RECT 29.750 223.850 30.050 224.760 ;
        RECT 33.430 223.850 33.730 224.760 ;
        RECT 37.110 223.850 37.410 224.760 ;
        RECT 40.790 223.850 41.090 224.760 ;
        RECT 44.470 223.850 44.770 224.760 ;
        RECT 48.150 223.850 48.450 224.760 ;
        RECT 51.830 223.850 52.130 224.760 ;
        RECT 55.510 223.850 55.810 224.760 ;
        RECT 59.190 223.850 59.490 224.760 ;
        RECT 62.870 223.850 63.170 224.760 ;
        RECT 66.550 223.850 66.850 224.760 ;
        RECT 70.230 223.850 70.530 224.760 ;
        RECT 73.910 223.850 74.210 224.760 ;
        RECT 77.590 223.850 77.890 224.760 ;
        RECT 81.270 223.850 81.570 224.760 ;
        RECT 84.950 223.850 85.250 224.760 ;
        RECT 88.630 223.850 88.930 224.760 ;
        RECT 2.850 223.550 88.930 223.850 ;
        RECT 49.650 220.760 49.950 223.550 ;
        RECT 2.500 63.450 33.650 64.950 ;
        RECT 50.500 44.550 105.970 46.050 ;
        RECT 99.910 31.140 101.410 44.550 ;
        RECT 99.910 27.120 101.450 31.140 ;
        RECT 99.950 10.550 101.450 27.120 ;
        RECT 152.495 8.700 153.705 8.705 ;
        RECT 156.410 8.700 157.310 31.750 ;
        RECT 152.495 7.500 157.310 8.700 ;
        RECT 152.495 7.495 153.705 7.500 ;
        RECT 156.410 1.000 157.310 7.500 ;
  END
END tt_um_mos_bandgap
END LIBRARY

