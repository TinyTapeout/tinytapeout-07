VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_nurirfansyah_alits02
  CLASS BLOCK ;
  FOREIGN tt_um_nurirfansyah_alits02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.810000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.405000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.405000 ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.810000 ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    ANTENNADIFFAREA 0.261000 ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    ANTENNADIFFAREA 0.261000 ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.135000 ;
    ANTENNADIFFAREA 5.690100 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 75.130 60.000 76.630 61.650 ;
        RECT 77.930 60.000 79.430 61.650 ;
        RECT 80.730 60.000 82.230 61.650 ;
        RECT 83.530 60.000 85.030 61.650 ;
        RECT 86.330 60.000 87.830 61.650 ;
        RECT 89.130 60.000 90.630 61.650 ;
        RECT 76.600 45.910 89.440 46.860 ;
        RECT 76.610 44.590 89.440 45.910 ;
      LAYER pwell ;
        RECT 76.610 42.230 89.440 44.280 ;
        RECT 84.460 41.900 84.820 42.230 ;
        RECT 86.450 42.210 86.620 42.230 ;
      LAYER nwell ;
        RECT 127.850 24.000 129.350 25.650 ;
        RECT 130.650 24.000 132.150 25.650 ;
        RECT 133.450 24.000 134.950 25.650 ;
        RECT 136.250 24.000 137.750 25.650 ;
        RECT 139.050 24.000 140.550 25.650 ;
        RECT 141.850 24.000 143.350 25.650 ;
      LAYER li1 ;
        RECT 75.330 61.100 75.880 61.400 ;
        RECT 76.080 61.000 76.630 61.950 ;
        RECT 78.130 61.100 79.230 61.400 ;
        RECT 80.930 61.100 81.480 61.400 ;
        RECT 75.330 59.200 75.730 60.850 ;
        RECT 76.030 60.150 76.430 60.750 ;
        RECT 78.130 60.300 78.530 61.100 ;
        RECT 80.930 61.000 81.330 61.100 ;
        RECT 81.680 61.000 82.230 61.950 ;
        RECT 83.730 61.100 84.830 61.400 ;
        RECT 86.530 61.100 87.080 61.400 ;
        RECT 76.030 59.750 76.630 60.150 ;
        RECT 77.930 59.850 78.580 60.100 ;
        RECT 76.030 59.200 76.430 59.750 ;
        RECT 75.330 58.550 75.880 58.850 ;
        RECT 76.080 58.000 76.630 58.950 ;
        RECT 78.130 58.850 78.530 59.650 ;
        RECT 78.830 59.200 79.230 60.750 ;
        RECT 80.930 59.200 81.330 60.750 ;
        RECT 81.630 60.150 82.030 60.750 ;
        RECT 83.730 60.300 84.130 61.100 ;
        RECT 86.530 61.000 86.930 61.100 ;
        RECT 87.280 61.000 87.830 61.950 ;
        RECT 89.330 61.100 90.430 61.400 ;
        RECT 81.630 59.750 82.230 60.150 ;
        RECT 83.530 59.850 84.180 60.100 ;
        RECT 81.630 59.200 82.030 59.750 ;
        RECT 78.130 58.550 79.230 58.850 ;
        RECT 80.930 58.550 81.480 58.850 ;
        RECT 81.680 58.000 82.230 58.950 ;
        RECT 83.730 58.850 84.130 59.650 ;
        RECT 84.430 59.200 84.830 60.750 ;
        RECT 86.530 59.200 86.930 60.750 ;
        RECT 87.230 60.150 87.630 60.750 ;
        RECT 89.330 60.300 89.730 61.100 ;
        RECT 87.230 59.750 87.830 60.150 ;
        RECT 89.130 59.850 89.780 60.100 ;
        RECT 87.230 59.200 87.630 59.750 ;
        RECT 83.730 58.550 84.830 58.850 ;
        RECT 86.530 58.550 87.080 58.850 ;
        RECT 87.280 58.000 87.830 58.950 ;
        RECT 89.330 58.850 89.730 59.650 ;
        RECT 90.030 59.200 90.430 60.750 ;
        RECT 89.330 58.550 90.430 58.850 ;
        RECT 77.170 45.440 77.500 46.660 ;
        RECT 78.480 45.440 78.810 46.660 ;
        RECT 79.390 45.950 79.720 46.660 ;
        RECT 76.705 45.290 76.875 45.300 ;
        RECT 76.700 44.560 76.880 45.290 ;
        RECT 77.090 45.270 77.580 45.440 ;
        RECT 77.170 45.260 77.500 45.270 ;
        RECT 77.090 44.830 77.580 45.000 ;
        RECT 78.015 44.970 78.185 45.300 ;
        RECT 78.400 45.270 78.890 45.440 ;
        RECT 78.400 44.830 78.890 45.000 ;
        RECT 79.470 44.900 79.640 45.950 ;
        RECT 79.910 45.700 80.080 46.660 ;
        RECT 80.780 46.190 84.220 46.360 ;
        RECT 80.780 45.775 80.950 46.190 ;
        RECT 80.700 45.605 81.030 45.775 ;
        RECT 82.970 45.600 83.310 45.840 ;
        RECT 84.050 45.775 84.220 46.190 ;
        RECT 83.970 45.605 84.300 45.775 ;
        RECT 86.010 45.700 86.180 46.660 ;
        RECT 86.360 45.950 86.690 46.660 ;
        RECT 84.050 45.600 84.220 45.605 ;
        RECT 76.700 44.380 78.200 44.560 ;
        RECT 76.750 42.400 76.920 44.050 ;
        RECT 77.090 44.020 77.580 44.190 ;
        RECT 78.020 43.800 78.200 44.380 ;
        RECT 79.420 44.340 79.700 44.670 ;
        RECT 78.400 44.020 78.890 44.190 ;
        RECT 77.090 43.580 77.580 43.750 ;
        RECT 78.400 43.580 78.890 43.750 ;
        RECT 79.470 43.630 79.640 44.120 ;
        RECT 79.910 43.630 80.080 45.390 ;
        RECT 80.560 44.590 80.730 45.390 ;
        RECT 80.550 44.420 80.730 44.590 ;
        RECT 80.560 43.630 80.730 44.420 ;
        RECT 81.000 44.610 81.170 45.390 ;
        RECT 81.650 44.900 81.820 45.390 ;
        RECT 81.000 44.280 81.590 44.610 ;
        RECT 81.000 43.630 81.170 44.280 ;
        RECT 81.650 44.110 81.820 44.120 ;
        RECT 81.500 43.630 81.820 44.110 ;
        RECT 82.090 43.630 82.260 45.390 ;
        RECT 82.740 44.900 82.910 45.390 ;
        RECT 82.570 43.630 82.910 44.120 ;
        RECT 83.180 43.630 83.350 45.390 ;
        RECT 83.830 44.040 84.000 45.390 ;
        RECT 84.270 44.590 84.440 45.390 ;
        RECT 84.260 44.420 84.450 44.590 ;
        RECT 83.520 43.630 84.000 44.040 ;
        RECT 84.270 43.630 84.440 44.420 ;
        RECT 78.020 43.190 78.200 43.520 ;
        RECT 78.400 43.140 78.890 43.310 ;
        RECT 80.700 43.290 81.030 43.460 ;
        RECT 79.910 42.600 80.080 43.170 ;
        RECT 80.780 42.800 80.950 43.290 ;
        RECT 81.500 43.080 81.670 43.630 ;
        RECT 81.880 43.260 82.220 43.440 ;
        RECT 82.570 43.080 82.740 43.630 ;
        RECT 83.520 43.440 83.690 43.630 ;
        RECT 82.970 43.260 83.690 43.440 ;
        RECT 84.060 43.260 84.400 43.440 ;
        RECT 81.500 42.910 82.740 43.080 ;
        RECT 80.780 42.740 81.020 42.800 ;
        RECT 84.140 42.740 84.320 43.260 ;
        RECT 80.780 42.570 84.320 42.740 ;
        RECT 84.920 42.400 85.090 45.390 ;
        RECT 85.360 44.890 85.530 45.390 ;
        RECT 85.330 44.340 85.520 44.670 ;
        RECT 85.360 42.910 85.530 44.120 ;
        RECT 86.010 43.630 86.180 45.390 ;
        RECT 86.450 44.900 86.620 45.950 ;
        RECT 87.220 45.440 87.550 46.660 ;
        RECT 88.540 45.440 88.870 46.660 ;
        RECT 87.140 45.270 87.630 45.440 ;
        RECT 87.140 44.830 87.630 45.000 ;
        RECT 87.845 44.970 88.015 45.300 ;
        RECT 88.460 45.270 88.950 45.440 ;
        RECT 88.460 44.830 88.950 45.000 ;
        RECT 86.390 44.340 86.670 44.670 ;
        RECT 89.160 44.620 89.340 45.300 ;
        RECT 87.820 44.440 89.340 44.620 ;
        RECT 86.010 42.600 86.180 43.170 ;
        RECT 86.450 42.910 86.620 44.120 ;
        RECT 87.140 44.020 87.630 44.190 ;
        RECT 87.820 43.810 88.000 44.440 ;
        RECT 88.460 44.020 88.950 44.190 ;
        RECT 87.140 43.580 87.630 43.750 ;
        RECT 88.460 43.580 88.950 43.750 ;
        RECT 87.140 43.140 87.630 43.310 ;
        RECT 87.820 43.190 88.000 43.520 ;
        RECT 89.120 42.400 89.290 44.050 ;
        RECT 76.750 42.230 89.290 42.400 ;
        RECT 128.050 25.100 128.600 25.400 ;
        RECT 128.800 25.000 129.350 25.950 ;
        RECT 130.850 25.100 131.950 25.400 ;
        RECT 133.650 25.100 134.200 25.400 ;
        RECT 128.050 23.200 128.450 24.850 ;
        RECT 128.750 24.150 129.150 24.750 ;
        RECT 130.850 24.300 131.250 25.100 ;
        RECT 133.650 25.000 134.050 25.100 ;
        RECT 134.400 25.000 134.950 25.950 ;
        RECT 136.450 25.100 137.550 25.400 ;
        RECT 139.250 25.100 139.800 25.400 ;
        RECT 128.750 23.750 129.350 24.150 ;
        RECT 130.650 23.850 131.300 24.100 ;
        RECT 128.750 23.200 129.150 23.750 ;
        RECT 128.050 22.550 128.600 22.850 ;
        RECT 128.800 22.000 129.350 22.950 ;
        RECT 130.850 22.850 131.250 23.650 ;
        RECT 131.550 23.200 131.950 24.750 ;
        RECT 133.650 23.200 134.050 24.750 ;
        RECT 134.350 24.150 134.750 24.750 ;
        RECT 136.450 24.300 136.850 25.100 ;
        RECT 139.250 25.000 139.650 25.100 ;
        RECT 140.000 25.000 140.550 25.950 ;
        RECT 142.050 25.100 143.150 25.400 ;
        RECT 134.350 23.750 134.950 24.150 ;
        RECT 136.250 23.850 136.900 24.100 ;
        RECT 134.350 23.200 134.750 23.750 ;
        RECT 130.850 22.550 131.950 22.850 ;
        RECT 133.650 22.550 134.200 22.850 ;
        RECT 134.400 22.000 134.950 22.950 ;
        RECT 136.450 22.850 136.850 23.650 ;
        RECT 137.150 23.200 137.550 24.750 ;
        RECT 139.250 23.200 139.650 24.750 ;
        RECT 139.950 24.150 140.350 24.750 ;
        RECT 142.050 24.300 142.450 25.100 ;
        RECT 139.950 23.750 140.550 24.150 ;
        RECT 141.850 23.850 142.500 24.100 ;
        RECT 139.950 23.200 140.350 23.750 ;
        RECT 136.450 22.550 137.550 22.850 ;
        RECT 139.250 22.550 139.800 22.850 ;
        RECT 140.000 22.000 140.550 22.950 ;
        RECT 142.050 22.850 142.450 23.650 ;
        RECT 142.750 23.200 143.150 24.750 ;
        RECT 142.050 22.550 143.150 22.850 ;
      LAYER met1 ;
        RECT 60.400 63.755 62.200 64.100 ;
        RECT 60.400 63.045 93.755 63.755 ;
        RECT 60.400 62.450 62.200 63.045 ;
        RECT 70.800 61.550 87.830 61.950 ;
        RECT 93.065 61.700 93.735 63.045 ;
        RECT 70.800 40.250 71.800 61.550 ;
        RECT 92.100 61.400 93.750 61.700 ;
        RECT 73.400 61.370 93.750 61.400 ;
        RECT 73.390 61.000 93.750 61.370 ;
        RECT 73.390 57.740 74.390 61.000 ;
        RECT 75.330 60.350 90.430 60.750 ;
        RECT 75.330 59.600 75.730 60.350 ;
        RECT 90.030 60.200 90.430 60.350 ;
        RECT 76.030 59.750 78.580 60.200 ;
        RECT 78.830 59.750 81.330 60.200 ;
        RECT 81.630 59.750 84.180 60.200 ;
        RECT 84.430 59.750 86.930 60.200 ;
        RECT 87.230 59.750 89.780 60.200 ;
        RECT 90.030 59.700 96.650 60.200 ;
        RECT 90.030 59.600 90.430 59.700 ;
        RECT 75.330 59.200 90.430 59.600 ;
        RECT 75.330 58.550 90.430 58.950 ;
        RECT 75.450 58.010 75.820 58.550 ;
        RECT 76.080 58.000 87.830 58.400 ;
        RECT 87.380 57.860 87.730 58.000 ;
        RECT 73.390 56.740 74.400 57.740 ;
        RECT 87.380 57.500 87.740 57.860 ;
        RECT 73.400 47.360 74.400 56.740 ;
        RECT 89.140 51.950 90.430 58.550 ;
        RECT 96.160 58.100 96.640 59.700 ;
        RECT 73.400 46.660 76.550 47.360 ;
        RECT 73.400 46.360 89.410 46.660 ;
        RECT 79.910 46.020 85.530 46.190 ;
        RECT 73.320 45.300 76.550 45.630 ;
        RECT 73.320 44.970 76.960 45.300 ;
        RECT 77.110 45.240 77.560 45.470 ;
        RECT 73.320 44.630 76.550 44.970 ;
        RECT 77.110 44.800 77.560 45.030 ;
        RECT 77.840 44.970 78.260 45.300 ;
        RECT 78.420 45.240 78.870 45.470 ;
        RECT 79.910 45.370 80.080 46.020 ;
        RECT 82.330 45.810 82.690 45.880 ;
        RECT 80.700 45.540 81.030 45.810 ;
        RECT 81.620 45.550 82.690 45.810 ;
        RECT 77.170 44.220 77.500 44.800 ;
        RECT 77.110 44.190 77.560 44.220 ;
        RECT 77.840 44.190 78.020 44.970 ;
        RECT 78.420 44.800 78.870 45.030 ;
        RECT 79.440 44.920 79.670 45.370 ;
        RECT 79.880 44.920 80.110 45.370 ;
        RECT 80.530 44.920 80.760 45.370 ;
        RECT 80.970 44.920 81.200 45.370 ;
        RECT 81.620 44.920 81.850 45.550 ;
        RECT 82.490 45.370 82.690 45.550 ;
        RECT 82.970 45.540 83.310 46.020 ;
        RECT 83.970 45.780 84.300 45.810 ;
        RECT 84.470 45.780 84.830 45.880 ;
        RECT 83.970 45.600 84.830 45.780 ;
        RECT 83.970 45.540 84.300 45.600 ;
        RECT 84.470 45.520 84.830 45.600 ;
        RECT 85.360 45.370 85.530 46.020 ;
        RECT 82.060 44.920 82.290 45.370 ;
        RECT 82.490 44.920 82.940 45.370 ;
        RECT 83.150 44.920 83.380 45.370 ;
        RECT 83.800 44.920 84.030 45.370 ;
        RECT 84.240 44.920 84.470 45.370 ;
        RECT 84.890 44.920 85.120 45.370 ;
        RECT 85.330 44.920 85.560 45.370 ;
        RECT 85.980 44.920 86.210 45.370 ;
        RECT 86.420 44.920 86.650 45.370 ;
        RECT 87.160 45.240 87.610 45.470 ;
        RECT 87.820 45.280 88.170 45.300 ;
        RECT 87.160 44.800 87.610 45.030 ;
        RECT 87.815 44.990 88.170 45.280 ;
        RECT 88.480 45.240 88.930 45.470 ;
        RECT 89.400 45.300 90.500 45.700 ;
        RECT 87.820 44.970 88.170 44.990 ;
        RECT 78.480 44.590 78.810 44.800 ;
        RECT 79.440 44.590 79.680 44.670 ;
        RECT 80.520 44.590 80.760 44.670 ;
        RECT 82.240 44.620 82.600 44.690 ;
        RECT 78.480 44.420 80.760 44.590 ;
        RECT 78.480 44.220 78.810 44.420 ;
        RECT 79.440 44.340 79.680 44.420 ;
        RECT 80.520 44.340 80.760 44.420 ;
        RECT 82.030 44.390 82.600 44.620 ;
        RECT 82.240 44.330 82.600 44.390 ;
        RECT 82.840 44.330 83.380 44.690 ;
        RECT 85.270 44.630 85.550 44.650 ;
        RECT 86.390 44.630 86.650 44.660 ;
        RECT 87.220 44.630 87.550 44.800 ;
        RECT 84.200 44.400 87.550 44.630 ;
        RECT 84.200 44.390 85.550 44.400 ;
        RECT 85.270 44.360 85.550 44.390 ;
        RECT 86.390 44.370 86.650 44.400 ;
        RECT 87.220 44.220 87.550 44.400 ;
        RECT 76.670 43.720 76.970 44.050 ;
        RECT 77.110 44.020 78.020 44.190 ;
        RECT 77.110 43.990 77.560 44.020 ;
        RECT 77.110 43.550 77.560 43.780 ;
        RECT 75.500 42.230 76.550 42.310 ;
        RECT 77.110 42.230 77.550 43.550 ;
        RECT 77.840 43.520 78.020 44.020 ;
        RECT 78.420 43.990 78.870 44.220 ;
        RECT 78.420 43.550 78.870 43.780 ;
        RECT 77.840 43.190 78.280 43.520 ;
        RECT 78.420 42.230 78.870 43.340 ;
        RECT 79.440 42.230 79.670 44.110 ;
        RECT 79.880 43.650 80.110 44.100 ;
        RECT 80.530 43.650 80.760 44.100 ;
        RECT 80.970 43.650 81.200 44.100 ;
        RECT 81.620 43.650 81.850 44.100 ;
        RECT 82.060 43.650 82.290 44.100 ;
        RECT 82.710 43.650 82.940 44.100 ;
        RECT 83.150 43.650 83.380 44.100 ;
        RECT 83.800 43.650 84.030 44.100 ;
        RECT 84.240 43.650 84.470 44.100 ;
        RECT 84.890 43.650 85.120 44.100 ;
        RECT 85.330 43.650 85.560 44.100 ;
        RECT 85.980 43.650 86.210 44.100 ;
        RECT 86.420 43.650 86.650 44.100 ;
        RECT 87.160 43.990 87.610 44.220 ;
        RECT 88.000 44.190 88.170 44.970 ;
        RECT 88.480 44.800 88.930 45.030 ;
        RECT 89.080 44.970 90.500 45.300 ;
        RECT 88.540 44.220 88.870 44.800 ;
        RECT 89.400 44.550 90.500 44.970 ;
        RECT 88.480 44.190 88.930 44.220 ;
        RECT 88.000 44.020 88.930 44.190 ;
        RECT 80.700 43.180 81.030 43.510 ;
        RECT 81.880 43.440 82.220 43.500 ;
        RECT 86.010 43.440 86.180 43.650 ;
        RECT 87.160 43.550 87.610 43.780 ;
        RECT 88.000 43.520 88.170 44.020 ;
        RECT 88.480 43.990 88.930 44.020 ;
        RECT 81.880 43.260 86.180 43.440 ;
        RECT 81.880 43.190 82.220 43.260 ;
        RECT 79.850 42.670 80.140 43.090 ;
        RECT 79.910 42.230 80.080 42.670 ;
        RECT 80.750 42.540 81.110 42.900 ;
        RECT 81.470 42.880 81.700 43.140 ;
        RECT 86.450 43.110 86.620 43.140 ;
        RECT 85.330 43.080 85.560 43.110 ;
        RECT 85.300 42.900 85.590 43.080 ;
        RECT 85.330 42.880 85.560 42.900 ;
        RECT 81.500 42.230 81.670 42.880 ;
        RECT 85.360 42.230 85.530 42.880 ;
        RECT 85.950 42.680 86.240 43.100 ;
        RECT 86.420 42.880 86.650 43.110 ;
        RECT 86.010 42.230 86.180 42.680 ;
        RECT 86.450 42.230 86.620 42.880 ;
        RECT 87.160 42.230 87.610 43.340 ;
        RECT 87.790 43.190 88.170 43.520 ;
        RECT 88.480 42.230 88.930 43.780 ;
        RECT 89.070 43.720 89.370 44.050 ;
        RECT 75.500 41.930 89.410 42.230 ;
        RECT 75.500 41.230 76.550 41.930 ;
        RECT 81.410 40.250 82.410 41.750 ;
        RECT 70.800 39.250 82.410 40.250 ;
        RECT 83.030 40.250 84.030 41.740 ;
        RECT 91.510 40.250 92.510 57.860 ;
        RECT 95.700 56.850 97.000 58.100 ;
        RECT 83.030 39.250 92.510 40.250 ;
        RECT 80.550 31.750 82.100 39.250 ;
        RECT 85.000 36.500 86.400 39.250 ;
        RECT 85.000 34.850 86.800 36.500 ;
        RECT 73.320 27.550 74.380 28.550 ;
        RECT 101.770 27.550 102.830 28.550 ;
        RECT 73.350 7.800 74.350 27.550 ;
        RECT 101.800 10.220 102.800 27.550 ;
        RECT 109.150 25.400 115.950 25.650 ;
        RECT 128.050 25.550 147.400 25.950 ;
        RECT 109.150 25.000 143.150 25.400 ;
        RECT 109.150 24.800 115.950 25.000 ;
        RECT 128.050 24.350 143.150 24.750 ;
        RECT 128.050 23.600 128.450 24.350 ;
        RECT 142.750 24.200 143.150 24.350 ;
        RECT 143.900 24.200 144.650 24.300 ;
        RECT 128.750 23.750 131.300 24.200 ;
        RECT 131.550 23.750 134.050 24.200 ;
        RECT 134.350 23.750 136.900 24.200 ;
        RECT 137.150 23.750 139.650 24.200 ;
        RECT 139.950 23.750 142.500 24.200 ;
        RECT 142.750 23.700 144.650 24.200 ;
        RECT 142.750 23.600 143.150 23.700 ;
        RECT 128.050 23.200 143.150 23.600 ;
        RECT 143.900 23.550 144.650 23.700 ;
        RECT 125.650 22.400 126.700 22.600 ;
        RECT 128.050 22.550 143.150 22.950 ;
        RECT 125.650 22.000 140.550 22.400 ;
        RECT 125.650 21.900 126.700 22.000 ;
        RECT 141.750 15.950 143.150 22.550 ;
        RECT 146.550 22.200 147.400 25.550 ;
        RECT 73.350 6.800 139.200 7.800 ;
        RECT 138.200 5.450 139.200 6.800 ;
        RECT 137.750 3.550 139.650 5.450 ;
      LAYER met2 ;
        RECT 0.250 62.450 62.200 64.100 ;
        RECT 76.530 59.750 78.030 60.200 ;
        RECT 82.130 59.750 83.630 60.200 ;
        RECT 87.730 59.750 89.230 60.200 ;
        RECT 75.450 57.350 75.820 58.370 ;
        RECT 87.380 57.500 92.510 57.860 ;
        RECT 73.350 27.520 74.350 45.660 ;
        RECT 75.450 41.240 76.540 57.350 ;
        RECT 89.140 51.950 90.430 57.050 ;
        RECT 95.700 56.850 97.000 58.100 ;
        RECT 80.170 46.330 80.530 46.690 ;
        RECT 82.330 46.330 82.690 46.690 ;
        RECT 80.270 42.800 80.440 46.330 ;
        RECT 82.430 45.880 82.600 46.330 ;
        RECT 82.330 45.520 82.690 45.880 ;
        RECT 84.470 45.520 84.830 45.880 ;
        RECT 89.400 45.630 90.500 45.700 ;
        RECT 82.240 44.330 82.600 44.690 ;
        RECT 82.840 44.330 83.200 44.690 ;
        RECT 80.750 42.800 81.110 42.900 ;
        RECT 80.270 42.630 81.110 42.800 ;
        RECT 80.750 42.540 81.110 42.630 ;
        RECT 82.240 41.750 82.410 44.330 ;
        RECT 82.050 41.390 82.410 41.750 ;
        RECT 83.030 41.740 83.200 44.330 ;
        RECT 84.560 42.260 84.730 45.520 ;
        RECT 89.400 44.630 102.800 45.630 ;
        RECT 89.400 44.550 90.500 44.630 ;
        RECT 84.460 41.900 84.820 42.260 ;
        RECT 83.030 41.380 83.390 41.740 ;
        RECT 85.000 34.850 86.800 36.500 ;
        RECT 80.550 31.750 82.100 33.350 ;
        RECT 101.800 27.520 102.800 44.630 ;
        RECT 0.700 23.950 116.150 25.950 ;
        RECT 129.250 23.750 130.750 24.200 ;
        RECT 134.850 23.750 136.350 24.200 ;
        RECT 140.450 23.750 141.950 24.200 ;
        RECT 143.900 23.550 157.450 24.350 ;
        RECT 125.650 21.900 126.700 22.600 ;
        RECT 146.450 22.200 147.500 23.100 ;
        RECT 141.850 18.850 143.150 21.050 ;
        RECT 48.550 15.950 143.150 18.850 ;
        RECT 101.770 10.250 102.830 11.250 ;
        RECT 101.800 5.050 102.800 10.250 ;
        RECT 112.050 5.050 126.650 5.250 ;
        RECT 137.750 5.150 139.650 5.450 ;
        RECT 101.800 4.150 126.650 5.050 ;
        RECT 101.800 4.050 114.950 4.150 ;
        RECT 133.950 4.100 147.750 5.150 ;
        RECT 137.750 3.550 139.650 4.100 ;
      LAYER met3 ;
        RECT 0.400 62.450 3.050 64.100 ;
        RECT 71.530 62.650 81.980 73.100 ;
        RECT 83.580 62.700 94.030 73.150 ;
        RECT 76.530 59.750 78.030 62.650 ;
        RECT 82.130 57.250 83.630 60.200 ;
        RECT 87.730 59.750 89.230 62.700 ;
        RECT 76.930 46.850 87.330 57.250 ;
        RECT 89.140 51.950 90.430 57.050 ;
        RECT 85.000 34.850 86.800 36.500 ;
        RECT 89.650 34.875 91.700 35.100 ;
        RECT 95.475 34.875 97.125 58.325 ;
        RECT 80.550 31.750 82.100 33.350 ;
        RECT 89.650 33.225 97.125 34.875 ;
        RECT 0.700 23.950 2.700 25.950 ;
        RECT 48.550 15.950 51.000 18.850 ;
        RECT 89.650 11.400 91.300 33.225 ;
        RECT 124.250 26.650 134.700 37.100 ;
        RECT 136.300 26.700 146.750 37.150 ;
        RECT 129.250 23.750 130.750 26.650 ;
        RECT 125.700 22.600 126.550 22.800 ;
        RECT 125.650 21.900 126.700 22.600 ;
        RECT 112.200 2.350 113.300 5.500 ;
        RECT 125.700 4.150 126.550 21.900 ;
        RECT 134.850 21.250 136.350 24.200 ;
        RECT 140.450 23.750 141.950 26.700 ;
        RECT 129.650 10.850 140.050 21.250 ;
        RECT 141.750 15.950 143.150 21.050 ;
        RECT 112.100 1.450 113.350 2.350 ;
        RECT 134.200 2.200 135.300 5.300 ;
        RECT 146.550 5.150 147.400 23.100 ;
        RECT 146.500 4.100 147.600 5.150 ;
        RECT 134.200 1.450 135.400 2.200 ;
        RECT 156.300 1.450 157.300 24.450 ;
      LAYER met4 ;
        RECT 3.800 224.100 59.740 224.760 ;
        RECT 49.000 220.760 50.500 224.100 ;
        RECT 71.880 67.500 76.630 67.550 ;
        RECT 0.400 62.450 1.000 64.100 ;
        RECT 2.500 62.450 3.050 64.100 ;
        RECT 71.880 63.000 93.780 67.500 ;
        RECT 71.880 62.950 76.630 63.000 ;
        RECT 81.980 57.050 86.980 63.000 ;
        RECT 81.930 54.000 90.430 57.050 ;
        RECT 50.500 52.550 90.430 54.000 ;
        RECT 81.930 51.950 90.430 52.550 ;
        RECT 81.930 51.900 87.130 51.950 ;
        RECT 85.000 34.850 86.800 36.500 ;
        RECT 80.550 31.750 82.100 33.350 ;
        RECT 0.700 23.950 1.000 25.950 ;
        RECT 2.500 23.950 2.700 25.950 ;
        RECT 81.025 21.125 82.075 31.750 ;
        RECT 62.075 20.075 82.075 21.125 ;
        RECT 48.550 15.950 49.000 18.850 ;
        RECT 50.500 15.950 51.000 18.850 ;
        RECT 62.075 2.050 63.125 20.075 ;
        RECT 67.975 13.520 69.025 13.525 ;
        RECT 85.220 13.520 86.270 34.850 ;
        RECT 124.600 31.500 129.350 31.550 ;
        RECT 124.600 27.000 146.500 31.500 ;
        RECT 124.600 26.950 129.350 27.000 ;
        RECT 134.700 21.050 139.700 27.000 ;
        RECT 134.650 15.950 143.150 21.050 ;
        RECT 134.650 15.900 139.850 15.950 ;
        RECT 67.975 12.485 86.270 13.520 ;
        RECT 67.975 2.050 69.025 12.485 ;
        RECT 85.220 12.475 86.270 12.485 ;
        RECT 90.005 2.050 91.045 14.470 ;
        RECT 45.750 1.000 63.175 2.050 ;
        RECT 67.900 1.000 69.200 2.050 ;
        RECT 90.000 1.000 91.300 2.050 ;
        RECT 112.100 1.450 113.350 2.350 ;
        RECT 134.200 1.450 135.350 2.200 ;
        RECT 156.300 1.450 157.450 2.300 ;
        RECT 112.250 1.000 113.150 1.450 ;
        RECT 134.330 1.000 135.230 1.450 ;
        RECT 156.410 1.000 157.310 1.450 ;
  END
END tt_um_nurirfansyah_alits02
END LIBRARY

